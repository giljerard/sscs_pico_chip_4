magic
tech sky130A
magscale 1 2
timestamp 1637083665
<< poly >>
rect -285 912 285 928
rect -285 878 -269 912
rect 269 878 285 912
rect -285 855 285 878
rect -285 -878 285 -855
rect -285 -912 -269 -878
rect 269 -912 285 -878
rect -285 -928 285 -912
<< polycont >>
rect -269 878 269 912
rect -269 -912 269 -878
<< npolyres >>
rect -285 -855 285 855
<< locali >>
rect -285 878 -269 912
rect 269 878 285 912
rect -285 -912 -269 -878
rect 269 -912 285 -878
<< viali >>
rect -269 878 269 912
rect -269 872 269 878
rect -269 -878 269 -872
rect -269 -912 269 -878
<< metal1 >>
rect -281 912 281 918
rect -281 872 -269 912
rect 269 872 281 912
rect -281 866 281 872
rect -281 -872 281 -866
rect -281 -912 -269 -872
rect 269 -912 281 -872
rect -281 -918 281 -912
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string parameters w 2.85 l 8.55 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 144.6 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
