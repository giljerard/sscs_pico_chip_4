magic
tech sky130A
magscale 1 2
timestamp 1636523469
<< nwell >>
rect 6634 2516 8002 8010
<< pwell >>
rect 4308 2542 5666 8036
<< pmoslvt >>
rect 6854 7614 7854 7814
rect 6854 7356 7854 7556
rect 6854 7098 7854 7298
rect 6854 6840 7854 7040
rect 6854 6582 7854 6782
rect 6854 6324 7854 6524
rect 6854 6066 7854 6266
rect 6854 5808 7854 6008
rect 6854 5550 7854 5750
rect 6854 5292 7854 5492
rect 6854 5034 7854 5234
rect 6854 4776 7854 4976
rect 6854 4518 7854 4718
rect 6854 4260 7854 4460
rect 6854 4002 7854 4202
rect 6854 3744 7854 3944
rect 6854 3486 7854 3686
rect 6854 3228 7854 3428
rect 6854 2970 7854 3170
rect 6854 2712 7854 2912
<< nmoslvt >>
rect 4456 7640 5456 7840
rect 4456 7382 5456 7582
rect 4456 7124 5456 7324
rect 4456 6866 5456 7066
rect 4456 6608 5456 6808
rect 4456 6350 5456 6550
rect 4456 6092 5456 6292
rect 4456 5834 5456 6034
rect 4456 5576 5456 5776
rect 4456 5318 5456 5518
rect 4456 5060 5456 5260
rect 4456 4802 5456 5002
rect 4456 4544 5456 4744
rect 4456 4286 5456 4486
rect 4456 4028 5456 4228
rect 4456 3770 5456 3970
rect 4456 3512 5456 3712
rect 4456 3254 5456 3454
rect 4456 2996 5456 3196
rect 4456 2738 5456 2938
<< ndiff >>
rect 4456 7886 5456 7898
rect 4456 7852 4468 7886
rect 5444 7852 5456 7886
rect 4456 7840 5456 7852
rect 4456 7628 5456 7640
rect 4456 7594 4468 7628
rect 5444 7594 5456 7628
rect 4456 7582 5456 7594
rect 4456 7370 5456 7382
rect 4456 7336 4468 7370
rect 5444 7336 5456 7370
rect 4456 7324 5456 7336
rect 4456 7112 5456 7124
rect 4456 7078 4468 7112
rect 5444 7078 5456 7112
rect 4456 7066 5456 7078
rect 4456 6854 5456 6866
rect 4456 6820 4468 6854
rect 5444 6820 5456 6854
rect 4456 6808 5456 6820
rect 4456 6596 5456 6608
rect 4456 6562 4468 6596
rect 5444 6562 5456 6596
rect 4456 6550 5456 6562
rect 4456 6338 5456 6350
rect 4456 6304 4468 6338
rect 5444 6304 5456 6338
rect 4456 6292 5456 6304
rect 4456 6080 5456 6092
rect 4456 6046 4468 6080
rect 5444 6046 5456 6080
rect 4456 6034 5456 6046
rect 4456 5822 5456 5834
rect 4456 5788 4468 5822
rect 5444 5788 5456 5822
rect 4456 5776 5456 5788
rect 4456 5564 5456 5576
rect 4456 5530 4468 5564
rect 5444 5530 5456 5564
rect 4456 5518 5456 5530
rect 4456 5306 5456 5318
rect 4456 5272 4468 5306
rect 5444 5272 5456 5306
rect 4456 5260 5456 5272
rect 4456 5048 5456 5060
rect 4456 5014 4468 5048
rect 5444 5014 5456 5048
rect 4456 5002 5456 5014
rect 4456 4790 5456 4802
rect 4456 4756 4468 4790
rect 5444 4756 5456 4790
rect 4456 4744 5456 4756
rect 4456 4532 5456 4544
rect 4456 4498 4468 4532
rect 5444 4498 5456 4532
rect 4456 4486 5456 4498
rect 4456 4274 5456 4286
rect 4456 4240 4468 4274
rect 5444 4240 5456 4274
rect 4456 4228 5456 4240
rect 4456 4016 5456 4028
rect 4456 3982 4468 4016
rect 5444 3982 5456 4016
rect 4456 3970 5456 3982
rect 4456 3758 5456 3770
rect 4456 3724 4468 3758
rect 5444 3724 5456 3758
rect 4456 3712 5456 3724
rect 4456 3500 5456 3512
rect 4456 3466 4468 3500
rect 5444 3466 5456 3500
rect 4456 3454 5456 3466
rect 4456 3242 5456 3254
rect 4456 3208 4468 3242
rect 5444 3208 5456 3242
rect 4456 3196 5456 3208
rect 4456 2984 5456 2996
rect 4456 2950 4468 2984
rect 5444 2950 5456 2984
rect 4456 2938 5456 2950
rect 4456 2726 5456 2738
rect 4456 2692 4468 2726
rect 5444 2692 5456 2726
rect 4456 2680 5456 2692
<< pdiff >>
rect 6854 7860 7854 7872
rect 6854 7826 6866 7860
rect 7842 7826 7854 7860
rect 6854 7814 7854 7826
rect 6854 7602 7854 7614
rect 6854 7568 6866 7602
rect 7842 7568 7854 7602
rect 6854 7556 7854 7568
rect 6854 7344 7854 7356
rect 6854 7310 6866 7344
rect 7842 7310 7854 7344
rect 6854 7298 7854 7310
rect 6854 7086 7854 7098
rect 6854 7052 6866 7086
rect 7842 7052 7854 7086
rect 6854 7040 7854 7052
rect 6854 6828 7854 6840
rect 6854 6794 6866 6828
rect 7842 6794 7854 6828
rect 6854 6782 7854 6794
rect 6854 6570 7854 6582
rect 6854 6536 6866 6570
rect 7842 6536 7854 6570
rect 6854 6524 7854 6536
rect 6854 6312 7854 6324
rect 6854 6278 6866 6312
rect 7842 6278 7854 6312
rect 6854 6266 7854 6278
rect 6854 6054 7854 6066
rect 6854 6020 6866 6054
rect 7842 6020 7854 6054
rect 6854 6008 7854 6020
rect 6854 5796 7854 5808
rect 6854 5762 6866 5796
rect 7842 5762 7854 5796
rect 6854 5750 7854 5762
rect 6854 5538 7854 5550
rect 6854 5504 6866 5538
rect 7842 5504 7854 5538
rect 6854 5492 7854 5504
rect 6854 5280 7854 5292
rect 6854 5246 6866 5280
rect 7842 5246 7854 5280
rect 6854 5234 7854 5246
rect 6854 5022 7854 5034
rect 6854 4988 6866 5022
rect 7842 4988 7854 5022
rect 6854 4976 7854 4988
rect 6854 4764 7854 4776
rect 6854 4730 6866 4764
rect 7842 4730 7854 4764
rect 6854 4718 7854 4730
rect 6854 4506 7854 4518
rect 6854 4472 6866 4506
rect 7842 4472 7854 4506
rect 6854 4460 7854 4472
rect 6854 4248 7854 4260
rect 6854 4214 6866 4248
rect 7842 4214 7854 4248
rect 6854 4202 7854 4214
rect 6854 3990 7854 4002
rect 6854 3956 6866 3990
rect 7842 3956 7854 3990
rect 6854 3944 7854 3956
rect 6854 3732 7854 3744
rect 6854 3698 6866 3732
rect 7842 3698 7854 3732
rect 6854 3686 7854 3698
rect 6854 3474 7854 3486
rect 6854 3440 6866 3474
rect 7842 3440 7854 3474
rect 6854 3428 7854 3440
rect 6854 3216 7854 3228
rect 6854 3182 6866 3216
rect 7842 3182 7854 3216
rect 6854 3170 7854 3182
rect 6854 2958 7854 2970
rect 6854 2924 6866 2958
rect 7842 2924 7854 2958
rect 6854 2912 7854 2924
rect 6854 2700 7854 2712
rect 6854 2666 6866 2700
rect 7842 2666 7854 2700
rect 6854 2654 7854 2666
<< ndiffc >>
rect 4468 7852 5444 7886
rect 4468 7594 5444 7628
rect 4468 7336 5444 7370
rect 4468 7078 5444 7112
rect 4468 6820 5444 6854
rect 4468 6562 5444 6596
rect 4468 6304 5444 6338
rect 4468 6046 5444 6080
rect 4468 5788 5444 5822
rect 4468 5530 5444 5564
rect 4468 5272 5444 5306
rect 4468 5014 5444 5048
rect 4468 4756 5444 4790
rect 4468 4498 5444 4532
rect 4468 4240 5444 4274
rect 4468 3982 5444 4016
rect 4468 3724 5444 3758
rect 4468 3466 5444 3500
rect 4468 3208 5444 3242
rect 4468 2950 5444 2984
rect 4468 2692 5444 2726
<< pdiffc >>
rect 6866 7826 7842 7860
rect 6866 7568 7842 7602
rect 6866 7310 7842 7344
rect 6866 7052 7842 7086
rect 6866 6794 7842 6828
rect 6866 6536 7842 6570
rect 6866 6278 7842 6312
rect 6866 6020 7842 6054
rect 6866 5762 7842 5796
rect 6866 5504 7842 5538
rect 6866 5246 7842 5280
rect 6866 4988 7842 5022
rect 6866 4730 7842 4764
rect 6866 4472 7842 4506
rect 6866 4214 7842 4248
rect 6866 3956 7842 3990
rect 6866 3698 7842 3732
rect 6866 3440 7842 3474
rect 6866 3182 7842 3216
rect 6866 2924 7842 2958
rect 6866 2666 7842 2700
<< psubdiff >>
rect 4344 7966 4440 8000
rect 5534 7966 5630 8000
rect 4344 7904 4378 7966
rect 5596 7904 5630 7966
rect 4344 2612 4378 2674
rect 5596 2612 5630 2674
rect 4344 2578 4440 2612
rect 5534 2578 5630 2612
<< nsubdiff >>
rect 6670 7940 6767 7974
rect 7869 7940 7966 7974
rect 6670 7878 6704 7940
rect 7932 7878 7966 7940
rect 6670 2586 6704 2648
rect 7932 2586 7966 2648
rect 6670 2552 6767 2586
rect 7869 2552 7966 2586
<< psubdiffcont >>
rect 4440 7966 5534 8000
rect 4344 2674 4378 7904
rect 5596 2674 5630 7904
rect 4440 2578 5534 2612
<< nsubdiffcont >>
rect 6767 7940 7869 7974
rect 6670 2648 6704 7878
rect 7932 2648 7966 7878
rect 6767 2552 7869 2586
<< poly >>
rect 4430 7640 4456 7840
rect 5456 7824 5544 7840
rect 5456 7656 5494 7824
rect 5528 7656 5544 7824
rect 5456 7640 5544 7656
rect 4430 7382 4456 7582
rect 5456 7566 5544 7582
rect 5456 7398 5494 7566
rect 5528 7398 5544 7566
rect 5456 7382 5544 7398
rect 4430 7124 4456 7324
rect 5456 7308 5544 7324
rect 5456 7140 5494 7308
rect 5528 7140 5544 7308
rect 5456 7124 5544 7140
rect 4430 6866 4456 7066
rect 5456 7050 5544 7066
rect 5456 6882 5494 7050
rect 5528 6882 5544 7050
rect 5456 6866 5544 6882
rect 4430 6608 4456 6808
rect 5456 6792 5544 6808
rect 5456 6624 5494 6792
rect 5528 6624 5544 6792
rect 5456 6608 5544 6624
rect 4430 6350 4456 6550
rect 5456 6534 5544 6550
rect 5456 6366 5494 6534
rect 5528 6366 5544 6534
rect 5456 6350 5544 6366
rect 4430 6092 4456 6292
rect 5456 6276 5544 6292
rect 5456 6108 5494 6276
rect 5528 6108 5544 6276
rect 5456 6092 5544 6108
rect 4430 5834 4456 6034
rect 5456 6018 5544 6034
rect 5456 5850 5494 6018
rect 5528 5850 5544 6018
rect 5456 5834 5544 5850
rect 4430 5576 4456 5776
rect 5456 5760 5544 5776
rect 5456 5592 5494 5760
rect 5528 5592 5544 5760
rect 5456 5576 5544 5592
rect 4430 5318 4456 5518
rect 5456 5502 5544 5518
rect 5456 5334 5494 5502
rect 5528 5334 5544 5502
rect 5456 5318 5544 5334
rect 4430 5060 4456 5260
rect 5456 5244 5544 5260
rect 5456 5076 5494 5244
rect 5528 5076 5544 5244
rect 5456 5060 5544 5076
rect 4430 4802 4456 5002
rect 5456 4986 5544 5002
rect 5456 4818 5494 4986
rect 5528 4818 5544 4986
rect 5456 4802 5544 4818
rect 4430 4544 4456 4744
rect 5456 4728 5544 4744
rect 5456 4560 5494 4728
rect 5528 4560 5544 4728
rect 5456 4544 5544 4560
rect 4430 4286 4456 4486
rect 5456 4470 5544 4486
rect 5456 4302 5494 4470
rect 5528 4302 5544 4470
rect 5456 4286 5544 4302
rect 4430 4028 4456 4228
rect 5456 4212 5544 4228
rect 5456 4044 5494 4212
rect 5528 4044 5544 4212
rect 5456 4028 5544 4044
rect 4430 3770 4456 3970
rect 5456 3954 5544 3970
rect 5456 3786 5494 3954
rect 5528 3786 5544 3954
rect 5456 3770 5544 3786
rect 4430 3512 4456 3712
rect 5456 3696 5544 3712
rect 5456 3528 5494 3696
rect 5528 3528 5544 3696
rect 5456 3512 5544 3528
rect 4430 3254 4456 3454
rect 5456 3438 5544 3454
rect 5456 3270 5494 3438
rect 5528 3270 5544 3438
rect 5456 3254 5544 3270
rect 4430 2996 4456 3196
rect 5456 3180 5544 3196
rect 5456 3012 5494 3180
rect 5528 3012 5544 3180
rect 5456 2996 5544 3012
rect 4430 2738 4456 2938
rect 5456 2922 5544 2938
rect 5456 2754 5494 2922
rect 5528 2754 5544 2922
rect 5456 2738 5544 2754
rect 6757 7798 6854 7814
rect 6757 7630 6773 7798
rect 6807 7630 6854 7798
rect 6757 7614 6854 7630
rect 7854 7614 7880 7814
rect 6757 7540 6854 7556
rect 6757 7372 6773 7540
rect 6807 7372 6854 7540
rect 6757 7356 6854 7372
rect 7854 7356 7880 7556
rect 6757 7282 6854 7298
rect 6757 7114 6773 7282
rect 6807 7114 6854 7282
rect 6757 7098 6854 7114
rect 7854 7098 7880 7298
rect 6757 7024 6854 7040
rect 6757 6856 6773 7024
rect 6807 6856 6854 7024
rect 6757 6840 6854 6856
rect 7854 6840 7880 7040
rect 6757 6766 6854 6782
rect 6757 6598 6773 6766
rect 6807 6598 6854 6766
rect 6757 6582 6854 6598
rect 7854 6582 7880 6782
rect 6757 6508 6854 6524
rect 6757 6340 6773 6508
rect 6807 6340 6854 6508
rect 6757 6324 6854 6340
rect 7854 6324 7880 6524
rect 6757 6250 6854 6266
rect 6757 6082 6773 6250
rect 6807 6082 6854 6250
rect 6757 6066 6854 6082
rect 7854 6066 7880 6266
rect 6757 5992 6854 6008
rect 6757 5824 6773 5992
rect 6807 5824 6854 5992
rect 6757 5808 6854 5824
rect 7854 5808 7880 6008
rect 6757 5734 6854 5750
rect 6757 5566 6773 5734
rect 6807 5566 6854 5734
rect 6757 5550 6854 5566
rect 7854 5550 7880 5750
rect 6757 5476 6854 5492
rect 6757 5308 6773 5476
rect 6807 5308 6854 5476
rect 6757 5292 6854 5308
rect 7854 5292 7880 5492
rect 6757 5218 6854 5234
rect 6757 5050 6773 5218
rect 6807 5050 6854 5218
rect 6757 5034 6854 5050
rect 7854 5034 7880 5234
rect 6757 4960 6854 4976
rect 6757 4792 6773 4960
rect 6807 4792 6854 4960
rect 6757 4776 6854 4792
rect 7854 4776 7880 4976
rect 6757 4702 6854 4718
rect 6757 4534 6773 4702
rect 6807 4534 6854 4702
rect 6757 4518 6854 4534
rect 7854 4518 7880 4718
rect 6757 4444 6854 4460
rect 6757 4276 6773 4444
rect 6807 4276 6854 4444
rect 6757 4260 6854 4276
rect 7854 4260 7880 4460
rect 6757 4186 6854 4202
rect 6757 4018 6773 4186
rect 6807 4018 6854 4186
rect 6757 4002 6854 4018
rect 7854 4002 7880 4202
rect 6757 3928 6854 3944
rect 6757 3760 6773 3928
rect 6807 3760 6854 3928
rect 6757 3744 6854 3760
rect 7854 3744 7880 3944
rect 6757 3670 6854 3686
rect 6757 3502 6773 3670
rect 6807 3502 6854 3670
rect 6757 3486 6854 3502
rect 7854 3486 7880 3686
rect 6757 3412 6854 3428
rect 6757 3244 6773 3412
rect 6807 3244 6854 3412
rect 6757 3228 6854 3244
rect 7854 3228 7880 3428
rect 6757 3154 6854 3170
rect 6757 2986 6773 3154
rect 6807 2986 6854 3154
rect 6757 2970 6854 2986
rect 7854 2970 7880 3170
rect 6757 2896 6854 2912
rect 6757 2728 6773 2896
rect 6807 2728 6854 2896
rect 6757 2712 6854 2728
rect 7854 2712 7880 2912
<< polycont >>
rect 5494 7656 5528 7824
rect 5494 7398 5528 7566
rect 5494 7140 5528 7308
rect 5494 6882 5528 7050
rect 5494 6624 5528 6792
rect 5494 6366 5528 6534
rect 5494 6108 5528 6276
rect 5494 5850 5528 6018
rect 5494 5592 5528 5760
rect 5494 5334 5528 5502
rect 5494 5076 5528 5244
rect 5494 4818 5528 4986
rect 5494 4560 5528 4728
rect 5494 4302 5528 4470
rect 5494 4044 5528 4212
rect 5494 3786 5528 3954
rect 5494 3528 5528 3696
rect 5494 3270 5528 3438
rect 5494 3012 5528 3180
rect 5494 2754 5528 2922
rect 6773 7630 6807 7798
rect 6773 7372 6807 7540
rect 6773 7114 6807 7282
rect 6773 6856 6807 7024
rect 6773 6598 6807 6766
rect 6773 6340 6807 6508
rect 6773 6082 6807 6250
rect 6773 5824 6807 5992
rect 6773 5566 6807 5734
rect 6773 5308 6807 5476
rect 6773 5050 6807 5218
rect 6773 4792 6807 4960
rect 6773 4534 6807 4702
rect 6773 4276 6807 4444
rect 6773 4018 6807 4186
rect 6773 3760 6807 3928
rect 6773 3502 6807 3670
rect 6773 3244 6807 3412
rect 6773 2986 6807 3154
rect 6773 2728 6807 2896
<< locali >>
rect 4344 7966 4440 8000
rect 5534 7966 5630 8000
rect 5596 7904 5630 7966
rect 4452 7852 4468 7886
rect 5444 7852 5460 7886
rect 5494 7824 5528 7888
rect 5494 7628 5528 7656
rect 4452 7594 4468 7628
rect 5444 7594 5528 7628
rect 5494 7566 5528 7594
rect 4452 7336 4468 7370
rect 5444 7336 5460 7370
rect 5494 7308 5528 7398
rect 5494 7112 5528 7140
rect 4452 7078 4468 7112
rect 5444 7078 5528 7112
rect 5494 7050 5528 7078
rect 4452 6820 4468 6854
rect 5444 6820 5460 6854
rect 5494 6792 5528 6882
rect 5494 6596 5528 6624
rect 4452 6562 4468 6596
rect 5444 6562 5528 6596
rect 5494 6534 5528 6562
rect 4452 6304 4468 6338
rect 5444 6304 5460 6338
rect 5494 6276 5528 6366
rect 5494 6080 5528 6108
rect 4452 6046 4468 6080
rect 5444 6046 5528 6080
rect 5494 6018 5528 6046
rect 4452 5788 4468 5822
rect 5444 5788 5460 5822
rect 5494 5760 5528 5850
rect 5494 5564 5528 5592
rect 4452 5530 4468 5564
rect 5444 5530 5528 5564
rect 5494 5502 5528 5530
rect 4452 5272 4468 5306
rect 5444 5272 5460 5306
rect 5494 5244 5528 5334
rect 5494 5048 5528 5076
rect 4452 5014 4468 5048
rect 5444 5014 5528 5048
rect 5494 4986 5528 5014
rect 4452 4756 4468 4790
rect 5444 4756 5460 4790
rect 5494 4728 5528 4818
rect 5494 4532 5528 4560
rect 4452 4498 4468 4532
rect 5444 4498 5528 4532
rect 5494 4470 5528 4498
rect 4452 4240 4468 4274
rect 5444 4240 5460 4274
rect 5494 4212 5528 4302
rect 5494 4016 5528 4044
rect 4452 3982 4468 4016
rect 5444 3982 5528 4016
rect 5494 3954 5528 3982
rect 4452 3724 4468 3758
rect 5444 3724 5460 3758
rect 5494 3696 5528 3786
rect 5494 3500 5528 3528
rect 4452 3466 4468 3500
rect 5444 3466 5528 3500
rect 5494 3438 5528 3466
rect 4452 3208 4468 3242
rect 5444 3208 5460 3242
rect 5494 3180 5528 3270
rect 5494 2984 5528 3012
rect 4452 2950 4468 2984
rect 5444 2950 5528 2984
rect 5494 2922 5528 2950
rect 4452 2692 4468 2726
rect 5444 2692 5460 2726
rect 5494 2691 5528 2754
rect 5596 2612 5630 2674
rect 4344 2578 4440 2612
rect 5534 2578 5630 2612
rect 6670 7940 6767 7974
rect 7869 7940 7966 7974
rect 6670 7878 6704 7940
rect 6773 7798 6807 7860
rect 6850 7826 6866 7860
rect 7842 7826 7858 7860
rect 6773 7602 6807 7630
rect 6773 7568 6866 7602
rect 7842 7568 7858 7602
rect 6773 7540 6807 7568
rect 6773 7282 6807 7372
rect 6850 7310 6866 7344
rect 7842 7310 7858 7344
rect 6773 7086 6807 7114
rect 6773 7052 6866 7086
rect 7842 7052 7858 7086
rect 6773 7024 6807 7052
rect 6773 6766 6807 6856
rect 6850 6794 6866 6828
rect 7842 6794 7858 6828
rect 6773 6570 6807 6598
rect 6773 6536 6866 6570
rect 7842 6536 7858 6570
rect 6773 6508 6807 6536
rect 6773 6250 6807 6340
rect 6850 6278 6866 6312
rect 7842 6278 7858 6312
rect 6773 6054 6807 6082
rect 6773 6020 6866 6054
rect 7842 6020 7858 6054
rect 6773 5992 6807 6020
rect 6773 5734 6807 5824
rect 6850 5762 6866 5796
rect 7842 5762 7858 5796
rect 6773 5538 6807 5566
rect 6773 5504 6866 5538
rect 7842 5504 7858 5538
rect 6773 5476 6807 5504
rect 6773 5218 6807 5308
rect 6850 5246 6866 5280
rect 7842 5246 7858 5280
rect 6773 5022 6807 5050
rect 6773 4988 6866 5022
rect 7842 4988 7858 5022
rect 6773 4960 6807 4988
rect 6773 4702 6807 4792
rect 6850 4730 6866 4764
rect 7842 4730 7858 4764
rect 6773 4506 6807 4534
rect 6773 4472 6866 4506
rect 7842 4472 7858 4506
rect 6773 4444 6807 4472
rect 6773 4186 6807 4276
rect 6850 4214 6866 4248
rect 7842 4214 7858 4248
rect 6773 3990 6807 4018
rect 6773 3956 6866 3990
rect 7842 3956 7858 3990
rect 6773 3928 6807 3956
rect 6773 3670 6807 3760
rect 6850 3698 6866 3732
rect 7842 3698 7858 3732
rect 6773 3474 6807 3502
rect 6773 3440 6866 3474
rect 7842 3440 7858 3474
rect 6773 3412 6807 3440
rect 6773 3154 6807 3244
rect 6850 3182 6866 3216
rect 7842 3182 7858 3216
rect 6773 2958 6807 2986
rect 6773 2924 6866 2958
rect 7842 2924 7858 2958
rect 6773 2896 6807 2924
rect 6773 2666 6807 2728
rect 6850 2666 6866 2700
rect 7842 2666 7858 2700
rect 6670 2586 6704 2648
rect 6670 2552 6767 2586
rect 7869 2552 7966 2586
<< viali >>
rect 4500 7966 5474 8000
rect 4344 7904 4378 7966
rect 4344 2674 4378 7904
rect 4468 7852 5444 7886
rect 5494 7698 5528 7782
rect 4468 7594 5444 7628
rect 5494 7440 5528 7524
rect 4468 7336 5444 7370
rect 5494 7182 5528 7266
rect 4468 7078 5444 7112
rect 5494 6924 5528 7008
rect 4468 6820 5444 6854
rect 5494 6666 5528 6750
rect 4468 6562 5444 6596
rect 5494 6408 5528 6492
rect 4468 6304 5444 6338
rect 5494 6150 5528 6234
rect 4468 6046 5444 6080
rect 5494 5892 5528 5976
rect 4468 5788 5444 5822
rect 5494 5634 5528 5718
rect 4468 5530 5444 5564
rect 5494 5376 5528 5460
rect 4468 5272 5444 5306
rect 5494 5118 5528 5202
rect 4468 5014 5444 5048
rect 5494 4860 5528 4944
rect 4468 4756 5444 4790
rect 5494 4602 5528 4686
rect 4468 4498 5444 4532
rect 5494 4344 5528 4428
rect 4468 4240 5444 4274
rect 5494 4086 5528 4170
rect 4468 3982 5444 4016
rect 5494 3828 5528 3912
rect 4468 3724 5444 3758
rect 5494 3570 5528 3654
rect 4468 3466 5444 3500
rect 5494 3312 5528 3396
rect 4468 3208 5444 3242
rect 5494 3054 5528 3138
rect 4468 2950 5444 2984
rect 5494 2796 5528 2880
rect 4468 2692 5444 2726
rect 4344 2612 4378 2674
rect 4500 2578 5474 2612
rect 6827 7940 7809 7974
rect 7932 7878 7966 7940
rect 6866 7826 7842 7860
rect 6773 7672 6807 7756
rect 6866 7568 7842 7602
rect 6773 7414 6807 7498
rect 6866 7310 7842 7344
rect 6773 7156 6807 7240
rect 6866 7052 7842 7086
rect 6773 6898 6807 6982
rect 6866 6794 7842 6828
rect 6773 6640 6807 6724
rect 6866 6536 7842 6570
rect 6773 6382 6807 6466
rect 6866 6278 7842 6312
rect 6773 6124 6807 6208
rect 6866 6020 7842 6054
rect 6773 5866 6807 5950
rect 6866 5762 7842 5796
rect 6773 5608 6807 5692
rect 6866 5504 7842 5538
rect 6773 5350 6807 5434
rect 6866 5246 7842 5280
rect 6773 5092 6807 5176
rect 6866 4988 7842 5022
rect 6773 4834 6807 4918
rect 6866 4730 7842 4764
rect 6773 4576 6807 4660
rect 6866 4472 7842 4506
rect 6773 4318 6807 4402
rect 6866 4214 7842 4248
rect 6773 4060 6807 4144
rect 6866 3956 7842 3990
rect 6773 3802 6807 3886
rect 6866 3698 7842 3732
rect 6773 3544 6807 3628
rect 6866 3440 7842 3474
rect 6773 3286 6807 3370
rect 6866 3182 7842 3216
rect 6773 3028 6807 3112
rect 6866 2924 7842 2958
rect 6773 2770 6807 2854
rect 6866 2666 7842 2700
rect 7932 2648 7966 7878
rect 7932 2586 7966 2648
rect 6827 2552 7809 2586
<< metal1 >>
rect 4117 8000 5486 8006
rect 4117 7966 4500 8000
rect 5474 7966 5486 8000
rect 4117 2612 4344 7966
rect 4378 7960 5486 7966
rect 4378 7628 4418 7960
rect 5600 7892 5875 8036
rect 4456 7886 5875 7892
rect 4456 7852 4468 7886
rect 5444 7852 5875 7886
rect 4456 7846 5875 7852
rect 5488 7782 5534 7794
rect 5488 7698 5494 7782
rect 5528 7698 5534 7782
rect 5488 7686 5534 7698
rect 4456 7628 5456 7634
rect 4378 7594 4468 7628
rect 5444 7594 5456 7628
rect 4378 7112 4418 7594
rect 4456 7588 5456 7594
rect 5488 7524 5534 7536
rect 5488 7440 5494 7524
rect 5528 7440 5534 7524
rect 5488 7428 5534 7440
rect 5600 7376 5875 7846
rect 4456 7370 5875 7376
rect 4456 7336 4468 7370
rect 5444 7336 5875 7370
rect 4456 7330 5875 7336
rect 5488 7266 5534 7278
rect 5488 7182 5494 7266
rect 5528 7182 5534 7266
rect 5488 7170 5534 7182
rect 4456 7112 5456 7118
rect 4378 7078 4468 7112
rect 5444 7078 5456 7112
rect 4378 6596 4418 7078
rect 4456 7072 5456 7078
rect 5488 7008 5534 7020
rect 5488 6924 5494 7008
rect 5528 6924 5534 7008
rect 5488 6912 5534 6924
rect 5600 6860 5875 7330
rect 4456 6854 5875 6860
rect 4456 6820 4468 6854
rect 5444 6820 5875 6854
rect 4456 6814 5875 6820
rect 5488 6750 5534 6762
rect 5488 6666 5494 6750
rect 5528 6666 5534 6750
rect 5488 6654 5534 6666
rect 4456 6596 5456 6602
rect 4378 6562 4468 6596
rect 5444 6562 5456 6596
rect 4378 6080 4418 6562
rect 4456 6556 5456 6562
rect 5488 6492 5534 6504
rect 5488 6408 5494 6492
rect 5528 6408 5534 6492
rect 5488 6396 5534 6408
rect 5600 6344 5875 6814
rect 4456 6338 5875 6344
rect 4456 6304 4468 6338
rect 5444 6304 5875 6338
rect 4456 6298 5875 6304
rect 5488 6234 5534 6246
rect 5488 6150 5494 6234
rect 5528 6150 5534 6234
rect 5488 6138 5534 6150
rect 4456 6080 5456 6086
rect 4378 6046 4468 6080
rect 5444 6046 5456 6080
rect 4378 5564 4418 6046
rect 4456 6040 5456 6046
rect 5488 5976 5534 5988
rect 5488 5892 5494 5976
rect 5528 5892 5534 5976
rect 5488 5880 5534 5892
rect 5600 5828 5875 6298
rect 4456 5822 5875 5828
rect 4456 5788 4468 5822
rect 5444 5788 5875 5822
rect 4456 5782 5875 5788
rect 5488 5718 5534 5730
rect 5488 5634 5494 5718
rect 5528 5634 5534 5718
rect 5488 5622 5534 5634
rect 4456 5564 5456 5570
rect 4378 5530 4468 5564
rect 5444 5530 5456 5564
rect 4378 5048 4418 5530
rect 4456 5524 5456 5530
rect 5488 5460 5534 5472
rect 5488 5376 5494 5460
rect 5528 5376 5534 5460
rect 5488 5364 5534 5376
rect 5600 5312 5875 5782
rect 4456 5306 5875 5312
rect 4456 5272 4468 5306
rect 5444 5272 5875 5306
rect 4456 5266 5875 5272
rect 5488 5202 5534 5214
rect 5488 5118 5494 5202
rect 5528 5118 5534 5202
rect 5488 5106 5534 5118
rect 4456 5048 5456 5054
rect 4378 5014 4468 5048
rect 5444 5014 5456 5048
rect 4378 4532 4418 5014
rect 4456 5008 5456 5014
rect 5488 4944 5534 4956
rect 5488 4860 5494 4944
rect 5528 4860 5534 4944
rect 5488 4848 5534 4860
rect 5600 4796 5875 5266
rect 4456 4790 5875 4796
rect 4456 4756 4468 4790
rect 5444 4756 5875 4790
rect 4456 4750 5875 4756
rect 5488 4686 5534 4698
rect 5488 4602 5494 4686
rect 5528 4602 5534 4686
rect 5488 4590 5534 4602
rect 4456 4532 5456 4538
rect 4378 4498 4468 4532
rect 5444 4498 5456 4532
rect 4378 4016 4418 4498
rect 4456 4492 5456 4498
rect 5488 4428 5534 4440
rect 5488 4344 5494 4428
rect 5528 4344 5534 4428
rect 5488 4332 5534 4344
rect 5600 4280 5875 4750
rect 4456 4274 5875 4280
rect 4456 4240 4468 4274
rect 5444 4240 5875 4274
rect 4456 4234 5875 4240
rect 5488 4170 5534 4182
rect 5488 4086 5494 4170
rect 5528 4086 5534 4170
rect 5488 4074 5534 4086
rect 4456 4016 5456 4022
rect 4378 3982 4468 4016
rect 5444 3982 5456 4016
rect 4378 3500 4418 3982
rect 4456 3976 5456 3982
rect 5488 3912 5534 3924
rect 5488 3828 5494 3912
rect 5528 3828 5534 3912
rect 5488 3816 5534 3828
rect 5600 3764 5875 4234
rect 4456 3758 5875 3764
rect 4456 3724 4468 3758
rect 5444 3724 5875 3758
rect 4456 3718 5875 3724
rect 5488 3654 5534 3666
rect 5488 3570 5494 3654
rect 5528 3570 5534 3654
rect 5488 3558 5534 3570
rect 4456 3500 5456 3506
rect 4378 3466 4468 3500
rect 5444 3466 5456 3500
rect 4378 2984 4418 3466
rect 4456 3460 5456 3466
rect 5488 3396 5534 3408
rect 5488 3312 5494 3396
rect 5528 3312 5534 3396
rect 5488 3300 5534 3312
rect 5600 3248 5875 3718
rect 4456 3242 5875 3248
rect 4456 3208 4468 3242
rect 5444 3208 5875 3242
rect 4456 3202 5875 3208
rect 5488 3138 5534 3150
rect 5488 3054 5494 3138
rect 5528 3054 5534 3138
rect 5488 3042 5534 3054
rect 4456 2984 5456 2990
rect 4378 2950 4468 2984
rect 5444 2950 5456 2984
rect 4378 2618 4418 2950
rect 4456 2944 5456 2950
rect 5488 2880 5534 2892
rect 5488 2796 5494 2880
rect 5528 2796 5534 2880
rect 5488 2784 5534 2796
rect 5600 2732 5875 3202
rect 4456 2726 5875 2732
rect 4456 2692 4468 2726
rect 5444 2692 5875 2726
rect 4456 2686 5875 2692
rect 4378 2612 5486 2618
rect 4117 2578 4500 2612
rect 5474 2578 5486 2612
rect 4117 2572 5486 2578
rect 5600 2542 5875 2686
rect 6454 7866 6729 8010
rect 6815 7974 8227 7980
rect 6815 7940 6827 7974
rect 7809 7940 8227 7974
rect 6815 7934 7932 7940
rect 6454 7860 7854 7866
rect 6454 7826 6866 7860
rect 7842 7826 7854 7860
rect 6454 7820 7854 7826
rect 6454 7350 6729 7820
rect 6767 7756 6813 7768
rect 6767 7672 6773 7756
rect 6807 7672 6813 7756
rect 6767 7660 6813 7672
rect 7926 7608 7932 7934
rect 6854 7602 7932 7608
rect 6854 7568 6866 7602
rect 7842 7568 7932 7602
rect 6854 7562 7932 7568
rect 6767 7498 6813 7510
rect 6767 7414 6773 7498
rect 6807 7414 6813 7498
rect 6767 7402 6813 7414
rect 6454 7344 7854 7350
rect 6454 7310 6866 7344
rect 7842 7310 7854 7344
rect 6454 7304 7854 7310
rect 6454 6834 6729 7304
rect 6767 7240 6813 7252
rect 6767 7156 6773 7240
rect 6807 7156 6813 7240
rect 6767 7144 6813 7156
rect 7926 7092 7932 7562
rect 6854 7086 7932 7092
rect 6854 7052 6866 7086
rect 7842 7052 7932 7086
rect 6854 7046 7932 7052
rect 6767 6982 6813 6994
rect 6767 6898 6773 6982
rect 6807 6898 6813 6982
rect 6767 6886 6813 6898
rect 6454 6828 7854 6834
rect 6454 6794 6866 6828
rect 7842 6794 7854 6828
rect 6454 6788 7854 6794
rect 6454 6318 6729 6788
rect 6767 6724 6813 6736
rect 6767 6640 6773 6724
rect 6807 6640 6813 6724
rect 6767 6628 6813 6640
rect 7926 6576 7932 7046
rect 6854 6570 7932 6576
rect 6854 6536 6866 6570
rect 7842 6536 7932 6570
rect 6854 6530 7932 6536
rect 6767 6466 6813 6478
rect 6767 6382 6773 6466
rect 6807 6382 6813 6466
rect 6767 6370 6813 6382
rect 6454 6312 7854 6318
rect 6454 6278 6866 6312
rect 7842 6278 7854 6312
rect 6454 6272 7854 6278
rect 6454 5802 6729 6272
rect 6767 6208 6813 6220
rect 6767 6124 6773 6208
rect 6807 6124 6813 6208
rect 6767 6112 6813 6124
rect 7926 6060 7932 6530
rect 6854 6054 7932 6060
rect 6854 6020 6866 6054
rect 7842 6020 7932 6054
rect 6854 6014 7932 6020
rect 6767 5950 6813 5962
rect 6767 5866 6773 5950
rect 6807 5866 6813 5950
rect 6767 5854 6813 5866
rect 6454 5796 7854 5802
rect 6454 5762 6866 5796
rect 7842 5762 7854 5796
rect 6454 5756 7854 5762
rect 6454 5286 6729 5756
rect 6767 5692 6813 5704
rect 6767 5608 6773 5692
rect 6807 5608 6813 5692
rect 6767 5596 6813 5608
rect 7926 5544 7932 6014
rect 6854 5538 7932 5544
rect 6854 5504 6866 5538
rect 7842 5504 7932 5538
rect 6854 5498 7932 5504
rect 6767 5434 6813 5446
rect 6767 5350 6773 5434
rect 6807 5350 6813 5434
rect 6767 5338 6813 5350
rect 6454 5280 7854 5286
rect 6454 5246 6866 5280
rect 7842 5246 7854 5280
rect 6454 5240 7854 5246
rect 6454 4770 6729 5240
rect 6767 5176 6813 5188
rect 6767 5092 6773 5176
rect 6807 5092 6813 5176
rect 6767 5080 6813 5092
rect 7926 5028 7932 5498
rect 6854 5022 7932 5028
rect 6854 4988 6866 5022
rect 7842 4988 7932 5022
rect 6854 4982 7932 4988
rect 6767 4918 6813 4930
rect 6767 4834 6773 4918
rect 6807 4834 6813 4918
rect 6767 4822 6813 4834
rect 6454 4764 7854 4770
rect 6454 4730 6866 4764
rect 7842 4730 7854 4764
rect 6454 4724 7854 4730
rect 6454 4254 6729 4724
rect 6767 4660 6813 4672
rect 6767 4576 6773 4660
rect 6807 4576 6813 4660
rect 6767 4564 6813 4576
rect 7926 4512 7932 4982
rect 6854 4506 7932 4512
rect 6854 4472 6866 4506
rect 7842 4472 7932 4506
rect 6854 4466 7932 4472
rect 6767 4402 6813 4414
rect 6767 4318 6773 4402
rect 6807 4318 6813 4402
rect 6767 4306 6813 4318
rect 6454 4248 7854 4254
rect 6454 4214 6866 4248
rect 7842 4214 7854 4248
rect 6454 4208 7854 4214
rect 6454 3738 6729 4208
rect 6767 4144 6813 4156
rect 6767 4060 6773 4144
rect 6807 4060 6813 4144
rect 6767 4048 6813 4060
rect 7926 3996 7932 4466
rect 6854 3990 7932 3996
rect 6854 3956 6866 3990
rect 7842 3956 7932 3990
rect 6854 3950 7932 3956
rect 6767 3886 6813 3898
rect 6767 3802 6773 3886
rect 6807 3802 6813 3886
rect 6767 3790 6813 3802
rect 6454 3732 7854 3738
rect 6454 3698 6866 3732
rect 7842 3698 7854 3732
rect 6454 3692 7854 3698
rect 6454 3222 6729 3692
rect 6767 3628 6813 3640
rect 6767 3544 6773 3628
rect 6807 3544 6813 3628
rect 6767 3532 6813 3544
rect 7926 3480 7932 3950
rect 6854 3474 7932 3480
rect 6854 3440 6866 3474
rect 7842 3440 7932 3474
rect 6854 3434 7932 3440
rect 6767 3370 6813 3382
rect 6767 3286 6773 3370
rect 6807 3286 6813 3370
rect 6767 3274 6813 3286
rect 6454 3216 7854 3222
rect 6454 3182 6866 3216
rect 7842 3182 7854 3216
rect 6454 3176 7854 3182
rect 6454 2706 6729 3176
rect 6767 3112 6813 3124
rect 6767 3028 6773 3112
rect 6807 3028 6813 3112
rect 6767 3016 6813 3028
rect 7926 2964 7932 3434
rect 6854 2958 7932 2964
rect 6854 2924 6866 2958
rect 7842 2924 7932 2958
rect 6854 2918 7932 2924
rect 6767 2854 6813 2866
rect 6767 2770 6773 2854
rect 6807 2770 6813 2854
rect 6767 2758 6813 2770
rect 6454 2700 7854 2706
rect 6454 2666 6866 2700
rect 7842 2666 7854 2700
rect 6454 2660 7854 2666
rect 6454 2516 6729 2660
rect 7926 2592 7932 2918
rect 6815 2586 7932 2592
rect 7966 2586 8227 7940
rect 6815 2552 6827 2586
rect 7809 2552 8227 2586
rect 6815 2546 8227 2552
<< labels >>
rlabel metal1 4226 5114 4226 5114 7 GND
port 3 n
rlabel metal1 8128 5180 8128 5180 1 VDD
port 1 n
rlabel metal1 6546 5216 6546 5216 1 clamped
port 2 n
<< end >>
