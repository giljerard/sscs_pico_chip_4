magic
tech sky130A
timestamp 1636526374
<< metal3 >>
rect 30770 1630 53370 7225
rect 30770 1510 30835 1630
rect 30955 1510 31000 1630
rect 31120 1510 31165 1630
rect 31285 1510 31330 1630
rect 31450 1510 31495 1630
rect 31615 1510 31660 1630
rect 31780 1510 31825 1630
rect 31945 1510 31990 1630
rect 32110 1510 32155 1630
rect 32275 1510 32320 1630
rect 32440 1510 32485 1630
rect 32605 1510 32650 1630
rect 32770 1510 32815 1630
rect 32935 1510 32980 1630
rect 33100 1510 33145 1630
rect 33265 1510 33310 1630
rect 33430 1510 33475 1630
rect 33595 1510 33640 1630
rect 33760 1510 33805 1630
rect 33925 1510 33970 1630
rect 34090 1510 34135 1630
rect 34255 1510 34300 1630
rect 34420 1510 34465 1630
rect 34585 1510 34630 1630
rect 34750 1510 34795 1630
rect 34915 1510 34960 1630
rect 35080 1510 35125 1630
rect 35245 1510 35290 1630
rect 35410 1510 35455 1630
rect 35575 1510 35620 1630
rect 35740 1510 35785 1630
rect 35905 1510 35950 1630
rect 36070 1510 36115 1630
rect 36235 1510 36525 1630
rect 36645 1510 36690 1630
rect 36810 1510 36855 1630
rect 36975 1510 37020 1630
rect 37140 1510 37185 1630
rect 37305 1510 37350 1630
rect 37470 1510 37515 1630
rect 37635 1510 37680 1630
rect 37800 1510 37845 1630
rect 37965 1510 38010 1630
rect 38130 1510 38175 1630
rect 38295 1510 38340 1630
rect 38460 1510 38505 1630
rect 38625 1510 38670 1630
rect 38790 1510 38835 1630
rect 38955 1510 39000 1630
rect 39120 1510 39165 1630
rect 39285 1510 39330 1630
rect 39450 1510 39495 1630
rect 39615 1510 39660 1630
rect 39780 1510 39825 1630
rect 39945 1510 39990 1630
rect 40110 1510 40155 1630
rect 40275 1510 40320 1630
rect 40440 1510 40485 1630
rect 40605 1510 40650 1630
rect 40770 1510 40815 1630
rect 40935 1510 40980 1630
rect 41100 1510 41145 1630
rect 41265 1510 41310 1630
rect 41430 1510 41475 1630
rect 41595 1510 41640 1630
rect 41760 1510 41805 1630
rect 41925 1510 42215 1630
rect 42335 1510 42380 1630
rect 42500 1510 42545 1630
rect 42665 1510 42710 1630
rect 42830 1510 42875 1630
rect 42995 1510 43040 1630
rect 43160 1510 43205 1630
rect 43325 1510 43370 1630
rect 43490 1510 43535 1630
rect 43655 1510 43700 1630
rect 43820 1510 43865 1630
rect 43985 1510 44030 1630
rect 44150 1510 44195 1630
rect 44315 1510 44360 1630
rect 44480 1510 44525 1630
rect 44645 1510 44690 1630
rect 44810 1510 44855 1630
rect 44975 1510 45020 1630
rect 45140 1510 45185 1630
rect 45305 1510 45350 1630
rect 45470 1510 45515 1630
rect 45635 1510 45680 1630
rect 45800 1510 45845 1630
rect 45965 1510 46010 1630
rect 46130 1510 46175 1630
rect 46295 1510 46340 1630
rect 46460 1510 46505 1630
rect 46625 1510 46670 1630
rect 46790 1510 46835 1630
rect 46955 1510 47000 1630
rect 47120 1510 47165 1630
rect 47285 1510 47330 1630
rect 47450 1510 47495 1630
rect 47615 1510 47905 1630
rect 48025 1510 48070 1630
rect 48190 1510 48235 1630
rect 48355 1510 48400 1630
rect 48520 1510 48565 1630
rect 48685 1510 48730 1630
rect 48850 1510 48895 1630
rect 49015 1510 49060 1630
rect 49180 1510 49225 1630
rect 49345 1510 49390 1630
rect 49510 1510 49555 1630
rect 49675 1510 49720 1630
rect 49840 1510 49885 1630
rect 50005 1510 50050 1630
rect 50170 1510 50215 1630
rect 50335 1510 50380 1630
rect 50500 1510 50545 1630
rect 50665 1510 50710 1630
rect 50830 1510 50875 1630
rect 50995 1510 51040 1630
rect 51160 1510 51205 1630
rect 51325 1510 51370 1630
rect 51490 1510 51535 1630
rect 51655 1510 51700 1630
rect 51820 1510 51865 1630
rect 51985 1510 52030 1630
rect 52150 1510 52195 1630
rect 52315 1510 52360 1630
rect 52480 1510 52525 1630
rect 52645 1510 52690 1630
rect 52810 1510 52855 1630
rect 52975 1510 53020 1630
rect 53140 1510 53185 1630
rect 53305 1510 53370 1630
rect 30770 -9840 53370 1510
rect 30770 -9960 30835 -9840
rect 30955 -9960 31000 -9840
rect 31120 -9960 31165 -9840
rect 31285 -9960 31330 -9840
rect 31450 -9960 31495 -9840
rect 31615 -9960 31660 -9840
rect 31780 -9960 31825 -9840
rect 31945 -9960 31990 -9840
rect 32110 -9960 32155 -9840
rect 32275 -9960 32320 -9840
rect 32440 -9960 32485 -9840
rect 32605 -9960 32650 -9840
rect 32770 -9960 32815 -9840
rect 32935 -9960 32980 -9840
rect 33100 -9960 33145 -9840
rect 33265 -9960 33310 -9840
rect 33430 -9960 33475 -9840
rect 33595 -9960 33640 -9840
rect 33760 -9960 33805 -9840
rect 33925 -9960 33970 -9840
rect 34090 -9960 34135 -9840
rect 34255 -9960 34300 -9840
rect 34420 -9960 34465 -9840
rect 34585 -9960 34630 -9840
rect 34750 -9960 34795 -9840
rect 34915 -9960 34960 -9840
rect 35080 -9960 35125 -9840
rect 35245 -9960 35290 -9840
rect 35410 -9960 35455 -9840
rect 35575 -9960 35620 -9840
rect 35740 -9960 35785 -9840
rect 35905 -9960 35950 -9840
rect 36070 -9960 36115 -9840
rect 36235 -9960 36525 -9840
rect 36645 -9960 36690 -9840
rect 36810 -9960 36855 -9840
rect 36975 -9960 37020 -9840
rect 37140 -9960 37185 -9840
rect 37305 -9960 37350 -9840
rect 37470 -9960 37515 -9840
rect 37635 -9960 37680 -9840
rect 37800 -9960 37845 -9840
rect 37965 -9960 38010 -9840
rect 38130 -9960 38175 -9840
rect 38295 -9960 38340 -9840
rect 38460 -9960 38505 -9840
rect 38625 -9960 38670 -9840
rect 38790 -9960 38835 -9840
rect 38955 -9960 39000 -9840
rect 39120 -9960 39165 -9840
rect 39285 -9960 39330 -9840
rect 39450 -9960 39495 -9840
rect 39615 -9960 39660 -9840
rect 39780 -9960 39825 -9840
rect 39945 -9960 39990 -9840
rect 40110 -9960 40155 -9840
rect 40275 -9960 40320 -9840
rect 40440 -9960 40485 -9840
rect 40605 -9960 40650 -9840
rect 40770 -9960 40815 -9840
rect 40935 -9960 40980 -9840
rect 41100 -9960 41145 -9840
rect 41265 -9960 41310 -9840
rect 41430 -9960 41475 -9840
rect 41595 -9960 41640 -9840
rect 41760 -9960 41805 -9840
rect 41925 -9960 42215 -9840
rect 42335 -9960 42380 -9840
rect 42500 -9960 42545 -9840
rect 42665 -9960 42710 -9840
rect 42830 -9960 42875 -9840
rect 42995 -9960 43040 -9840
rect 43160 -9960 43205 -9840
rect 43325 -9960 43370 -9840
rect 43490 -9960 43535 -9840
rect 43655 -9960 43700 -9840
rect 43820 -9960 43865 -9840
rect 43985 -9960 44030 -9840
rect 44150 -9960 44195 -9840
rect 44315 -9960 44360 -9840
rect 44480 -9960 44525 -9840
rect 44645 -9960 44690 -9840
rect 44810 -9960 44855 -9840
rect 44975 -9960 45020 -9840
rect 45140 -9960 45185 -9840
rect 45305 -9960 45350 -9840
rect 45470 -9960 45515 -9840
rect 45635 -9960 45680 -9840
rect 45800 -9960 45845 -9840
rect 45965 -9960 46010 -9840
rect 46130 -9960 46175 -9840
rect 46295 -9960 46340 -9840
rect 46460 -9960 46505 -9840
rect 46625 -9960 46670 -9840
rect 46790 -9960 46835 -9840
rect 46955 -9960 47000 -9840
rect 47120 -9960 47165 -9840
rect 47285 -9960 47330 -9840
rect 47450 -9960 47495 -9840
rect 47615 -9960 47905 -9840
rect 48025 -9960 48070 -9840
rect 48190 -9960 48235 -9840
rect 48355 -9960 48400 -9840
rect 48520 -9960 48565 -9840
rect 48685 -9960 48730 -9840
rect 48850 -9960 48895 -9840
rect 49015 -9960 49060 -9840
rect 49180 -9960 49225 -9840
rect 49345 -9960 49390 -9840
rect 49510 -9960 49555 -9840
rect 49675 -9960 49720 -9840
rect 49840 -9960 49885 -9840
rect 50005 -9960 50050 -9840
rect 50170 -9960 50215 -9840
rect 50335 -9960 50380 -9840
rect 50500 -9960 50545 -9840
rect 50665 -9960 50710 -9840
rect 50830 -9960 50875 -9840
rect 50995 -9960 51040 -9840
rect 51160 -9960 51205 -9840
rect 51325 -9960 51370 -9840
rect 51490 -9960 51535 -9840
rect 51655 -9960 51700 -9840
rect 51820 -9960 51865 -9840
rect 51985 -9960 52030 -9840
rect 52150 -9960 52195 -9840
rect 52315 -9960 52360 -9840
rect 52480 -9960 52525 -9840
rect 52645 -9960 52690 -9840
rect 52810 -9960 52855 -9840
rect 52975 -9960 53020 -9840
rect 53140 -9960 53185 -9840
rect 53305 -9960 53370 -9840
rect 30770 -15555 53370 -9960
<< via3 >>
rect 30835 1510 30955 1630
rect 31000 1510 31120 1630
rect 31165 1510 31285 1630
rect 31330 1510 31450 1630
rect 31495 1510 31615 1630
rect 31660 1510 31780 1630
rect 31825 1510 31945 1630
rect 31990 1510 32110 1630
rect 32155 1510 32275 1630
rect 32320 1510 32440 1630
rect 32485 1510 32605 1630
rect 32650 1510 32770 1630
rect 32815 1510 32935 1630
rect 32980 1510 33100 1630
rect 33145 1510 33265 1630
rect 33310 1510 33430 1630
rect 33475 1510 33595 1630
rect 33640 1510 33760 1630
rect 33805 1510 33925 1630
rect 33970 1510 34090 1630
rect 34135 1510 34255 1630
rect 34300 1510 34420 1630
rect 34465 1510 34585 1630
rect 34630 1510 34750 1630
rect 34795 1510 34915 1630
rect 34960 1510 35080 1630
rect 35125 1510 35245 1630
rect 35290 1510 35410 1630
rect 35455 1510 35575 1630
rect 35620 1510 35740 1630
rect 35785 1510 35905 1630
rect 35950 1510 36070 1630
rect 36115 1510 36235 1630
rect 36525 1510 36645 1630
rect 36690 1510 36810 1630
rect 36855 1510 36975 1630
rect 37020 1510 37140 1630
rect 37185 1510 37305 1630
rect 37350 1510 37470 1630
rect 37515 1510 37635 1630
rect 37680 1510 37800 1630
rect 37845 1510 37965 1630
rect 38010 1510 38130 1630
rect 38175 1510 38295 1630
rect 38340 1510 38460 1630
rect 38505 1510 38625 1630
rect 38670 1510 38790 1630
rect 38835 1510 38955 1630
rect 39000 1510 39120 1630
rect 39165 1510 39285 1630
rect 39330 1510 39450 1630
rect 39495 1510 39615 1630
rect 39660 1510 39780 1630
rect 39825 1510 39945 1630
rect 39990 1510 40110 1630
rect 40155 1510 40275 1630
rect 40320 1510 40440 1630
rect 40485 1510 40605 1630
rect 40650 1510 40770 1630
rect 40815 1510 40935 1630
rect 40980 1510 41100 1630
rect 41145 1510 41265 1630
rect 41310 1510 41430 1630
rect 41475 1510 41595 1630
rect 41640 1510 41760 1630
rect 41805 1510 41925 1630
rect 42215 1510 42335 1630
rect 42380 1510 42500 1630
rect 42545 1510 42665 1630
rect 42710 1510 42830 1630
rect 42875 1510 42995 1630
rect 43040 1510 43160 1630
rect 43205 1510 43325 1630
rect 43370 1510 43490 1630
rect 43535 1510 43655 1630
rect 43700 1510 43820 1630
rect 43865 1510 43985 1630
rect 44030 1510 44150 1630
rect 44195 1510 44315 1630
rect 44360 1510 44480 1630
rect 44525 1510 44645 1630
rect 44690 1510 44810 1630
rect 44855 1510 44975 1630
rect 45020 1510 45140 1630
rect 45185 1510 45305 1630
rect 45350 1510 45470 1630
rect 45515 1510 45635 1630
rect 45680 1510 45800 1630
rect 45845 1510 45965 1630
rect 46010 1510 46130 1630
rect 46175 1510 46295 1630
rect 46340 1510 46460 1630
rect 46505 1510 46625 1630
rect 46670 1510 46790 1630
rect 46835 1510 46955 1630
rect 47000 1510 47120 1630
rect 47165 1510 47285 1630
rect 47330 1510 47450 1630
rect 47495 1510 47615 1630
rect 47905 1510 48025 1630
rect 48070 1510 48190 1630
rect 48235 1510 48355 1630
rect 48400 1510 48520 1630
rect 48565 1510 48685 1630
rect 48730 1510 48850 1630
rect 48895 1510 49015 1630
rect 49060 1510 49180 1630
rect 49225 1510 49345 1630
rect 49390 1510 49510 1630
rect 49555 1510 49675 1630
rect 49720 1510 49840 1630
rect 49885 1510 50005 1630
rect 50050 1510 50170 1630
rect 50215 1510 50335 1630
rect 50380 1510 50500 1630
rect 50545 1510 50665 1630
rect 50710 1510 50830 1630
rect 50875 1510 50995 1630
rect 51040 1510 51160 1630
rect 51205 1510 51325 1630
rect 51370 1510 51490 1630
rect 51535 1510 51655 1630
rect 51700 1510 51820 1630
rect 51865 1510 51985 1630
rect 52030 1510 52150 1630
rect 52195 1510 52315 1630
rect 52360 1510 52480 1630
rect 52525 1510 52645 1630
rect 52690 1510 52810 1630
rect 52855 1510 52975 1630
rect 53020 1510 53140 1630
rect 53185 1510 53305 1630
rect 30835 -9960 30955 -9840
rect 31000 -9960 31120 -9840
rect 31165 -9960 31285 -9840
rect 31330 -9960 31450 -9840
rect 31495 -9960 31615 -9840
rect 31660 -9960 31780 -9840
rect 31825 -9960 31945 -9840
rect 31990 -9960 32110 -9840
rect 32155 -9960 32275 -9840
rect 32320 -9960 32440 -9840
rect 32485 -9960 32605 -9840
rect 32650 -9960 32770 -9840
rect 32815 -9960 32935 -9840
rect 32980 -9960 33100 -9840
rect 33145 -9960 33265 -9840
rect 33310 -9960 33430 -9840
rect 33475 -9960 33595 -9840
rect 33640 -9960 33760 -9840
rect 33805 -9960 33925 -9840
rect 33970 -9960 34090 -9840
rect 34135 -9960 34255 -9840
rect 34300 -9960 34420 -9840
rect 34465 -9960 34585 -9840
rect 34630 -9960 34750 -9840
rect 34795 -9960 34915 -9840
rect 34960 -9960 35080 -9840
rect 35125 -9960 35245 -9840
rect 35290 -9960 35410 -9840
rect 35455 -9960 35575 -9840
rect 35620 -9960 35740 -9840
rect 35785 -9960 35905 -9840
rect 35950 -9960 36070 -9840
rect 36115 -9960 36235 -9840
rect 36525 -9960 36645 -9840
rect 36690 -9960 36810 -9840
rect 36855 -9960 36975 -9840
rect 37020 -9960 37140 -9840
rect 37185 -9960 37305 -9840
rect 37350 -9960 37470 -9840
rect 37515 -9960 37635 -9840
rect 37680 -9960 37800 -9840
rect 37845 -9960 37965 -9840
rect 38010 -9960 38130 -9840
rect 38175 -9960 38295 -9840
rect 38340 -9960 38460 -9840
rect 38505 -9960 38625 -9840
rect 38670 -9960 38790 -9840
rect 38835 -9960 38955 -9840
rect 39000 -9960 39120 -9840
rect 39165 -9960 39285 -9840
rect 39330 -9960 39450 -9840
rect 39495 -9960 39615 -9840
rect 39660 -9960 39780 -9840
rect 39825 -9960 39945 -9840
rect 39990 -9960 40110 -9840
rect 40155 -9960 40275 -9840
rect 40320 -9960 40440 -9840
rect 40485 -9960 40605 -9840
rect 40650 -9960 40770 -9840
rect 40815 -9960 40935 -9840
rect 40980 -9960 41100 -9840
rect 41145 -9960 41265 -9840
rect 41310 -9960 41430 -9840
rect 41475 -9960 41595 -9840
rect 41640 -9960 41760 -9840
rect 41805 -9960 41925 -9840
rect 42215 -9960 42335 -9840
rect 42380 -9960 42500 -9840
rect 42545 -9960 42665 -9840
rect 42710 -9960 42830 -9840
rect 42875 -9960 42995 -9840
rect 43040 -9960 43160 -9840
rect 43205 -9960 43325 -9840
rect 43370 -9960 43490 -9840
rect 43535 -9960 43655 -9840
rect 43700 -9960 43820 -9840
rect 43865 -9960 43985 -9840
rect 44030 -9960 44150 -9840
rect 44195 -9960 44315 -9840
rect 44360 -9960 44480 -9840
rect 44525 -9960 44645 -9840
rect 44690 -9960 44810 -9840
rect 44855 -9960 44975 -9840
rect 45020 -9960 45140 -9840
rect 45185 -9960 45305 -9840
rect 45350 -9960 45470 -9840
rect 45515 -9960 45635 -9840
rect 45680 -9960 45800 -9840
rect 45845 -9960 45965 -9840
rect 46010 -9960 46130 -9840
rect 46175 -9960 46295 -9840
rect 46340 -9960 46460 -9840
rect 46505 -9960 46625 -9840
rect 46670 -9960 46790 -9840
rect 46835 -9960 46955 -9840
rect 47000 -9960 47120 -9840
rect 47165 -9960 47285 -9840
rect 47330 -9960 47450 -9840
rect 47495 -9960 47615 -9840
rect 47905 -9960 48025 -9840
rect 48070 -9960 48190 -9840
rect 48235 -9960 48355 -9840
rect 48400 -9960 48520 -9840
rect 48565 -9960 48685 -9840
rect 48730 -9960 48850 -9840
rect 48895 -9960 49015 -9840
rect 49060 -9960 49180 -9840
rect 49225 -9960 49345 -9840
rect 49390 -9960 49510 -9840
rect 49555 -9960 49675 -9840
rect 49720 -9960 49840 -9840
rect 49885 -9960 50005 -9840
rect 50050 -9960 50170 -9840
rect 50215 -9960 50335 -9840
rect 50380 -9960 50500 -9840
rect 50545 -9960 50665 -9840
rect 50710 -9960 50830 -9840
rect 50875 -9960 50995 -9840
rect 51040 -9960 51160 -9840
rect 51205 -9960 51325 -9840
rect 51370 -9960 51490 -9840
rect 51535 -9960 51655 -9840
rect 51700 -9960 51820 -9840
rect 51865 -9960 51985 -9840
rect 52030 -9960 52150 -9840
rect 52195 -9960 52315 -9840
rect 52360 -9960 52480 -9840
rect 52525 -9960 52645 -9840
rect 52690 -9960 52810 -9840
rect 52855 -9960 52975 -9840
rect 53020 -9960 53140 -9840
rect 53185 -9960 53305 -9840
<< mimcap >>
rect 30785 7200 36285 7210
rect 30785 7080 30795 7200
rect 30915 7080 30960 7200
rect 31080 7080 31125 7200
rect 31245 7080 31290 7200
rect 31410 7080 31465 7200
rect 31585 7080 31630 7200
rect 31750 7080 31795 7200
rect 31915 7080 31960 7200
rect 32080 7080 32135 7200
rect 32255 7080 32300 7200
rect 32420 7080 32465 7200
rect 32585 7080 32630 7200
rect 32750 7080 32805 7200
rect 32925 7080 32970 7200
rect 33090 7080 33135 7200
rect 33255 7080 33300 7200
rect 33420 7080 33475 7200
rect 33595 7080 33640 7200
rect 33760 7080 33805 7200
rect 33925 7080 33970 7200
rect 34090 7080 34145 7200
rect 34265 7080 34310 7200
rect 34430 7080 34475 7200
rect 34595 7080 34640 7200
rect 34760 7080 34815 7200
rect 34935 7080 34980 7200
rect 35100 7080 35145 7200
rect 35265 7080 35310 7200
rect 35430 7080 35485 7200
rect 35605 7080 35650 7200
rect 35770 7080 35815 7200
rect 35935 7080 35980 7200
rect 36100 7080 36155 7200
rect 36275 7080 36285 7200
rect 30785 7025 36285 7080
rect 30785 6905 30795 7025
rect 30915 6905 30960 7025
rect 31080 6905 31125 7025
rect 31245 6905 31290 7025
rect 31410 6905 31465 7025
rect 31585 6905 31630 7025
rect 31750 6905 31795 7025
rect 31915 6905 31960 7025
rect 32080 6905 32135 7025
rect 32255 6905 32300 7025
rect 32420 6905 32465 7025
rect 32585 6905 32630 7025
rect 32750 6905 32805 7025
rect 32925 6905 32970 7025
rect 33090 6905 33135 7025
rect 33255 6905 33300 7025
rect 33420 6905 33475 7025
rect 33595 6905 33640 7025
rect 33760 6905 33805 7025
rect 33925 6905 33970 7025
rect 34090 6905 34145 7025
rect 34265 6905 34310 7025
rect 34430 6905 34475 7025
rect 34595 6905 34640 7025
rect 34760 6905 34815 7025
rect 34935 6905 34980 7025
rect 35100 6905 35145 7025
rect 35265 6905 35310 7025
rect 35430 6905 35485 7025
rect 35605 6905 35650 7025
rect 35770 6905 35815 7025
rect 35935 6905 35980 7025
rect 36100 6905 36155 7025
rect 36275 6905 36285 7025
rect 30785 6860 36285 6905
rect 30785 6740 30795 6860
rect 30915 6740 30960 6860
rect 31080 6740 31125 6860
rect 31245 6740 31290 6860
rect 31410 6740 31465 6860
rect 31585 6740 31630 6860
rect 31750 6740 31795 6860
rect 31915 6740 31960 6860
rect 32080 6740 32135 6860
rect 32255 6740 32300 6860
rect 32420 6740 32465 6860
rect 32585 6740 32630 6860
rect 32750 6740 32805 6860
rect 32925 6740 32970 6860
rect 33090 6740 33135 6860
rect 33255 6740 33300 6860
rect 33420 6740 33475 6860
rect 33595 6740 33640 6860
rect 33760 6740 33805 6860
rect 33925 6740 33970 6860
rect 34090 6740 34145 6860
rect 34265 6740 34310 6860
rect 34430 6740 34475 6860
rect 34595 6740 34640 6860
rect 34760 6740 34815 6860
rect 34935 6740 34980 6860
rect 35100 6740 35145 6860
rect 35265 6740 35310 6860
rect 35430 6740 35485 6860
rect 35605 6740 35650 6860
rect 35770 6740 35815 6860
rect 35935 6740 35980 6860
rect 36100 6740 36155 6860
rect 36275 6740 36285 6860
rect 30785 6695 36285 6740
rect 30785 6575 30795 6695
rect 30915 6575 30960 6695
rect 31080 6575 31125 6695
rect 31245 6575 31290 6695
rect 31410 6575 31465 6695
rect 31585 6575 31630 6695
rect 31750 6575 31795 6695
rect 31915 6575 31960 6695
rect 32080 6575 32135 6695
rect 32255 6575 32300 6695
rect 32420 6575 32465 6695
rect 32585 6575 32630 6695
rect 32750 6575 32805 6695
rect 32925 6575 32970 6695
rect 33090 6575 33135 6695
rect 33255 6575 33300 6695
rect 33420 6575 33475 6695
rect 33595 6575 33640 6695
rect 33760 6575 33805 6695
rect 33925 6575 33970 6695
rect 34090 6575 34145 6695
rect 34265 6575 34310 6695
rect 34430 6575 34475 6695
rect 34595 6575 34640 6695
rect 34760 6575 34815 6695
rect 34935 6575 34980 6695
rect 35100 6575 35145 6695
rect 35265 6575 35310 6695
rect 35430 6575 35485 6695
rect 35605 6575 35650 6695
rect 35770 6575 35815 6695
rect 35935 6575 35980 6695
rect 36100 6575 36155 6695
rect 36275 6575 36285 6695
rect 30785 6530 36285 6575
rect 30785 6410 30795 6530
rect 30915 6410 30960 6530
rect 31080 6410 31125 6530
rect 31245 6410 31290 6530
rect 31410 6410 31465 6530
rect 31585 6410 31630 6530
rect 31750 6410 31795 6530
rect 31915 6410 31960 6530
rect 32080 6410 32135 6530
rect 32255 6410 32300 6530
rect 32420 6410 32465 6530
rect 32585 6410 32630 6530
rect 32750 6410 32805 6530
rect 32925 6410 32970 6530
rect 33090 6410 33135 6530
rect 33255 6410 33300 6530
rect 33420 6410 33475 6530
rect 33595 6410 33640 6530
rect 33760 6410 33805 6530
rect 33925 6410 33970 6530
rect 34090 6410 34145 6530
rect 34265 6410 34310 6530
rect 34430 6410 34475 6530
rect 34595 6410 34640 6530
rect 34760 6410 34815 6530
rect 34935 6410 34980 6530
rect 35100 6410 35145 6530
rect 35265 6410 35310 6530
rect 35430 6410 35485 6530
rect 35605 6410 35650 6530
rect 35770 6410 35815 6530
rect 35935 6410 35980 6530
rect 36100 6410 36155 6530
rect 36275 6410 36285 6530
rect 30785 6355 36285 6410
rect 30785 6235 30795 6355
rect 30915 6235 30960 6355
rect 31080 6235 31125 6355
rect 31245 6235 31290 6355
rect 31410 6235 31465 6355
rect 31585 6235 31630 6355
rect 31750 6235 31795 6355
rect 31915 6235 31960 6355
rect 32080 6235 32135 6355
rect 32255 6235 32300 6355
rect 32420 6235 32465 6355
rect 32585 6235 32630 6355
rect 32750 6235 32805 6355
rect 32925 6235 32970 6355
rect 33090 6235 33135 6355
rect 33255 6235 33300 6355
rect 33420 6235 33475 6355
rect 33595 6235 33640 6355
rect 33760 6235 33805 6355
rect 33925 6235 33970 6355
rect 34090 6235 34145 6355
rect 34265 6235 34310 6355
rect 34430 6235 34475 6355
rect 34595 6235 34640 6355
rect 34760 6235 34815 6355
rect 34935 6235 34980 6355
rect 35100 6235 35145 6355
rect 35265 6235 35310 6355
rect 35430 6235 35485 6355
rect 35605 6235 35650 6355
rect 35770 6235 35815 6355
rect 35935 6235 35980 6355
rect 36100 6235 36155 6355
rect 36275 6235 36285 6355
rect 30785 6190 36285 6235
rect 30785 6070 30795 6190
rect 30915 6070 30960 6190
rect 31080 6070 31125 6190
rect 31245 6070 31290 6190
rect 31410 6070 31465 6190
rect 31585 6070 31630 6190
rect 31750 6070 31795 6190
rect 31915 6070 31960 6190
rect 32080 6070 32135 6190
rect 32255 6070 32300 6190
rect 32420 6070 32465 6190
rect 32585 6070 32630 6190
rect 32750 6070 32805 6190
rect 32925 6070 32970 6190
rect 33090 6070 33135 6190
rect 33255 6070 33300 6190
rect 33420 6070 33475 6190
rect 33595 6070 33640 6190
rect 33760 6070 33805 6190
rect 33925 6070 33970 6190
rect 34090 6070 34145 6190
rect 34265 6070 34310 6190
rect 34430 6070 34475 6190
rect 34595 6070 34640 6190
rect 34760 6070 34815 6190
rect 34935 6070 34980 6190
rect 35100 6070 35145 6190
rect 35265 6070 35310 6190
rect 35430 6070 35485 6190
rect 35605 6070 35650 6190
rect 35770 6070 35815 6190
rect 35935 6070 35980 6190
rect 36100 6070 36155 6190
rect 36275 6070 36285 6190
rect 30785 6025 36285 6070
rect 30785 5905 30795 6025
rect 30915 5905 30960 6025
rect 31080 5905 31125 6025
rect 31245 5905 31290 6025
rect 31410 5905 31465 6025
rect 31585 5905 31630 6025
rect 31750 5905 31795 6025
rect 31915 5905 31960 6025
rect 32080 5905 32135 6025
rect 32255 5905 32300 6025
rect 32420 5905 32465 6025
rect 32585 5905 32630 6025
rect 32750 5905 32805 6025
rect 32925 5905 32970 6025
rect 33090 5905 33135 6025
rect 33255 5905 33300 6025
rect 33420 5905 33475 6025
rect 33595 5905 33640 6025
rect 33760 5905 33805 6025
rect 33925 5905 33970 6025
rect 34090 5905 34145 6025
rect 34265 5905 34310 6025
rect 34430 5905 34475 6025
rect 34595 5905 34640 6025
rect 34760 5905 34815 6025
rect 34935 5905 34980 6025
rect 35100 5905 35145 6025
rect 35265 5905 35310 6025
rect 35430 5905 35485 6025
rect 35605 5905 35650 6025
rect 35770 5905 35815 6025
rect 35935 5905 35980 6025
rect 36100 5905 36155 6025
rect 36275 5905 36285 6025
rect 30785 5860 36285 5905
rect 30785 5740 30795 5860
rect 30915 5740 30960 5860
rect 31080 5740 31125 5860
rect 31245 5740 31290 5860
rect 31410 5740 31465 5860
rect 31585 5740 31630 5860
rect 31750 5740 31795 5860
rect 31915 5740 31960 5860
rect 32080 5740 32135 5860
rect 32255 5740 32300 5860
rect 32420 5740 32465 5860
rect 32585 5740 32630 5860
rect 32750 5740 32805 5860
rect 32925 5740 32970 5860
rect 33090 5740 33135 5860
rect 33255 5740 33300 5860
rect 33420 5740 33475 5860
rect 33595 5740 33640 5860
rect 33760 5740 33805 5860
rect 33925 5740 33970 5860
rect 34090 5740 34145 5860
rect 34265 5740 34310 5860
rect 34430 5740 34475 5860
rect 34595 5740 34640 5860
rect 34760 5740 34815 5860
rect 34935 5740 34980 5860
rect 35100 5740 35145 5860
rect 35265 5740 35310 5860
rect 35430 5740 35485 5860
rect 35605 5740 35650 5860
rect 35770 5740 35815 5860
rect 35935 5740 35980 5860
rect 36100 5740 36155 5860
rect 36275 5740 36285 5860
rect 30785 5685 36285 5740
rect 30785 5565 30795 5685
rect 30915 5565 30960 5685
rect 31080 5565 31125 5685
rect 31245 5565 31290 5685
rect 31410 5565 31465 5685
rect 31585 5565 31630 5685
rect 31750 5565 31795 5685
rect 31915 5565 31960 5685
rect 32080 5565 32135 5685
rect 32255 5565 32300 5685
rect 32420 5565 32465 5685
rect 32585 5565 32630 5685
rect 32750 5565 32805 5685
rect 32925 5565 32970 5685
rect 33090 5565 33135 5685
rect 33255 5565 33300 5685
rect 33420 5565 33475 5685
rect 33595 5565 33640 5685
rect 33760 5565 33805 5685
rect 33925 5565 33970 5685
rect 34090 5565 34145 5685
rect 34265 5565 34310 5685
rect 34430 5565 34475 5685
rect 34595 5565 34640 5685
rect 34760 5565 34815 5685
rect 34935 5565 34980 5685
rect 35100 5565 35145 5685
rect 35265 5565 35310 5685
rect 35430 5565 35485 5685
rect 35605 5565 35650 5685
rect 35770 5565 35815 5685
rect 35935 5565 35980 5685
rect 36100 5565 36155 5685
rect 36275 5565 36285 5685
rect 30785 5520 36285 5565
rect 30785 5400 30795 5520
rect 30915 5400 30960 5520
rect 31080 5400 31125 5520
rect 31245 5400 31290 5520
rect 31410 5400 31465 5520
rect 31585 5400 31630 5520
rect 31750 5400 31795 5520
rect 31915 5400 31960 5520
rect 32080 5400 32135 5520
rect 32255 5400 32300 5520
rect 32420 5400 32465 5520
rect 32585 5400 32630 5520
rect 32750 5400 32805 5520
rect 32925 5400 32970 5520
rect 33090 5400 33135 5520
rect 33255 5400 33300 5520
rect 33420 5400 33475 5520
rect 33595 5400 33640 5520
rect 33760 5400 33805 5520
rect 33925 5400 33970 5520
rect 34090 5400 34145 5520
rect 34265 5400 34310 5520
rect 34430 5400 34475 5520
rect 34595 5400 34640 5520
rect 34760 5400 34815 5520
rect 34935 5400 34980 5520
rect 35100 5400 35145 5520
rect 35265 5400 35310 5520
rect 35430 5400 35485 5520
rect 35605 5400 35650 5520
rect 35770 5400 35815 5520
rect 35935 5400 35980 5520
rect 36100 5400 36155 5520
rect 36275 5400 36285 5520
rect 30785 5355 36285 5400
rect 30785 5235 30795 5355
rect 30915 5235 30960 5355
rect 31080 5235 31125 5355
rect 31245 5235 31290 5355
rect 31410 5235 31465 5355
rect 31585 5235 31630 5355
rect 31750 5235 31795 5355
rect 31915 5235 31960 5355
rect 32080 5235 32135 5355
rect 32255 5235 32300 5355
rect 32420 5235 32465 5355
rect 32585 5235 32630 5355
rect 32750 5235 32805 5355
rect 32925 5235 32970 5355
rect 33090 5235 33135 5355
rect 33255 5235 33300 5355
rect 33420 5235 33475 5355
rect 33595 5235 33640 5355
rect 33760 5235 33805 5355
rect 33925 5235 33970 5355
rect 34090 5235 34145 5355
rect 34265 5235 34310 5355
rect 34430 5235 34475 5355
rect 34595 5235 34640 5355
rect 34760 5235 34815 5355
rect 34935 5235 34980 5355
rect 35100 5235 35145 5355
rect 35265 5235 35310 5355
rect 35430 5235 35485 5355
rect 35605 5235 35650 5355
rect 35770 5235 35815 5355
rect 35935 5235 35980 5355
rect 36100 5235 36155 5355
rect 36275 5235 36285 5355
rect 30785 5190 36285 5235
rect 30785 5070 30795 5190
rect 30915 5070 30960 5190
rect 31080 5070 31125 5190
rect 31245 5070 31290 5190
rect 31410 5070 31465 5190
rect 31585 5070 31630 5190
rect 31750 5070 31795 5190
rect 31915 5070 31960 5190
rect 32080 5070 32135 5190
rect 32255 5070 32300 5190
rect 32420 5070 32465 5190
rect 32585 5070 32630 5190
rect 32750 5070 32805 5190
rect 32925 5070 32970 5190
rect 33090 5070 33135 5190
rect 33255 5070 33300 5190
rect 33420 5070 33475 5190
rect 33595 5070 33640 5190
rect 33760 5070 33805 5190
rect 33925 5070 33970 5190
rect 34090 5070 34145 5190
rect 34265 5070 34310 5190
rect 34430 5070 34475 5190
rect 34595 5070 34640 5190
rect 34760 5070 34815 5190
rect 34935 5070 34980 5190
rect 35100 5070 35145 5190
rect 35265 5070 35310 5190
rect 35430 5070 35485 5190
rect 35605 5070 35650 5190
rect 35770 5070 35815 5190
rect 35935 5070 35980 5190
rect 36100 5070 36155 5190
rect 36275 5070 36285 5190
rect 30785 5015 36285 5070
rect 30785 4895 30795 5015
rect 30915 4895 30960 5015
rect 31080 4895 31125 5015
rect 31245 4895 31290 5015
rect 31410 4895 31465 5015
rect 31585 4895 31630 5015
rect 31750 4895 31795 5015
rect 31915 4895 31960 5015
rect 32080 4895 32135 5015
rect 32255 4895 32300 5015
rect 32420 4895 32465 5015
rect 32585 4895 32630 5015
rect 32750 4895 32805 5015
rect 32925 4895 32970 5015
rect 33090 4895 33135 5015
rect 33255 4895 33300 5015
rect 33420 4895 33475 5015
rect 33595 4895 33640 5015
rect 33760 4895 33805 5015
rect 33925 4895 33970 5015
rect 34090 4895 34145 5015
rect 34265 4895 34310 5015
rect 34430 4895 34475 5015
rect 34595 4895 34640 5015
rect 34760 4895 34815 5015
rect 34935 4895 34980 5015
rect 35100 4895 35145 5015
rect 35265 4895 35310 5015
rect 35430 4895 35485 5015
rect 35605 4895 35650 5015
rect 35770 4895 35815 5015
rect 35935 4895 35980 5015
rect 36100 4895 36155 5015
rect 36275 4895 36285 5015
rect 30785 4850 36285 4895
rect 30785 4730 30795 4850
rect 30915 4730 30960 4850
rect 31080 4730 31125 4850
rect 31245 4730 31290 4850
rect 31410 4730 31465 4850
rect 31585 4730 31630 4850
rect 31750 4730 31795 4850
rect 31915 4730 31960 4850
rect 32080 4730 32135 4850
rect 32255 4730 32300 4850
rect 32420 4730 32465 4850
rect 32585 4730 32630 4850
rect 32750 4730 32805 4850
rect 32925 4730 32970 4850
rect 33090 4730 33135 4850
rect 33255 4730 33300 4850
rect 33420 4730 33475 4850
rect 33595 4730 33640 4850
rect 33760 4730 33805 4850
rect 33925 4730 33970 4850
rect 34090 4730 34145 4850
rect 34265 4730 34310 4850
rect 34430 4730 34475 4850
rect 34595 4730 34640 4850
rect 34760 4730 34815 4850
rect 34935 4730 34980 4850
rect 35100 4730 35145 4850
rect 35265 4730 35310 4850
rect 35430 4730 35485 4850
rect 35605 4730 35650 4850
rect 35770 4730 35815 4850
rect 35935 4730 35980 4850
rect 36100 4730 36155 4850
rect 36275 4730 36285 4850
rect 30785 4685 36285 4730
rect 30785 4565 30795 4685
rect 30915 4565 30960 4685
rect 31080 4565 31125 4685
rect 31245 4565 31290 4685
rect 31410 4565 31465 4685
rect 31585 4565 31630 4685
rect 31750 4565 31795 4685
rect 31915 4565 31960 4685
rect 32080 4565 32135 4685
rect 32255 4565 32300 4685
rect 32420 4565 32465 4685
rect 32585 4565 32630 4685
rect 32750 4565 32805 4685
rect 32925 4565 32970 4685
rect 33090 4565 33135 4685
rect 33255 4565 33300 4685
rect 33420 4565 33475 4685
rect 33595 4565 33640 4685
rect 33760 4565 33805 4685
rect 33925 4565 33970 4685
rect 34090 4565 34145 4685
rect 34265 4565 34310 4685
rect 34430 4565 34475 4685
rect 34595 4565 34640 4685
rect 34760 4565 34815 4685
rect 34935 4565 34980 4685
rect 35100 4565 35145 4685
rect 35265 4565 35310 4685
rect 35430 4565 35485 4685
rect 35605 4565 35650 4685
rect 35770 4565 35815 4685
rect 35935 4565 35980 4685
rect 36100 4565 36155 4685
rect 36275 4565 36285 4685
rect 30785 4520 36285 4565
rect 30785 4400 30795 4520
rect 30915 4400 30960 4520
rect 31080 4400 31125 4520
rect 31245 4400 31290 4520
rect 31410 4400 31465 4520
rect 31585 4400 31630 4520
rect 31750 4400 31795 4520
rect 31915 4400 31960 4520
rect 32080 4400 32135 4520
rect 32255 4400 32300 4520
rect 32420 4400 32465 4520
rect 32585 4400 32630 4520
rect 32750 4400 32805 4520
rect 32925 4400 32970 4520
rect 33090 4400 33135 4520
rect 33255 4400 33300 4520
rect 33420 4400 33475 4520
rect 33595 4400 33640 4520
rect 33760 4400 33805 4520
rect 33925 4400 33970 4520
rect 34090 4400 34145 4520
rect 34265 4400 34310 4520
rect 34430 4400 34475 4520
rect 34595 4400 34640 4520
rect 34760 4400 34815 4520
rect 34935 4400 34980 4520
rect 35100 4400 35145 4520
rect 35265 4400 35310 4520
rect 35430 4400 35485 4520
rect 35605 4400 35650 4520
rect 35770 4400 35815 4520
rect 35935 4400 35980 4520
rect 36100 4400 36155 4520
rect 36275 4400 36285 4520
rect 30785 4345 36285 4400
rect 30785 4225 30795 4345
rect 30915 4225 30960 4345
rect 31080 4225 31125 4345
rect 31245 4225 31290 4345
rect 31410 4225 31465 4345
rect 31585 4225 31630 4345
rect 31750 4225 31795 4345
rect 31915 4225 31960 4345
rect 32080 4225 32135 4345
rect 32255 4225 32300 4345
rect 32420 4225 32465 4345
rect 32585 4225 32630 4345
rect 32750 4225 32805 4345
rect 32925 4225 32970 4345
rect 33090 4225 33135 4345
rect 33255 4225 33300 4345
rect 33420 4225 33475 4345
rect 33595 4225 33640 4345
rect 33760 4225 33805 4345
rect 33925 4225 33970 4345
rect 34090 4225 34145 4345
rect 34265 4225 34310 4345
rect 34430 4225 34475 4345
rect 34595 4225 34640 4345
rect 34760 4225 34815 4345
rect 34935 4225 34980 4345
rect 35100 4225 35145 4345
rect 35265 4225 35310 4345
rect 35430 4225 35485 4345
rect 35605 4225 35650 4345
rect 35770 4225 35815 4345
rect 35935 4225 35980 4345
rect 36100 4225 36155 4345
rect 36275 4225 36285 4345
rect 30785 4180 36285 4225
rect 30785 4060 30795 4180
rect 30915 4060 30960 4180
rect 31080 4060 31125 4180
rect 31245 4060 31290 4180
rect 31410 4060 31465 4180
rect 31585 4060 31630 4180
rect 31750 4060 31795 4180
rect 31915 4060 31960 4180
rect 32080 4060 32135 4180
rect 32255 4060 32300 4180
rect 32420 4060 32465 4180
rect 32585 4060 32630 4180
rect 32750 4060 32805 4180
rect 32925 4060 32970 4180
rect 33090 4060 33135 4180
rect 33255 4060 33300 4180
rect 33420 4060 33475 4180
rect 33595 4060 33640 4180
rect 33760 4060 33805 4180
rect 33925 4060 33970 4180
rect 34090 4060 34145 4180
rect 34265 4060 34310 4180
rect 34430 4060 34475 4180
rect 34595 4060 34640 4180
rect 34760 4060 34815 4180
rect 34935 4060 34980 4180
rect 35100 4060 35145 4180
rect 35265 4060 35310 4180
rect 35430 4060 35485 4180
rect 35605 4060 35650 4180
rect 35770 4060 35815 4180
rect 35935 4060 35980 4180
rect 36100 4060 36155 4180
rect 36275 4060 36285 4180
rect 30785 4015 36285 4060
rect 30785 3895 30795 4015
rect 30915 3895 30960 4015
rect 31080 3895 31125 4015
rect 31245 3895 31290 4015
rect 31410 3895 31465 4015
rect 31585 3895 31630 4015
rect 31750 3895 31795 4015
rect 31915 3895 31960 4015
rect 32080 3895 32135 4015
rect 32255 3895 32300 4015
rect 32420 3895 32465 4015
rect 32585 3895 32630 4015
rect 32750 3895 32805 4015
rect 32925 3895 32970 4015
rect 33090 3895 33135 4015
rect 33255 3895 33300 4015
rect 33420 3895 33475 4015
rect 33595 3895 33640 4015
rect 33760 3895 33805 4015
rect 33925 3895 33970 4015
rect 34090 3895 34145 4015
rect 34265 3895 34310 4015
rect 34430 3895 34475 4015
rect 34595 3895 34640 4015
rect 34760 3895 34815 4015
rect 34935 3895 34980 4015
rect 35100 3895 35145 4015
rect 35265 3895 35310 4015
rect 35430 3895 35485 4015
rect 35605 3895 35650 4015
rect 35770 3895 35815 4015
rect 35935 3895 35980 4015
rect 36100 3895 36155 4015
rect 36275 3895 36285 4015
rect 30785 3850 36285 3895
rect 30785 3730 30795 3850
rect 30915 3730 30960 3850
rect 31080 3730 31125 3850
rect 31245 3730 31290 3850
rect 31410 3730 31465 3850
rect 31585 3730 31630 3850
rect 31750 3730 31795 3850
rect 31915 3730 31960 3850
rect 32080 3730 32135 3850
rect 32255 3730 32300 3850
rect 32420 3730 32465 3850
rect 32585 3730 32630 3850
rect 32750 3730 32805 3850
rect 32925 3730 32970 3850
rect 33090 3730 33135 3850
rect 33255 3730 33300 3850
rect 33420 3730 33475 3850
rect 33595 3730 33640 3850
rect 33760 3730 33805 3850
rect 33925 3730 33970 3850
rect 34090 3730 34145 3850
rect 34265 3730 34310 3850
rect 34430 3730 34475 3850
rect 34595 3730 34640 3850
rect 34760 3730 34815 3850
rect 34935 3730 34980 3850
rect 35100 3730 35145 3850
rect 35265 3730 35310 3850
rect 35430 3730 35485 3850
rect 35605 3730 35650 3850
rect 35770 3730 35815 3850
rect 35935 3730 35980 3850
rect 36100 3730 36155 3850
rect 36275 3730 36285 3850
rect 30785 3675 36285 3730
rect 30785 3555 30795 3675
rect 30915 3555 30960 3675
rect 31080 3555 31125 3675
rect 31245 3555 31290 3675
rect 31410 3555 31465 3675
rect 31585 3555 31630 3675
rect 31750 3555 31795 3675
rect 31915 3555 31960 3675
rect 32080 3555 32135 3675
rect 32255 3555 32300 3675
rect 32420 3555 32465 3675
rect 32585 3555 32630 3675
rect 32750 3555 32805 3675
rect 32925 3555 32970 3675
rect 33090 3555 33135 3675
rect 33255 3555 33300 3675
rect 33420 3555 33475 3675
rect 33595 3555 33640 3675
rect 33760 3555 33805 3675
rect 33925 3555 33970 3675
rect 34090 3555 34145 3675
rect 34265 3555 34310 3675
rect 34430 3555 34475 3675
rect 34595 3555 34640 3675
rect 34760 3555 34815 3675
rect 34935 3555 34980 3675
rect 35100 3555 35145 3675
rect 35265 3555 35310 3675
rect 35430 3555 35485 3675
rect 35605 3555 35650 3675
rect 35770 3555 35815 3675
rect 35935 3555 35980 3675
rect 36100 3555 36155 3675
rect 36275 3555 36285 3675
rect 30785 3510 36285 3555
rect 30785 3390 30795 3510
rect 30915 3390 30960 3510
rect 31080 3390 31125 3510
rect 31245 3390 31290 3510
rect 31410 3390 31465 3510
rect 31585 3390 31630 3510
rect 31750 3390 31795 3510
rect 31915 3390 31960 3510
rect 32080 3390 32135 3510
rect 32255 3390 32300 3510
rect 32420 3390 32465 3510
rect 32585 3390 32630 3510
rect 32750 3390 32805 3510
rect 32925 3390 32970 3510
rect 33090 3390 33135 3510
rect 33255 3390 33300 3510
rect 33420 3390 33475 3510
rect 33595 3390 33640 3510
rect 33760 3390 33805 3510
rect 33925 3390 33970 3510
rect 34090 3390 34145 3510
rect 34265 3390 34310 3510
rect 34430 3390 34475 3510
rect 34595 3390 34640 3510
rect 34760 3390 34815 3510
rect 34935 3390 34980 3510
rect 35100 3390 35145 3510
rect 35265 3390 35310 3510
rect 35430 3390 35485 3510
rect 35605 3390 35650 3510
rect 35770 3390 35815 3510
rect 35935 3390 35980 3510
rect 36100 3390 36155 3510
rect 36275 3390 36285 3510
rect 30785 3345 36285 3390
rect 30785 3225 30795 3345
rect 30915 3225 30960 3345
rect 31080 3225 31125 3345
rect 31245 3225 31290 3345
rect 31410 3225 31465 3345
rect 31585 3225 31630 3345
rect 31750 3225 31795 3345
rect 31915 3225 31960 3345
rect 32080 3225 32135 3345
rect 32255 3225 32300 3345
rect 32420 3225 32465 3345
rect 32585 3225 32630 3345
rect 32750 3225 32805 3345
rect 32925 3225 32970 3345
rect 33090 3225 33135 3345
rect 33255 3225 33300 3345
rect 33420 3225 33475 3345
rect 33595 3225 33640 3345
rect 33760 3225 33805 3345
rect 33925 3225 33970 3345
rect 34090 3225 34145 3345
rect 34265 3225 34310 3345
rect 34430 3225 34475 3345
rect 34595 3225 34640 3345
rect 34760 3225 34815 3345
rect 34935 3225 34980 3345
rect 35100 3225 35145 3345
rect 35265 3225 35310 3345
rect 35430 3225 35485 3345
rect 35605 3225 35650 3345
rect 35770 3225 35815 3345
rect 35935 3225 35980 3345
rect 36100 3225 36155 3345
rect 36275 3225 36285 3345
rect 30785 3180 36285 3225
rect 30785 3060 30795 3180
rect 30915 3060 30960 3180
rect 31080 3060 31125 3180
rect 31245 3060 31290 3180
rect 31410 3060 31465 3180
rect 31585 3060 31630 3180
rect 31750 3060 31795 3180
rect 31915 3060 31960 3180
rect 32080 3060 32135 3180
rect 32255 3060 32300 3180
rect 32420 3060 32465 3180
rect 32585 3060 32630 3180
rect 32750 3060 32805 3180
rect 32925 3060 32970 3180
rect 33090 3060 33135 3180
rect 33255 3060 33300 3180
rect 33420 3060 33475 3180
rect 33595 3060 33640 3180
rect 33760 3060 33805 3180
rect 33925 3060 33970 3180
rect 34090 3060 34145 3180
rect 34265 3060 34310 3180
rect 34430 3060 34475 3180
rect 34595 3060 34640 3180
rect 34760 3060 34815 3180
rect 34935 3060 34980 3180
rect 35100 3060 35145 3180
rect 35265 3060 35310 3180
rect 35430 3060 35485 3180
rect 35605 3060 35650 3180
rect 35770 3060 35815 3180
rect 35935 3060 35980 3180
rect 36100 3060 36155 3180
rect 36275 3060 36285 3180
rect 30785 3005 36285 3060
rect 30785 2885 30795 3005
rect 30915 2885 30960 3005
rect 31080 2885 31125 3005
rect 31245 2885 31290 3005
rect 31410 2885 31465 3005
rect 31585 2885 31630 3005
rect 31750 2885 31795 3005
rect 31915 2885 31960 3005
rect 32080 2885 32135 3005
rect 32255 2885 32300 3005
rect 32420 2885 32465 3005
rect 32585 2885 32630 3005
rect 32750 2885 32805 3005
rect 32925 2885 32970 3005
rect 33090 2885 33135 3005
rect 33255 2885 33300 3005
rect 33420 2885 33475 3005
rect 33595 2885 33640 3005
rect 33760 2885 33805 3005
rect 33925 2885 33970 3005
rect 34090 2885 34145 3005
rect 34265 2885 34310 3005
rect 34430 2885 34475 3005
rect 34595 2885 34640 3005
rect 34760 2885 34815 3005
rect 34935 2885 34980 3005
rect 35100 2885 35145 3005
rect 35265 2885 35310 3005
rect 35430 2885 35485 3005
rect 35605 2885 35650 3005
rect 35770 2885 35815 3005
rect 35935 2885 35980 3005
rect 36100 2885 36155 3005
rect 36275 2885 36285 3005
rect 30785 2840 36285 2885
rect 30785 2720 30795 2840
rect 30915 2720 30960 2840
rect 31080 2720 31125 2840
rect 31245 2720 31290 2840
rect 31410 2720 31465 2840
rect 31585 2720 31630 2840
rect 31750 2720 31795 2840
rect 31915 2720 31960 2840
rect 32080 2720 32135 2840
rect 32255 2720 32300 2840
rect 32420 2720 32465 2840
rect 32585 2720 32630 2840
rect 32750 2720 32805 2840
rect 32925 2720 32970 2840
rect 33090 2720 33135 2840
rect 33255 2720 33300 2840
rect 33420 2720 33475 2840
rect 33595 2720 33640 2840
rect 33760 2720 33805 2840
rect 33925 2720 33970 2840
rect 34090 2720 34145 2840
rect 34265 2720 34310 2840
rect 34430 2720 34475 2840
rect 34595 2720 34640 2840
rect 34760 2720 34815 2840
rect 34935 2720 34980 2840
rect 35100 2720 35145 2840
rect 35265 2720 35310 2840
rect 35430 2720 35485 2840
rect 35605 2720 35650 2840
rect 35770 2720 35815 2840
rect 35935 2720 35980 2840
rect 36100 2720 36155 2840
rect 36275 2720 36285 2840
rect 30785 2675 36285 2720
rect 30785 2555 30795 2675
rect 30915 2555 30960 2675
rect 31080 2555 31125 2675
rect 31245 2555 31290 2675
rect 31410 2555 31465 2675
rect 31585 2555 31630 2675
rect 31750 2555 31795 2675
rect 31915 2555 31960 2675
rect 32080 2555 32135 2675
rect 32255 2555 32300 2675
rect 32420 2555 32465 2675
rect 32585 2555 32630 2675
rect 32750 2555 32805 2675
rect 32925 2555 32970 2675
rect 33090 2555 33135 2675
rect 33255 2555 33300 2675
rect 33420 2555 33475 2675
rect 33595 2555 33640 2675
rect 33760 2555 33805 2675
rect 33925 2555 33970 2675
rect 34090 2555 34145 2675
rect 34265 2555 34310 2675
rect 34430 2555 34475 2675
rect 34595 2555 34640 2675
rect 34760 2555 34815 2675
rect 34935 2555 34980 2675
rect 35100 2555 35145 2675
rect 35265 2555 35310 2675
rect 35430 2555 35485 2675
rect 35605 2555 35650 2675
rect 35770 2555 35815 2675
rect 35935 2555 35980 2675
rect 36100 2555 36155 2675
rect 36275 2555 36285 2675
rect 30785 2510 36285 2555
rect 30785 2390 30795 2510
rect 30915 2390 30960 2510
rect 31080 2390 31125 2510
rect 31245 2390 31290 2510
rect 31410 2390 31465 2510
rect 31585 2390 31630 2510
rect 31750 2390 31795 2510
rect 31915 2390 31960 2510
rect 32080 2390 32135 2510
rect 32255 2390 32300 2510
rect 32420 2390 32465 2510
rect 32585 2390 32630 2510
rect 32750 2390 32805 2510
rect 32925 2390 32970 2510
rect 33090 2390 33135 2510
rect 33255 2390 33300 2510
rect 33420 2390 33475 2510
rect 33595 2390 33640 2510
rect 33760 2390 33805 2510
rect 33925 2390 33970 2510
rect 34090 2390 34145 2510
rect 34265 2390 34310 2510
rect 34430 2390 34475 2510
rect 34595 2390 34640 2510
rect 34760 2390 34815 2510
rect 34935 2390 34980 2510
rect 35100 2390 35145 2510
rect 35265 2390 35310 2510
rect 35430 2390 35485 2510
rect 35605 2390 35650 2510
rect 35770 2390 35815 2510
rect 35935 2390 35980 2510
rect 36100 2390 36155 2510
rect 36275 2390 36285 2510
rect 30785 2335 36285 2390
rect 30785 2215 30795 2335
rect 30915 2215 30960 2335
rect 31080 2215 31125 2335
rect 31245 2215 31290 2335
rect 31410 2215 31465 2335
rect 31585 2215 31630 2335
rect 31750 2215 31795 2335
rect 31915 2215 31960 2335
rect 32080 2215 32135 2335
rect 32255 2215 32300 2335
rect 32420 2215 32465 2335
rect 32585 2215 32630 2335
rect 32750 2215 32805 2335
rect 32925 2215 32970 2335
rect 33090 2215 33135 2335
rect 33255 2215 33300 2335
rect 33420 2215 33475 2335
rect 33595 2215 33640 2335
rect 33760 2215 33805 2335
rect 33925 2215 33970 2335
rect 34090 2215 34145 2335
rect 34265 2215 34310 2335
rect 34430 2215 34475 2335
rect 34595 2215 34640 2335
rect 34760 2215 34815 2335
rect 34935 2215 34980 2335
rect 35100 2215 35145 2335
rect 35265 2215 35310 2335
rect 35430 2215 35485 2335
rect 35605 2215 35650 2335
rect 35770 2215 35815 2335
rect 35935 2215 35980 2335
rect 36100 2215 36155 2335
rect 36275 2215 36285 2335
rect 30785 2170 36285 2215
rect 30785 2050 30795 2170
rect 30915 2050 30960 2170
rect 31080 2050 31125 2170
rect 31245 2050 31290 2170
rect 31410 2050 31465 2170
rect 31585 2050 31630 2170
rect 31750 2050 31795 2170
rect 31915 2050 31960 2170
rect 32080 2050 32135 2170
rect 32255 2050 32300 2170
rect 32420 2050 32465 2170
rect 32585 2050 32630 2170
rect 32750 2050 32805 2170
rect 32925 2050 32970 2170
rect 33090 2050 33135 2170
rect 33255 2050 33300 2170
rect 33420 2050 33475 2170
rect 33595 2050 33640 2170
rect 33760 2050 33805 2170
rect 33925 2050 33970 2170
rect 34090 2050 34145 2170
rect 34265 2050 34310 2170
rect 34430 2050 34475 2170
rect 34595 2050 34640 2170
rect 34760 2050 34815 2170
rect 34935 2050 34980 2170
rect 35100 2050 35145 2170
rect 35265 2050 35310 2170
rect 35430 2050 35485 2170
rect 35605 2050 35650 2170
rect 35770 2050 35815 2170
rect 35935 2050 35980 2170
rect 36100 2050 36155 2170
rect 36275 2050 36285 2170
rect 30785 2005 36285 2050
rect 30785 1885 30795 2005
rect 30915 1885 30960 2005
rect 31080 1885 31125 2005
rect 31245 1885 31290 2005
rect 31410 1885 31465 2005
rect 31585 1885 31630 2005
rect 31750 1885 31795 2005
rect 31915 1885 31960 2005
rect 32080 1885 32135 2005
rect 32255 1885 32300 2005
rect 32420 1885 32465 2005
rect 32585 1885 32630 2005
rect 32750 1885 32805 2005
rect 32925 1885 32970 2005
rect 33090 1885 33135 2005
rect 33255 1885 33300 2005
rect 33420 1885 33475 2005
rect 33595 1885 33640 2005
rect 33760 1885 33805 2005
rect 33925 1885 33970 2005
rect 34090 1885 34145 2005
rect 34265 1885 34310 2005
rect 34430 1885 34475 2005
rect 34595 1885 34640 2005
rect 34760 1885 34815 2005
rect 34935 1885 34980 2005
rect 35100 1885 35145 2005
rect 35265 1885 35310 2005
rect 35430 1885 35485 2005
rect 35605 1885 35650 2005
rect 35770 1885 35815 2005
rect 35935 1885 35980 2005
rect 36100 1885 36155 2005
rect 36275 1885 36285 2005
rect 30785 1840 36285 1885
rect 30785 1720 30795 1840
rect 30915 1720 30960 1840
rect 31080 1720 31125 1840
rect 31245 1720 31290 1840
rect 31410 1720 31465 1840
rect 31585 1720 31630 1840
rect 31750 1720 31795 1840
rect 31915 1720 31960 1840
rect 32080 1720 32135 1840
rect 32255 1720 32300 1840
rect 32420 1720 32465 1840
rect 32585 1720 32630 1840
rect 32750 1720 32805 1840
rect 32925 1720 32970 1840
rect 33090 1720 33135 1840
rect 33255 1720 33300 1840
rect 33420 1720 33475 1840
rect 33595 1720 33640 1840
rect 33760 1720 33805 1840
rect 33925 1720 33970 1840
rect 34090 1720 34145 1840
rect 34265 1720 34310 1840
rect 34430 1720 34475 1840
rect 34595 1720 34640 1840
rect 34760 1720 34815 1840
rect 34935 1720 34980 1840
rect 35100 1720 35145 1840
rect 35265 1720 35310 1840
rect 35430 1720 35485 1840
rect 35605 1720 35650 1840
rect 35770 1720 35815 1840
rect 35935 1720 35980 1840
rect 36100 1720 36155 1840
rect 36275 1720 36285 1840
rect 30785 1710 36285 1720
rect 36475 7200 41975 7210
rect 36475 7080 36485 7200
rect 36605 7080 36650 7200
rect 36770 7080 36815 7200
rect 36935 7080 36980 7200
rect 37100 7080 37155 7200
rect 37275 7080 37320 7200
rect 37440 7080 37485 7200
rect 37605 7080 37650 7200
rect 37770 7080 37825 7200
rect 37945 7080 37990 7200
rect 38110 7080 38155 7200
rect 38275 7080 38320 7200
rect 38440 7080 38495 7200
rect 38615 7080 38660 7200
rect 38780 7080 38825 7200
rect 38945 7080 38990 7200
rect 39110 7080 39165 7200
rect 39285 7080 39330 7200
rect 39450 7080 39495 7200
rect 39615 7080 39660 7200
rect 39780 7080 39835 7200
rect 39955 7080 40000 7200
rect 40120 7080 40165 7200
rect 40285 7080 40330 7200
rect 40450 7080 40505 7200
rect 40625 7080 40670 7200
rect 40790 7080 40835 7200
rect 40955 7080 41000 7200
rect 41120 7080 41175 7200
rect 41295 7080 41340 7200
rect 41460 7080 41505 7200
rect 41625 7080 41670 7200
rect 41790 7080 41845 7200
rect 41965 7080 41975 7200
rect 36475 7025 41975 7080
rect 36475 6905 36485 7025
rect 36605 6905 36650 7025
rect 36770 6905 36815 7025
rect 36935 6905 36980 7025
rect 37100 6905 37155 7025
rect 37275 6905 37320 7025
rect 37440 6905 37485 7025
rect 37605 6905 37650 7025
rect 37770 6905 37825 7025
rect 37945 6905 37990 7025
rect 38110 6905 38155 7025
rect 38275 6905 38320 7025
rect 38440 6905 38495 7025
rect 38615 6905 38660 7025
rect 38780 6905 38825 7025
rect 38945 6905 38990 7025
rect 39110 6905 39165 7025
rect 39285 6905 39330 7025
rect 39450 6905 39495 7025
rect 39615 6905 39660 7025
rect 39780 6905 39835 7025
rect 39955 6905 40000 7025
rect 40120 6905 40165 7025
rect 40285 6905 40330 7025
rect 40450 6905 40505 7025
rect 40625 6905 40670 7025
rect 40790 6905 40835 7025
rect 40955 6905 41000 7025
rect 41120 6905 41175 7025
rect 41295 6905 41340 7025
rect 41460 6905 41505 7025
rect 41625 6905 41670 7025
rect 41790 6905 41845 7025
rect 41965 6905 41975 7025
rect 36475 6860 41975 6905
rect 36475 6740 36485 6860
rect 36605 6740 36650 6860
rect 36770 6740 36815 6860
rect 36935 6740 36980 6860
rect 37100 6740 37155 6860
rect 37275 6740 37320 6860
rect 37440 6740 37485 6860
rect 37605 6740 37650 6860
rect 37770 6740 37825 6860
rect 37945 6740 37990 6860
rect 38110 6740 38155 6860
rect 38275 6740 38320 6860
rect 38440 6740 38495 6860
rect 38615 6740 38660 6860
rect 38780 6740 38825 6860
rect 38945 6740 38990 6860
rect 39110 6740 39165 6860
rect 39285 6740 39330 6860
rect 39450 6740 39495 6860
rect 39615 6740 39660 6860
rect 39780 6740 39835 6860
rect 39955 6740 40000 6860
rect 40120 6740 40165 6860
rect 40285 6740 40330 6860
rect 40450 6740 40505 6860
rect 40625 6740 40670 6860
rect 40790 6740 40835 6860
rect 40955 6740 41000 6860
rect 41120 6740 41175 6860
rect 41295 6740 41340 6860
rect 41460 6740 41505 6860
rect 41625 6740 41670 6860
rect 41790 6740 41845 6860
rect 41965 6740 41975 6860
rect 36475 6695 41975 6740
rect 36475 6575 36485 6695
rect 36605 6575 36650 6695
rect 36770 6575 36815 6695
rect 36935 6575 36980 6695
rect 37100 6575 37155 6695
rect 37275 6575 37320 6695
rect 37440 6575 37485 6695
rect 37605 6575 37650 6695
rect 37770 6575 37825 6695
rect 37945 6575 37990 6695
rect 38110 6575 38155 6695
rect 38275 6575 38320 6695
rect 38440 6575 38495 6695
rect 38615 6575 38660 6695
rect 38780 6575 38825 6695
rect 38945 6575 38990 6695
rect 39110 6575 39165 6695
rect 39285 6575 39330 6695
rect 39450 6575 39495 6695
rect 39615 6575 39660 6695
rect 39780 6575 39835 6695
rect 39955 6575 40000 6695
rect 40120 6575 40165 6695
rect 40285 6575 40330 6695
rect 40450 6575 40505 6695
rect 40625 6575 40670 6695
rect 40790 6575 40835 6695
rect 40955 6575 41000 6695
rect 41120 6575 41175 6695
rect 41295 6575 41340 6695
rect 41460 6575 41505 6695
rect 41625 6575 41670 6695
rect 41790 6575 41845 6695
rect 41965 6575 41975 6695
rect 36475 6530 41975 6575
rect 36475 6410 36485 6530
rect 36605 6410 36650 6530
rect 36770 6410 36815 6530
rect 36935 6410 36980 6530
rect 37100 6410 37155 6530
rect 37275 6410 37320 6530
rect 37440 6410 37485 6530
rect 37605 6410 37650 6530
rect 37770 6410 37825 6530
rect 37945 6410 37990 6530
rect 38110 6410 38155 6530
rect 38275 6410 38320 6530
rect 38440 6410 38495 6530
rect 38615 6410 38660 6530
rect 38780 6410 38825 6530
rect 38945 6410 38990 6530
rect 39110 6410 39165 6530
rect 39285 6410 39330 6530
rect 39450 6410 39495 6530
rect 39615 6410 39660 6530
rect 39780 6410 39835 6530
rect 39955 6410 40000 6530
rect 40120 6410 40165 6530
rect 40285 6410 40330 6530
rect 40450 6410 40505 6530
rect 40625 6410 40670 6530
rect 40790 6410 40835 6530
rect 40955 6410 41000 6530
rect 41120 6410 41175 6530
rect 41295 6410 41340 6530
rect 41460 6410 41505 6530
rect 41625 6410 41670 6530
rect 41790 6410 41845 6530
rect 41965 6410 41975 6530
rect 36475 6355 41975 6410
rect 36475 6235 36485 6355
rect 36605 6235 36650 6355
rect 36770 6235 36815 6355
rect 36935 6235 36980 6355
rect 37100 6235 37155 6355
rect 37275 6235 37320 6355
rect 37440 6235 37485 6355
rect 37605 6235 37650 6355
rect 37770 6235 37825 6355
rect 37945 6235 37990 6355
rect 38110 6235 38155 6355
rect 38275 6235 38320 6355
rect 38440 6235 38495 6355
rect 38615 6235 38660 6355
rect 38780 6235 38825 6355
rect 38945 6235 38990 6355
rect 39110 6235 39165 6355
rect 39285 6235 39330 6355
rect 39450 6235 39495 6355
rect 39615 6235 39660 6355
rect 39780 6235 39835 6355
rect 39955 6235 40000 6355
rect 40120 6235 40165 6355
rect 40285 6235 40330 6355
rect 40450 6235 40505 6355
rect 40625 6235 40670 6355
rect 40790 6235 40835 6355
rect 40955 6235 41000 6355
rect 41120 6235 41175 6355
rect 41295 6235 41340 6355
rect 41460 6235 41505 6355
rect 41625 6235 41670 6355
rect 41790 6235 41845 6355
rect 41965 6235 41975 6355
rect 36475 6190 41975 6235
rect 36475 6070 36485 6190
rect 36605 6070 36650 6190
rect 36770 6070 36815 6190
rect 36935 6070 36980 6190
rect 37100 6070 37155 6190
rect 37275 6070 37320 6190
rect 37440 6070 37485 6190
rect 37605 6070 37650 6190
rect 37770 6070 37825 6190
rect 37945 6070 37990 6190
rect 38110 6070 38155 6190
rect 38275 6070 38320 6190
rect 38440 6070 38495 6190
rect 38615 6070 38660 6190
rect 38780 6070 38825 6190
rect 38945 6070 38990 6190
rect 39110 6070 39165 6190
rect 39285 6070 39330 6190
rect 39450 6070 39495 6190
rect 39615 6070 39660 6190
rect 39780 6070 39835 6190
rect 39955 6070 40000 6190
rect 40120 6070 40165 6190
rect 40285 6070 40330 6190
rect 40450 6070 40505 6190
rect 40625 6070 40670 6190
rect 40790 6070 40835 6190
rect 40955 6070 41000 6190
rect 41120 6070 41175 6190
rect 41295 6070 41340 6190
rect 41460 6070 41505 6190
rect 41625 6070 41670 6190
rect 41790 6070 41845 6190
rect 41965 6070 41975 6190
rect 36475 6025 41975 6070
rect 36475 5905 36485 6025
rect 36605 5905 36650 6025
rect 36770 5905 36815 6025
rect 36935 5905 36980 6025
rect 37100 5905 37155 6025
rect 37275 5905 37320 6025
rect 37440 5905 37485 6025
rect 37605 5905 37650 6025
rect 37770 5905 37825 6025
rect 37945 5905 37990 6025
rect 38110 5905 38155 6025
rect 38275 5905 38320 6025
rect 38440 5905 38495 6025
rect 38615 5905 38660 6025
rect 38780 5905 38825 6025
rect 38945 5905 38990 6025
rect 39110 5905 39165 6025
rect 39285 5905 39330 6025
rect 39450 5905 39495 6025
rect 39615 5905 39660 6025
rect 39780 5905 39835 6025
rect 39955 5905 40000 6025
rect 40120 5905 40165 6025
rect 40285 5905 40330 6025
rect 40450 5905 40505 6025
rect 40625 5905 40670 6025
rect 40790 5905 40835 6025
rect 40955 5905 41000 6025
rect 41120 5905 41175 6025
rect 41295 5905 41340 6025
rect 41460 5905 41505 6025
rect 41625 5905 41670 6025
rect 41790 5905 41845 6025
rect 41965 5905 41975 6025
rect 36475 5860 41975 5905
rect 36475 5740 36485 5860
rect 36605 5740 36650 5860
rect 36770 5740 36815 5860
rect 36935 5740 36980 5860
rect 37100 5740 37155 5860
rect 37275 5740 37320 5860
rect 37440 5740 37485 5860
rect 37605 5740 37650 5860
rect 37770 5740 37825 5860
rect 37945 5740 37990 5860
rect 38110 5740 38155 5860
rect 38275 5740 38320 5860
rect 38440 5740 38495 5860
rect 38615 5740 38660 5860
rect 38780 5740 38825 5860
rect 38945 5740 38990 5860
rect 39110 5740 39165 5860
rect 39285 5740 39330 5860
rect 39450 5740 39495 5860
rect 39615 5740 39660 5860
rect 39780 5740 39835 5860
rect 39955 5740 40000 5860
rect 40120 5740 40165 5860
rect 40285 5740 40330 5860
rect 40450 5740 40505 5860
rect 40625 5740 40670 5860
rect 40790 5740 40835 5860
rect 40955 5740 41000 5860
rect 41120 5740 41175 5860
rect 41295 5740 41340 5860
rect 41460 5740 41505 5860
rect 41625 5740 41670 5860
rect 41790 5740 41845 5860
rect 41965 5740 41975 5860
rect 36475 5685 41975 5740
rect 36475 5565 36485 5685
rect 36605 5565 36650 5685
rect 36770 5565 36815 5685
rect 36935 5565 36980 5685
rect 37100 5565 37155 5685
rect 37275 5565 37320 5685
rect 37440 5565 37485 5685
rect 37605 5565 37650 5685
rect 37770 5565 37825 5685
rect 37945 5565 37990 5685
rect 38110 5565 38155 5685
rect 38275 5565 38320 5685
rect 38440 5565 38495 5685
rect 38615 5565 38660 5685
rect 38780 5565 38825 5685
rect 38945 5565 38990 5685
rect 39110 5565 39165 5685
rect 39285 5565 39330 5685
rect 39450 5565 39495 5685
rect 39615 5565 39660 5685
rect 39780 5565 39835 5685
rect 39955 5565 40000 5685
rect 40120 5565 40165 5685
rect 40285 5565 40330 5685
rect 40450 5565 40505 5685
rect 40625 5565 40670 5685
rect 40790 5565 40835 5685
rect 40955 5565 41000 5685
rect 41120 5565 41175 5685
rect 41295 5565 41340 5685
rect 41460 5565 41505 5685
rect 41625 5565 41670 5685
rect 41790 5565 41845 5685
rect 41965 5565 41975 5685
rect 36475 5520 41975 5565
rect 36475 5400 36485 5520
rect 36605 5400 36650 5520
rect 36770 5400 36815 5520
rect 36935 5400 36980 5520
rect 37100 5400 37155 5520
rect 37275 5400 37320 5520
rect 37440 5400 37485 5520
rect 37605 5400 37650 5520
rect 37770 5400 37825 5520
rect 37945 5400 37990 5520
rect 38110 5400 38155 5520
rect 38275 5400 38320 5520
rect 38440 5400 38495 5520
rect 38615 5400 38660 5520
rect 38780 5400 38825 5520
rect 38945 5400 38990 5520
rect 39110 5400 39165 5520
rect 39285 5400 39330 5520
rect 39450 5400 39495 5520
rect 39615 5400 39660 5520
rect 39780 5400 39835 5520
rect 39955 5400 40000 5520
rect 40120 5400 40165 5520
rect 40285 5400 40330 5520
rect 40450 5400 40505 5520
rect 40625 5400 40670 5520
rect 40790 5400 40835 5520
rect 40955 5400 41000 5520
rect 41120 5400 41175 5520
rect 41295 5400 41340 5520
rect 41460 5400 41505 5520
rect 41625 5400 41670 5520
rect 41790 5400 41845 5520
rect 41965 5400 41975 5520
rect 36475 5355 41975 5400
rect 36475 5235 36485 5355
rect 36605 5235 36650 5355
rect 36770 5235 36815 5355
rect 36935 5235 36980 5355
rect 37100 5235 37155 5355
rect 37275 5235 37320 5355
rect 37440 5235 37485 5355
rect 37605 5235 37650 5355
rect 37770 5235 37825 5355
rect 37945 5235 37990 5355
rect 38110 5235 38155 5355
rect 38275 5235 38320 5355
rect 38440 5235 38495 5355
rect 38615 5235 38660 5355
rect 38780 5235 38825 5355
rect 38945 5235 38990 5355
rect 39110 5235 39165 5355
rect 39285 5235 39330 5355
rect 39450 5235 39495 5355
rect 39615 5235 39660 5355
rect 39780 5235 39835 5355
rect 39955 5235 40000 5355
rect 40120 5235 40165 5355
rect 40285 5235 40330 5355
rect 40450 5235 40505 5355
rect 40625 5235 40670 5355
rect 40790 5235 40835 5355
rect 40955 5235 41000 5355
rect 41120 5235 41175 5355
rect 41295 5235 41340 5355
rect 41460 5235 41505 5355
rect 41625 5235 41670 5355
rect 41790 5235 41845 5355
rect 41965 5235 41975 5355
rect 36475 5190 41975 5235
rect 36475 5070 36485 5190
rect 36605 5070 36650 5190
rect 36770 5070 36815 5190
rect 36935 5070 36980 5190
rect 37100 5070 37155 5190
rect 37275 5070 37320 5190
rect 37440 5070 37485 5190
rect 37605 5070 37650 5190
rect 37770 5070 37825 5190
rect 37945 5070 37990 5190
rect 38110 5070 38155 5190
rect 38275 5070 38320 5190
rect 38440 5070 38495 5190
rect 38615 5070 38660 5190
rect 38780 5070 38825 5190
rect 38945 5070 38990 5190
rect 39110 5070 39165 5190
rect 39285 5070 39330 5190
rect 39450 5070 39495 5190
rect 39615 5070 39660 5190
rect 39780 5070 39835 5190
rect 39955 5070 40000 5190
rect 40120 5070 40165 5190
rect 40285 5070 40330 5190
rect 40450 5070 40505 5190
rect 40625 5070 40670 5190
rect 40790 5070 40835 5190
rect 40955 5070 41000 5190
rect 41120 5070 41175 5190
rect 41295 5070 41340 5190
rect 41460 5070 41505 5190
rect 41625 5070 41670 5190
rect 41790 5070 41845 5190
rect 41965 5070 41975 5190
rect 36475 5015 41975 5070
rect 36475 4895 36485 5015
rect 36605 4895 36650 5015
rect 36770 4895 36815 5015
rect 36935 4895 36980 5015
rect 37100 4895 37155 5015
rect 37275 4895 37320 5015
rect 37440 4895 37485 5015
rect 37605 4895 37650 5015
rect 37770 4895 37825 5015
rect 37945 4895 37990 5015
rect 38110 4895 38155 5015
rect 38275 4895 38320 5015
rect 38440 4895 38495 5015
rect 38615 4895 38660 5015
rect 38780 4895 38825 5015
rect 38945 4895 38990 5015
rect 39110 4895 39165 5015
rect 39285 4895 39330 5015
rect 39450 4895 39495 5015
rect 39615 4895 39660 5015
rect 39780 4895 39835 5015
rect 39955 4895 40000 5015
rect 40120 4895 40165 5015
rect 40285 4895 40330 5015
rect 40450 4895 40505 5015
rect 40625 4895 40670 5015
rect 40790 4895 40835 5015
rect 40955 4895 41000 5015
rect 41120 4895 41175 5015
rect 41295 4895 41340 5015
rect 41460 4895 41505 5015
rect 41625 4895 41670 5015
rect 41790 4895 41845 5015
rect 41965 4895 41975 5015
rect 36475 4850 41975 4895
rect 36475 4730 36485 4850
rect 36605 4730 36650 4850
rect 36770 4730 36815 4850
rect 36935 4730 36980 4850
rect 37100 4730 37155 4850
rect 37275 4730 37320 4850
rect 37440 4730 37485 4850
rect 37605 4730 37650 4850
rect 37770 4730 37825 4850
rect 37945 4730 37990 4850
rect 38110 4730 38155 4850
rect 38275 4730 38320 4850
rect 38440 4730 38495 4850
rect 38615 4730 38660 4850
rect 38780 4730 38825 4850
rect 38945 4730 38990 4850
rect 39110 4730 39165 4850
rect 39285 4730 39330 4850
rect 39450 4730 39495 4850
rect 39615 4730 39660 4850
rect 39780 4730 39835 4850
rect 39955 4730 40000 4850
rect 40120 4730 40165 4850
rect 40285 4730 40330 4850
rect 40450 4730 40505 4850
rect 40625 4730 40670 4850
rect 40790 4730 40835 4850
rect 40955 4730 41000 4850
rect 41120 4730 41175 4850
rect 41295 4730 41340 4850
rect 41460 4730 41505 4850
rect 41625 4730 41670 4850
rect 41790 4730 41845 4850
rect 41965 4730 41975 4850
rect 36475 4685 41975 4730
rect 36475 4565 36485 4685
rect 36605 4565 36650 4685
rect 36770 4565 36815 4685
rect 36935 4565 36980 4685
rect 37100 4565 37155 4685
rect 37275 4565 37320 4685
rect 37440 4565 37485 4685
rect 37605 4565 37650 4685
rect 37770 4565 37825 4685
rect 37945 4565 37990 4685
rect 38110 4565 38155 4685
rect 38275 4565 38320 4685
rect 38440 4565 38495 4685
rect 38615 4565 38660 4685
rect 38780 4565 38825 4685
rect 38945 4565 38990 4685
rect 39110 4565 39165 4685
rect 39285 4565 39330 4685
rect 39450 4565 39495 4685
rect 39615 4565 39660 4685
rect 39780 4565 39835 4685
rect 39955 4565 40000 4685
rect 40120 4565 40165 4685
rect 40285 4565 40330 4685
rect 40450 4565 40505 4685
rect 40625 4565 40670 4685
rect 40790 4565 40835 4685
rect 40955 4565 41000 4685
rect 41120 4565 41175 4685
rect 41295 4565 41340 4685
rect 41460 4565 41505 4685
rect 41625 4565 41670 4685
rect 41790 4565 41845 4685
rect 41965 4565 41975 4685
rect 36475 4520 41975 4565
rect 36475 4400 36485 4520
rect 36605 4400 36650 4520
rect 36770 4400 36815 4520
rect 36935 4400 36980 4520
rect 37100 4400 37155 4520
rect 37275 4400 37320 4520
rect 37440 4400 37485 4520
rect 37605 4400 37650 4520
rect 37770 4400 37825 4520
rect 37945 4400 37990 4520
rect 38110 4400 38155 4520
rect 38275 4400 38320 4520
rect 38440 4400 38495 4520
rect 38615 4400 38660 4520
rect 38780 4400 38825 4520
rect 38945 4400 38990 4520
rect 39110 4400 39165 4520
rect 39285 4400 39330 4520
rect 39450 4400 39495 4520
rect 39615 4400 39660 4520
rect 39780 4400 39835 4520
rect 39955 4400 40000 4520
rect 40120 4400 40165 4520
rect 40285 4400 40330 4520
rect 40450 4400 40505 4520
rect 40625 4400 40670 4520
rect 40790 4400 40835 4520
rect 40955 4400 41000 4520
rect 41120 4400 41175 4520
rect 41295 4400 41340 4520
rect 41460 4400 41505 4520
rect 41625 4400 41670 4520
rect 41790 4400 41845 4520
rect 41965 4400 41975 4520
rect 36475 4345 41975 4400
rect 36475 4225 36485 4345
rect 36605 4225 36650 4345
rect 36770 4225 36815 4345
rect 36935 4225 36980 4345
rect 37100 4225 37155 4345
rect 37275 4225 37320 4345
rect 37440 4225 37485 4345
rect 37605 4225 37650 4345
rect 37770 4225 37825 4345
rect 37945 4225 37990 4345
rect 38110 4225 38155 4345
rect 38275 4225 38320 4345
rect 38440 4225 38495 4345
rect 38615 4225 38660 4345
rect 38780 4225 38825 4345
rect 38945 4225 38990 4345
rect 39110 4225 39165 4345
rect 39285 4225 39330 4345
rect 39450 4225 39495 4345
rect 39615 4225 39660 4345
rect 39780 4225 39835 4345
rect 39955 4225 40000 4345
rect 40120 4225 40165 4345
rect 40285 4225 40330 4345
rect 40450 4225 40505 4345
rect 40625 4225 40670 4345
rect 40790 4225 40835 4345
rect 40955 4225 41000 4345
rect 41120 4225 41175 4345
rect 41295 4225 41340 4345
rect 41460 4225 41505 4345
rect 41625 4225 41670 4345
rect 41790 4225 41845 4345
rect 41965 4225 41975 4345
rect 36475 4180 41975 4225
rect 36475 4060 36485 4180
rect 36605 4060 36650 4180
rect 36770 4060 36815 4180
rect 36935 4060 36980 4180
rect 37100 4060 37155 4180
rect 37275 4060 37320 4180
rect 37440 4060 37485 4180
rect 37605 4060 37650 4180
rect 37770 4060 37825 4180
rect 37945 4060 37990 4180
rect 38110 4060 38155 4180
rect 38275 4060 38320 4180
rect 38440 4060 38495 4180
rect 38615 4060 38660 4180
rect 38780 4060 38825 4180
rect 38945 4060 38990 4180
rect 39110 4060 39165 4180
rect 39285 4060 39330 4180
rect 39450 4060 39495 4180
rect 39615 4060 39660 4180
rect 39780 4060 39835 4180
rect 39955 4060 40000 4180
rect 40120 4060 40165 4180
rect 40285 4060 40330 4180
rect 40450 4060 40505 4180
rect 40625 4060 40670 4180
rect 40790 4060 40835 4180
rect 40955 4060 41000 4180
rect 41120 4060 41175 4180
rect 41295 4060 41340 4180
rect 41460 4060 41505 4180
rect 41625 4060 41670 4180
rect 41790 4060 41845 4180
rect 41965 4060 41975 4180
rect 36475 4015 41975 4060
rect 36475 3895 36485 4015
rect 36605 3895 36650 4015
rect 36770 3895 36815 4015
rect 36935 3895 36980 4015
rect 37100 3895 37155 4015
rect 37275 3895 37320 4015
rect 37440 3895 37485 4015
rect 37605 3895 37650 4015
rect 37770 3895 37825 4015
rect 37945 3895 37990 4015
rect 38110 3895 38155 4015
rect 38275 3895 38320 4015
rect 38440 3895 38495 4015
rect 38615 3895 38660 4015
rect 38780 3895 38825 4015
rect 38945 3895 38990 4015
rect 39110 3895 39165 4015
rect 39285 3895 39330 4015
rect 39450 3895 39495 4015
rect 39615 3895 39660 4015
rect 39780 3895 39835 4015
rect 39955 3895 40000 4015
rect 40120 3895 40165 4015
rect 40285 3895 40330 4015
rect 40450 3895 40505 4015
rect 40625 3895 40670 4015
rect 40790 3895 40835 4015
rect 40955 3895 41000 4015
rect 41120 3895 41175 4015
rect 41295 3895 41340 4015
rect 41460 3895 41505 4015
rect 41625 3895 41670 4015
rect 41790 3895 41845 4015
rect 41965 3895 41975 4015
rect 36475 3850 41975 3895
rect 36475 3730 36485 3850
rect 36605 3730 36650 3850
rect 36770 3730 36815 3850
rect 36935 3730 36980 3850
rect 37100 3730 37155 3850
rect 37275 3730 37320 3850
rect 37440 3730 37485 3850
rect 37605 3730 37650 3850
rect 37770 3730 37825 3850
rect 37945 3730 37990 3850
rect 38110 3730 38155 3850
rect 38275 3730 38320 3850
rect 38440 3730 38495 3850
rect 38615 3730 38660 3850
rect 38780 3730 38825 3850
rect 38945 3730 38990 3850
rect 39110 3730 39165 3850
rect 39285 3730 39330 3850
rect 39450 3730 39495 3850
rect 39615 3730 39660 3850
rect 39780 3730 39835 3850
rect 39955 3730 40000 3850
rect 40120 3730 40165 3850
rect 40285 3730 40330 3850
rect 40450 3730 40505 3850
rect 40625 3730 40670 3850
rect 40790 3730 40835 3850
rect 40955 3730 41000 3850
rect 41120 3730 41175 3850
rect 41295 3730 41340 3850
rect 41460 3730 41505 3850
rect 41625 3730 41670 3850
rect 41790 3730 41845 3850
rect 41965 3730 41975 3850
rect 36475 3675 41975 3730
rect 36475 3555 36485 3675
rect 36605 3555 36650 3675
rect 36770 3555 36815 3675
rect 36935 3555 36980 3675
rect 37100 3555 37155 3675
rect 37275 3555 37320 3675
rect 37440 3555 37485 3675
rect 37605 3555 37650 3675
rect 37770 3555 37825 3675
rect 37945 3555 37990 3675
rect 38110 3555 38155 3675
rect 38275 3555 38320 3675
rect 38440 3555 38495 3675
rect 38615 3555 38660 3675
rect 38780 3555 38825 3675
rect 38945 3555 38990 3675
rect 39110 3555 39165 3675
rect 39285 3555 39330 3675
rect 39450 3555 39495 3675
rect 39615 3555 39660 3675
rect 39780 3555 39835 3675
rect 39955 3555 40000 3675
rect 40120 3555 40165 3675
rect 40285 3555 40330 3675
rect 40450 3555 40505 3675
rect 40625 3555 40670 3675
rect 40790 3555 40835 3675
rect 40955 3555 41000 3675
rect 41120 3555 41175 3675
rect 41295 3555 41340 3675
rect 41460 3555 41505 3675
rect 41625 3555 41670 3675
rect 41790 3555 41845 3675
rect 41965 3555 41975 3675
rect 36475 3510 41975 3555
rect 36475 3390 36485 3510
rect 36605 3390 36650 3510
rect 36770 3390 36815 3510
rect 36935 3390 36980 3510
rect 37100 3390 37155 3510
rect 37275 3390 37320 3510
rect 37440 3390 37485 3510
rect 37605 3390 37650 3510
rect 37770 3390 37825 3510
rect 37945 3390 37990 3510
rect 38110 3390 38155 3510
rect 38275 3390 38320 3510
rect 38440 3390 38495 3510
rect 38615 3390 38660 3510
rect 38780 3390 38825 3510
rect 38945 3390 38990 3510
rect 39110 3390 39165 3510
rect 39285 3390 39330 3510
rect 39450 3390 39495 3510
rect 39615 3390 39660 3510
rect 39780 3390 39835 3510
rect 39955 3390 40000 3510
rect 40120 3390 40165 3510
rect 40285 3390 40330 3510
rect 40450 3390 40505 3510
rect 40625 3390 40670 3510
rect 40790 3390 40835 3510
rect 40955 3390 41000 3510
rect 41120 3390 41175 3510
rect 41295 3390 41340 3510
rect 41460 3390 41505 3510
rect 41625 3390 41670 3510
rect 41790 3390 41845 3510
rect 41965 3390 41975 3510
rect 36475 3345 41975 3390
rect 36475 3225 36485 3345
rect 36605 3225 36650 3345
rect 36770 3225 36815 3345
rect 36935 3225 36980 3345
rect 37100 3225 37155 3345
rect 37275 3225 37320 3345
rect 37440 3225 37485 3345
rect 37605 3225 37650 3345
rect 37770 3225 37825 3345
rect 37945 3225 37990 3345
rect 38110 3225 38155 3345
rect 38275 3225 38320 3345
rect 38440 3225 38495 3345
rect 38615 3225 38660 3345
rect 38780 3225 38825 3345
rect 38945 3225 38990 3345
rect 39110 3225 39165 3345
rect 39285 3225 39330 3345
rect 39450 3225 39495 3345
rect 39615 3225 39660 3345
rect 39780 3225 39835 3345
rect 39955 3225 40000 3345
rect 40120 3225 40165 3345
rect 40285 3225 40330 3345
rect 40450 3225 40505 3345
rect 40625 3225 40670 3345
rect 40790 3225 40835 3345
rect 40955 3225 41000 3345
rect 41120 3225 41175 3345
rect 41295 3225 41340 3345
rect 41460 3225 41505 3345
rect 41625 3225 41670 3345
rect 41790 3225 41845 3345
rect 41965 3225 41975 3345
rect 36475 3180 41975 3225
rect 36475 3060 36485 3180
rect 36605 3060 36650 3180
rect 36770 3060 36815 3180
rect 36935 3060 36980 3180
rect 37100 3060 37155 3180
rect 37275 3060 37320 3180
rect 37440 3060 37485 3180
rect 37605 3060 37650 3180
rect 37770 3060 37825 3180
rect 37945 3060 37990 3180
rect 38110 3060 38155 3180
rect 38275 3060 38320 3180
rect 38440 3060 38495 3180
rect 38615 3060 38660 3180
rect 38780 3060 38825 3180
rect 38945 3060 38990 3180
rect 39110 3060 39165 3180
rect 39285 3060 39330 3180
rect 39450 3060 39495 3180
rect 39615 3060 39660 3180
rect 39780 3060 39835 3180
rect 39955 3060 40000 3180
rect 40120 3060 40165 3180
rect 40285 3060 40330 3180
rect 40450 3060 40505 3180
rect 40625 3060 40670 3180
rect 40790 3060 40835 3180
rect 40955 3060 41000 3180
rect 41120 3060 41175 3180
rect 41295 3060 41340 3180
rect 41460 3060 41505 3180
rect 41625 3060 41670 3180
rect 41790 3060 41845 3180
rect 41965 3060 41975 3180
rect 36475 3005 41975 3060
rect 36475 2885 36485 3005
rect 36605 2885 36650 3005
rect 36770 2885 36815 3005
rect 36935 2885 36980 3005
rect 37100 2885 37155 3005
rect 37275 2885 37320 3005
rect 37440 2885 37485 3005
rect 37605 2885 37650 3005
rect 37770 2885 37825 3005
rect 37945 2885 37990 3005
rect 38110 2885 38155 3005
rect 38275 2885 38320 3005
rect 38440 2885 38495 3005
rect 38615 2885 38660 3005
rect 38780 2885 38825 3005
rect 38945 2885 38990 3005
rect 39110 2885 39165 3005
rect 39285 2885 39330 3005
rect 39450 2885 39495 3005
rect 39615 2885 39660 3005
rect 39780 2885 39835 3005
rect 39955 2885 40000 3005
rect 40120 2885 40165 3005
rect 40285 2885 40330 3005
rect 40450 2885 40505 3005
rect 40625 2885 40670 3005
rect 40790 2885 40835 3005
rect 40955 2885 41000 3005
rect 41120 2885 41175 3005
rect 41295 2885 41340 3005
rect 41460 2885 41505 3005
rect 41625 2885 41670 3005
rect 41790 2885 41845 3005
rect 41965 2885 41975 3005
rect 36475 2840 41975 2885
rect 36475 2720 36485 2840
rect 36605 2720 36650 2840
rect 36770 2720 36815 2840
rect 36935 2720 36980 2840
rect 37100 2720 37155 2840
rect 37275 2720 37320 2840
rect 37440 2720 37485 2840
rect 37605 2720 37650 2840
rect 37770 2720 37825 2840
rect 37945 2720 37990 2840
rect 38110 2720 38155 2840
rect 38275 2720 38320 2840
rect 38440 2720 38495 2840
rect 38615 2720 38660 2840
rect 38780 2720 38825 2840
rect 38945 2720 38990 2840
rect 39110 2720 39165 2840
rect 39285 2720 39330 2840
rect 39450 2720 39495 2840
rect 39615 2720 39660 2840
rect 39780 2720 39835 2840
rect 39955 2720 40000 2840
rect 40120 2720 40165 2840
rect 40285 2720 40330 2840
rect 40450 2720 40505 2840
rect 40625 2720 40670 2840
rect 40790 2720 40835 2840
rect 40955 2720 41000 2840
rect 41120 2720 41175 2840
rect 41295 2720 41340 2840
rect 41460 2720 41505 2840
rect 41625 2720 41670 2840
rect 41790 2720 41845 2840
rect 41965 2720 41975 2840
rect 36475 2675 41975 2720
rect 36475 2555 36485 2675
rect 36605 2555 36650 2675
rect 36770 2555 36815 2675
rect 36935 2555 36980 2675
rect 37100 2555 37155 2675
rect 37275 2555 37320 2675
rect 37440 2555 37485 2675
rect 37605 2555 37650 2675
rect 37770 2555 37825 2675
rect 37945 2555 37990 2675
rect 38110 2555 38155 2675
rect 38275 2555 38320 2675
rect 38440 2555 38495 2675
rect 38615 2555 38660 2675
rect 38780 2555 38825 2675
rect 38945 2555 38990 2675
rect 39110 2555 39165 2675
rect 39285 2555 39330 2675
rect 39450 2555 39495 2675
rect 39615 2555 39660 2675
rect 39780 2555 39835 2675
rect 39955 2555 40000 2675
rect 40120 2555 40165 2675
rect 40285 2555 40330 2675
rect 40450 2555 40505 2675
rect 40625 2555 40670 2675
rect 40790 2555 40835 2675
rect 40955 2555 41000 2675
rect 41120 2555 41175 2675
rect 41295 2555 41340 2675
rect 41460 2555 41505 2675
rect 41625 2555 41670 2675
rect 41790 2555 41845 2675
rect 41965 2555 41975 2675
rect 36475 2510 41975 2555
rect 36475 2390 36485 2510
rect 36605 2390 36650 2510
rect 36770 2390 36815 2510
rect 36935 2390 36980 2510
rect 37100 2390 37155 2510
rect 37275 2390 37320 2510
rect 37440 2390 37485 2510
rect 37605 2390 37650 2510
rect 37770 2390 37825 2510
rect 37945 2390 37990 2510
rect 38110 2390 38155 2510
rect 38275 2390 38320 2510
rect 38440 2390 38495 2510
rect 38615 2390 38660 2510
rect 38780 2390 38825 2510
rect 38945 2390 38990 2510
rect 39110 2390 39165 2510
rect 39285 2390 39330 2510
rect 39450 2390 39495 2510
rect 39615 2390 39660 2510
rect 39780 2390 39835 2510
rect 39955 2390 40000 2510
rect 40120 2390 40165 2510
rect 40285 2390 40330 2510
rect 40450 2390 40505 2510
rect 40625 2390 40670 2510
rect 40790 2390 40835 2510
rect 40955 2390 41000 2510
rect 41120 2390 41175 2510
rect 41295 2390 41340 2510
rect 41460 2390 41505 2510
rect 41625 2390 41670 2510
rect 41790 2390 41845 2510
rect 41965 2390 41975 2510
rect 36475 2335 41975 2390
rect 36475 2215 36485 2335
rect 36605 2215 36650 2335
rect 36770 2215 36815 2335
rect 36935 2215 36980 2335
rect 37100 2215 37155 2335
rect 37275 2215 37320 2335
rect 37440 2215 37485 2335
rect 37605 2215 37650 2335
rect 37770 2215 37825 2335
rect 37945 2215 37990 2335
rect 38110 2215 38155 2335
rect 38275 2215 38320 2335
rect 38440 2215 38495 2335
rect 38615 2215 38660 2335
rect 38780 2215 38825 2335
rect 38945 2215 38990 2335
rect 39110 2215 39165 2335
rect 39285 2215 39330 2335
rect 39450 2215 39495 2335
rect 39615 2215 39660 2335
rect 39780 2215 39835 2335
rect 39955 2215 40000 2335
rect 40120 2215 40165 2335
rect 40285 2215 40330 2335
rect 40450 2215 40505 2335
rect 40625 2215 40670 2335
rect 40790 2215 40835 2335
rect 40955 2215 41000 2335
rect 41120 2215 41175 2335
rect 41295 2215 41340 2335
rect 41460 2215 41505 2335
rect 41625 2215 41670 2335
rect 41790 2215 41845 2335
rect 41965 2215 41975 2335
rect 36475 2170 41975 2215
rect 36475 2050 36485 2170
rect 36605 2050 36650 2170
rect 36770 2050 36815 2170
rect 36935 2050 36980 2170
rect 37100 2050 37155 2170
rect 37275 2050 37320 2170
rect 37440 2050 37485 2170
rect 37605 2050 37650 2170
rect 37770 2050 37825 2170
rect 37945 2050 37990 2170
rect 38110 2050 38155 2170
rect 38275 2050 38320 2170
rect 38440 2050 38495 2170
rect 38615 2050 38660 2170
rect 38780 2050 38825 2170
rect 38945 2050 38990 2170
rect 39110 2050 39165 2170
rect 39285 2050 39330 2170
rect 39450 2050 39495 2170
rect 39615 2050 39660 2170
rect 39780 2050 39835 2170
rect 39955 2050 40000 2170
rect 40120 2050 40165 2170
rect 40285 2050 40330 2170
rect 40450 2050 40505 2170
rect 40625 2050 40670 2170
rect 40790 2050 40835 2170
rect 40955 2050 41000 2170
rect 41120 2050 41175 2170
rect 41295 2050 41340 2170
rect 41460 2050 41505 2170
rect 41625 2050 41670 2170
rect 41790 2050 41845 2170
rect 41965 2050 41975 2170
rect 36475 2005 41975 2050
rect 36475 1885 36485 2005
rect 36605 1885 36650 2005
rect 36770 1885 36815 2005
rect 36935 1885 36980 2005
rect 37100 1885 37155 2005
rect 37275 1885 37320 2005
rect 37440 1885 37485 2005
rect 37605 1885 37650 2005
rect 37770 1885 37825 2005
rect 37945 1885 37990 2005
rect 38110 1885 38155 2005
rect 38275 1885 38320 2005
rect 38440 1885 38495 2005
rect 38615 1885 38660 2005
rect 38780 1885 38825 2005
rect 38945 1885 38990 2005
rect 39110 1885 39165 2005
rect 39285 1885 39330 2005
rect 39450 1885 39495 2005
rect 39615 1885 39660 2005
rect 39780 1885 39835 2005
rect 39955 1885 40000 2005
rect 40120 1885 40165 2005
rect 40285 1885 40330 2005
rect 40450 1885 40505 2005
rect 40625 1885 40670 2005
rect 40790 1885 40835 2005
rect 40955 1885 41000 2005
rect 41120 1885 41175 2005
rect 41295 1885 41340 2005
rect 41460 1885 41505 2005
rect 41625 1885 41670 2005
rect 41790 1885 41845 2005
rect 41965 1885 41975 2005
rect 36475 1840 41975 1885
rect 36475 1720 36485 1840
rect 36605 1720 36650 1840
rect 36770 1720 36815 1840
rect 36935 1720 36980 1840
rect 37100 1720 37155 1840
rect 37275 1720 37320 1840
rect 37440 1720 37485 1840
rect 37605 1720 37650 1840
rect 37770 1720 37825 1840
rect 37945 1720 37990 1840
rect 38110 1720 38155 1840
rect 38275 1720 38320 1840
rect 38440 1720 38495 1840
rect 38615 1720 38660 1840
rect 38780 1720 38825 1840
rect 38945 1720 38990 1840
rect 39110 1720 39165 1840
rect 39285 1720 39330 1840
rect 39450 1720 39495 1840
rect 39615 1720 39660 1840
rect 39780 1720 39835 1840
rect 39955 1720 40000 1840
rect 40120 1720 40165 1840
rect 40285 1720 40330 1840
rect 40450 1720 40505 1840
rect 40625 1720 40670 1840
rect 40790 1720 40835 1840
rect 40955 1720 41000 1840
rect 41120 1720 41175 1840
rect 41295 1720 41340 1840
rect 41460 1720 41505 1840
rect 41625 1720 41670 1840
rect 41790 1720 41845 1840
rect 41965 1720 41975 1840
rect 36475 1710 41975 1720
rect 42165 7200 47665 7210
rect 42165 7080 42175 7200
rect 42295 7080 42340 7200
rect 42460 7080 42505 7200
rect 42625 7080 42670 7200
rect 42790 7080 42845 7200
rect 42965 7080 43010 7200
rect 43130 7080 43175 7200
rect 43295 7080 43340 7200
rect 43460 7080 43515 7200
rect 43635 7080 43680 7200
rect 43800 7080 43845 7200
rect 43965 7080 44010 7200
rect 44130 7080 44185 7200
rect 44305 7080 44350 7200
rect 44470 7080 44515 7200
rect 44635 7080 44680 7200
rect 44800 7080 44855 7200
rect 44975 7080 45020 7200
rect 45140 7080 45185 7200
rect 45305 7080 45350 7200
rect 45470 7080 45525 7200
rect 45645 7080 45690 7200
rect 45810 7080 45855 7200
rect 45975 7080 46020 7200
rect 46140 7080 46195 7200
rect 46315 7080 46360 7200
rect 46480 7080 46525 7200
rect 46645 7080 46690 7200
rect 46810 7080 46865 7200
rect 46985 7080 47030 7200
rect 47150 7080 47195 7200
rect 47315 7080 47360 7200
rect 47480 7080 47535 7200
rect 47655 7080 47665 7200
rect 42165 7025 47665 7080
rect 42165 6905 42175 7025
rect 42295 6905 42340 7025
rect 42460 6905 42505 7025
rect 42625 6905 42670 7025
rect 42790 6905 42845 7025
rect 42965 6905 43010 7025
rect 43130 6905 43175 7025
rect 43295 6905 43340 7025
rect 43460 6905 43515 7025
rect 43635 6905 43680 7025
rect 43800 6905 43845 7025
rect 43965 6905 44010 7025
rect 44130 6905 44185 7025
rect 44305 6905 44350 7025
rect 44470 6905 44515 7025
rect 44635 6905 44680 7025
rect 44800 6905 44855 7025
rect 44975 6905 45020 7025
rect 45140 6905 45185 7025
rect 45305 6905 45350 7025
rect 45470 6905 45525 7025
rect 45645 6905 45690 7025
rect 45810 6905 45855 7025
rect 45975 6905 46020 7025
rect 46140 6905 46195 7025
rect 46315 6905 46360 7025
rect 46480 6905 46525 7025
rect 46645 6905 46690 7025
rect 46810 6905 46865 7025
rect 46985 6905 47030 7025
rect 47150 6905 47195 7025
rect 47315 6905 47360 7025
rect 47480 6905 47535 7025
rect 47655 6905 47665 7025
rect 42165 6860 47665 6905
rect 42165 6740 42175 6860
rect 42295 6740 42340 6860
rect 42460 6740 42505 6860
rect 42625 6740 42670 6860
rect 42790 6740 42845 6860
rect 42965 6740 43010 6860
rect 43130 6740 43175 6860
rect 43295 6740 43340 6860
rect 43460 6740 43515 6860
rect 43635 6740 43680 6860
rect 43800 6740 43845 6860
rect 43965 6740 44010 6860
rect 44130 6740 44185 6860
rect 44305 6740 44350 6860
rect 44470 6740 44515 6860
rect 44635 6740 44680 6860
rect 44800 6740 44855 6860
rect 44975 6740 45020 6860
rect 45140 6740 45185 6860
rect 45305 6740 45350 6860
rect 45470 6740 45525 6860
rect 45645 6740 45690 6860
rect 45810 6740 45855 6860
rect 45975 6740 46020 6860
rect 46140 6740 46195 6860
rect 46315 6740 46360 6860
rect 46480 6740 46525 6860
rect 46645 6740 46690 6860
rect 46810 6740 46865 6860
rect 46985 6740 47030 6860
rect 47150 6740 47195 6860
rect 47315 6740 47360 6860
rect 47480 6740 47535 6860
rect 47655 6740 47665 6860
rect 42165 6695 47665 6740
rect 42165 6575 42175 6695
rect 42295 6575 42340 6695
rect 42460 6575 42505 6695
rect 42625 6575 42670 6695
rect 42790 6575 42845 6695
rect 42965 6575 43010 6695
rect 43130 6575 43175 6695
rect 43295 6575 43340 6695
rect 43460 6575 43515 6695
rect 43635 6575 43680 6695
rect 43800 6575 43845 6695
rect 43965 6575 44010 6695
rect 44130 6575 44185 6695
rect 44305 6575 44350 6695
rect 44470 6575 44515 6695
rect 44635 6575 44680 6695
rect 44800 6575 44855 6695
rect 44975 6575 45020 6695
rect 45140 6575 45185 6695
rect 45305 6575 45350 6695
rect 45470 6575 45525 6695
rect 45645 6575 45690 6695
rect 45810 6575 45855 6695
rect 45975 6575 46020 6695
rect 46140 6575 46195 6695
rect 46315 6575 46360 6695
rect 46480 6575 46525 6695
rect 46645 6575 46690 6695
rect 46810 6575 46865 6695
rect 46985 6575 47030 6695
rect 47150 6575 47195 6695
rect 47315 6575 47360 6695
rect 47480 6575 47535 6695
rect 47655 6575 47665 6695
rect 42165 6530 47665 6575
rect 42165 6410 42175 6530
rect 42295 6410 42340 6530
rect 42460 6410 42505 6530
rect 42625 6410 42670 6530
rect 42790 6410 42845 6530
rect 42965 6410 43010 6530
rect 43130 6410 43175 6530
rect 43295 6410 43340 6530
rect 43460 6410 43515 6530
rect 43635 6410 43680 6530
rect 43800 6410 43845 6530
rect 43965 6410 44010 6530
rect 44130 6410 44185 6530
rect 44305 6410 44350 6530
rect 44470 6410 44515 6530
rect 44635 6410 44680 6530
rect 44800 6410 44855 6530
rect 44975 6410 45020 6530
rect 45140 6410 45185 6530
rect 45305 6410 45350 6530
rect 45470 6410 45525 6530
rect 45645 6410 45690 6530
rect 45810 6410 45855 6530
rect 45975 6410 46020 6530
rect 46140 6410 46195 6530
rect 46315 6410 46360 6530
rect 46480 6410 46525 6530
rect 46645 6410 46690 6530
rect 46810 6410 46865 6530
rect 46985 6410 47030 6530
rect 47150 6410 47195 6530
rect 47315 6410 47360 6530
rect 47480 6410 47535 6530
rect 47655 6410 47665 6530
rect 42165 6355 47665 6410
rect 42165 6235 42175 6355
rect 42295 6235 42340 6355
rect 42460 6235 42505 6355
rect 42625 6235 42670 6355
rect 42790 6235 42845 6355
rect 42965 6235 43010 6355
rect 43130 6235 43175 6355
rect 43295 6235 43340 6355
rect 43460 6235 43515 6355
rect 43635 6235 43680 6355
rect 43800 6235 43845 6355
rect 43965 6235 44010 6355
rect 44130 6235 44185 6355
rect 44305 6235 44350 6355
rect 44470 6235 44515 6355
rect 44635 6235 44680 6355
rect 44800 6235 44855 6355
rect 44975 6235 45020 6355
rect 45140 6235 45185 6355
rect 45305 6235 45350 6355
rect 45470 6235 45525 6355
rect 45645 6235 45690 6355
rect 45810 6235 45855 6355
rect 45975 6235 46020 6355
rect 46140 6235 46195 6355
rect 46315 6235 46360 6355
rect 46480 6235 46525 6355
rect 46645 6235 46690 6355
rect 46810 6235 46865 6355
rect 46985 6235 47030 6355
rect 47150 6235 47195 6355
rect 47315 6235 47360 6355
rect 47480 6235 47535 6355
rect 47655 6235 47665 6355
rect 42165 6190 47665 6235
rect 42165 6070 42175 6190
rect 42295 6070 42340 6190
rect 42460 6070 42505 6190
rect 42625 6070 42670 6190
rect 42790 6070 42845 6190
rect 42965 6070 43010 6190
rect 43130 6070 43175 6190
rect 43295 6070 43340 6190
rect 43460 6070 43515 6190
rect 43635 6070 43680 6190
rect 43800 6070 43845 6190
rect 43965 6070 44010 6190
rect 44130 6070 44185 6190
rect 44305 6070 44350 6190
rect 44470 6070 44515 6190
rect 44635 6070 44680 6190
rect 44800 6070 44855 6190
rect 44975 6070 45020 6190
rect 45140 6070 45185 6190
rect 45305 6070 45350 6190
rect 45470 6070 45525 6190
rect 45645 6070 45690 6190
rect 45810 6070 45855 6190
rect 45975 6070 46020 6190
rect 46140 6070 46195 6190
rect 46315 6070 46360 6190
rect 46480 6070 46525 6190
rect 46645 6070 46690 6190
rect 46810 6070 46865 6190
rect 46985 6070 47030 6190
rect 47150 6070 47195 6190
rect 47315 6070 47360 6190
rect 47480 6070 47535 6190
rect 47655 6070 47665 6190
rect 42165 6025 47665 6070
rect 42165 5905 42175 6025
rect 42295 5905 42340 6025
rect 42460 5905 42505 6025
rect 42625 5905 42670 6025
rect 42790 5905 42845 6025
rect 42965 5905 43010 6025
rect 43130 5905 43175 6025
rect 43295 5905 43340 6025
rect 43460 5905 43515 6025
rect 43635 5905 43680 6025
rect 43800 5905 43845 6025
rect 43965 5905 44010 6025
rect 44130 5905 44185 6025
rect 44305 5905 44350 6025
rect 44470 5905 44515 6025
rect 44635 5905 44680 6025
rect 44800 5905 44855 6025
rect 44975 5905 45020 6025
rect 45140 5905 45185 6025
rect 45305 5905 45350 6025
rect 45470 5905 45525 6025
rect 45645 5905 45690 6025
rect 45810 5905 45855 6025
rect 45975 5905 46020 6025
rect 46140 5905 46195 6025
rect 46315 5905 46360 6025
rect 46480 5905 46525 6025
rect 46645 5905 46690 6025
rect 46810 5905 46865 6025
rect 46985 5905 47030 6025
rect 47150 5905 47195 6025
rect 47315 5905 47360 6025
rect 47480 5905 47535 6025
rect 47655 5905 47665 6025
rect 42165 5860 47665 5905
rect 42165 5740 42175 5860
rect 42295 5740 42340 5860
rect 42460 5740 42505 5860
rect 42625 5740 42670 5860
rect 42790 5740 42845 5860
rect 42965 5740 43010 5860
rect 43130 5740 43175 5860
rect 43295 5740 43340 5860
rect 43460 5740 43515 5860
rect 43635 5740 43680 5860
rect 43800 5740 43845 5860
rect 43965 5740 44010 5860
rect 44130 5740 44185 5860
rect 44305 5740 44350 5860
rect 44470 5740 44515 5860
rect 44635 5740 44680 5860
rect 44800 5740 44855 5860
rect 44975 5740 45020 5860
rect 45140 5740 45185 5860
rect 45305 5740 45350 5860
rect 45470 5740 45525 5860
rect 45645 5740 45690 5860
rect 45810 5740 45855 5860
rect 45975 5740 46020 5860
rect 46140 5740 46195 5860
rect 46315 5740 46360 5860
rect 46480 5740 46525 5860
rect 46645 5740 46690 5860
rect 46810 5740 46865 5860
rect 46985 5740 47030 5860
rect 47150 5740 47195 5860
rect 47315 5740 47360 5860
rect 47480 5740 47535 5860
rect 47655 5740 47665 5860
rect 42165 5685 47665 5740
rect 42165 5565 42175 5685
rect 42295 5565 42340 5685
rect 42460 5565 42505 5685
rect 42625 5565 42670 5685
rect 42790 5565 42845 5685
rect 42965 5565 43010 5685
rect 43130 5565 43175 5685
rect 43295 5565 43340 5685
rect 43460 5565 43515 5685
rect 43635 5565 43680 5685
rect 43800 5565 43845 5685
rect 43965 5565 44010 5685
rect 44130 5565 44185 5685
rect 44305 5565 44350 5685
rect 44470 5565 44515 5685
rect 44635 5565 44680 5685
rect 44800 5565 44855 5685
rect 44975 5565 45020 5685
rect 45140 5565 45185 5685
rect 45305 5565 45350 5685
rect 45470 5565 45525 5685
rect 45645 5565 45690 5685
rect 45810 5565 45855 5685
rect 45975 5565 46020 5685
rect 46140 5565 46195 5685
rect 46315 5565 46360 5685
rect 46480 5565 46525 5685
rect 46645 5565 46690 5685
rect 46810 5565 46865 5685
rect 46985 5565 47030 5685
rect 47150 5565 47195 5685
rect 47315 5565 47360 5685
rect 47480 5565 47535 5685
rect 47655 5565 47665 5685
rect 42165 5520 47665 5565
rect 42165 5400 42175 5520
rect 42295 5400 42340 5520
rect 42460 5400 42505 5520
rect 42625 5400 42670 5520
rect 42790 5400 42845 5520
rect 42965 5400 43010 5520
rect 43130 5400 43175 5520
rect 43295 5400 43340 5520
rect 43460 5400 43515 5520
rect 43635 5400 43680 5520
rect 43800 5400 43845 5520
rect 43965 5400 44010 5520
rect 44130 5400 44185 5520
rect 44305 5400 44350 5520
rect 44470 5400 44515 5520
rect 44635 5400 44680 5520
rect 44800 5400 44855 5520
rect 44975 5400 45020 5520
rect 45140 5400 45185 5520
rect 45305 5400 45350 5520
rect 45470 5400 45525 5520
rect 45645 5400 45690 5520
rect 45810 5400 45855 5520
rect 45975 5400 46020 5520
rect 46140 5400 46195 5520
rect 46315 5400 46360 5520
rect 46480 5400 46525 5520
rect 46645 5400 46690 5520
rect 46810 5400 46865 5520
rect 46985 5400 47030 5520
rect 47150 5400 47195 5520
rect 47315 5400 47360 5520
rect 47480 5400 47535 5520
rect 47655 5400 47665 5520
rect 42165 5355 47665 5400
rect 42165 5235 42175 5355
rect 42295 5235 42340 5355
rect 42460 5235 42505 5355
rect 42625 5235 42670 5355
rect 42790 5235 42845 5355
rect 42965 5235 43010 5355
rect 43130 5235 43175 5355
rect 43295 5235 43340 5355
rect 43460 5235 43515 5355
rect 43635 5235 43680 5355
rect 43800 5235 43845 5355
rect 43965 5235 44010 5355
rect 44130 5235 44185 5355
rect 44305 5235 44350 5355
rect 44470 5235 44515 5355
rect 44635 5235 44680 5355
rect 44800 5235 44855 5355
rect 44975 5235 45020 5355
rect 45140 5235 45185 5355
rect 45305 5235 45350 5355
rect 45470 5235 45525 5355
rect 45645 5235 45690 5355
rect 45810 5235 45855 5355
rect 45975 5235 46020 5355
rect 46140 5235 46195 5355
rect 46315 5235 46360 5355
rect 46480 5235 46525 5355
rect 46645 5235 46690 5355
rect 46810 5235 46865 5355
rect 46985 5235 47030 5355
rect 47150 5235 47195 5355
rect 47315 5235 47360 5355
rect 47480 5235 47535 5355
rect 47655 5235 47665 5355
rect 42165 5190 47665 5235
rect 42165 5070 42175 5190
rect 42295 5070 42340 5190
rect 42460 5070 42505 5190
rect 42625 5070 42670 5190
rect 42790 5070 42845 5190
rect 42965 5070 43010 5190
rect 43130 5070 43175 5190
rect 43295 5070 43340 5190
rect 43460 5070 43515 5190
rect 43635 5070 43680 5190
rect 43800 5070 43845 5190
rect 43965 5070 44010 5190
rect 44130 5070 44185 5190
rect 44305 5070 44350 5190
rect 44470 5070 44515 5190
rect 44635 5070 44680 5190
rect 44800 5070 44855 5190
rect 44975 5070 45020 5190
rect 45140 5070 45185 5190
rect 45305 5070 45350 5190
rect 45470 5070 45525 5190
rect 45645 5070 45690 5190
rect 45810 5070 45855 5190
rect 45975 5070 46020 5190
rect 46140 5070 46195 5190
rect 46315 5070 46360 5190
rect 46480 5070 46525 5190
rect 46645 5070 46690 5190
rect 46810 5070 46865 5190
rect 46985 5070 47030 5190
rect 47150 5070 47195 5190
rect 47315 5070 47360 5190
rect 47480 5070 47535 5190
rect 47655 5070 47665 5190
rect 42165 5015 47665 5070
rect 42165 4895 42175 5015
rect 42295 4895 42340 5015
rect 42460 4895 42505 5015
rect 42625 4895 42670 5015
rect 42790 4895 42845 5015
rect 42965 4895 43010 5015
rect 43130 4895 43175 5015
rect 43295 4895 43340 5015
rect 43460 4895 43515 5015
rect 43635 4895 43680 5015
rect 43800 4895 43845 5015
rect 43965 4895 44010 5015
rect 44130 4895 44185 5015
rect 44305 4895 44350 5015
rect 44470 4895 44515 5015
rect 44635 4895 44680 5015
rect 44800 4895 44855 5015
rect 44975 4895 45020 5015
rect 45140 4895 45185 5015
rect 45305 4895 45350 5015
rect 45470 4895 45525 5015
rect 45645 4895 45690 5015
rect 45810 4895 45855 5015
rect 45975 4895 46020 5015
rect 46140 4895 46195 5015
rect 46315 4895 46360 5015
rect 46480 4895 46525 5015
rect 46645 4895 46690 5015
rect 46810 4895 46865 5015
rect 46985 4895 47030 5015
rect 47150 4895 47195 5015
rect 47315 4895 47360 5015
rect 47480 4895 47535 5015
rect 47655 4895 47665 5015
rect 42165 4850 47665 4895
rect 42165 4730 42175 4850
rect 42295 4730 42340 4850
rect 42460 4730 42505 4850
rect 42625 4730 42670 4850
rect 42790 4730 42845 4850
rect 42965 4730 43010 4850
rect 43130 4730 43175 4850
rect 43295 4730 43340 4850
rect 43460 4730 43515 4850
rect 43635 4730 43680 4850
rect 43800 4730 43845 4850
rect 43965 4730 44010 4850
rect 44130 4730 44185 4850
rect 44305 4730 44350 4850
rect 44470 4730 44515 4850
rect 44635 4730 44680 4850
rect 44800 4730 44855 4850
rect 44975 4730 45020 4850
rect 45140 4730 45185 4850
rect 45305 4730 45350 4850
rect 45470 4730 45525 4850
rect 45645 4730 45690 4850
rect 45810 4730 45855 4850
rect 45975 4730 46020 4850
rect 46140 4730 46195 4850
rect 46315 4730 46360 4850
rect 46480 4730 46525 4850
rect 46645 4730 46690 4850
rect 46810 4730 46865 4850
rect 46985 4730 47030 4850
rect 47150 4730 47195 4850
rect 47315 4730 47360 4850
rect 47480 4730 47535 4850
rect 47655 4730 47665 4850
rect 42165 4685 47665 4730
rect 42165 4565 42175 4685
rect 42295 4565 42340 4685
rect 42460 4565 42505 4685
rect 42625 4565 42670 4685
rect 42790 4565 42845 4685
rect 42965 4565 43010 4685
rect 43130 4565 43175 4685
rect 43295 4565 43340 4685
rect 43460 4565 43515 4685
rect 43635 4565 43680 4685
rect 43800 4565 43845 4685
rect 43965 4565 44010 4685
rect 44130 4565 44185 4685
rect 44305 4565 44350 4685
rect 44470 4565 44515 4685
rect 44635 4565 44680 4685
rect 44800 4565 44855 4685
rect 44975 4565 45020 4685
rect 45140 4565 45185 4685
rect 45305 4565 45350 4685
rect 45470 4565 45525 4685
rect 45645 4565 45690 4685
rect 45810 4565 45855 4685
rect 45975 4565 46020 4685
rect 46140 4565 46195 4685
rect 46315 4565 46360 4685
rect 46480 4565 46525 4685
rect 46645 4565 46690 4685
rect 46810 4565 46865 4685
rect 46985 4565 47030 4685
rect 47150 4565 47195 4685
rect 47315 4565 47360 4685
rect 47480 4565 47535 4685
rect 47655 4565 47665 4685
rect 42165 4520 47665 4565
rect 42165 4400 42175 4520
rect 42295 4400 42340 4520
rect 42460 4400 42505 4520
rect 42625 4400 42670 4520
rect 42790 4400 42845 4520
rect 42965 4400 43010 4520
rect 43130 4400 43175 4520
rect 43295 4400 43340 4520
rect 43460 4400 43515 4520
rect 43635 4400 43680 4520
rect 43800 4400 43845 4520
rect 43965 4400 44010 4520
rect 44130 4400 44185 4520
rect 44305 4400 44350 4520
rect 44470 4400 44515 4520
rect 44635 4400 44680 4520
rect 44800 4400 44855 4520
rect 44975 4400 45020 4520
rect 45140 4400 45185 4520
rect 45305 4400 45350 4520
rect 45470 4400 45525 4520
rect 45645 4400 45690 4520
rect 45810 4400 45855 4520
rect 45975 4400 46020 4520
rect 46140 4400 46195 4520
rect 46315 4400 46360 4520
rect 46480 4400 46525 4520
rect 46645 4400 46690 4520
rect 46810 4400 46865 4520
rect 46985 4400 47030 4520
rect 47150 4400 47195 4520
rect 47315 4400 47360 4520
rect 47480 4400 47535 4520
rect 47655 4400 47665 4520
rect 42165 4345 47665 4400
rect 42165 4225 42175 4345
rect 42295 4225 42340 4345
rect 42460 4225 42505 4345
rect 42625 4225 42670 4345
rect 42790 4225 42845 4345
rect 42965 4225 43010 4345
rect 43130 4225 43175 4345
rect 43295 4225 43340 4345
rect 43460 4225 43515 4345
rect 43635 4225 43680 4345
rect 43800 4225 43845 4345
rect 43965 4225 44010 4345
rect 44130 4225 44185 4345
rect 44305 4225 44350 4345
rect 44470 4225 44515 4345
rect 44635 4225 44680 4345
rect 44800 4225 44855 4345
rect 44975 4225 45020 4345
rect 45140 4225 45185 4345
rect 45305 4225 45350 4345
rect 45470 4225 45525 4345
rect 45645 4225 45690 4345
rect 45810 4225 45855 4345
rect 45975 4225 46020 4345
rect 46140 4225 46195 4345
rect 46315 4225 46360 4345
rect 46480 4225 46525 4345
rect 46645 4225 46690 4345
rect 46810 4225 46865 4345
rect 46985 4225 47030 4345
rect 47150 4225 47195 4345
rect 47315 4225 47360 4345
rect 47480 4225 47535 4345
rect 47655 4225 47665 4345
rect 42165 4180 47665 4225
rect 42165 4060 42175 4180
rect 42295 4060 42340 4180
rect 42460 4060 42505 4180
rect 42625 4060 42670 4180
rect 42790 4060 42845 4180
rect 42965 4060 43010 4180
rect 43130 4060 43175 4180
rect 43295 4060 43340 4180
rect 43460 4060 43515 4180
rect 43635 4060 43680 4180
rect 43800 4060 43845 4180
rect 43965 4060 44010 4180
rect 44130 4060 44185 4180
rect 44305 4060 44350 4180
rect 44470 4060 44515 4180
rect 44635 4060 44680 4180
rect 44800 4060 44855 4180
rect 44975 4060 45020 4180
rect 45140 4060 45185 4180
rect 45305 4060 45350 4180
rect 45470 4060 45525 4180
rect 45645 4060 45690 4180
rect 45810 4060 45855 4180
rect 45975 4060 46020 4180
rect 46140 4060 46195 4180
rect 46315 4060 46360 4180
rect 46480 4060 46525 4180
rect 46645 4060 46690 4180
rect 46810 4060 46865 4180
rect 46985 4060 47030 4180
rect 47150 4060 47195 4180
rect 47315 4060 47360 4180
rect 47480 4060 47535 4180
rect 47655 4060 47665 4180
rect 42165 4015 47665 4060
rect 42165 3895 42175 4015
rect 42295 3895 42340 4015
rect 42460 3895 42505 4015
rect 42625 3895 42670 4015
rect 42790 3895 42845 4015
rect 42965 3895 43010 4015
rect 43130 3895 43175 4015
rect 43295 3895 43340 4015
rect 43460 3895 43515 4015
rect 43635 3895 43680 4015
rect 43800 3895 43845 4015
rect 43965 3895 44010 4015
rect 44130 3895 44185 4015
rect 44305 3895 44350 4015
rect 44470 3895 44515 4015
rect 44635 3895 44680 4015
rect 44800 3895 44855 4015
rect 44975 3895 45020 4015
rect 45140 3895 45185 4015
rect 45305 3895 45350 4015
rect 45470 3895 45525 4015
rect 45645 3895 45690 4015
rect 45810 3895 45855 4015
rect 45975 3895 46020 4015
rect 46140 3895 46195 4015
rect 46315 3895 46360 4015
rect 46480 3895 46525 4015
rect 46645 3895 46690 4015
rect 46810 3895 46865 4015
rect 46985 3895 47030 4015
rect 47150 3895 47195 4015
rect 47315 3895 47360 4015
rect 47480 3895 47535 4015
rect 47655 3895 47665 4015
rect 42165 3850 47665 3895
rect 42165 3730 42175 3850
rect 42295 3730 42340 3850
rect 42460 3730 42505 3850
rect 42625 3730 42670 3850
rect 42790 3730 42845 3850
rect 42965 3730 43010 3850
rect 43130 3730 43175 3850
rect 43295 3730 43340 3850
rect 43460 3730 43515 3850
rect 43635 3730 43680 3850
rect 43800 3730 43845 3850
rect 43965 3730 44010 3850
rect 44130 3730 44185 3850
rect 44305 3730 44350 3850
rect 44470 3730 44515 3850
rect 44635 3730 44680 3850
rect 44800 3730 44855 3850
rect 44975 3730 45020 3850
rect 45140 3730 45185 3850
rect 45305 3730 45350 3850
rect 45470 3730 45525 3850
rect 45645 3730 45690 3850
rect 45810 3730 45855 3850
rect 45975 3730 46020 3850
rect 46140 3730 46195 3850
rect 46315 3730 46360 3850
rect 46480 3730 46525 3850
rect 46645 3730 46690 3850
rect 46810 3730 46865 3850
rect 46985 3730 47030 3850
rect 47150 3730 47195 3850
rect 47315 3730 47360 3850
rect 47480 3730 47535 3850
rect 47655 3730 47665 3850
rect 42165 3675 47665 3730
rect 42165 3555 42175 3675
rect 42295 3555 42340 3675
rect 42460 3555 42505 3675
rect 42625 3555 42670 3675
rect 42790 3555 42845 3675
rect 42965 3555 43010 3675
rect 43130 3555 43175 3675
rect 43295 3555 43340 3675
rect 43460 3555 43515 3675
rect 43635 3555 43680 3675
rect 43800 3555 43845 3675
rect 43965 3555 44010 3675
rect 44130 3555 44185 3675
rect 44305 3555 44350 3675
rect 44470 3555 44515 3675
rect 44635 3555 44680 3675
rect 44800 3555 44855 3675
rect 44975 3555 45020 3675
rect 45140 3555 45185 3675
rect 45305 3555 45350 3675
rect 45470 3555 45525 3675
rect 45645 3555 45690 3675
rect 45810 3555 45855 3675
rect 45975 3555 46020 3675
rect 46140 3555 46195 3675
rect 46315 3555 46360 3675
rect 46480 3555 46525 3675
rect 46645 3555 46690 3675
rect 46810 3555 46865 3675
rect 46985 3555 47030 3675
rect 47150 3555 47195 3675
rect 47315 3555 47360 3675
rect 47480 3555 47535 3675
rect 47655 3555 47665 3675
rect 42165 3510 47665 3555
rect 42165 3390 42175 3510
rect 42295 3390 42340 3510
rect 42460 3390 42505 3510
rect 42625 3390 42670 3510
rect 42790 3390 42845 3510
rect 42965 3390 43010 3510
rect 43130 3390 43175 3510
rect 43295 3390 43340 3510
rect 43460 3390 43515 3510
rect 43635 3390 43680 3510
rect 43800 3390 43845 3510
rect 43965 3390 44010 3510
rect 44130 3390 44185 3510
rect 44305 3390 44350 3510
rect 44470 3390 44515 3510
rect 44635 3390 44680 3510
rect 44800 3390 44855 3510
rect 44975 3390 45020 3510
rect 45140 3390 45185 3510
rect 45305 3390 45350 3510
rect 45470 3390 45525 3510
rect 45645 3390 45690 3510
rect 45810 3390 45855 3510
rect 45975 3390 46020 3510
rect 46140 3390 46195 3510
rect 46315 3390 46360 3510
rect 46480 3390 46525 3510
rect 46645 3390 46690 3510
rect 46810 3390 46865 3510
rect 46985 3390 47030 3510
rect 47150 3390 47195 3510
rect 47315 3390 47360 3510
rect 47480 3390 47535 3510
rect 47655 3390 47665 3510
rect 42165 3345 47665 3390
rect 42165 3225 42175 3345
rect 42295 3225 42340 3345
rect 42460 3225 42505 3345
rect 42625 3225 42670 3345
rect 42790 3225 42845 3345
rect 42965 3225 43010 3345
rect 43130 3225 43175 3345
rect 43295 3225 43340 3345
rect 43460 3225 43515 3345
rect 43635 3225 43680 3345
rect 43800 3225 43845 3345
rect 43965 3225 44010 3345
rect 44130 3225 44185 3345
rect 44305 3225 44350 3345
rect 44470 3225 44515 3345
rect 44635 3225 44680 3345
rect 44800 3225 44855 3345
rect 44975 3225 45020 3345
rect 45140 3225 45185 3345
rect 45305 3225 45350 3345
rect 45470 3225 45525 3345
rect 45645 3225 45690 3345
rect 45810 3225 45855 3345
rect 45975 3225 46020 3345
rect 46140 3225 46195 3345
rect 46315 3225 46360 3345
rect 46480 3225 46525 3345
rect 46645 3225 46690 3345
rect 46810 3225 46865 3345
rect 46985 3225 47030 3345
rect 47150 3225 47195 3345
rect 47315 3225 47360 3345
rect 47480 3225 47535 3345
rect 47655 3225 47665 3345
rect 42165 3180 47665 3225
rect 42165 3060 42175 3180
rect 42295 3060 42340 3180
rect 42460 3060 42505 3180
rect 42625 3060 42670 3180
rect 42790 3060 42845 3180
rect 42965 3060 43010 3180
rect 43130 3060 43175 3180
rect 43295 3060 43340 3180
rect 43460 3060 43515 3180
rect 43635 3060 43680 3180
rect 43800 3060 43845 3180
rect 43965 3060 44010 3180
rect 44130 3060 44185 3180
rect 44305 3060 44350 3180
rect 44470 3060 44515 3180
rect 44635 3060 44680 3180
rect 44800 3060 44855 3180
rect 44975 3060 45020 3180
rect 45140 3060 45185 3180
rect 45305 3060 45350 3180
rect 45470 3060 45525 3180
rect 45645 3060 45690 3180
rect 45810 3060 45855 3180
rect 45975 3060 46020 3180
rect 46140 3060 46195 3180
rect 46315 3060 46360 3180
rect 46480 3060 46525 3180
rect 46645 3060 46690 3180
rect 46810 3060 46865 3180
rect 46985 3060 47030 3180
rect 47150 3060 47195 3180
rect 47315 3060 47360 3180
rect 47480 3060 47535 3180
rect 47655 3060 47665 3180
rect 42165 3005 47665 3060
rect 42165 2885 42175 3005
rect 42295 2885 42340 3005
rect 42460 2885 42505 3005
rect 42625 2885 42670 3005
rect 42790 2885 42845 3005
rect 42965 2885 43010 3005
rect 43130 2885 43175 3005
rect 43295 2885 43340 3005
rect 43460 2885 43515 3005
rect 43635 2885 43680 3005
rect 43800 2885 43845 3005
rect 43965 2885 44010 3005
rect 44130 2885 44185 3005
rect 44305 2885 44350 3005
rect 44470 2885 44515 3005
rect 44635 2885 44680 3005
rect 44800 2885 44855 3005
rect 44975 2885 45020 3005
rect 45140 2885 45185 3005
rect 45305 2885 45350 3005
rect 45470 2885 45525 3005
rect 45645 2885 45690 3005
rect 45810 2885 45855 3005
rect 45975 2885 46020 3005
rect 46140 2885 46195 3005
rect 46315 2885 46360 3005
rect 46480 2885 46525 3005
rect 46645 2885 46690 3005
rect 46810 2885 46865 3005
rect 46985 2885 47030 3005
rect 47150 2885 47195 3005
rect 47315 2885 47360 3005
rect 47480 2885 47535 3005
rect 47655 2885 47665 3005
rect 42165 2840 47665 2885
rect 42165 2720 42175 2840
rect 42295 2720 42340 2840
rect 42460 2720 42505 2840
rect 42625 2720 42670 2840
rect 42790 2720 42845 2840
rect 42965 2720 43010 2840
rect 43130 2720 43175 2840
rect 43295 2720 43340 2840
rect 43460 2720 43515 2840
rect 43635 2720 43680 2840
rect 43800 2720 43845 2840
rect 43965 2720 44010 2840
rect 44130 2720 44185 2840
rect 44305 2720 44350 2840
rect 44470 2720 44515 2840
rect 44635 2720 44680 2840
rect 44800 2720 44855 2840
rect 44975 2720 45020 2840
rect 45140 2720 45185 2840
rect 45305 2720 45350 2840
rect 45470 2720 45525 2840
rect 45645 2720 45690 2840
rect 45810 2720 45855 2840
rect 45975 2720 46020 2840
rect 46140 2720 46195 2840
rect 46315 2720 46360 2840
rect 46480 2720 46525 2840
rect 46645 2720 46690 2840
rect 46810 2720 46865 2840
rect 46985 2720 47030 2840
rect 47150 2720 47195 2840
rect 47315 2720 47360 2840
rect 47480 2720 47535 2840
rect 47655 2720 47665 2840
rect 42165 2675 47665 2720
rect 42165 2555 42175 2675
rect 42295 2555 42340 2675
rect 42460 2555 42505 2675
rect 42625 2555 42670 2675
rect 42790 2555 42845 2675
rect 42965 2555 43010 2675
rect 43130 2555 43175 2675
rect 43295 2555 43340 2675
rect 43460 2555 43515 2675
rect 43635 2555 43680 2675
rect 43800 2555 43845 2675
rect 43965 2555 44010 2675
rect 44130 2555 44185 2675
rect 44305 2555 44350 2675
rect 44470 2555 44515 2675
rect 44635 2555 44680 2675
rect 44800 2555 44855 2675
rect 44975 2555 45020 2675
rect 45140 2555 45185 2675
rect 45305 2555 45350 2675
rect 45470 2555 45525 2675
rect 45645 2555 45690 2675
rect 45810 2555 45855 2675
rect 45975 2555 46020 2675
rect 46140 2555 46195 2675
rect 46315 2555 46360 2675
rect 46480 2555 46525 2675
rect 46645 2555 46690 2675
rect 46810 2555 46865 2675
rect 46985 2555 47030 2675
rect 47150 2555 47195 2675
rect 47315 2555 47360 2675
rect 47480 2555 47535 2675
rect 47655 2555 47665 2675
rect 42165 2510 47665 2555
rect 42165 2390 42175 2510
rect 42295 2390 42340 2510
rect 42460 2390 42505 2510
rect 42625 2390 42670 2510
rect 42790 2390 42845 2510
rect 42965 2390 43010 2510
rect 43130 2390 43175 2510
rect 43295 2390 43340 2510
rect 43460 2390 43515 2510
rect 43635 2390 43680 2510
rect 43800 2390 43845 2510
rect 43965 2390 44010 2510
rect 44130 2390 44185 2510
rect 44305 2390 44350 2510
rect 44470 2390 44515 2510
rect 44635 2390 44680 2510
rect 44800 2390 44855 2510
rect 44975 2390 45020 2510
rect 45140 2390 45185 2510
rect 45305 2390 45350 2510
rect 45470 2390 45525 2510
rect 45645 2390 45690 2510
rect 45810 2390 45855 2510
rect 45975 2390 46020 2510
rect 46140 2390 46195 2510
rect 46315 2390 46360 2510
rect 46480 2390 46525 2510
rect 46645 2390 46690 2510
rect 46810 2390 46865 2510
rect 46985 2390 47030 2510
rect 47150 2390 47195 2510
rect 47315 2390 47360 2510
rect 47480 2390 47535 2510
rect 47655 2390 47665 2510
rect 42165 2335 47665 2390
rect 42165 2215 42175 2335
rect 42295 2215 42340 2335
rect 42460 2215 42505 2335
rect 42625 2215 42670 2335
rect 42790 2215 42845 2335
rect 42965 2215 43010 2335
rect 43130 2215 43175 2335
rect 43295 2215 43340 2335
rect 43460 2215 43515 2335
rect 43635 2215 43680 2335
rect 43800 2215 43845 2335
rect 43965 2215 44010 2335
rect 44130 2215 44185 2335
rect 44305 2215 44350 2335
rect 44470 2215 44515 2335
rect 44635 2215 44680 2335
rect 44800 2215 44855 2335
rect 44975 2215 45020 2335
rect 45140 2215 45185 2335
rect 45305 2215 45350 2335
rect 45470 2215 45525 2335
rect 45645 2215 45690 2335
rect 45810 2215 45855 2335
rect 45975 2215 46020 2335
rect 46140 2215 46195 2335
rect 46315 2215 46360 2335
rect 46480 2215 46525 2335
rect 46645 2215 46690 2335
rect 46810 2215 46865 2335
rect 46985 2215 47030 2335
rect 47150 2215 47195 2335
rect 47315 2215 47360 2335
rect 47480 2215 47535 2335
rect 47655 2215 47665 2335
rect 42165 2170 47665 2215
rect 42165 2050 42175 2170
rect 42295 2050 42340 2170
rect 42460 2050 42505 2170
rect 42625 2050 42670 2170
rect 42790 2050 42845 2170
rect 42965 2050 43010 2170
rect 43130 2050 43175 2170
rect 43295 2050 43340 2170
rect 43460 2050 43515 2170
rect 43635 2050 43680 2170
rect 43800 2050 43845 2170
rect 43965 2050 44010 2170
rect 44130 2050 44185 2170
rect 44305 2050 44350 2170
rect 44470 2050 44515 2170
rect 44635 2050 44680 2170
rect 44800 2050 44855 2170
rect 44975 2050 45020 2170
rect 45140 2050 45185 2170
rect 45305 2050 45350 2170
rect 45470 2050 45525 2170
rect 45645 2050 45690 2170
rect 45810 2050 45855 2170
rect 45975 2050 46020 2170
rect 46140 2050 46195 2170
rect 46315 2050 46360 2170
rect 46480 2050 46525 2170
rect 46645 2050 46690 2170
rect 46810 2050 46865 2170
rect 46985 2050 47030 2170
rect 47150 2050 47195 2170
rect 47315 2050 47360 2170
rect 47480 2050 47535 2170
rect 47655 2050 47665 2170
rect 42165 2005 47665 2050
rect 42165 1885 42175 2005
rect 42295 1885 42340 2005
rect 42460 1885 42505 2005
rect 42625 1885 42670 2005
rect 42790 1885 42845 2005
rect 42965 1885 43010 2005
rect 43130 1885 43175 2005
rect 43295 1885 43340 2005
rect 43460 1885 43515 2005
rect 43635 1885 43680 2005
rect 43800 1885 43845 2005
rect 43965 1885 44010 2005
rect 44130 1885 44185 2005
rect 44305 1885 44350 2005
rect 44470 1885 44515 2005
rect 44635 1885 44680 2005
rect 44800 1885 44855 2005
rect 44975 1885 45020 2005
rect 45140 1885 45185 2005
rect 45305 1885 45350 2005
rect 45470 1885 45525 2005
rect 45645 1885 45690 2005
rect 45810 1885 45855 2005
rect 45975 1885 46020 2005
rect 46140 1885 46195 2005
rect 46315 1885 46360 2005
rect 46480 1885 46525 2005
rect 46645 1885 46690 2005
rect 46810 1885 46865 2005
rect 46985 1885 47030 2005
rect 47150 1885 47195 2005
rect 47315 1885 47360 2005
rect 47480 1885 47535 2005
rect 47655 1885 47665 2005
rect 42165 1840 47665 1885
rect 42165 1720 42175 1840
rect 42295 1720 42340 1840
rect 42460 1720 42505 1840
rect 42625 1720 42670 1840
rect 42790 1720 42845 1840
rect 42965 1720 43010 1840
rect 43130 1720 43175 1840
rect 43295 1720 43340 1840
rect 43460 1720 43515 1840
rect 43635 1720 43680 1840
rect 43800 1720 43845 1840
rect 43965 1720 44010 1840
rect 44130 1720 44185 1840
rect 44305 1720 44350 1840
rect 44470 1720 44515 1840
rect 44635 1720 44680 1840
rect 44800 1720 44855 1840
rect 44975 1720 45020 1840
rect 45140 1720 45185 1840
rect 45305 1720 45350 1840
rect 45470 1720 45525 1840
rect 45645 1720 45690 1840
rect 45810 1720 45855 1840
rect 45975 1720 46020 1840
rect 46140 1720 46195 1840
rect 46315 1720 46360 1840
rect 46480 1720 46525 1840
rect 46645 1720 46690 1840
rect 46810 1720 46865 1840
rect 46985 1720 47030 1840
rect 47150 1720 47195 1840
rect 47315 1720 47360 1840
rect 47480 1720 47535 1840
rect 47655 1720 47665 1840
rect 42165 1710 47665 1720
rect 47855 7200 53355 7210
rect 47855 7080 47865 7200
rect 47985 7080 48030 7200
rect 48150 7080 48195 7200
rect 48315 7080 48360 7200
rect 48480 7080 48535 7200
rect 48655 7080 48700 7200
rect 48820 7080 48865 7200
rect 48985 7080 49030 7200
rect 49150 7080 49205 7200
rect 49325 7080 49370 7200
rect 49490 7080 49535 7200
rect 49655 7080 49700 7200
rect 49820 7080 49875 7200
rect 49995 7080 50040 7200
rect 50160 7080 50205 7200
rect 50325 7080 50370 7200
rect 50490 7080 50545 7200
rect 50665 7080 50710 7200
rect 50830 7080 50875 7200
rect 50995 7080 51040 7200
rect 51160 7080 51215 7200
rect 51335 7080 51380 7200
rect 51500 7080 51545 7200
rect 51665 7080 51710 7200
rect 51830 7080 51885 7200
rect 52005 7080 52050 7200
rect 52170 7080 52215 7200
rect 52335 7080 52380 7200
rect 52500 7080 52555 7200
rect 52675 7080 52720 7200
rect 52840 7080 52885 7200
rect 53005 7080 53050 7200
rect 53170 7080 53225 7200
rect 53345 7080 53355 7200
rect 47855 7025 53355 7080
rect 47855 6905 47865 7025
rect 47985 6905 48030 7025
rect 48150 6905 48195 7025
rect 48315 6905 48360 7025
rect 48480 6905 48535 7025
rect 48655 6905 48700 7025
rect 48820 6905 48865 7025
rect 48985 6905 49030 7025
rect 49150 6905 49205 7025
rect 49325 6905 49370 7025
rect 49490 6905 49535 7025
rect 49655 6905 49700 7025
rect 49820 6905 49875 7025
rect 49995 6905 50040 7025
rect 50160 6905 50205 7025
rect 50325 6905 50370 7025
rect 50490 6905 50545 7025
rect 50665 6905 50710 7025
rect 50830 6905 50875 7025
rect 50995 6905 51040 7025
rect 51160 6905 51215 7025
rect 51335 6905 51380 7025
rect 51500 6905 51545 7025
rect 51665 6905 51710 7025
rect 51830 6905 51885 7025
rect 52005 6905 52050 7025
rect 52170 6905 52215 7025
rect 52335 6905 52380 7025
rect 52500 6905 52555 7025
rect 52675 6905 52720 7025
rect 52840 6905 52885 7025
rect 53005 6905 53050 7025
rect 53170 6905 53225 7025
rect 53345 6905 53355 7025
rect 47855 6860 53355 6905
rect 47855 6740 47865 6860
rect 47985 6740 48030 6860
rect 48150 6740 48195 6860
rect 48315 6740 48360 6860
rect 48480 6740 48535 6860
rect 48655 6740 48700 6860
rect 48820 6740 48865 6860
rect 48985 6740 49030 6860
rect 49150 6740 49205 6860
rect 49325 6740 49370 6860
rect 49490 6740 49535 6860
rect 49655 6740 49700 6860
rect 49820 6740 49875 6860
rect 49995 6740 50040 6860
rect 50160 6740 50205 6860
rect 50325 6740 50370 6860
rect 50490 6740 50545 6860
rect 50665 6740 50710 6860
rect 50830 6740 50875 6860
rect 50995 6740 51040 6860
rect 51160 6740 51215 6860
rect 51335 6740 51380 6860
rect 51500 6740 51545 6860
rect 51665 6740 51710 6860
rect 51830 6740 51885 6860
rect 52005 6740 52050 6860
rect 52170 6740 52215 6860
rect 52335 6740 52380 6860
rect 52500 6740 52555 6860
rect 52675 6740 52720 6860
rect 52840 6740 52885 6860
rect 53005 6740 53050 6860
rect 53170 6740 53225 6860
rect 53345 6740 53355 6860
rect 47855 6695 53355 6740
rect 47855 6575 47865 6695
rect 47985 6575 48030 6695
rect 48150 6575 48195 6695
rect 48315 6575 48360 6695
rect 48480 6575 48535 6695
rect 48655 6575 48700 6695
rect 48820 6575 48865 6695
rect 48985 6575 49030 6695
rect 49150 6575 49205 6695
rect 49325 6575 49370 6695
rect 49490 6575 49535 6695
rect 49655 6575 49700 6695
rect 49820 6575 49875 6695
rect 49995 6575 50040 6695
rect 50160 6575 50205 6695
rect 50325 6575 50370 6695
rect 50490 6575 50545 6695
rect 50665 6575 50710 6695
rect 50830 6575 50875 6695
rect 50995 6575 51040 6695
rect 51160 6575 51215 6695
rect 51335 6575 51380 6695
rect 51500 6575 51545 6695
rect 51665 6575 51710 6695
rect 51830 6575 51885 6695
rect 52005 6575 52050 6695
rect 52170 6575 52215 6695
rect 52335 6575 52380 6695
rect 52500 6575 52555 6695
rect 52675 6575 52720 6695
rect 52840 6575 52885 6695
rect 53005 6575 53050 6695
rect 53170 6575 53225 6695
rect 53345 6575 53355 6695
rect 47855 6530 53355 6575
rect 47855 6410 47865 6530
rect 47985 6410 48030 6530
rect 48150 6410 48195 6530
rect 48315 6410 48360 6530
rect 48480 6410 48535 6530
rect 48655 6410 48700 6530
rect 48820 6410 48865 6530
rect 48985 6410 49030 6530
rect 49150 6410 49205 6530
rect 49325 6410 49370 6530
rect 49490 6410 49535 6530
rect 49655 6410 49700 6530
rect 49820 6410 49875 6530
rect 49995 6410 50040 6530
rect 50160 6410 50205 6530
rect 50325 6410 50370 6530
rect 50490 6410 50545 6530
rect 50665 6410 50710 6530
rect 50830 6410 50875 6530
rect 50995 6410 51040 6530
rect 51160 6410 51215 6530
rect 51335 6410 51380 6530
rect 51500 6410 51545 6530
rect 51665 6410 51710 6530
rect 51830 6410 51885 6530
rect 52005 6410 52050 6530
rect 52170 6410 52215 6530
rect 52335 6410 52380 6530
rect 52500 6410 52555 6530
rect 52675 6410 52720 6530
rect 52840 6410 52885 6530
rect 53005 6410 53050 6530
rect 53170 6410 53225 6530
rect 53345 6410 53355 6530
rect 47855 6355 53355 6410
rect 47855 6235 47865 6355
rect 47985 6235 48030 6355
rect 48150 6235 48195 6355
rect 48315 6235 48360 6355
rect 48480 6235 48535 6355
rect 48655 6235 48700 6355
rect 48820 6235 48865 6355
rect 48985 6235 49030 6355
rect 49150 6235 49205 6355
rect 49325 6235 49370 6355
rect 49490 6235 49535 6355
rect 49655 6235 49700 6355
rect 49820 6235 49875 6355
rect 49995 6235 50040 6355
rect 50160 6235 50205 6355
rect 50325 6235 50370 6355
rect 50490 6235 50545 6355
rect 50665 6235 50710 6355
rect 50830 6235 50875 6355
rect 50995 6235 51040 6355
rect 51160 6235 51215 6355
rect 51335 6235 51380 6355
rect 51500 6235 51545 6355
rect 51665 6235 51710 6355
rect 51830 6235 51885 6355
rect 52005 6235 52050 6355
rect 52170 6235 52215 6355
rect 52335 6235 52380 6355
rect 52500 6235 52555 6355
rect 52675 6235 52720 6355
rect 52840 6235 52885 6355
rect 53005 6235 53050 6355
rect 53170 6235 53225 6355
rect 53345 6235 53355 6355
rect 47855 6190 53355 6235
rect 47855 6070 47865 6190
rect 47985 6070 48030 6190
rect 48150 6070 48195 6190
rect 48315 6070 48360 6190
rect 48480 6070 48535 6190
rect 48655 6070 48700 6190
rect 48820 6070 48865 6190
rect 48985 6070 49030 6190
rect 49150 6070 49205 6190
rect 49325 6070 49370 6190
rect 49490 6070 49535 6190
rect 49655 6070 49700 6190
rect 49820 6070 49875 6190
rect 49995 6070 50040 6190
rect 50160 6070 50205 6190
rect 50325 6070 50370 6190
rect 50490 6070 50545 6190
rect 50665 6070 50710 6190
rect 50830 6070 50875 6190
rect 50995 6070 51040 6190
rect 51160 6070 51215 6190
rect 51335 6070 51380 6190
rect 51500 6070 51545 6190
rect 51665 6070 51710 6190
rect 51830 6070 51885 6190
rect 52005 6070 52050 6190
rect 52170 6070 52215 6190
rect 52335 6070 52380 6190
rect 52500 6070 52555 6190
rect 52675 6070 52720 6190
rect 52840 6070 52885 6190
rect 53005 6070 53050 6190
rect 53170 6070 53225 6190
rect 53345 6070 53355 6190
rect 47855 6025 53355 6070
rect 47855 5905 47865 6025
rect 47985 5905 48030 6025
rect 48150 5905 48195 6025
rect 48315 5905 48360 6025
rect 48480 5905 48535 6025
rect 48655 5905 48700 6025
rect 48820 5905 48865 6025
rect 48985 5905 49030 6025
rect 49150 5905 49205 6025
rect 49325 5905 49370 6025
rect 49490 5905 49535 6025
rect 49655 5905 49700 6025
rect 49820 5905 49875 6025
rect 49995 5905 50040 6025
rect 50160 5905 50205 6025
rect 50325 5905 50370 6025
rect 50490 5905 50545 6025
rect 50665 5905 50710 6025
rect 50830 5905 50875 6025
rect 50995 5905 51040 6025
rect 51160 5905 51215 6025
rect 51335 5905 51380 6025
rect 51500 5905 51545 6025
rect 51665 5905 51710 6025
rect 51830 5905 51885 6025
rect 52005 5905 52050 6025
rect 52170 5905 52215 6025
rect 52335 5905 52380 6025
rect 52500 5905 52555 6025
rect 52675 5905 52720 6025
rect 52840 5905 52885 6025
rect 53005 5905 53050 6025
rect 53170 5905 53225 6025
rect 53345 5905 53355 6025
rect 47855 5860 53355 5905
rect 47855 5740 47865 5860
rect 47985 5740 48030 5860
rect 48150 5740 48195 5860
rect 48315 5740 48360 5860
rect 48480 5740 48535 5860
rect 48655 5740 48700 5860
rect 48820 5740 48865 5860
rect 48985 5740 49030 5860
rect 49150 5740 49205 5860
rect 49325 5740 49370 5860
rect 49490 5740 49535 5860
rect 49655 5740 49700 5860
rect 49820 5740 49875 5860
rect 49995 5740 50040 5860
rect 50160 5740 50205 5860
rect 50325 5740 50370 5860
rect 50490 5740 50545 5860
rect 50665 5740 50710 5860
rect 50830 5740 50875 5860
rect 50995 5740 51040 5860
rect 51160 5740 51215 5860
rect 51335 5740 51380 5860
rect 51500 5740 51545 5860
rect 51665 5740 51710 5860
rect 51830 5740 51885 5860
rect 52005 5740 52050 5860
rect 52170 5740 52215 5860
rect 52335 5740 52380 5860
rect 52500 5740 52555 5860
rect 52675 5740 52720 5860
rect 52840 5740 52885 5860
rect 53005 5740 53050 5860
rect 53170 5740 53225 5860
rect 53345 5740 53355 5860
rect 47855 5685 53355 5740
rect 47855 5565 47865 5685
rect 47985 5565 48030 5685
rect 48150 5565 48195 5685
rect 48315 5565 48360 5685
rect 48480 5565 48535 5685
rect 48655 5565 48700 5685
rect 48820 5565 48865 5685
rect 48985 5565 49030 5685
rect 49150 5565 49205 5685
rect 49325 5565 49370 5685
rect 49490 5565 49535 5685
rect 49655 5565 49700 5685
rect 49820 5565 49875 5685
rect 49995 5565 50040 5685
rect 50160 5565 50205 5685
rect 50325 5565 50370 5685
rect 50490 5565 50545 5685
rect 50665 5565 50710 5685
rect 50830 5565 50875 5685
rect 50995 5565 51040 5685
rect 51160 5565 51215 5685
rect 51335 5565 51380 5685
rect 51500 5565 51545 5685
rect 51665 5565 51710 5685
rect 51830 5565 51885 5685
rect 52005 5565 52050 5685
rect 52170 5565 52215 5685
rect 52335 5565 52380 5685
rect 52500 5565 52555 5685
rect 52675 5565 52720 5685
rect 52840 5565 52885 5685
rect 53005 5565 53050 5685
rect 53170 5565 53225 5685
rect 53345 5565 53355 5685
rect 47855 5520 53355 5565
rect 47855 5400 47865 5520
rect 47985 5400 48030 5520
rect 48150 5400 48195 5520
rect 48315 5400 48360 5520
rect 48480 5400 48535 5520
rect 48655 5400 48700 5520
rect 48820 5400 48865 5520
rect 48985 5400 49030 5520
rect 49150 5400 49205 5520
rect 49325 5400 49370 5520
rect 49490 5400 49535 5520
rect 49655 5400 49700 5520
rect 49820 5400 49875 5520
rect 49995 5400 50040 5520
rect 50160 5400 50205 5520
rect 50325 5400 50370 5520
rect 50490 5400 50545 5520
rect 50665 5400 50710 5520
rect 50830 5400 50875 5520
rect 50995 5400 51040 5520
rect 51160 5400 51215 5520
rect 51335 5400 51380 5520
rect 51500 5400 51545 5520
rect 51665 5400 51710 5520
rect 51830 5400 51885 5520
rect 52005 5400 52050 5520
rect 52170 5400 52215 5520
rect 52335 5400 52380 5520
rect 52500 5400 52555 5520
rect 52675 5400 52720 5520
rect 52840 5400 52885 5520
rect 53005 5400 53050 5520
rect 53170 5400 53225 5520
rect 53345 5400 53355 5520
rect 47855 5355 53355 5400
rect 47855 5235 47865 5355
rect 47985 5235 48030 5355
rect 48150 5235 48195 5355
rect 48315 5235 48360 5355
rect 48480 5235 48535 5355
rect 48655 5235 48700 5355
rect 48820 5235 48865 5355
rect 48985 5235 49030 5355
rect 49150 5235 49205 5355
rect 49325 5235 49370 5355
rect 49490 5235 49535 5355
rect 49655 5235 49700 5355
rect 49820 5235 49875 5355
rect 49995 5235 50040 5355
rect 50160 5235 50205 5355
rect 50325 5235 50370 5355
rect 50490 5235 50545 5355
rect 50665 5235 50710 5355
rect 50830 5235 50875 5355
rect 50995 5235 51040 5355
rect 51160 5235 51215 5355
rect 51335 5235 51380 5355
rect 51500 5235 51545 5355
rect 51665 5235 51710 5355
rect 51830 5235 51885 5355
rect 52005 5235 52050 5355
rect 52170 5235 52215 5355
rect 52335 5235 52380 5355
rect 52500 5235 52555 5355
rect 52675 5235 52720 5355
rect 52840 5235 52885 5355
rect 53005 5235 53050 5355
rect 53170 5235 53225 5355
rect 53345 5235 53355 5355
rect 47855 5190 53355 5235
rect 47855 5070 47865 5190
rect 47985 5070 48030 5190
rect 48150 5070 48195 5190
rect 48315 5070 48360 5190
rect 48480 5070 48535 5190
rect 48655 5070 48700 5190
rect 48820 5070 48865 5190
rect 48985 5070 49030 5190
rect 49150 5070 49205 5190
rect 49325 5070 49370 5190
rect 49490 5070 49535 5190
rect 49655 5070 49700 5190
rect 49820 5070 49875 5190
rect 49995 5070 50040 5190
rect 50160 5070 50205 5190
rect 50325 5070 50370 5190
rect 50490 5070 50545 5190
rect 50665 5070 50710 5190
rect 50830 5070 50875 5190
rect 50995 5070 51040 5190
rect 51160 5070 51215 5190
rect 51335 5070 51380 5190
rect 51500 5070 51545 5190
rect 51665 5070 51710 5190
rect 51830 5070 51885 5190
rect 52005 5070 52050 5190
rect 52170 5070 52215 5190
rect 52335 5070 52380 5190
rect 52500 5070 52555 5190
rect 52675 5070 52720 5190
rect 52840 5070 52885 5190
rect 53005 5070 53050 5190
rect 53170 5070 53225 5190
rect 53345 5070 53355 5190
rect 47855 5015 53355 5070
rect 47855 4895 47865 5015
rect 47985 4895 48030 5015
rect 48150 4895 48195 5015
rect 48315 4895 48360 5015
rect 48480 4895 48535 5015
rect 48655 4895 48700 5015
rect 48820 4895 48865 5015
rect 48985 4895 49030 5015
rect 49150 4895 49205 5015
rect 49325 4895 49370 5015
rect 49490 4895 49535 5015
rect 49655 4895 49700 5015
rect 49820 4895 49875 5015
rect 49995 4895 50040 5015
rect 50160 4895 50205 5015
rect 50325 4895 50370 5015
rect 50490 4895 50545 5015
rect 50665 4895 50710 5015
rect 50830 4895 50875 5015
rect 50995 4895 51040 5015
rect 51160 4895 51215 5015
rect 51335 4895 51380 5015
rect 51500 4895 51545 5015
rect 51665 4895 51710 5015
rect 51830 4895 51885 5015
rect 52005 4895 52050 5015
rect 52170 4895 52215 5015
rect 52335 4895 52380 5015
rect 52500 4895 52555 5015
rect 52675 4895 52720 5015
rect 52840 4895 52885 5015
rect 53005 4895 53050 5015
rect 53170 4895 53225 5015
rect 53345 4895 53355 5015
rect 47855 4850 53355 4895
rect 47855 4730 47865 4850
rect 47985 4730 48030 4850
rect 48150 4730 48195 4850
rect 48315 4730 48360 4850
rect 48480 4730 48535 4850
rect 48655 4730 48700 4850
rect 48820 4730 48865 4850
rect 48985 4730 49030 4850
rect 49150 4730 49205 4850
rect 49325 4730 49370 4850
rect 49490 4730 49535 4850
rect 49655 4730 49700 4850
rect 49820 4730 49875 4850
rect 49995 4730 50040 4850
rect 50160 4730 50205 4850
rect 50325 4730 50370 4850
rect 50490 4730 50545 4850
rect 50665 4730 50710 4850
rect 50830 4730 50875 4850
rect 50995 4730 51040 4850
rect 51160 4730 51215 4850
rect 51335 4730 51380 4850
rect 51500 4730 51545 4850
rect 51665 4730 51710 4850
rect 51830 4730 51885 4850
rect 52005 4730 52050 4850
rect 52170 4730 52215 4850
rect 52335 4730 52380 4850
rect 52500 4730 52555 4850
rect 52675 4730 52720 4850
rect 52840 4730 52885 4850
rect 53005 4730 53050 4850
rect 53170 4730 53225 4850
rect 53345 4730 53355 4850
rect 47855 4685 53355 4730
rect 47855 4565 47865 4685
rect 47985 4565 48030 4685
rect 48150 4565 48195 4685
rect 48315 4565 48360 4685
rect 48480 4565 48535 4685
rect 48655 4565 48700 4685
rect 48820 4565 48865 4685
rect 48985 4565 49030 4685
rect 49150 4565 49205 4685
rect 49325 4565 49370 4685
rect 49490 4565 49535 4685
rect 49655 4565 49700 4685
rect 49820 4565 49875 4685
rect 49995 4565 50040 4685
rect 50160 4565 50205 4685
rect 50325 4565 50370 4685
rect 50490 4565 50545 4685
rect 50665 4565 50710 4685
rect 50830 4565 50875 4685
rect 50995 4565 51040 4685
rect 51160 4565 51215 4685
rect 51335 4565 51380 4685
rect 51500 4565 51545 4685
rect 51665 4565 51710 4685
rect 51830 4565 51885 4685
rect 52005 4565 52050 4685
rect 52170 4565 52215 4685
rect 52335 4565 52380 4685
rect 52500 4565 52555 4685
rect 52675 4565 52720 4685
rect 52840 4565 52885 4685
rect 53005 4565 53050 4685
rect 53170 4565 53225 4685
rect 53345 4565 53355 4685
rect 47855 4520 53355 4565
rect 47855 4400 47865 4520
rect 47985 4400 48030 4520
rect 48150 4400 48195 4520
rect 48315 4400 48360 4520
rect 48480 4400 48535 4520
rect 48655 4400 48700 4520
rect 48820 4400 48865 4520
rect 48985 4400 49030 4520
rect 49150 4400 49205 4520
rect 49325 4400 49370 4520
rect 49490 4400 49535 4520
rect 49655 4400 49700 4520
rect 49820 4400 49875 4520
rect 49995 4400 50040 4520
rect 50160 4400 50205 4520
rect 50325 4400 50370 4520
rect 50490 4400 50545 4520
rect 50665 4400 50710 4520
rect 50830 4400 50875 4520
rect 50995 4400 51040 4520
rect 51160 4400 51215 4520
rect 51335 4400 51380 4520
rect 51500 4400 51545 4520
rect 51665 4400 51710 4520
rect 51830 4400 51885 4520
rect 52005 4400 52050 4520
rect 52170 4400 52215 4520
rect 52335 4400 52380 4520
rect 52500 4400 52555 4520
rect 52675 4400 52720 4520
rect 52840 4400 52885 4520
rect 53005 4400 53050 4520
rect 53170 4400 53225 4520
rect 53345 4400 53355 4520
rect 47855 4345 53355 4400
rect 47855 4225 47865 4345
rect 47985 4225 48030 4345
rect 48150 4225 48195 4345
rect 48315 4225 48360 4345
rect 48480 4225 48535 4345
rect 48655 4225 48700 4345
rect 48820 4225 48865 4345
rect 48985 4225 49030 4345
rect 49150 4225 49205 4345
rect 49325 4225 49370 4345
rect 49490 4225 49535 4345
rect 49655 4225 49700 4345
rect 49820 4225 49875 4345
rect 49995 4225 50040 4345
rect 50160 4225 50205 4345
rect 50325 4225 50370 4345
rect 50490 4225 50545 4345
rect 50665 4225 50710 4345
rect 50830 4225 50875 4345
rect 50995 4225 51040 4345
rect 51160 4225 51215 4345
rect 51335 4225 51380 4345
rect 51500 4225 51545 4345
rect 51665 4225 51710 4345
rect 51830 4225 51885 4345
rect 52005 4225 52050 4345
rect 52170 4225 52215 4345
rect 52335 4225 52380 4345
rect 52500 4225 52555 4345
rect 52675 4225 52720 4345
rect 52840 4225 52885 4345
rect 53005 4225 53050 4345
rect 53170 4225 53225 4345
rect 53345 4225 53355 4345
rect 47855 4180 53355 4225
rect 47855 4060 47865 4180
rect 47985 4060 48030 4180
rect 48150 4060 48195 4180
rect 48315 4060 48360 4180
rect 48480 4060 48535 4180
rect 48655 4060 48700 4180
rect 48820 4060 48865 4180
rect 48985 4060 49030 4180
rect 49150 4060 49205 4180
rect 49325 4060 49370 4180
rect 49490 4060 49535 4180
rect 49655 4060 49700 4180
rect 49820 4060 49875 4180
rect 49995 4060 50040 4180
rect 50160 4060 50205 4180
rect 50325 4060 50370 4180
rect 50490 4060 50545 4180
rect 50665 4060 50710 4180
rect 50830 4060 50875 4180
rect 50995 4060 51040 4180
rect 51160 4060 51215 4180
rect 51335 4060 51380 4180
rect 51500 4060 51545 4180
rect 51665 4060 51710 4180
rect 51830 4060 51885 4180
rect 52005 4060 52050 4180
rect 52170 4060 52215 4180
rect 52335 4060 52380 4180
rect 52500 4060 52555 4180
rect 52675 4060 52720 4180
rect 52840 4060 52885 4180
rect 53005 4060 53050 4180
rect 53170 4060 53225 4180
rect 53345 4060 53355 4180
rect 47855 4015 53355 4060
rect 47855 3895 47865 4015
rect 47985 3895 48030 4015
rect 48150 3895 48195 4015
rect 48315 3895 48360 4015
rect 48480 3895 48535 4015
rect 48655 3895 48700 4015
rect 48820 3895 48865 4015
rect 48985 3895 49030 4015
rect 49150 3895 49205 4015
rect 49325 3895 49370 4015
rect 49490 3895 49535 4015
rect 49655 3895 49700 4015
rect 49820 3895 49875 4015
rect 49995 3895 50040 4015
rect 50160 3895 50205 4015
rect 50325 3895 50370 4015
rect 50490 3895 50545 4015
rect 50665 3895 50710 4015
rect 50830 3895 50875 4015
rect 50995 3895 51040 4015
rect 51160 3895 51215 4015
rect 51335 3895 51380 4015
rect 51500 3895 51545 4015
rect 51665 3895 51710 4015
rect 51830 3895 51885 4015
rect 52005 3895 52050 4015
rect 52170 3895 52215 4015
rect 52335 3895 52380 4015
rect 52500 3895 52555 4015
rect 52675 3895 52720 4015
rect 52840 3895 52885 4015
rect 53005 3895 53050 4015
rect 53170 3895 53225 4015
rect 53345 3895 53355 4015
rect 47855 3850 53355 3895
rect 47855 3730 47865 3850
rect 47985 3730 48030 3850
rect 48150 3730 48195 3850
rect 48315 3730 48360 3850
rect 48480 3730 48535 3850
rect 48655 3730 48700 3850
rect 48820 3730 48865 3850
rect 48985 3730 49030 3850
rect 49150 3730 49205 3850
rect 49325 3730 49370 3850
rect 49490 3730 49535 3850
rect 49655 3730 49700 3850
rect 49820 3730 49875 3850
rect 49995 3730 50040 3850
rect 50160 3730 50205 3850
rect 50325 3730 50370 3850
rect 50490 3730 50545 3850
rect 50665 3730 50710 3850
rect 50830 3730 50875 3850
rect 50995 3730 51040 3850
rect 51160 3730 51215 3850
rect 51335 3730 51380 3850
rect 51500 3730 51545 3850
rect 51665 3730 51710 3850
rect 51830 3730 51885 3850
rect 52005 3730 52050 3850
rect 52170 3730 52215 3850
rect 52335 3730 52380 3850
rect 52500 3730 52555 3850
rect 52675 3730 52720 3850
rect 52840 3730 52885 3850
rect 53005 3730 53050 3850
rect 53170 3730 53225 3850
rect 53345 3730 53355 3850
rect 47855 3675 53355 3730
rect 47855 3555 47865 3675
rect 47985 3555 48030 3675
rect 48150 3555 48195 3675
rect 48315 3555 48360 3675
rect 48480 3555 48535 3675
rect 48655 3555 48700 3675
rect 48820 3555 48865 3675
rect 48985 3555 49030 3675
rect 49150 3555 49205 3675
rect 49325 3555 49370 3675
rect 49490 3555 49535 3675
rect 49655 3555 49700 3675
rect 49820 3555 49875 3675
rect 49995 3555 50040 3675
rect 50160 3555 50205 3675
rect 50325 3555 50370 3675
rect 50490 3555 50545 3675
rect 50665 3555 50710 3675
rect 50830 3555 50875 3675
rect 50995 3555 51040 3675
rect 51160 3555 51215 3675
rect 51335 3555 51380 3675
rect 51500 3555 51545 3675
rect 51665 3555 51710 3675
rect 51830 3555 51885 3675
rect 52005 3555 52050 3675
rect 52170 3555 52215 3675
rect 52335 3555 52380 3675
rect 52500 3555 52555 3675
rect 52675 3555 52720 3675
rect 52840 3555 52885 3675
rect 53005 3555 53050 3675
rect 53170 3555 53225 3675
rect 53345 3555 53355 3675
rect 47855 3510 53355 3555
rect 47855 3390 47865 3510
rect 47985 3390 48030 3510
rect 48150 3390 48195 3510
rect 48315 3390 48360 3510
rect 48480 3390 48535 3510
rect 48655 3390 48700 3510
rect 48820 3390 48865 3510
rect 48985 3390 49030 3510
rect 49150 3390 49205 3510
rect 49325 3390 49370 3510
rect 49490 3390 49535 3510
rect 49655 3390 49700 3510
rect 49820 3390 49875 3510
rect 49995 3390 50040 3510
rect 50160 3390 50205 3510
rect 50325 3390 50370 3510
rect 50490 3390 50545 3510
rect 50665 3390 50710 3510
rect 50830 3390 50875 3510
rect 50995 3390 51040 3510
rect 51160 3390 51215 3510
rect 51335 3390 51380 3510
rect 51500 3390 51545 3510
rect 51665 3390 51710 3510
rect 51830 3390 51885 3510
rect 52005 3390 52050 3510
rect 52170 3390 52215 3510
rect 52335 3390 52380 3510
rect 52500 3390 52555 3510
rect 52675 3390 52720 3510
rect 52840 3390 52885 3510
rect 53005 3390 53050 3510
rect 53170 3390 53225 3510
rect 53345 3390 53355 3510
rect 47855 3345 53355 3390
rect 47855 3225 47865 3345
rect 47985 3225 48030 3345
rect 48150 3225 48195 3345
rect 48315 3225 48360 3345
rect 48480 3225 48535 3345
rect 48655 3225 48700 3345
rect 48820 3225 48865 3345
rect 48985 3225 49030 3345
rect 49150 3225 49205 3345
rect 49325 3225 49370 3345
rect 49490 3225 49535 3345
rect 49655 3225 49700 3345
rect 49820 3225 49875 3345
rect 49995 3225 50040 3345
rect 50160 3225 50205 3345
rect 50325 3225 50370 3345
rect 50490 3225 50545 3345
rect 50665 3225 50710 3345
rect 50830 3225 50875 3345
rect 50995 3225 51040 3345
rect 51160 3225 51215 3345
rect 51335 3225 51380 3345
rect 51500 3225 51545 3345
rect 51665 3225 51710 3345
rect 51830 3225 51885 3345
rect 52005 3225 52050 3345
rect 52170 3225 52215 3345
rect 52335 3225 52380 3345
rect 52500 3225 52555 3345
rect 52675 3225 52720 3345
rect 52840 3225 52885 3345
rect 53005 3225 53050 3345
rect 53170 3225 53225 3345
rect 53345 3225 53355 3345
rect 47855 3180 53355 3225
rect 47855 3060 47865 3180
rect 47985 3060 48030 3180
rect 48150 3060 48195 3180
rect 48315 3060 48360 3180
rect 48480 3060 48535 3180
rect 48655 3060 48700 3180
rect 48820 3060 48865 3180
rect 48985 3060 49030 3180
rect 49150 3060 49205 3180
rect 49325 3060 49370 3180
rect 49490 3060 49535 3180
rect 49655 3060 49700 3180
rect 49820 3060 49875 3180
rect 49995 3060 50040 3180
rect 50160 3060 50205 3180
rect 50325 3060 50370 3180
rect 50490 3060 50545 3180
rect 50665 3060 50710 3180
rect 50830 3060 50875 3180
rect 50995 3060 51040 3180
rect 51160 3060 51215 3180
rect 51335 3060 51380 3180
rect 51500 3060 51545 3180
rect 51665 3060 51710 3180
rect 51830 3060 51885 3180
rect 52005 3060 52050 3180
rect 52170 3060 52215 3180
rect 52335 3060 52380 3180
rect 52500 3060 52555 3180
rect 52675 3060 52720 3180
rect 52840 3060 52885 3180
rect 53005 3060 53050 3180
rect 53170 3060 53225 3180
rect 53345 3060 53355 3180
rect 47855 3005 53355 3060
rect 47855 2885 47865 3005
rect 47985 2885 48030 3005
rect 48150 2885 48195 3005
rect 48315 2885 48360 3005
rect 48480 2885 48535 3005
rect 48655 2885 48700 3005
rect 48820 2885 48865 3005
rect 48985 2885 49030 3005
rect 49150 2885 49205 3005
rect 49325 2885 49370 3005
rect 49490 2885 49535 3005
rect 49655 2885 49700 3005
rect 49820 2885 49875 3005
rect 49995 2885 50040 3005
rect 50160 2885 50205 3005
rect 50325 2885 50370 3005
rect 50490 2885 50545 3005
rect 50665 2885 50710 3005
rect 50830 2885 50875 3005
rect 50995 2885 51040 3005
rect 51160 2885 51215 3005
rect 51335 2885 51380 3005
rect 51500 2885 51545 3005
rect 51665 2885 51710 3005
rect 51830 2885 51885 3005
rect 52005 2885 52050 3005
rect 52170 2885 52215 3005
rect 52335 2885 52380 3005
rect 52500 2885 52555 3005
rect 52675 2885 52720 3005
rect 52840 2885 52885 3005
rect 53005 2885 53050 3005
rect 53170 2885 53225 3005
rect 53345 2885 53355 3005
rect 47855 2840 53355 2885
rect 47855 2720 47865 2840
rect 47985 2720 48030 2840
rect 48150 2720 48195 2840
rect 48315 2720 48360 2840
rect 48480 2720 48535 2840
rect 48655 2720 48700 2840
rect 48820 2720 48865 2840
rect 48985 2720 49030 2840
rect 49150 2720 49205 2840
rect 49325 2720 49370 2840
rect 49490 2720 49535 2840
rect 49655 2720 49700 2840
rect 49820 2720 49875 2840
rect 49995 2720 50040 2840
rect 50160 2720 50205 2840
rect 50325 2720 50370 2840
rect 50490 2720 50545 2840
rect 50665 2720 50710 2840
rect 50830 2720 50875 2840
rect 50995 2720 51040 2840
rect 51160 2720 51215 2840
rect 51335 2720 51380 2840
rect 51500 2720 51545 2840
rect 51665 2720 51710 2840
rect 51830 2720 51885 2840
rect 52005 2720 52050 2840
rect 52170 2720 52215 2840
rect 52335 2720 52380 2840
rect 52500 2720 52555 2840
rect 52675 2720 52720 2840
rect 52840 2720 52885 2840
rect 53005 2720 53050 2840
rect 53170 2720 53225 2840
rect 53345 2720 53355 2840
rect 47855 2675 53355 2720
rect 47855 2555 47865 2675
rect 47985 2555 48030 2675
rect 48150 2555 48195 2675
rect 48315 2555 48360 2675
rect 48480 2555 48535 2675
rect 48655 2555 48700 2675
rect 48820 2555 48865 2675
rect 48985 2555 49030 2675
rect 49150 2555 49205 2675
rect 49325 2555 49370 2675
rect 49490 2555 49535 2675
rect 49655 2555 49700 2675
rect 49820 2555 49875 2675
rect 49995 2555 50040 2675
rect 50160 2555 50205 2675
rect 50325 2555 50370 2675
rect 50490 2555 50545 2675
rect 50665 2555 50710 2675
rect 50830 2555 50875 2675
rect 50995 2555 51040 2675
rect 51160 2555 51215 2675
rect 51335 2555 51380 2675
rect 51500 2555 51545 2675
rect 51665 2555 51710 2675
rect 51830 2555 51885 2675
rect 52005 2555 52050 2675
rect 52170 2555 52215 2675
rect 52335 2555 52380 2675
rect 52500 2555 52555 2675
rect 52675 2555 52720 2675
rect 52840 2555 52885 2675
rect 53005 2555 53050 2675
rect 53170 2555 53225 2675
rect 53345 2555 53355 2675
rect 47855 2510 53355 2555
rect 47855 2390 47865 2510
rect 47985 2390 48030 2510
rect 48150 2390 48195 2510
rect 48315 2390 48360 2510
rect 48480 2390 48535 2510
rect 48655 2390 48700 2510
rect 48820 2390 48865 2510
rect 48985 2390 49030 2510
rect 49150 2390 49205 2510
rect 49325 2390 49370 2510
rect 49490 2390 49535 2510
rect 49655 2390 49700 2510
rect 49820 2390 49875 2510
rect 49995 2390 50040 2510
rect 50160 2390 50205 2510
rect 50325 2390 50370 2510
rect 50490 2390 50545 2510
rect 50665 2390 50710 2510
rect 50830 2390 50875 2510
rect 50995 2390 51040 2510
rect 51160 2390 51215 2510
rect 51335 2390 51380 2510
rect 51500 2390 51545 2510
rect 51665 2390 51710 2510
rect 51830 2390 51885 2510
rect 52005 2390 52050 2510
rect 52170 2390 52215 2510
rect 52335 2390 52380 2510
rect 52500 2390 52555 2510
rect 52675 2390 52720 2510
rect 52840 2390 52885 2510
rect 53005 2390 53050 2510
rect 53170 2390 53225 2510
rect 53345 2390 53355 2510
rect 47855 2335 53355 2390
rect 47855 2215 47865 2335
rect 47985 2215 48030 2335
rect 48150 2215 48195 2335
rect 48315 2215 48360 2335
rect 48480 2215 48535 2335
rect 48655 2215 48700 2335
rect 48820 2215 48865 2335
rect 48985 2215 49030 2335
rect 49150 2215 49205 2335
rect 49325 2215 49370 2335
rect 49490 2215 49535 2335
rect 49655 2215 49700 2335
rect 49820 2215 49875 2335
rect 49995 2215 50040 2335
rect 50160 2215 50205 2335
rect 50325 2215 50370 2335
rect 50490 2215 50545 2335
rect 50665 2215 50710 2335
rect 50830 2215 50875 2335
rect 50995 2215 51040 2335
rect 51160 2215 51215 2335
rect 51335 2215 51380 2335
rect 51500 2215 51545 2335
rect 51665 2215 51710 2335
rect 51830 2215 51885 2335
rect 52005 2215 52050 2335
rect 52170 2215 52215 2335
rect 52335 2215 52380 2335
rect 52500 2215 52555 2335
rect 52675 2215 52720 2335
rect 52840 2215 52885 2335
rect 53005 2215 53050 2335
rect 53170 2215 53225 2335
rect 53345 2215 53355 2335
rect 47855 2170 53355 2215
rect 47855 2050 47865 2170
rect 47985 2050 48030 2170
rect 48150 2050 48195 2170
rect 48315 2050 48360 2170
rect 48480 2050 48535 2170
rect 48655 2050 48700 2170
rect 48820 2050 48865 2170
rect 48985 2050 49030 2170
rect 49150 2050 49205 2170
rect 49325 2050 49370 2170
rect 49490 2050 49535 2170
rect 49655 2050 49700 2170
rect 49820 2050 49875 2170
rect 49995 2050 50040 2170
rect 50160 2050 50205 2170
rect 50325 2050 50370 2170
rect 50490 2050 50545 2170
rect 50665 2050 50710 2170
rect 50830 2050 50875 2170
rect 50995 2050 51040 2170
rect 51160 2050 51215 2170
rect 51335 2050 51380 2170
rect 51500 2050 51545 2170
rect 51665 2050 51710 2170
rect 51830 2050 51885 2170
rect 52005 2050 52050 2170
rect 52170 2050 52215 2170
rect 52335 2050 52380 2170
rect 52500 2050 52555 2170
rect 52675 2050 52720 2170
rect 52840 2050 52885 2170
rect 53005 2050 53050 2170
rect 53170 2050 53225 2170
rect 53345 2050 53355 2170
rect 47855 2005 53355 2050
rect 47855 1885 47865 2005
rect 47985 1885 48030 2005
rect 48150 1885 48195 2005
rect 48315 1885 48360 2005
rect 48480 1885 48535 2005
rect 48655 1885 48700 2005
rect 48820 1885 48865 2005
rect 48985 1885 49030 2005
rect 49150 1885 49205 2005
rect 49325 1885 49370 2005
rect 49490 1885 49535 2005
rect 49655 1885 49700 2005
rect 49820 1885 49875 2005
rect 49995 1885 50040 2005
rect 50160 1885 50205 2005
rect 50325 1885 50370 2005
rect 50490 1885 50545 2005
rect 50665 1885 50710 2005
rect 50830 1885 50875 2005
rect 50995 1885 51040 2005
rect 51160 1885 51215 2005
rect 51335 1885 51380 2005
rect 51500 1885 51545 2005
rect 51665 1885 51710 2005
rect 51830 1885 51885 2005
rect 52005 1885 52050 2005
rect 52170 1885 52215 2005
rect 52335 1885 52380 2005
rect 52500 1885 52555 2005
rect 52675 1885 52720 2005
rect 52840 1885 52885 2005
rect 53005 1885 53050 2005
rect 53170 1885 53225 2005
rect 53345 1885 53355 2005
rect 47855 1840 53355 1885
rect 47855 1720 47865 1840
rect 47985 1720 48030 1840
rect 48150 1720 48195 1840
rect 48315 1720 48360 1840
rect 48480 1720 48535 1840
rect 48655 1720 48700 1840
rect 48820 1720 48865 1840
rect 48985 1720 49030 1840
rect 49150 1720 49205 1840
rect 49325 1720 49370 1840
rect 49490 1720 49535 1840
rect 49655 1720 49700 1840
rect 49820 1720 49875 1840
rect 49995 1720 50040 1840
rect 50160 1720 50205 1840
rect 50325 1720 50370 1840
rect 50490 1720 50545 1840
rect 50665 1720 50710 1840
rect 50830 1720 50875 1840
rect 50995 1720 51040 1840
rect 51160 1720 51215 1840
rect 51335 1720 51380 1840
rect 51500 1720 51545 1840
rect 51665 1720 51710 1840
rect 51830 1720 51885 1840
rect 52005 1720 52050 1840
rect 52170 1720 52215 1840
rect 52335 1720 52380 1840
rect 52500 1720 52555 1840
rect 52675 1720 52720 1840
rect 52840 1720 52885 1840
rect 53005 1720 53050 1840
rect 53170 1720 53225 1840
rect 53345 1720 53355 1840
rect 47855 1710 53355 1720
rect 30785 1420 36285 1430
rect 30785 1300 30795 1420
rect 30915 1300 30970 1420
rect 31090 1300 31135 1420
rect 31255 1300 31300 1420
rect 31420 1300 31465 1420
rect 31585 1300 31640 1420
rect 31760 1300 31805 1420
rect 31925 1300 31970 1420
rect 32090 1300 32135 1420
rect 32255 1300 32310 1420
rect 32430 1300 32475 1420
rect 32595 1300 32640 1420
rect 32760 1300 32805 1420
rect 32925 1300 32980 1420
rect 33100 1300 33145 1420
rect 33265 1300 33310 1420
rect 33430 1300 33475 1420
rect 33595 1300 33650 1420
rect 33770 1300 33815 1420
rect 33935 1300 33980 1420
rect 34100 1300 34145 1420
rect 34265 1300 34320 1420
rect 34440 1300 34485 1420
rect 34605 1300 34650 1420
rect 34770 1300 34815 1420
rect 34935 1300 34990 1420
rect 35110 1300 35155 1420
rect 35275 1300 35320 1420
rect 35440 1300 35485 1420
rect 35605 1300 35660 1420
rect 35780 1300 35825 1420
rect 35945 1300 35990 1420
rect 36110 1300 36155 1420
rect 36275 1300 36285 1420
rect 30785 1255 36285 1300
rect 30785 1135 30795 1255
rect 30915 1135 30970 1255
rect 31090 1135 31135 1255
rect 31255 1135 31300 1255
rect 31420 1135 31465 1255
rect 31585 1135 31640 1255
rect 31760 1135 31805 1255
rect 31925 1135 31970 1255
rect 32090 1135 32135 1255
rect 32255 1135 32310 1255
rect 32430 1135 32475 1255
rect 32595 1135 32640 1255
rect 32760 1135 32805 1255
rect 32925 1135 32980 1255
rect 33100 1135 33145 1255
rect 33265 1135 33310 1255
rect 33430 1135 33475 1255
rect 33595 1135 33650 1255
rect 33770 1135 33815 1255
rect 33935 1135 33980 1255
rect 34100 1135 34145 1255
rect 34265 1135 34320 1255
rect 34440 1135 34485 1255
rect 34605 1135 34650 1255
rect 34770 1135 34815 1255
rect 34935 1135 34990 1255
rect 35110 1135 35155 1255
rect 35275 1135 35320 1255
rect 35440 1135 35485 1255
rect 35605 1135 35660 1255
rect 35780 1135 35825 1255
rect 35945 1135 35990 1255
rect 36110 1135 36155 1255
rect 36275 1135 36285 1255
rect 30785 1090 36285 1135
rect 30785 970 30795 1090
rect 30915 970 30970 1090
rect 31090 970 31135 1090
rect 31255 970 31300 1090
rect 31420 970 31465 1090
rect 31585 970 31640 1090
rect 31760 970 31805 1090
rect 31925 970 31970 1090
rect 32090 970 32135 1090
rect 32255 970 32310 1090
rect 32430 970 32475 1090
rect 32595 970 32640 1090
rect 32760 970 32805 1090
rect 32925 970 32980 1090
rect 33100 970 33145 1090
rect 33265 970 33310 1090
rect 33430 970 33475 1090
rect 33595 970 33650 1090
rect 33770 970 33815 1090
rect 33935 970 33980 1090
rect 34100 970 34145 1090
rect 34265 970 34320 1090
rect 34440 970 34485 1090
rect 34605 970 34650 1090
rect 34770 970 34815 1090
rect 34935 970 34990 1090
rect 35110 970 35155 1090
rect 35275 970 35320 1090
rect 35440 970 35485 1090
rect 35605 970 35660 1090
rect 35780 970 35825 1090
rect 35945 970 35990 1090
rect 36110 970 36155 1090
rect 36275 970 36285 1090
rect 30785 925 36285 970
rect 30785 805 30795 925
rect 30915 805 30970 925
rect 31090 805 31135 925
rect 31255 805 31300 925
rect 31420 805 31465 925
rect 31585 805 31640 925
rect 31760 805 31805 925
rect 31925 805 31970 925
rect 32090 805 32135 925
rect 32255 805 32310 925
rect 32430 805 32475 925
rect 32595 805 32640 925
rect 32760 805 32805 925
rect 32925 805 32980 925
rect 33100 805 33145 925
rect 33265 805 33310 925
rect 33430 805 33475 925
rect 33595 805 33650 925
rect 33770 805 33815 925
rect 33935 805 33980 925
rect 34100 805 34145 925
rect 34265 805 34320 925
rect 34440 805 34485 925
rect 34605 805 34650 925
rect 34770 805 34815 925
rect 34935 805 34990 925
rect 35110 805 35155 925
rect 35275 805 35320 925
rect 35440 805 35485 925
rect 35605 805 35660 925
rect 35780 805 35825 925
rect 35945 805 35990 925
rect 36110 805 36155 925
rect 36275 805 36285 925
rect 30785 750 36285 805
rect 30785 630 30795 750
rect 30915 630 30970 750
rect 31090 630 31135 750
rect 31255 630 31300 750
rect 31420 630 31465 750
rect 31585 630 31640 750
rect 31760 630 31805 750
rect 31925 630 31970 750
rect 32090 630 32135 750
rect 32255 630 32310 750
rect 32430 630 32475 750
rect 32595 630 32640 750
rect 32760 630 32805 750
rect 32925 630 32980 750
rect 33100 630 33145 750
rect 33265 630 33310 750
rect 33430 630 33475 750
rect 33595 630 33650 750
rect 33770 630 33815 750
rect 33935 630 33980 750
rect 34100 630 34145 750
rect 34265 630 34320 750
rect 34440 630 34485 750
rect 34605 630 34650 750
rect 34770 630 34815 750
rect 34935 630 34990 750
rect 35110 630 35155 750
rect 35275 630 35320 750
rect 35440 630 35485 750
rect 35605 630 35660 750
rect 35780 630 35825 750
rect 35945 630 35990 750
rect 36110 630 36155 750
rect 36275 630 36285 750
rect 30785 585 36285 630
rect 30785 465 30795 585
rect 30915 465 30970 585
rect 31090 465 31135 585
rect 31255 465 31300 585
rect 31420 465 31465 585
rect 31585 465 31640 585
rect 31760 465 31805 585
rect 31925 465 31970 585
rect 32090 465 32135 585
rect 32255 465 32310 585
rect 32430 465 32475 585
rect 32595 465 32640 585
rect 32760 465 32805 585
rect 32925 465 32980 585
rect 33100 465 33145 585
rect 33265 465 33310 585
rect 33430 465 33475 585
rect 33595 465 33650 585
rect 33770 465 33815 585
rect 33935 465 33980 585
rect 34100 465 34145 585
rect 34265 465 34320 585
rect 34440 465 34485 585
rect 34605 465 34650 585
rect 34770 465 34815 585
rect 34935 465 34990 585
rect 35110 465 35155 585
rect 35275 465 35320 585
rect 35440 465 35485 585
rect 35605 465 35660 585
rect 35780 465 35825 585
rect 35945 465 35990 585
rect 36110 465 36155 585
rect 36275 465 36285 585
rect 30785 420 36285 465
rect 30785 300 30795 420
rect 30915 300 30970 420
rect 31090 300 31135 420
rect 31255 300 31300 420
rect 31420 300 31465 420
rect 31585 300 31640 420
rect 31760 300 31805 420
rect 31925 300 31970 420
rect 32090 300 32135 420
rect 32255 300 32310 420
rect 32430 300 32475 420
rect 32595 300 32640 420
rect 32760 300 32805 420
rect 32925 300 32980 420
rect 33100 300 33145 420
rect 33265 300 33310 420
rect 33430 300 33475 420
rect 33595 300 33650 420
rect 33770 300 33815 420
rect 33935 300 33980 420
rect 34100 300 34145 420
rect 34265 300 34320 420
rect 34440 300 34485 420
rect 34605 300 34650 420
rect 34770 300 34815 420
rect 34935 300 34990 420
rect 35110 300 35155 420
rect 35275 300 35320 420
rect 35440 300 35485 420
rect 35605 300 35660 420
rect 35780 300 35825 420
rect 35945 300 35990 420
rect 36110 300 36155 420
rect 36275 300 36285 420
rect 30785 255 36285 300
rect 30785 135 30795 255
rect 30915 135 30970 255
rect 31090 135 31135 255
rect 31255 135 31300 255
rect 31420 135 31465 255
rect 31585 135 31640 255
rect 31760 135 31805 255
rect 31925 135 31970 255
rect 32090 135 32135 255
rect 32255 135 32310 255
rect 32430 135 32475 255
rect 32595 135 32640 255
rect 32760 135 32805 255
rect 32925 135 32980 255
rect 33100 135 33145 255
rect 33265 135 33310 255
rect 33430 135 33475 255
rect 33595 135 33650 255
rect 33770 135 33815 255
rect 33935 135 33980 255
rect 34100 135 34145 255
rect 34265 135 34320 255
rect 34440 135 34485 255
rect 34605 135 34650 255
rect 34770 135 34815 255
rect 34935 135 34990 255
rect 35110 135 35155 255
rect 35275 135 35320 255
rect 35440 135 35485 255
rect 35605 135 35660 255
rect 35780 135 35825 255
rect 35945 135 35990 255
rect 36110 135 36155 255
rect 36275 135 36285 255
rect 30785 80 36285 135
rect 30785 -40 30795 80
rect 30915 -40 30970 80
rect 31090 -40 31135 80
rect 31255 -40 31300 80
rect 31420 -40 31465 80
rect 31585 -40 31640 80
rect 31760 -40 31805 80
rect 31925 -40 31970 80
rect 32090 -40 32135 80
rect 32255 -40 32310 80
rect 32430 -40 32475 80
rect 32595 -40 32640 80
rect 32760 -40 32805 80
rect 32925 -40 32980 80
rect 33100 -40 33145 80
rect 33265 -40 33310 80
rect 33430 -40 33475 80
rect 33595 -40 33650 80
rect 33770 -40 33815 80
rect 33935 -40 33980 80
rect 34100 -40 34145 80
rect 34265 -40 34320 80
rect 34440 -40 34485 80
rect 34605 -40 34650 80
rect 34770 -40 34815 80
rect 34935 -40 34990 80
rect 35110 -40 35155 80
rect 35275 -40 35320 80
rect 35440 -40 35485 80
rect 35605 -40 35660 80
rect 35780 -40 35825 80
rect 35945 -40 35990 80
rect 36110 -40 36155 80
rect 36275 -40 36285 80
rect 30785 -85 36285 -40
rect 30785 -205 30795 -85
rect 30915 -205 30970 -85
rect 31090 -205 31135 -85
rect 31255 -205 31300 -85
rect 31420 -205 31465 -85
rect 31585 -205 31640 -85
rect 31760 -205 31805 -85
rect 31925 -205 31970 -85
rect 32090 -205 32135 -85
rect 32255 -205 32310 -85
rect 32430 -205 32475 -85
rect 32595 -205 32640 -85
rect 32760 -205 32805 -85
rect 32925 -205 32980 -85
rect 33100 -205 33145 -85
rect 33265 -205 33310 -85
rect 33430 -205 33475 -85
rect 33595 -205 33650 -85
rect 33770 -205 33815 -85
rect 33935 -205 33980 -85
rect 34100 -205 34145 -85
rect 34265 -205 34320 -85
rect 34440 -205 34485 -85
rect 34605 -205 34650 -85
rect 34770 -205 34815 -85
rect 34935 -205 34990 -85
rect 35110 -205 35155 -85
rect 35275 -205 35320 -85
rect 35440 -205 35485 -85
rect 35605 -205 35660 -85
rect 35780 -205 35825 -85
rect 35945 -205 35990 -85
rect 36110 -205 36155 -85
rect 36275 -205 36285 -85
rect 30785 -250 36285 -205
rect 30785 -370 30795 -250
rect 30915 -370 30970 -250
rect 31090 -370 31135 -250
rect 31255 -370 31300 -250
rect 31420 -370 31465 -250
rect 31585 -370 31640 -250
rect 31760 -370 31805 -250
rect 31925 -370 31970 -250
rect 32090 -370 32135 -250
rect 32255 -370 32310 -250
rect 32430 -370 32475 -250
rect 32595 -370 32640 -250
rect 32760 -370 32805 -250
rect 32925 -370 32980 -250
rect 33100 -370 33145 -250
rect 33265 -370 33310 -250
rect 33430 -370 33475 -250
rect 33595 -370 33650 -250
rect 33770 -370 33815 -250
rect 33935 -370 33980 -250
rect 34100 -370 34145 -250
rect 34265 -370 34320 -250
rect 34440 -370 34485 -250
rect 34605 -370 34650 -250
rect 34770 -370 34815 -250
rect 34935 -370 34990 -250
rect 35110 -370 35155 -250
rect 35275 -370 35320 -250
rect 35440 -370 35485 -250
rect 35605 -370 35660 -250
rect 35780 -370 35825 -250
rect 35945 -370 35990 -250
rect 36110 -370 36155 -250
rect 36275 -370 36285 -250
rect 30785 -415 36285 -370
rect 30785 -535 30795 -415
rect 30915 -535 30970 -415
rect 31090 -535 31135 -415
rect 31255 -535 31300 -415
rect 31420 -535 31465 -415
rect 31585 -535 31640 -415
rect 31760 -535 31805 -415
rect 31925 -535 31970 -415
rect 32090 -535 32135 -415
rect 32255 -535 32310 -415
rect 32430 -535 32475 -415
rect 32595 -535 32640 -415
rect 32760 -535 32805 -415
rect 32925 -535 32980 -415
rect 33100 -535 33145 -415
rect 33265 -535 33310 -415
rect 33430 -535 33475 -415
rect 33595 -535 33650 -415
rect 33770 -535 33815 -415
rect 33935 -535 33980 -415
rect 34100 -535 34145 -415
rect 34265 -535 34320 -415
rect 34440 -535 34485 -415
rect 34605 -535 34650 -415
rect 34770 -535 34815 -415
rect 34935 -535 34990 -415
rect 35110 -535 35155 -415
rect 35275 -535 35320 -415
rect 35440 -535 35485 -415
rect 35605 -535 35660 -415
rect 35780 -535 35825 -415
rect 35945 -535 35990 -415
rect 36110 -535 36155 -415
rect 36275 -535 36285 -415
rect 30785 -590 36285 -535
rect 30785 -710 30795 -590
rect 30915 -710 30970 -590
rect 31090 -710 31135 -590
rect 31255 -710 31300 -590
rect 31420 -710 31465 -590
rect 31585 -710 31640 -590
rect 31760 -710 31805 -590
rect 31925 -710 31970 -590
rect 32090 -710 32135 -590
rect 32255 -710 32310 -590
rect 32430 -710 32475 -590
rect 32595 -710 32640 -590
rect 32760 -710 32805 -590
rect 32925 -710 32980 -590
rect 33100 -710 33145 -590
rect 33265 -710 33310 -590
rect 33430 -710 33475 -590
rect 33595 -710 33650 -590
rect 33770 -710 33815 -590
rect 33935 -710 33980 -590
rect 34100 -710 34145 -590
rect 34265 -710 34320 -590
rect 34440 -710 34485 -590
rect 34605 -710 34650 -590
rect 34770 -710 34815 -590
rect 34935 -710 34990 -590
rect 35110 -710 35155 -590
rect 35275 -710 35320 -590
rect 35440 -710 35485 -590
rect 35605 -710 35660 -590
rect 35780 -710 35825 -590
rect 35945 -710 35990 -590
rect 36110 -710 36155 -590
rect 36275 -710 36285 -590
rect 30785 -755 36285 -710
rect 30785 -875 30795 -755
rect 30915 -875 30970 -755
rect 31090 -875 31135 -755
rect 31255 -875 31300 -755
rect 31420 -875 31465 -755
rect 31585 -875 31640 -755
rect 31760 -875 31805 -755
rect 31925 -875 31970 -755
rect 32090 -875 32135 -755
rect 32255 -875 32310 -755
rect 32430 -875 32475 -755
rect 32595 -875 32640 -755
rect 32760 -875 32805 -755
rect 32925 -875 32980 -755
rect 33100 -875 33145 -755
rect 33265 -875 33310 -755
rect 33430 -875 33475 -755
rect 33595 -875 33650 -755
rect 33770 -875 33815 -755
rect 33935 -875 33980 -755
rect 34100 -875 34145 -755
rect 34265 -875 34320 -755
rect 34440 -875 34485 -755
rect 34605 -875 34650 -755
rect 34770 -875 34815 -755
rect 34935 -875 34990 -755
rect 35110 -875 35155 -755
rect 35275 -875 35320 -755
rect 35440 -875 35485 -755
rect 35605 -875 35660 -755
rect 35780 -875 35825 -755
rect 35945 -875 35990 -755
rect 36110 -875 36155 -755
rect 36275 -875 36285 -755
rect 30785 -920 36285 -875
rect 30785 -1040 30795 -920
rect 30915 -1040 30970 -920
rect 31090 -1040 31135 -920
rect 31255 -1040 31300 -920
rect 31420 -1040 31465 -920
rect 31585 -1040 31640 -920
rect 31760 -1040 31805 -920
rect 31925 -1040 31970 -920
rect 32090 -1040 32135 -920
rect 32255 -1040 32310 -920
rect 32430 -1040 32475 -920
rect 32595 -1040 32640 -920
rect 32760 -1040 32805 -920
rect 32925 -1040 32980 -920
rect 33100 -1040 33145 -920
rect 33265 -1040 33310 -920
rect 33430 -1040 33475 -920
rect 33595 -1040 33650 -920
rect 33770 -1040 33815 -920
rect 33935 -1040 33980 -920
rect 34100 -1040 34145 -920
rect 34265 -1040 34320 -920
rect 34440 -1040 34485 -920
rect 34605 -1040 34650 -920
rect 34770 -1040 34815 -920
rect 34935 -1040 34990 -920
rect 35110 -1040 35155 -920
rect 35275 -1040 35320 -920
rect 35440 -1040 35485 -920
rect 35605 -1040 35660 -920
rect 35780 -1040 35825 -920
rect 35945 -1040 35990 -920
rect 36110 -1040 36155 -920
rect 36275 -1040 36285 -920
rect 30785 -1085 36285 -1040
rect 30785 -1205 30795 -1085
rect 30915 -1205 30970 -1085
rect 31090 -1205 31135 -1085
rect 31255 -1205 31300 -1085
rect 31420 -1205 31465 -1085
rect 31585 -1205 31640 -1085
rect 31760 -1205 31805 -1085
rect 31925 -1205 31970 -1085
rect 32090 -1205 32135 -1085
rect 32255 -1205 32310 -1085
rect 32430 -1205 32475 -1085
rect 32595 -1205 32640 -1085
rect 32760 -1205 32805 -1085
rect 32925 -1205 32980 -1085
rect 33100 -1205 33145 -1085
rect 33265 -1205 33310 -1085
rect 33430 -1205 33475 -1085
rect 33595 -1205 33650 -1085
rect 33770 -1205 33815 -1085
rect 33935 -1205 33980 -1085
rect 34100 -1205 34145 -1085
rect 34265 -1205 34320 -1085
rect 34440 -1205 34485 -1085
rect 34605 -1205 34650 -1085
rect 34770 -1205 34815 -1085
rect 34935 -1205 34990 -1085
rect 35110 -1205 35155 -1085
rect 35275 -1205 35320 -1085
rect 35440 -1205 35485 -1085
rect 35605 -1205 35660 -1085
rect 35780 -1205 35825 -1085
rect 35945 -1205 35990 -1085
rect 36110 -1205 36155 -1085
rect 36275 -1205 36285 -1085
rect 30785 -1260 36285 -1205
rect 30785 -1380 30795 -1260
rect 30915 -1380 30970 -1260
rect 31090 -1380 31135 -1260
rect 31255 -1380 31300 -1260
rect 31420 -1380 31465 -1260
rect 31585 -1380 31640 -1260
rect 31760 -1380 31805 -1260
rect 31925 -1380 31970 -1260
rect 32090 -1380 32135 -1260
rect 32255 -1380 32310 -1260
rect 32430 -1380 32475 -1260
rect 32595 -1380 32640 -1260
rect 32760 -1380 32805 -1260
rect 32925 -1380 32980 -1260
rect 33100 -1380 33145 -1260
rect 33265 -1380 33310 -1260
rect 33430 -1380 33475 -1260
rect 33595 -1380 33650 -1260
rect 33770 -1380 33815 -1260
rect 33935 -1380 33980 -1260
rect 34100 -1380 34145 -1260
rect 34265 -1380 34320 -1260
rect 34440 -1380 34485 -1260
rect 34605 -1380 34650 -1260
rect 34770 -1380 34815 -1260
rect 34935 -1380 34990 -1260
rect 35110 -1380 35155 -1260
rect 35275 -1380 35320 -1260
rect 35440 -1380 35485 -1260
rect 35605 -1380 35660 -1260
rect 35780 -1380 35825 -1260
rect 35945 -1380 35990 -1260
rect 36110 -1380 36155 -1260
rect 36275 -1380 36285 -1260
rect 30785 -1425 36285 -1380
rect 30785 -1545 30795 -1425
rect 30915 -1545 30970 -1425
rect 31090 -1545 31135 -1425
rect 31255 -1545 31300 -1425
rect 31420 -1545 31465 -1425
rect 31585 -1545 31640 -1425
rect 31760 -1545 31805 -1425
rect 31925 -1545 31970 -1425
rect 32090 -1545 32135 -1425
rect 32255 -1545 32310 -1425
rect 32430 -1545 32475 -1425
rect 32595 -1545 32640 -1425
rect 32760 -1545 32805 -1425
rect 32925 -1545 32980 -1425
rect 33100 -1545 33145 -1425
rect 33265 -1545 33310 -1425
rect 33430 -1545 33475 -1425
rect 33595 -1545 33650 -1425
rect 33770 -1545 33815 -1425
rect 33935 -1545 33980 -1425
rect 34100 -1545 34145 -1425
rect 34265 -1545 34320 -1425
rect 34440 -1545 34485 -1425
rect 34605 -1545 34650 -1425
rect 34770 -1545 34815 -1425
rect 34935 -1545 34990 -1425
rect 35110 -1545 35155 -1425
rect 35275 -1545 35320 -1425
rect 35440 -1545 35485 -1425
rect 35605 -1545 35660 -1425
rect 35780 -1545 35825 -1425
rect 35945 -1545 35990 -1425
rect 36110 -1545 36155 -1425
rect 36275 -1545 36285 -1425
rect 30785 -1590 36285 -1545
rect 30785 -1710 30795 -1590
rect 30915 -1710 30970 -1590
rect 31090 -1710 31135 -1590
rect 31255 -1710 31300 -1590
rect 31420 -1710 31465 -1590
rect 31585 -1710 31640 -1590
rect 31760 -1710 31805 -1590
rect 31925 -1710 31970 -1590
rect 32090 -1710 32135 -1590
rect 32255 -1710 32310 -1590
rect 32430 -1710 32475 -1590
rect 32595 -1710 32640 -1590
rect 32760 -1710 32805 -1590
rect 32925 -1710 32980 -1590
rect 33100 -1710 33145 -1590
rect 33265 -1710 33310 -1590
rect 33430 -1710 33475 -1590
rect 33595 -1710 33650 -1590
rect 33770 -1710 33815 -1590
rect 33935 -1710 33980 -1590
rect 34100 -1710 34145 -1590
rect 34265 -1710 34320 -1590
rect 34440 -1710 34485 -1590
rect 34605 -1710 34650 -1590
rect 34770 -1710 34815 -1590
rect 34935 -1710 34990 -1590
rect 35110 -1710 35155 -1590
rect 35275 -1710 35320 -1590
rect 35440 -1710 35485 -1590
rect 35605 -1710 35660 -1590
rect 35780 -1710 35825 -1590
rect 35945 -1710 35990 -1590
rect 36110 -1710 36155 -1590
rect 36275 -1710 36285 -1590
rect 30785 -1755 36285 -1710
rect 30785 -1875 30795 -1755
rect 30915 -1875 30970 -1755
rect 31090 -1875 31135 -1755
rect 31255 -1875 31300 -1755
rect 31420 -1875 31465 -1755
rect 31585 -1875 31640 -1755
rect 31760 -1875 31805 -1755
rect 31925 -1875 31970 -1755
rect 32090 -1875 32135 -1755
rect 32255 -1875 32310 -1755
rect 32430 -1875 32475 -1755
rect 32595 -1875 32640 -1755
rect 32760 -1875 32805 -1755
rect 32925 -1875 32980 -1755
rect 33100 -1875 33145 -1755
rect 33265 -1875 33310 -1755
rect 33430 -1875 33475 -1755
rect 33595 -1875 33650 -1755
rect 33770 -1875 33815 -1755
rect 33935 -1875 33980 -1755
rect 34100 -1875 34145 -1755
rect 34265 -1875 34320 -1755
rect 34440 -1875 34485 -1755
rect 34605 -1875 34650 -1755
rect 34770 -1875 34815 -1755
rect 34935 -1875 34990 -1755
rect 35110 -1875 35155 -1755
rect 35275 -1875 35320 -1755
rect 35440 -1875 35485 -1755
rect 35605 -1875 35660 -1755
rect 35780 -1875 35825 -1755
rect 35945 -1875 35990 -1755
rect 36110 -1875 36155 -1755
rect 36275 -1875 36285 -1755
rect 30785 -1930 36285 -1875
rect 30785 -2050 30795 -1930
rect 30915 -2050 30970 -1930
rect 31090 -2050 31135 -1930
rect 31255 -2050 31300 -1930
rect 31420 -2050 31465 -1930
rect 31585 -2050 31640 -1930
rect 31760 -2050 31805 -1930
rect 31925 -2050 31970 -1930
rect 32090 -2050 32135 -1930
rect 32255 -2050 32310 -1930
rect 32430 -2050 32475 -1930
rect 32595 -2050 32640 -1930
rect 32760 -2050 32805 -1930
rect 32925 -2050 32980 -1930
rect 33100 -2050 33145 -1930
rect 33265 -2050 33310 -1930
rect 33430 -2050 33475 -1930
rect 33595 -2050 33650 -1930
rect 33770 -2050 33815 -1930
rect 33935 -2050 33980 -1930
rect 34100 -2050 34145 -1930
rect 34265 -2050 34320 -1930
rect 34440 -2050 34485 -1930
rect 34605 -2050 34650 -1930
rect 34770 -2050 34815 -1930
rect 34935 -2050 34990 -1930
rect 35110 -2050 35155 -1930
rect 35275 -2050 35320 -1930
rect 35440 -2050 35485 -1930
rect 35605 -2050 35660 -1930
rect 35780 -2050 35825 -1930
rect 35945 -2050 35990 -1930
rect 36110 -2050 36155 -1930
rect 36275 -2050 36285 -1930
rect 30785 -2095 36285 -2050
rect 30785 -2215 30795 -2095
rect 30915 -2215 30970 -2095
rect 31090 -2215 31135 -2095
rect 31255 -2215 31300 -2095
rect 31420 -2215 31465 -2095
rect 31585 -2215 31640 -2095
rect 31760 -2215 31805 -2095
rect 31925 -2215 31970 -2095
rect 32090 -2215 32135 -2095
rect 32255 -2215 32310 -2095
rect 32430 -2215 32475 -2095
rect 32595 -2215 32640 -2095
rect 32760 -2215 32805 -2095
rect 32925 -2215 32980 -2095
rect 33100 -2215 33145 -2095
rect 33265 -2215 33310 -2095
rect 33430 -2215 33475 -2095
rect 33595 -2215 33650 -2095
rect 33770 -2215 33815 -2095
rect 33935 -2215 33980 -2095
rect 34100 -2215 34145 -2095
rect 34265 -2215 34320 -2095
rect 34440 -2215 34485 -2095
rect 34605 -2215 34650 -2095
rect 34770 -2215 34815 -2095
rect 34935 -2215 34990 -2095
rect 35110 -2215 35155 -2095
rect 35275 -2215 35320 -2095
rect 35440 -2215 35485 -2095
rect 35605 -2215 35660 -2095
rect 35780 -2215 35825 -2095
rect 35945 -2215 35990 -2095
rect 36110 -2215 36155 -2095
rect 36275 -2215 36285 -2095
rect 30785 -2260 36285 -2215
rect 30785 -2380 30795 -2260
rect 30915 -2380 30970 -2260
rect 31090 -2380 31135 -2260
rect 31255 -2380 31300 -2260
rect 31420 -2380 31465 -2260
rect 31585 -2380 31640 -2260
rect 31760 -2380 31805 -2260
rect 31925 -2380 31970 -2260
rect 32090 -2380 32135 -2260
rect 32255 -2380 32310 -2260
rect 32430 -2380 32475 -2260
rect 32595 -2380 32640 -2260
rect 32760 -2380 32805 -2260
rect 32925 -2380 32980 -2260
rect 33100 -2380 33145 -2260
rect 33265 -2380 33310 -2260
rect 33430 -2380 33475 -2260
rect 33595 -2380 33650 -2260
rect 33770 -2380 33815 -2260
rect 33935 -2380 33980 -2260
rect 34100 -2380 34145 -2260
rect 34265 -2380 34320 -2260
rect 34440 -2380 34485 -2260
rect 34605 -2380 34650 -2260
rect 34770 -2380 34815 -2260
rect 34935 -2380 34990 -2260
rect 35110 -2380 35155 -2260
rect 35275 -2380 35320 -2260
rect 35440 -2380 35485 -2260
rect 35605 -2380 35660 -2260
rect 35780 -2380 35825 -2260
rect 35945 -2380 35990 -2260
rect 36110 -2380 36155 -2260
rect 36275 -2380 36285 -2260
rect 30785 -2425 36285 -2380
rect 30785 -2545 30795 -2425
rect 30915 -2545 30970 -2425
rect 31090 -2545 31135 -2425
rect 31255 -2545 31300 -2425
rect 31420 -2545 31465 -2425
rect 31585 -2545 31640 -2425
rect 31760 -2545 31805 -2425
rect 31925 -2545 31970 -2425
rect 32090 -2545 32135 -2425
rect 32255 -2545 32310 -2425
rect 32430 -2545 32475 -2425
rect 32595 -2545 32640 -2425
rect 32760 -2545 32805 -2425
rect 32925 -2545 32980 -2425
rect 33100 -2545 33145 -2425
rect 33265 -2545 33310 -2425
rect 33430 -2545 33475 -2425
rect 33595 -2545 33650 -2425
rect 33770 -2545 33815 -2425
rect 33935 -2545 33980 -2425
rect 34100 -2545 34145 -2425
rect 34265 -2545 34320 -2425
rect 34440 -2545 34485 -2425
rect 34605 -2545 34650 -2425
rect 34770 -2545 34815 -2425
rect 34935 -2545 34990 -2425
rect 35110 -2545 35155 -2425
rect 35275 -2545 35320 -2425
rect 35440 -2545 35485 -2425
rect 35605 -2545 35660 -2425
rect 35780 -2545 35825 -2425
rect 35945 -2545 35990 -2425
rect 36110 -2545 36155 -2425
rect 36275 -2545 36285 -2425
rect 30785 -2600 36285 -2545
rect 30785 -2720 30795 -2600
rect 30915 -2720 30970 -2600
rect 31090 -2720 31135 -2600
rect 31255 -2720 31300 -2600
rect 31420 -2720 31465 -2600
rect 31585 -2720 31640 -2600
rect 31760 -2720 31805 -2600
rect 31925 -2720 31970 -2600
rect 32090 -2720 32135 -2600
rect 32255 -2720 32310 -2600
rect 32430 -2720 32475 -2600
rect 32595 -2720 32640 -2600
rect 32760 -2720 32805 -2600
rect 32925 -2720 32980 -2600
rect 33100 -2720 33145 -2600
rect 33265 -2720 33310 -2600
rect 33430 -2720 33475 -2600
rect 33595 -2720 33650 -2600
rect 33770 -2720 33815 -2600
rect 33935 -2720 33980 -2600
rect 34100 -2720 34145 -2600
rect 34265 -2720 34320 -2600
rect 34440 -2720 34485 -2600
rect 34605 -2720 34650 -2600
rect 34770 -2720 34815 -2600
rect 34935 -2720 34990 -2600
rect 35110 -2720 35155 -2600
rect 35275 -2720 35320 -2600
rect 35440 -2720 35485 -2600
rect 35605 -2720 35660 -2600
rect 35780 -2720 35825 -2600
rect 35945 -2720 35990 -2600
rect 36110 -2720 36155 -2600
rect 36275 -2720 36285 -2600
rect 30785 -2765 36285 -2720
rect 30785 -2885 30795 -2765
rect 30915 -2885 30970 -2765
rect 31090 -2885 31135 -2765
rect 31255 -2885 31300 -2765
rect 31420 -2885 31465 -2765
rect 31585 -2885 31640 -2765
rect 31760 -2885 31805 -2765
rect 31925 -2885 31970 -2765
rect 32090 -2885 32135 -2765
rect 32255 -2885 32310 -2765
rect 32430 -2885 32475 -2765
rect 32595 -2885 32640 -2765
rect 32760 -2885 32805 -2765
rect 32925 -2885 32980 -2765
rect 33100 -2885 33145 -2765
rect 33265 -2885 33310 -2765
rect 33430 -2885 33475 -2765
rect 33595 -2885 33650 -2765
rect 33770 -2885 33815 -2765
rect 33935 -2885 33980 -2765
rect 34100 -2885 34145 -2765
rect 34265 -2885 34320 -2765
rect 34440 -2885 34485 -2765
rect 34605 -2885 34650 -2765
rect 34770 -2885 34815 -2765
rect 34935 -2885 34990 -2765
rect 35110 -2885 35155 -2765
rect 35275 -2885 35320 -2765
rect 35440 -2885 35485 -2765
rect 35605 -2885 35660 -2765
rect 35780 -2885 35825 -2765
rect 35945 -2885 35990 -2765
rect 36110 -2885 36155 -2765
rect 36275 -2885 36285 -2765
rect 30785 -2930 36285 -2885
rect 30785 -3050 30795 -2930
rect 30915 -3050 30970 -2930
rect 31090 -3050 31135 -2930
rect 31255 -3050 31300 -2930
rect 31420 -3050 31465 -2930
rect 31585 -3050 31640 -2930
rect 31760 -3050 31805 -2930
rect 31925 -3050 31970 -2930
rect 32090 -3050 32135 -2930
rect 32255 -3050 32310 -2930
rect 32430 -3050 32475 -2930
rect 32595 -3050 32640 -2930
rect 32760 -3050 32805 -2930
rect 32925 -3050 32980 -2930
rect 33100 -3050 33145 -2930
rect 33265 -3050 33310 -2930
rect 33430 -3050 33475 -2930
rect 33595 -3050 33650 -2930
rect 33770 -3050 33815 -2930
rect 33935 -3050 33980 -2930
rect 34100 -3050 34145 -2930
rect 34265 -3050 34320 -2930
rect 34440 -3050 34485 -2930
rect 34605 -3050 34650 -2930
rect 34770 -3050 34815 -2930
rect 34935 -3050 34990 -2930
rect 35110 -3050 35155 -2930
rect 35275 -3050 35320 -2930
rect 35440 -3050 35485 -2930
rect 35605 -3050 35660 -2930
rect 35780 -3050 35825 -2930
rect 35945 -3050 35990 -2930
rect 36110 -3050 36155 -2930
rect 36275 -3050 36285 -2930
rect 30785 -3095 36285 -3050
rect 30785 -3215 30795 -3095
rect 30915 -3215 30970 -3095
rect 31090 -3215 31135 -3095
rect 31255 -3215 31300 -3095
rect 31420 -3215 31465 -3095
rect 31585 -3215 31640 -3095
rect 31760 -3215 31805 -3095
rect 31925 -3215 31970 -3095
rect 32090 -3215 32135 -3095
rect 32255 -3215 32310 -3095
rect 32430 -3215 32475 -3095
rect 32595 -3215 32640 -3095
rect 32760 -3215 32805 -3095
rect 32925 -3215 32980 -3095
rect 33100 -3215 33145 -3095
rect 33265 -3215 33310 -3095
rect 33430 -3215 33475 -3095
rect 33595 -3215 33650 -3095
rect 33770 -3215 33815 -3095
rect 33935 -3215 33980 -3095
rect 34100 -3215 34145 -3095
rect 34265 -3215 34320 -3095
rect 34440 -3215 34485 -3095
rect 34605 -3215 34650 -3095
rect 34770 -3215 34815 -3095
rect 34935 -3215 34990 -3095
rect 35110 -3215 35155 -3095
rect 35275 -3215 35320 -3095
rect 35440 -3215 35485 -3095
rect 35605 -3215 35660 -3095
rect 35780 -3215 35825 -3095
rect 35945 -3215 35990 -3095
rect 36110 -3215 36155 -3095
rect 36275 -3215 36285 -3095
rect 30785 -3270 36285 -3215
rect 30785 -3390 30795 -3270
rect 30915 -3390 30970 -3270
rect 31090 -3390 31135 -3270
rect 31255 -3390 31300 -3270
rect 31420 -3390 31465 -3270
rect 31585 -3390 31640 -3270
rect 31760 -3390 31805 -3270
rect 31925 -3390 31970 -3270
rect 32090 -3390 32135 -3270
rect 32255 -3390 32310 -3270
rect 32430 -3390 32475 -3270
rect 32595 -3390 32640 -3270
rect 32760 -3390 32805 -3270
rect 32925 -3390 32980 -3270
rect 33100 -3390 33145 -3270
rect 33265 -3390 33310 -3270
rect 33430 -3390 33475 -3270
rect 33595 -3390 33650 -3270
rect 33770 -3390 33815 -3270
rect 33935 -3390 33980 -3270
rect 34100 -3390 34145 -3270
rect 34265 -3390 34320 -3270
rect 34440 -3390 34485 -3270
rect 34605 -3390 34650 -3270
rect 34770 -3390 34815 -3270
rect 34935 -3390 34990 -3270
rect 35110 -3390 35155 -3270
rect 35275 -3390 35320 -3270
rect 35440 -3390 35485 -3270
rect 35605 -3390 35660 -3270
rect 35780 -3390 35825 -3270
rect 35945 -3390 35990 -3270
rect 36110 -3390 36155 -3270
rect 36275 -3390 36285 -3270
rect 30785 -3435 36285 -3390
rect 30785 -3555 30795 -3435
rect 30915 -3555 30970 -3435
rect 31090 -3555 31135 -3435
rect 31255 -3555 31300 -3435
rect 31420 -3555 31465 -3435
rect 31585 -3555 31640 -3435
rect 31760 -3555 31805 -3435
rect 31925 -3555 31970 -3435
rect 32090 -3555 32135 -3435
rect 32255 -3555 32310 -3435
rect 32430 -3555 32475 -3435
rect 32595 -3555 32640 -3435
rect 32760 -3555 32805 -3435
rect 32925 -3555 32980 -3435
rect 33100 -3555 33145 -3435
rect 33265 -3555 33310 -3435
rect 33430 -3555 33475 -3435
rect 33595 -3555 33650 -3435
rect 33770 -3555 33815 -3435
rect 33935 -3555 33980 -3435
rect 34100 -3555 34145 -3435
rect 34265 -3555 34320 -3435
rect 34440 -3555 34485 -3435
rect 34605 -3555 34650 -3435
rect 34770 -3555 34815 -3435
rect 34935 -3555 34990 -3435
rect 35110 -3555 35155 -3435
rect 35275 -3555 35320 -3435
rect 35440 -3555 35485 -3435
rect 35605 -3555 35660 -3435
rect 35780 -3555 35825 -3435
rect 35945 -3555 35990 -3435
rect 36110 -3555 36155 -3435
rect 36275 -3555 36285 -3435
rect 30785 -3600 36285 -3555
rect 30785 -3720 30795 -3600
rect 30915 -3720 30970 -3600
rect 31090 -3720 31135 -3600
rect 31255 -3720 31300 -3600
rect 31420 -3720 31465 -3600
rect 31585 -3720 31640 -3600
rect 31760 -3720 31805 -3600
rect 31925 -3720 31970 -3600
rect 32090 -3720 32135 -3600
rect 32255 -3720 32310 -3600
rect 32430 -3720 32475 -3600
rect 32595 -3720 32640 -3600
rect 32760 -3720 32805 -3600
rect 32925 -3720 32980 -3600
rect 33100 -3720 33145 -3600
rect 33265 -3720 33310 -3600
rect 33430 -3720 33475 -3600
rect 33595 -3720 33650 -3600
rect 33770 -3720 33815 -3600
rect 33935 -3720 33980 -3600
rect 34100 -3720 34145 -3600
rect 34265 -3720 34320 -3600
rect 34440 -3720 34485 -3600
rect 34605 -3720 34650 -3600
rect 34770 -3720 34815 -3600
rect 34935 -3720 34990 -3600
rect 35110 -3720 35155 -3600
rect 35275 -3720 35320 -3600
rect 35440 -3720 35485 -3600
rect 35605 -3720 35660 -3600
rect 35780 -3720 35825 -3600
rect 35945 -3720 35990 -3600
rect 36110 -3720 36155 -3600
rect 36275 -3720 36285 -3600
rect 30785 -3765 36285 -3720
rect 30785 -3885 30795 -3765
rect 30915 -3885 30970 -3765
rect 31090 -3885 31135 -3765
rect 31255 -3885 31300 -3765
rect 31420 -3885 31465 -3765
rect 31585 -3885 31640 -3765
rect 31760 -3885 31805 -3765
rect 31925 -3885 31970 -3765
rect 32090 -3885 32135 -3765
rect 32255 -3885 32310 -3765
rect 32430 -3885 32475 -3765
rect 32595 -3885 32640 -3765
rect 32760 -3885 32805 -3765
rect 32925 -3885 32980 -3765
rect 33100 -3885 33145 -3765
rect 33265 -3885 33310 -3765
rect 33430 -3885 33475 -3765
rect 33595 -3885 33650 -3765
rect 33770 -3885 33815 -3765
rect 33935 -3885 33980 -3765
rect 34100 -3885 34145 -3765
rect 34265 -3885 34320 -3765
rect 34440 -3885 34485 -3765
rect 34605 -3885 34650 -3765
rect 34770 -3885 34815 -3765
rect 34935 -3885 34990 -3765
rect 35110 -3885 35155 -3765
rect 35275 -3885 35320 -3765
rect 35440 -3885 35485 -3765
rect 35605 -3885 35660 -3765
rect 35780 -3885 35825 -3765
rect 35945 -3885 35990 -3765
rect 36110 -3885 36155 -3765
rect 36275 -3885 36285 -3765
rect 30785 -3940 36285 -3885
rect 30785 -4060 30795 -3940
rect 30915 -4060 30970 -3940
rect 31090 -4060 31135 -3940
rect 31255 -4060 31300 -3940
rect 31420 -4060 31465 -3940
rect 31585 -4060 31640 -3940
rect 31760 -4060 31805 -3940
rect 31925 -4060 31970 -3940
rect 32090 -4060 32135 -3940
rect 32255 -4060 32310 -3940
rect 32430 -4060 32475 -3940
rect 32595 -4060 32640 -3940
rect 32760 -4060 32805 -3940
rect 32925 -4060 32980 -3940
rect 33100 -4060 33145 -3940
rect 33265 -4060 33310 -3940
rect 33430 -4060 33475 -3940
rect 33595 -4060 33650 -3940
rect 33770 -4060 33815 -3940
rect 33935 -4060 33980 -3940
rect 34100 -4060 34145 -3940
rect 34265 -4060 34320 -3940
rect 34440 -4060 34485 -3940
rect 34605 -4060 34650 -3940
rect 34770 -4060 34815 -3940
rect 34935 -4060 34990 -3940
rect 35110 -4060 35155 -3940
rect 35275 -4060 35320 -3940
rect 35440 -4060 35485 -3940
rect 35605 -4060 35660 -3940
rect 35780 -4060 35825 -3940
rect 35945 -4060 35990 -3940
rect 36110 -4060 36155 -3940
rect 36275 -4060 36285 -3940
rect 30785 -4070 36285 -4060
rect 36475 1420 41975 1430
rect 36475 1300 36485 1420
rect 36605 1300 36660 1420
rect 36780 1300 36825 1420
rect 36945 1300 36990 1420
rect 37110 1300 37155 1420
rect 37275 1300 37330 1420
rect 37450 1300 37495 1420
rect 37615 1300 37660 1420
rect 37780 1300 37825 1420
rect 37945 1300 38000 1420
rect 38120 1300 38165 1420
rect 38285 1300 38330 1420
rect 38450 1300 38495 1420
rect 38615 1300 38670 1420
rect 38790 1300 38835 1420
rect 38955 1300 39000 1420
rect 39120 1300 39165 1420
rect 39285 1300 39340 1420
rect 39460 1300 39505 1420
rect 39625 1300 39670 1420
rect 39790 1300 39835 1420
rect 39955 1300 40010 1420
rect 40130 1300 40175 1420
rect 40295 1300 40340 1420
rect 40460 1300 40505 1420
rect 40625 1300 40680 1420
rect 40800 1300 40845 1420
rect 40965 1300 41010 1420
rect 41130 1300 41175 1420
rect 41295 1300 41350 1420
rect 41470 1300 41515 1420
rect 41635 1300 41680 1420
rect 41800 1300 41845 1420
rect 41965 1300 41975 1420
rect 36475 1255 41975 1300
rect 36475 1135 36485 1255
rect 36605 1135 36660 1255
rect 36780 1135 36825 1255
rect 36945 1135 36990 1255
rect 37110 1135 37155 1255
rect 37275 1135 37330 1255
rect 37450 1135 37495 1255
rect 37615 1135 37660 1255
rect 37780 1135 37825 1255
rect 37945 1135 38000 1255
rect 38120 1135 38165 1255
rect 38285 1135 38330 1255
rect 38450 1135 38495 1255
rect 38615 1135 38670 1255
rect 38790 1135 38835 1255
rect 38955 1135 39000 1255
rect 39120 1135 39165 1255
rect 39285 1135 39340 1255
rect 39460 1135 39505 1255
rect 39625 1135 39670 1255
rect 39790 1135 39835 1255
rect 39955 1135 40010 1255
rect 40130 1135 40175 1255
rect 40295 1135 40340 1255
rect 40460 1135 40505 1255
rect 40625 1135 40680 1255
rect 40800 1135 40845 1255
rect 40965 1135 41010 1255
rect 41130 1135 41175 1255
rect 41295 1135 41350 1255
rect 41470 1135 41515 1255
rect 41635 1135 41680 1255
rect 41800 1135 41845 1255
rect 41965 1135 41975 1255
rect 36475 1090 41975 1135
rect 36475 970 36485 1090
rect 36605 970 36660 1090
rect 36780 970 36825 1090
rect 36945 970 36990 1090
rect 37110 970 37155 1090
rect 37275 970 37330 1090
rect 37450 970 37495 1090
rect 37615 970 37660 1090
rect 37780 970 37825 1090
rect 37945 970 38000 1090
rect 38120 970 38165 1090
rect 38285 970 38330 1090
rect 38450 970 38495 1090
rect 38615 970 38670 1090
rect 38790 970 38835 1090
rect 38955 970 39000 1090
rect 39120 970 39165 1090
rect 39285 970 39340 1090
rect 39460 970 39505 1090
rect 39625 970 39670 1090
rect 39790 970 39835 1090
rect 39955 970 40010 1090
rect 40130 970 40175 1090
rect 40295 970 40340 1090
rect 40460 970 40505 1090
rect 40625 970 40680 1090
rect 40800 970 40845 1090
rect 40965 970 41010 1090
rect 41130 970 41175 1090
rect 41295 970 41350 1090
rect 41470 970 41515 1090
rect 41635 970 41680 1090
rect 41800 970 41845 1090
rect 41965 970 41975 1090
rect 36475 925 41975 970
rect 36475 805 36485 925
rect 36605 805 36660 925
rect 36780 805 36825 925
rect 36945 805 36990 925
rect 37110 805 37155 925
rect 37275 805 37330 925
rect 37450 805 37495 925
rect 37615 805 37660 925
rect 37780 805 37825 925
rect 37945 805 38000 925
rect 38120 805 38165 925
rect 38285 805 38330 925
rect 38450 805 38495 925
rect 38615 805 38670 925
rect 38790 805 38835 925
rect 38955 805 39000 925
rect 39120 805 39165 925
rect 39285 805 39340 925
rect 39460 805 39505 925
rect 39625 805 39670 925
rect 39790 805 39835 925
rect 39955 805 40010 925
rect 40130 805 40175 925
rect 40295 805 40340 925
rect 40460 805 40505 925
rect 40625 805 40680 925
rect 40800 805 40845 925
rect 40965 805 41010 925
rect 41130 805 41175 925
rect 41295 805 41350 925
rect 41470 805 41515 925
rect 41635 805 41680 925
rect 41800 805 41845 925
rect 41965 805 41975 925
rect 36475 750 41975 805
rect 36475 630 36485 750
rect 36605 630 36660 750
rect 36780 630 36825 750
rect 36945 630 36990 750
rect 37110 630 37155 750
rect 37275 630 37330 750
rect 37450 630 37495 750
rect 37615 630 37660 750
rect 37780 630 37825 750
rect 37945 630 38000 750
rect 38120 630 38165 750
rect 38285 630 38330 750
rect 38450 630 38495 750
rect 38615 630 38670 750
rect 38790 630 38835 750
rect 38955 630 39000 750
rect 39120 630 39165 750
rect 39285 630 39340 750
rect 39460 630 39505 750
rect 39625 630 39670 750
rect 39790 630 39835 750
rect 39955 630 40010 750
rect 40130 630 40175 750
rect 40295 630 40340 750
rect 40460 630 40505 750
rect 40625 630 40680 750
rect 40800 630 40845 750
rect 40965 630 41010 750
rect 41130 630 41175 750
rect 41295 630 41350 750
rect 41470 630 41515 750
rect 41635 630 41680 750
rect 41800 630 41845 750
rect 41965 630 41975 750
rect 36475 585 41975 630
rect 36475 465 36485 585
rect 36605 465 36660 585
rect 36780 465 36825 585
rect 36945 465 36990 585
rect 37110 465 37155 585
rect 37275 465 37330 585
rect 37450 465 37495 585
rect 37615 465 37660 585
rect 37780 465 37825 585
rect 37945 465 38000 585
rect 38120 465 38165 585
rect 38285 465 38330 585
rect 38450 465 38495 585
rect 38615 465 38670 585
rect 38790 465 38835 585
rect 38955 465 39000 585
rect 39120 465 39165 585
rect 39285 465 39340 585
rect 39460 465 39505 585
rect 39625 465 39670 585
rect 39790 465 39835 585
rect 39955 465 40010 585
rect 40130 465 40175 585
rect 40295 465 40340 585
rect 40460 465 40505 585
rect 40625 465 40680 585
rect 40800 465 40845 585
rect 40965 465 41010 585
rect 41130 465 41175 585
rect 41295 465 41350 585
rect 41470 465 41515 585
rect 41635 465 41680 585
rect 41800 465 41845 585
rect 41965 465 41975 585
rect 36475 420 41975 465
rect 36475 300 36485 420
rect 36605 300 36660 420
rect 36780 300 36825 420
rect 36945 300 36990 420
rect 37110 300 37155 420
rect 37275 300 37330 420
rect 37450 300 37495 420
rect 37615 300 37660 420
rect 37780 300 37825 420
rect 37945 300 38000 420
rect 38120 300 38165 420
rect 38285 300 38330 420
rect 38450 300 38495 420
rect 38615 300 38670 420
rect 38790 300 38835 420
rect 38955 300 39000 420
rect 39120 300 39165 420
rect 39285 300 39340 420
rect 39460 300 39505 420
rect 39625 300 39670 420
rect 39790 300 39835 420
rect 39955 300 40010 420
rect 40130 300 40175 420
rect 40295 300 40340 420
rect 40460 300 40505 420
rect 40625 300 40680 420
rect 40800 300 40845 420
rect 40965 300 41010 420
rect 41130 300 41175 420
rect 41295 300 41350 420
rect 41470 300 41515 420
rect 41635 300 41680 420
rect 41800 300 41845 420
rect 41965 300 41975 420
rect 36475 255 41975 300
rect 36475 135 36485 255
rect 36605 135 36660 255
rect 36780 135 36825 255
rect 36945 135 36990 255
rect 37110 135 37155 255
rect 37275 135 37330 255
rect 37450 135 37495 255
rect 37615 135 37660 255
rect 37780 135 37825 255
rect 37945 135 38000 255
rect 38120 135 38165 255
rect 38285 135 38330 255
rect 38450 135 38495 255
rect 38615 135 38670 255
rect 38790 135 38835 255
rect 38955 135 39000 255
rect 39120 135 39165 255
rect 39285 135 39340 255
rect 39460 135 39505 255
rect 39625 135 39670 255
rect 39790 135 39835 255
rect 39955 135 40010 255
rect 40130 135 40175 255
rect 40295 135 40340 255
rect 40460 135 40505 255
rect 40625 135 40680 255
rect 40800 135 40845 255
rect 40965 135 41010 255
rect 41130 135 41175 255
rect 41295 135 41350 255
rect 41470 135 41515 255
rect 41635 135 41680 255
rect 41800 135 41845 255
rect 41965 135 41975 255
rect 36475 80 41975 135
rect 36475 -40 36485 80
rect 36605 -40 36660 80
rect 36780 -40 36825 80
rect 36945 -40 36990 80
rect 37110 -40 37155 80
rect 37275 -40 37330 80
rect 37450 -40 37495 80
rect 37615 -40 37660 80
rect 37780 -40 37825 80
rect 37945 -40 38000 80
rect 38120 -40 38165 80
rect 38285 -40 38330 80
rect 38450 -40 38495 80
rect 38615 -40 38670 80
rect 38790 -40 38835 80
rect 38955 -40 39000 80
rect 39120 -40 39165 80
rect 39285 -40 39340 80
rect 39460 -40 39505 80
rect 39625 -40 39670 80
rect 39790 -40 39835 80
rect 39955 -40 40010 80
rect 40130 -40 40175 80
rect 40295 -40 40340 80
rect 40460 -40 40505 80
rect 40625 -40 40680 80
rect 40800 -40 40845 80
rect 40965 -40 41010 80
rect 41130 -40 41175 80
rect 41295 -40 41350 80
rect 41470 -40 41515 80
rect 41635 -40 41680 80
rect 41800 -40 41845 80
rect 41965 -40 41975 80
rect 36475 -85 41975 -40
rect 36475 -205 36485 -85
rect 36605 -205 36660 -85
rect 36780 -205 36825 -85
rect 36945 -205 36990 -85
rect 37110 -205 37155 -85
rect 37275 -205 37330 -85
rect 37450 -205 37495 -85
rect 37615 -205 37660 -85
rect 37780 -205 37825 -85
rect 37945 -205 38000 -85
rect 38120 -205 38165 -85
rect 38285 -205 38330 -85
rect 38450 -205 38495 -85
rect 38615 -205 38670 -85
rect 38790 -205 38835 -85
rect 38955 -205 39000 -85
rect 39120 -205 39165 -85
rect 39285 -205 39340 -85
rect 39460 -205 39505 -85
rect 39625 -205 39670 -85
rect 39790 -205 39835 -85
rect 39955 -205 40010 -85
rect 40130 -205 40175 -85
rect 40295 -205 40340 -85
rect 40460 -205 40505 -85
rect 40625 -205 40680 -85
rect 40800 -205 40845 -85
rect 40965 -205 41010 -85
rect 41130 -205 41175 -85
rect 41295 -205 41350 -85
rect 41470 -205 41515 -85
rect 41635 -205 41680 -85
rect 41800 -205 41845 -85
rect 41965 -205 41975 -85
rect 36475 -250 41975 -205
rect 36475 -370 36485 -250
rect 36605 -370 36660 -250
rect 36780 -370 36825 -250
rect 36945 -370 36990 -250
rect 37110 -370 37155 -250
rect 37275 -370 37330 -250
rect 37450 -370 37495 -250
rect 37615 -370 37660 -250
rect 37780 -370 37825 -250
rect 37945 -370 38000 -250
rect 38120 -370 38165 -250
rect 38285 -370 38330 -250
rect 38450 -370 38495 -250
rect 38615 -370 38670 -250
rect 38790 -370 38835 -250
rect 38955 -370 39000 -250
rect 39120 -370 39165 -250
rect 39285 -370 39340 -250
rect 39460 -370 39505 -250
rect 39625 -370 39670 -250
rect 39790 -370 39835 -250
rect 39955 -370 40010 -250
rect 40130 -370 40175 -250
rect 40295 -370 40340 -250
rect 40460 -370 40505 -250
rect 40625 -370 40680 -250
rect 40800 -370 40845 -250
rect 40965 -370 41010 -250
rect 41130 -370 41175 -250
rect 41295 -370 41350 -250
rect 41470 -370 41515 -250
rect 41635 -370 41680 -250
rect 41800 -370 41845 -250
rect 41965 -370 41975 -250
rect 36475 -415 41975 -370
rect 36475 -535 36485 -415
rect 36605 -535 36660 -415
rect 36780 -535 36825 -415
rect 36945 -535 36990 -415
rect 37110 -535 37155 -415
rect 37275 -535 37330 -415
rect 37450 -535 37495 -415
rect 37615 -535 37660 -415
rect 37780 -535 37825 -415
rect 37945 -535 38000 -415
rect 38120 -535 38165 -415
rect 38285 -535 38330 -415
rect 38450 -535 38495 -415
rect 38615 -535 38670 -415
rect 38790 -535 38835 -415
rect 38955 -535 39000 -415
rect 39120 -535 39165 -415
rect 39285 -535 39340 -415
rect 39460 -535 39505 -415
rect 39625 -535 39670 -415
rect 39790 -535 39835 -415
rect 39955 -535 40010 -415
rect 40130 -535 40175 -415
rect 40295 -535 40340 -415
rect 40460 -535 40505 -415
rect 40625 -535 40680 -415
rect 40800 -535 40845 -415
rect 40965 -535 41010 -415
rect 41130 -535 41175 -415
rect 41295 -535 41350 -415
rect 41470 -535 41515 -415
rect 41635 -535 41680 -415
rect 41800 -535 41845 -415
rect 41965 -535 41975 -415
rect 36475 -590 41975 -535
rect 36475 -710 36485 -590
rect 36605 -710 36660 -590
rect 36780 -710 36825 -590
rect 36945 -710 36990 -590
rect 37110 -710 37155 -590
rect 37275 -710 37330 -590
rect 37450 -710 37495 -590
rect 37615 -710 37660 -590
rect 37780 -710 37825 -590
rect 37945 -710 38000 -590
rect 38120 -710 38165 -590
rect 38285 -710 38330 -590
rect 38450 -710 38495 -590
rect 38615 -710 38670 -590
rect 38790 -710 38835 -590
rect 38955 -710 39000 -590
rect 39120 -710 39165 -590
rect 39285 -710 39340 -590
rect 39460 -710 39505 -590
rect 39625 -710 39670 -590
rect 39790 -710 39835 -590
rect 39955 -710 40010 -590
rect 40130 -710 40175 -590
rect 40295 -710 40340 -590
rect 40460 -710 40505 -590
rect 40625 -710 40680 -590
rect 40800 -710 40845 -590
rect 40965 -710 41010 -590
rect 41130 -710 41175 -590
rect 41295 -710 41350 -590
rect 41470 -710 41515 -590
rect 41635 -710 41680 -590
rect 41800 -710 41845 -590
rect 41965 -710 41975 -590
rect 36475 -755 41975 -710
rect 36475 -875 36485 -755
rect 36605 -875 36660 -755
rect 36780 -875 36825 -755
rect 36945 -875 36990 -755
rect 37110 -875 37155 -755
rect 37275 -875 37330 -755
rect 37450 -875 37495 -755
rect 37615 -875 37660 -755
rect 37780 -875 37825 -755
rect 37945 -875 38000 -755
rect 38120 -875 38165 -755
rect 38285 -875 38330 -755
rect 38450 -875 38495 -755
rect 38615 -875 38670 -755
rect 38790 -875 38835 -755
rect 38955 -875 39000 -755
rect 39120 -875 39165 -755
rect 39285 -875 39340 -755
rect 39460 -875 39505 -755
rect 39625 -875 39670 -755
rect 39790 -875 39835 -755
rect 39955 -875 40010 -755
rect 40130 -875 40175 -755
rect 40295 -875 40340 -755
rect 40460 -875 40505 -755
rect 40625 -875 40680 -755
rect 40800 -875 40845 -755
rect 40965 -875 41010 -755
rect 41130 -875 41175 -755
rect 41295 -875 41350 -755
rect 41470 -875 41515 -755
rect 41635 -875 41680 -755
rect 41800 -875 41845 -755
rect 41965 -875 41975 -755
rect 36475 -920 41975 -875
rect 36475 -1040 36485 -920
rect 36605 -1040 36660 -920
rect 36780 -1040 36825 -920
rect 36945 -1040 36990 -920
rect 37110 -1040 37155 -920
rect 37275 -1040 37330 -920
rect 37450 -1040 37495 -920
rect 37615 -1040 37660 -920
rect 37780 -1040 37825 -920
rect 37945 -1040 38000 -920
rect 38120 -1040 38165 -920
rect 38285 -1040 38330 -920
rect 38450 -1040 38495 -920
rect 38615 -1040 38670 -920
rect 38790 -1040 38835 -920
rect 38955 -1040 39000 -920
rect 39120 -1040 39165 -920
rect 39285 -1040 39340 -920
rect 39460 -1040 39505 -920
rect 39625 -1040 39670 -920
rect 39790 -1040 39835 -920
rect 39955 -1040 40010 -920
rect 40130 -1040 40175 -920
rect 40295 -1040 40340 -920
rect 40460 -1040 40505 -920
rect 40625 -1040 40680 -920
rect 40800 -1040 40845 -920
rect 40965 -1040 41010 -920
rect 41130 -1040 41175 -920
rect 41295 -1040 41350 -920
rect 41470 -1040 41515 -920
rect 41635 -1040 41680 -920
rect 41800 -1040 41845 -920
rect 41965 -1040 41975 -920
rect 36475 -1085 41975 -1040
rect 36475 -1205 36485 -1085
rect 36605 -1205 36660 -1085
rect 36780 -1205 36825 -1085
rect 36945 -1205 36990 -1085
rect 37110 -1205 37155 -1085
rect 37275 -1205 37330 -1085
rect 37450 -1205 37495 -1085
rect 37615 -1205 37660 -1085
rect 37780 -1205 37825 -1085
rect 37945 -1205 38000 -1085
rect 38120 -1205 38165 -1085
rect 38285 -1205 38330 -1085
rect 38450 -1205 38495 -1085
rect 38615 -1205 38670 -1085
rect 38790 -1205 38835 -1085
rect 38955 -1205 39000 -1085
rect 39120 -1205 39165 -1085
rect 39285 -1205 39340 -1085
rect 39460 -1205 39505 -1085
rect 39625 -1205 39670 -1085
rect 39790 -1205 39835 -1085
rect 39955 -1205 40010 -1085
rect 40130 -1205 40175 -1085
rect 40295 -1205 40340 -1085
rect 40460 -1205 40505 -1085
rect 40625 -1205 40680 -1085
rect 40800 -1205 40845 -1085
rect 40965 -1205 41010 -1085
rect 41130 -1205 41175 -1085
rect 41295 -1205 41350 -1085
rect 41470 -1205 41515 -1085
rect 41635 -1205 41680 -1085
rect 41800 -1205 41845 -1085
rect 41965 -1205 41975 -1085
rect 36475 -1260 41975 -1205
rect 36475 -1380 36485 -1260
rect 36605 -1380 36660 -1260
rect 36780 -1380 36825 -1260
rect 36945 -1380 36990 -1260
rect 37110 -1380 37155 -1260
rect 37275 -1380 37330 -1260
rect 37450 -1380 37495 -1260
rect 37615 -1380 37660 -1260
rect 37780 -1380 37825 -1260
rect 37945 -1380 38000 -1260
rect 38120 -1380 38165 -1260
rect 38285 -1380 38330 -1260
rect 38450 -1380 38495 -1260
rect 38615 -1380 38670 -1260
rect 38790 -1380 38835 -1260
rect 38955 -1380 39000 -1260
rect 39120 -1380 39165 -1260
rect 39285 -1380 39340 -1260
rect 39460 -1380 39505 -1260
rect 39625 -1380 39670 -1260
rect 39790 -1380 39835 -1260
rect 39955 -1380 40010 -1260
rect 40130 -1380 40175 -1260
rect 40295 -1380 40340 -1260
rect 40460 -1380 40505 -1260
rect 40625 -1380 40680 -1260
rect 40800 -1380 40845 -1260
rect 40965 -1380 41010 -1260
rect 41130 -1380 41175 -1260
rect 41295 -1380 41350 -1260
rect 41470 -1380 41515 -1260
rect 41635 -1380 41680 -1260
rect 41800 -1380 41845 -1260
rect 41965 -1380 41975 -1260
rect 36475 -1425 41975 -1380
rect 36475 -1545 36485 -1425
rect 36605 -1545 36660 -1425
rect 36780 -1545 36825 -1425
rect 36945 -1545 36990 -1425
rect 37110 -1545 37155 -1425
rect 37275 -1545 37330 -1425
rect 37450 -1545 37495 -1425
rect 37615 -1545 37660 -1425
rect 37780 -1545 37825 -1425
rect 37945 -1545 38000 -1425
rect 38120 -1545 38165 -1425
rect 38285 -1545 38330 -1425
rect 38450 -1545 38495 -1425
rect 38615 -1545 38670 -1425
rect 38790 -1545 38835 -1425
rect 38955 -1545 39000 -1425
rect 39120 -1545 39165 -1425
rect 39285 -1545 39340 -1425
rect 39460 -1545 39505 -1425
rect 39625 -1545 39670 -1425
rect 39790 -1545 39835 -1425
rect 39955 -1545 40010 -1425
rect 40130 -1545 40175 -1425
rect 40295 -1545 40340 -1425
rect 40460 -1545 40505 -1425
rect 40625 -1545 40680 -1425
rect 40800 -1545 40845 -1425
rect 40965 -1545 41010 -1425
rect 41130 -1545 41175 -1425
rect 41295 -1545 41350 -1425
rect 41470 -1545 41515 -1425
rect 41635 -1545 41680 -1425
rect 41800 -1545 41845 -1425
rect 41965 -1545 41975 -1425
rect 36475 -1590 41975 -1545
rect 36475 -1710 36485 -1590
rect 36605 -1710 36660 -1590
rect 36780 -1710 36825 -1590
rect 36945 -1710 36990 -1590
rect 37110 -1710 37155 -1590
rect 37275 -1710 37330 -1590
rect 37450 -1710 37495 -1590
rect 37615 -1710 37660 -1590
rect 37780 -1710 37825 -1590
rect 37945 -1710 38000 -1590
rect 38120 -1710 38165 -1590
rect 38285 -1710 38330 -1590
rect 38450 -1710 38495 -1590
rect 38615 -1710 38670 -1590
rect 38790 -1710 38835 -1590
rect 38955 -1710 39000 -1590
rect 39120 -1710 39165 -1590
rect 39285 -1710 39340 -1590
rect 39460 -1710 39505 -1590
rect 39625 -1710 39670 -1590
rect 39790 -1710 39835 -1590
rect 39955 -1710 40010 -1590
rect 40130 -1710 40175 -1590
rect 40295 -1710 40340 -1590
rect 40460 -1710 40505 -1590
rect 40625 -1710 40680 -1590
rect 40800 -1710 40845 -1590
rect 40965 -1710 41010 -1590
rect 41130 -1710 41175 -1590
rect 41295 -1710 41350 -1590
rect 41470 -1710 41515 -1590
rect 41635 -1710 41680 -1590
rect 41800 -1710 41845 -1590
rect 41965 -1710 41975 -1590
rect 36475 -1755 41975 -1710
rect 36475 -1875 36485 -1755
rect 36605 -1875 36660 -1755
rect 36780 -1875 36825 -1755
rect 36945 -1875 36990 -1755
rect 37110 -1875 37155 -1755
rect 37275 -1875 37330 -1755
rect 37450 -1875 37495 -1755
rect 37615 -1875 37660 -1755
rect 37780 -1875 37825 -1755
rect 37945 -1875 38000 -1755
rect 38120 -1875 38165 -1755
rect 38285 -1875 38330 -1755
rect 38450 -1875 38495 -1755
rect 38615 -1875 38670 -1755
rect 38790 -1875 38835 -1755
rect 38955 -1875 39000 -1755
rect 39120 -1875 39165 -1755
rect 39285 -1875 39340 -1755
rect 39460 -1875 39505 -1755
rect 39625 -1875 39670 -1755
rect 39790 -1875 39835 -1755
rect 39955 -1875 40010 -1755
rect 40130 -1875 40175 -1755
rect 40295 -1875 40340 -1755
rect 40460 -1875 40505 -1755
rect 40625 -1875 40680 -1755
rect 40800 -1875 40845 -1755
rect 40965 -1875 41010 -1755
rect 41130 -1875 41175 -1755
rect 41295 -1875 41350 -1755
rect 41470 -1875 41515 -1755
rect 41635 -1875 41680 -1755
rect 41800 -1875 41845 -1755
rect 41965 -1875 41975 -1755
rect 36475 -1930 41975 -1875
rect 36475 -2050 36485 -1930
rect 36605 -2050 36660 -1930
rect 36780 -2050 36825 -1930
rect 36945 -2050 36990 -1930
rect 37110 -2050 37155 -1930
rect 37275 -2050 37330 -1930
rect 37450 -2050 37495 -1930
rect 37615 -2050 37660 -1930
rect 37780 -2050 37825 -1930
rect 37945 -2050 38000 -1930
rect 38120 -2050 38165 -1930
rect 38285 -2050 38330 -1930
rect 38450 -2050 38495 -1930
rect 38615 -2050 38670 -1930
rect 38790 -2050 38835 -1930
rect 38955 -2050 39000 -1930
rect 39120 -2050 39165 -1930
rect 39285 -2050 39340 -1930
rect 39460 -2050 39505 -1930
rect 39625 -2050 39670 -1930
rect 39790 -2050 39835 -1930
rect 39955 -2050 40010 -1930
rect 40130 -2050 40175 -1930
rect 40295 -2050 40340 -1930
rect 40460 -2050 40505 -1930
rect 40625 -2050 40680 -1930
rect 40800 -2050 40845 -1930
rect 40965 -2050 41010 -1930
rect 41130 -2050 41175 -1930
rect 41295 -2050 41350 -1930
rect 41470 -2050 41515 -1930
rect 41635 -2050 41680 -1930
rect 41800 -2050 41845 -1930
rect 41965 -2050 41975 -1930
rect 36475 -2095 41975 -2050
rect 36475 -2215 36485 -2095
rect 36605 -2215 36660 -2095
rect 36780 -2215 36825 -2095
rect 36945 -2215 36990 -2095
rect 37110 -2215 37155 -2095
rect 37275 -2215 37330 -2095
rect 37450 -2215 37495 -2095
rect 37615 -2215 37660 -2095
rect 37780 -2215 37825 -2095
rect 37945 -2215 38000 -2095
rect 38120 -2215 38165 -2095
rect 38285 -2215 38330 -2095
rect 38450 -2215 38495 -2095
rect 38615 -2215 38670 -2095
rect 38790 -2215 38835 -2095
rect 38955 -2215 39000 -2095
rect 39120 -2215 39165 -2095
rect 39285 -2215 39340 -2095
rect 39460 -2215 39505 -2095
rect 39625 -2215 39670 -2095
rect 39790 -2215 39835 -2095
rect 39955 -2215 40010 -2095
rect 40130 -2215 40175 -2095
rect 40295 -2215 40340 -2095
rect 40460 -2215 40505 -2095
rect 40625 -2215 40680 -2095
rect 40800 -2215 40845 -2095
rect 40965 -2215 41010 -2095
rect 41130 -2215 41175 -2095
rect 41295 -2215 41350 -2095
rect 41470 -2215 41515 -2095
rect 41635 -2215 41680 -2095
rect 41800 -2215 41845 -2095
rect 41965 -2215 41975 -2095
rect 36475 -2260 41975 -2215
rect 36475 -2380 36485 -2260
rect 36605 -2380 36660 -2260
rect 36780 -2380 36825 -2260
rect 36945 -2380 36990 -2260
rect 37110 -2380 37155 -2260
rect 37275 -2380 37330 -2260
rect 37450 -2380 37495 -2260
rect 37615 -2380 37660 -2260
rect 37780 -2380 37825 -2260
rect 37945 -2380 38000 -2260
rect 38120 -2380 38165 -2260
rect 38285 -2380 38330 -2260
rect 38450 -2380 38495 -2260
rect 38615 -2380 38670 -2260
rect 38790 -2380 38835 -2260
rect 38955 -2380 39000 -2260
rect 39120 -2380 39165 -2260
rect 39285 -2380 39340 -2260
rect 39460 -2380 39505 -2260
rect 39625 -2380 39670 -2260
rect 39790 -2380 39835 -2260
rect 39955 -2380 40010 -2260
rect 40130 -2380 40175 -2260
rect 40295 -2380 40340 -2260
rect 40460 -2380 40505 -2260
rect 40625 -2380 40680 -2260
rect 40800 -2380 40845 -2260
rect 40965 -2380 41010 -2260
rect 41130 -2380 41175 -2260
rect 41295 -2380 41350 -2260
rect 41470 -2380 41515 -2260
rect 41635 -2380 41680 -2260
rect 41800 -2380 41845 -2260
rect 41965 -2380 41975 -2260
rect 36475 -2425 41975 -2380
rect 36475 -2545 36485 -2425
rect 36605 -2545 36660 -2425
rect 36780 -2545 36825 -2425
rect 36945 -2545 36990 -2425
rect 37110 -2545 37155 -2425
rect 37275 -2545 37330 -2425
rect 37450 -2545 37495 -2425
rect 37615 -2545 37660 -2425
rect 37780 -2545 37825 -2425
rect 37945 -2545 38000 -2425
rect 38120 -2545 38165 -2425
rect 38285 -2545 38330 -2425
rect 38450 -2545 38495 -2425
rect 38615 -2545 38670 -2425
rect 38790 -2545 38835 -2425
rect 38955 -2545 39000 -2425
rect 39120 -2545 39165 -2425
rect 39285 -2545 39340 -2425
rect 39460 -2545 39505 -2425
rect 39625 -2545 39670 -2425
rect 39790 -2545 39835 -2425
rect 39955 -2545 40010 -2425
rect 40130 -2545 40175 -2425
rect 40295 -2545 40340 -2425
rect 40460 -2545 40505 -2425
rect 40625 -2545 40680 -2425
rect 40800 -2545 40845 -2425
rect 40965 -2545 41010 -2425
rect 41130 -2545 41175 -2425
rect 41295 -2545 41350 -2425
rect 41470 -2545 41515 -2425
rect 41635 -2545 41680 -2425
rect 41800 -2545 41845 -2425
rect 41965 -2545 41975 -2425
rect 36475 -2600 41975 -2545
rect 36475 -2720 36485 -2600
rect 36605 -2720 36660 -2600
rect 36780 -2720 36825 -2600
rect 36945 -2720 36990 -2600
rect 37110 -2720 37155 -2600
rect 37275 -2720 37330 -2600
rect 37450 -2720 37495 -2600
rect 37615 -2720 37660 -2600
rect 37780 -2720 37825 -2600
rect 37945 -2720 38000 -2600
rect 38120 -2720 38165 -2600
rect 38285 -2720 38330 -2600
rect 38450 -2720 38495 -2600
rect 38615 -2720 38670 -2600
rect 38790 -2720 38835 -2600
rect 38955 -2720 39000 -2600
rect 39120 -2720 39165 -2600
rect 39285 -2720 39340 -2600
rect 39460 -2720 39505 -2600
rect 39625 -2720 39670 -2600
rect 39790 -2720 39835 -2600
rect 39955 -2720 40010 -2600
rect 40130 -2720 40175 -2600
rect 40295 -2720 40340 -2600
rect 40460 -2720 40505 -2600
rect 40625 -2720 40680 -2600
rect 40800 -2720 40845 -2600
rect 40965 -2720 41010 -2600
rect 41130 -2720 41175 -2600
rect 41295 -2720 41350 -2600
rect 41470 -2720 41515 -2600
rect 41635 -2720 41680 -2600
rect 41800 -2720 41845 -2600
rect 41965 -2720 41975 -2600
rect 36475 -2765 41975 -2720
rect 36475 -2885 36485 -2765
rect 36605 -2885 36660 -2765
rect 36780 -2885 36825 -2765
rect 36945 -2885 36990 -2765
rect 37110 -2885 37155 -2765
rect 37275 -2885 37330 -2765
rect 37450 -2885 37495 -2765
rect 37615 -2885 37660 -2765
rect 37780 -2885 37825 -2765
rect 37945 -2885 38000 -2765
rect 38120 -2885 38165 -2765
rect 38285 -2885 38330 -2765
rect 38450 -2885 38495 -2765
rect 38615 -2885 38670 -2765
rect 38790 -2885 38835 -2765
rect 38955 -2885 39000 -2765
rect 39120 -2885 39165 -2765
rect 39285 -2885 39340 -2765
rect 39460 -2885 39505 -2765
rect 39625 -2885 39670 -2765
rect 39790 -2885 39835 -2765
rect 39955 -2885 40010 -2765
rect 40130 -2885 40175 -2765
rect 40295 -2885 40340 -2765
rect 40460 -2885 40505 -2765
rect 40625 -2885 40680 -2765
rect 40800 -2885 40845 -2765
rect 40965 -2885 41010 -2765
rect 41130 -2885 41175 -2765
rect 41295 -2885 41350 -2765
rect 41470 -2885 41515 -2765
rect 41635 -2885 41680 -2765
rect 41800 -2885 41845 -2765
rect 41965 -2885 41975 -2765
rect 36475 -2930 41975 -2885
rect 36475 -3050 36485 -2930
rect 36605 -3050 36660 -2930
rect 36780 -3050 36825 -2930
rect 36945 -3050 36990 -2930
rect 37110 -3050 37155 -2930
rect 37275 -3050 37330 -2930
rect 37450 -3050 37495 -2930
rect 37615 -3050 37660 -2930
rect 37780 -3050 37825 -2930
rect 37945 -3050 38000 -2930
rect 38120 -3050 38165 -2930
rect 38285 -3050 38330 -2930
rect 38450 -3050 38495 -2930
rect 38615 -3050 38670 -2930
rect 38790 -3050 38835 -2930
rect 38955 -3050 39000 -2930
rect 39120 -3050 39165 -2930
rect 39285 -3050 39340 -2930
rect 39460 -3050 39505 -2930
rect 39625 -3050 39670 -2930
rect 39790 -3050 39835 -2930
rect 39955 -3050 40010 -2930
rect 40130 -3050 40175 -2930
rect 40295 -3050 40340 -2930
rect 40460 -3050 40505 -2930
rect 40625 -3050 40680 -2930
rect 40800 -3050 40845 -2930
rect 40965 -3050 41010 -2930
rect 41130 -3050 41175 -2930
rect 41295 -3050 41350 -2930
rect 41470 -3050 41515 -2930
rect 41635 -3050 41680 -2930
rect 41800 -3050 41845 -2930
rect 41965 -3050 41975 -2930
rect 36475 -3095 41975 -3050
rect 36475 -3215 36485 -3095
rect 36605 -3215 36660 -3095
rect 36780 -3215 36825 -3095
rect 36945 -3215 36990 -3095
rect 37110 -3215 37155 -3095
rect 37275 -3215 37330 -3095
rect 37450 -3215 37495 -3095
rect 37615 -3215 37660 -3095
rect 37780 -3215 37825 -3095
rect 37945 -3215 38000 -3095
rect 38120 -3215 38165 -3095
rect 38285 -3215 38330 -3095
rect 38450 -3215 38495 -3095
rect 38615 -3215 38670 -3095
rect 38790 -3215 38835 -3095
rect 38955 -3215 39000 -3095
rect 39120 -3215 39165 -3095
rect 39285 -3215 39340 -3095
rect 39460 -3215 39505 -3095
rect 39625 -3215 39670 -3095
rect 39790 -3215 39835 -3095
rect 39955 -3215 40010 -3095
rect 40130 -3215 40175 -3095
rect 40295 -3215 40340 -3095
rect 40460 -3215 40505 -3095
rect 40625 -3215 40680 -3095
rect 40800 -3215 40845 -3095
rect 40965 -3215 41010 -3095
rect 41130 -3215 41175 -3095
rect 41295 -3215 41350 -3095
rect 41470 -3215 41515 -3095
rect 41635 -3215 41680 -3095
rect 41800 -3215 41845 -3095
rect 41965 -3215 41975 -3095
rect 36475 -3270 41975 -3215
rect 36475 -3390 36485 -3270
rect 36605 -3390 36660 -3270
rect 36780 -3390 36825 -3270
rect 36945 -3390 36990 -3270
rect 37110 -3390 37155 -3270
rect 37275 -3390 37330 -3270
rect 37450 -3390 37495 -3270
rect 37615 -3390 37660 -3270
rect 37780 -3390 37825 -3270
rect 37945 -3390 38000 -3270
rect 38120 -3390 38165 -3270
rect 38285 -3390 38330 -3270
rect 38450 -3390 38495 -3270
rect 38615 -3390 38670 -3270
rect 38790 -3390 38835 -3270
rect 38955 -3390 39000 -3270
rect 39120 -3390 39165 -3270
rect 39285 -3390 39340 -3270
rect 39460 -3390 39505 -3270
rect 39625 -3390 39670 -3270
rect 39790 -3390 39835 -3270
rect 39955 -3390 40010 -3270
rect 40130 -3390 40175 -3270
rect 40295 -3390 40340 -3270
rect 40460 -3390 40505 -3270
rect 40625 -3390 40680 -3270
rect 40800 -3390 40845 -3270
rect 40965 -3390 41010 -3270
rect 41130 -3390 41175 -3270
rect 41295 -3390 41350 -3270
rect 41470 -3390 41515 -3270
rect 41635 -3390 41680 -3270
rect 41800 -3390 41845 -3270
rect 41965 -3390 41975 -3270
rect 36475 -3435 41975 -3390
rect 36475 -3555 36485 -3435
rect 36605 -3555 36660 -3435
rect 36780 -3555 36825 -3435
rect 36945 -3555 36990 -3435
rect 37110 -3555 37155 -3435
rect 37275 -3555 37330 -3435
rect 37450 -3555 37495 -3435
rect 37615 -3555 37660 -3435
rect 37780 -3555 37825 -3435
rect 37945 -3555 38000 -3435
rect 38120 -3555 38165 -3435
rect 38285 -3555 38330 -3435
rect 38450 -3555 38495 -3435
rect 38615 -3555 38670 -3435
rect 38790 -3555 38835 -3435
rect 38955 -3555 39000 -3435
rect 39120 -3555 39165 -3435
rect 39285 -3555 39340 -3435
rect 39460 -3555 39505 -3435
rect 39625 -3555 39670 -3435
rect 39790 -3555 39835 -3435
rect 39955 -3555 40010 -3435
rect 40130 -3555 40175 -3435
rect 40295 -3555 40340 -3435
rect 40460 -3555 40505 -3435
rect 40625 -3555 40680 -3435
rect 40800 -3555 40845 -3435
rect 40965 -3555 41010 -3435
rect 41130 -3555 41175 -3435
rect 41295 -3555 41350 -3435
rect 41470 -3555 41515 -3435
rect 41635 -3555 41680 -3435
rect 41800 -3555 41845 -3435
rect 41965 -3555 41975 -3435
rect 36475 -3600 41975 -3555
rect 36475 -3720 36485 -3600
rect 36605 -3720 36660 -3600
rect 36780 -3720 36825 -3600
rect 36945 -3720 36990 -3600
rect 37110 -3720 37155 -3600
rect 37275 -3720 37330 -3600
rect 37450 -3720 37495 -3600
rect 37615 -3720 37660 -3600
rect 37780 -3720 37825 -3600
rect 37945 -3720 38000 -3600
rect 38120 -3720 38165 -3600
rect 38285 -3720 38330 -3600
rect 38450 -3720 38495 -3600
rect 38615 -3720 38670 -3600
rect 38790 -3720 38835 -3600
rect 38955 -3720 39000 -3600
rect 39120 -3720 39165 -3600
rect 39285 -3720 39340 -3600
rect 39460 -3720 39505 -3600
rect 39625 -3720 39670 -3600
rect 39790 -3720 39835 -3600
rect 39955 -3720 40010 -3600
rect 40130 -3720 40175 -3600
rect 40295 -3720 40340 -3600
rect 40460 -3720 40505 -3600
rect 40625 -3720 40680 -3600
rect 40800 -3720 40845 -3600
rect 40965 -3720 41010 -3600
rect 41130 -3720 41175 -3600
rect 41295 -3720 41350 -3600
rect 41470 -3720 41515 -3600
rect 41635 -3720 41680 -3600
rect 41800 -3720 41845 -3600
rect 41965 -3720 41975 -3600
rect 36475 -3765 41975 -3720
rect 36475 -3885 36485 -3765
rect 36605 -3885 36660 -3765
rect 36780 -3885 36825 -3765
rect 36945 -3885 36990 -3765
rect 37110 -3885 37155 -3765
rect 37275 -3885 37330 -3765
rect 37450 -3885 37495 -3765
rect 37615 -3885 37660 -3765
rect 37780 -3885 37825 -3765
rect 37945 -3885 38000 -3765
rect 38120 -3885 38165 -3765
rect 38285 -3885 38330 -3765
rect 38450 -3885 38495 -3765
rect 38615 -3885 38670 -3765
rect 38790 -3885 38835 -3765
rect 38955 -3885 39000 -3765
rect 39120 -3885 39165 -3765
rect 39285 -3885 39340 -3765
rect 39460 -3885 39505 -3765
rect 39625 -3885 39670 -3765
rect 39790 -3885 39835 -3765
rect 39955 -3885 40010 -3765
rect 40130 -3885 40175 -3765
rect 40295 -3885 40340 -3765
rect 40460 -3885 40505 -3765
rect 40625 -3885 40680 -3765
rect 40800 -3885 40845 -3765
rect 40965 -3885 41010 -3765
rect 41130 -3885 41175 -3765
rect 41295 -3885 41350 -3765
rect 41470 -3885 41515 -3765
rect 41635 -3885 41680 -3765
rect 41800 -3885 41845 -3765
rect 41965 -3885 41975 -3765
rect 36475 -3940 41975 -3885
rect 36475 -4060 36485 -3940
rect 36605 -4060 36660 -3940
rect 36780 -4060 36825 -3940
rect 36945 -4060 36990 -3940
rect 37110 -4060 37155 -3940
rect 37275 -4060 37330 -3940
rect 37450 -4060 37495 -3940
rect 37615 -4060 37660 -3940
rect 37780 -4060 37825 -3940
rect 37945 -4060 38000 -3940
rect 38120 -4060 38165 -3940
rect 38285 -4060 38330 -3940
rect 38450 -4060 38495 -3940
rect 38615 -4060 38670 -3940
rect 38790 -4060 38835 -3940
rect 38955 -4060 39000 -3940
rect 39120 -4060 39165 -3940
rect 39285 -4060 39340 -3940
rect 39460 -4060 39505 -3940
rect 39625 -4060 39670 -3940
rect 39790 -4060 39835 -3940
rect 39955 -4060 40010 -3940
rect 40130 -4060 40175 -3940
rect 40295 -4060 40340 -3940
rect 40460 -4060 40505 -3940
rect 40625 -4060 40680 -3940
rect 40800 -4060 40845 -3940
rect 40965 -4060 41010 -3940
rect 41130 -4060 41175 -3940
rect 41295 -4060 41350 -3940
rect 41470 -4060 41515 -3940
rect 41635 -4060 41680 -3940
rect 41800 -4060 41845 -3940
rect 41965 -4060 41975 -3940
rect 36475 -4070 41975 -4060
rect 42165 1420 47665 1430
rect 42165 1300 42175 1420
rect 42295 1300 42350 1420
rect 42470 1300 42515 1420
rect 42635 1300 42680 1420
rect 42800 1300 42845 1420
rect 42965 1300 43020 1420
rect 43140 1300 43185 1420
rect 43305 1300 43350 1420
rect 43470 1300 43515 1420
rect 43635 1300 43690 1420
rect 43810 1300 43855 1420
rect 43975 1300 44020 1420
rect 44140 1300 44185 1420
rect 44305 1300 44360 1420
rect 44480 1300 44525 1420
rect 44645 1300 44690 1420
rect 44810 1300 44855 1420
rect 44975 1300 45030 1420
rect 45150 1300 45195 1420
rect 45315 1300 45360 1420
rect 45480 1300 45525 1420
rect 45645 1300 45700 1420
rect 45820 1300 45865 1420
rect 45985 1300 46030 1420
rect 46150 1300 46195 1420
rect 46315 1300 46370 1420
rect 46490 1300 46535 1420
rect 46655 1300 46700 1420
rect 46820 1300 46865 1420
rect 46985 1300 47040 1420
rect 47160 1300 47205 1420
rect 47325 1300 47370 1420
rect 47490 1300 47535 1420
rect 47655 1300 47665 1420
rect 42165 1255 47665 1300
rect 42165 1135 42175 1255
rect 42295 1135 42350 1255
rect 42470 1135 42515 1255
rect 42635 1135 42680 1255
rect 42800 1135 42845 1255
rect 42965 1135 43020 1255
rect 43140 1135 43185 1255
rect 43305 1135 43350 1255
rect 43470 1135 43515 1255
rect 43635 1135 43690 1255
rect 43810 1135 43855 1255
rect 43975 1135 44020 1255
rect 44140 1135 44185 1255
rect 44305 1135 44360 1255
rect 44480 1135 44525 1255
rect 44645 1135 44690 1255
rect 44810 1135 44855 1255
rect 44975 1135 45030 1255
rect 45150 1135 45195 1255
rect 45315 1135 45360 1255
rect 45480 1135 45525 1255
rect 45645 1135 45700 1255
rect 45820 1135 45865 1255
rect 45985 1135 46030 1255
rect 46150 1135 46195 1255
rect 46315 1135 46370 1255
rect 46490 1135 46535 1255
rect 46655 1135 46700 1255
rect 46820 1135 46865 1255
rect 46985 1135 47040 1255
rect 47160 1135 47205 1255
rect 47325 1135 47370 1255
rect 47490 1135 47535 1255
rect 47655 1135 47665 1255
rect 42165 1090 47665 1135
rect 42165 970 42175 1090
rect 42295 970 42350 1090
rect 42470 970 42515 1090
rect 42635 970 42680 1090
rect 42800 970 42845 1090
rect 42965 970 43020 1090
rect 43140 970 43185 1090
rect 43305 970 43350 1090
rect 43470 970 43515 1090
rect 43635 970 43690 1090
rect 43810 970 43855 1090
rect 43975 970 44020 1090
rect 44140 970 44185 1090
rect 44305 970 44360 1090
rect 44480 970 44525 1090
rect 44645 970 44690 1090
rect 44810 970 44855 1090
rect 44975 970 45030 1090
rect 45150 970 45195 1090
rect 45315 970 45360 1090
rect 45480 970 45525 1090
rect 45645 970 45700 1090
rect 45820 970 45865 1090
rect 45985 970 46030 1090
rect 46150 970 46195 1090
rect 46315 970 46370 1090
rect 46490 970 46535 1090
rect 46655 970 46700 1090
rect 46820 970 46865 1090
rect 46985 970 47040 1090
rect 47160 970 47205 1090
rect 47325 970 47370 1090
rect 47490 970 47535 1090
rect 47655 970 47665 1090
rect 42165 925 47665 970
rect 42165 805 42175 925
rect 42295 805 42350 925
rect 42470 805 42515 925
rect 42635 805 42680 925
rect 42800 805 42845 925
rect 42965 805 43020 925
rect 43140 805 43185 925
rect 43305 805 43350 925
rect 43470 805 43515 925
rect 43635 805 43690 925
rect 43810 805 43855 925
rect 43975 805 44020 925
rect 44140 805 44185 925
rect 44305 805 44360 925
rect 44480 805 44525 925
rect 44645 805 44690 925
rect 44810 805 44855 925
rect 44975 805 45030 925
rect 45150 805 45195 925
rect 45315 805 45360 925
rect 45480 805 45525 925
rect 45645 805 45700 925
rect 45820 805 45865 925
rect 45985 805 46030 925
rect 46150 805 46195 925
rect 46315 805 46370 925
rect 46490 805 46535 925
rect 46655 805 46700 925
rect 46820 805 46865 925
rect 46985 805 47040 925
rect 47160 805 47205 925
rect 47325 805 47370 925
rect 47490 805 47535 925
rect 47655 805 47665 925
rect 42165 750 47665 805
rect 42165 630 42175 750
rect 42295 630 42350 750
rect 42470 630 42515 750
rect 42635 630 42680 750
rect 42800 630 42845 750
rect 42965 630 43020 750
rect 43140 630 43185 750
rect 43305 630 43350 750
rect 43470 630 43515 750
rect 43635 630 43690 750
rect 43810 630 43855 750
rect 43975 630 44020 750
rect 44140 630 44185 750
rect 44305 630 44360 750
rect 44480 630 44525 750
rect 44645 630 44690 750
rect 44810 630 44855 750
rect 44975 630 45030 750
rect 45150 630 45195 750
rect 45315 630 45360 750
rect 45480 630 45525 750
rect 45645 630 45700 750
rect 45820 630 45865 750
rect 45985 630 46030 750
rect 46150 630 46195 750
rect 46315 630 46370 750
rect 46490 630 46535 750
rect 46655 630 46700 750
rect 46820 630 46865 750
rect 46985 630 47040 750
rect 47160 630 47205 750
rect 47325 630 47370 750
rect 47490 630 47535 750
rect 47655 630 47665 750
rect 42165 585 47665 630
rect 42165 465 42175 585
rect 42295 465 42350 585
rect 42470 465 42515 585
rect 42635 465 42680 585
rect 42800 465 42845 585
rect 42965 465 43020 585
rect 43140 465 43185 585
rect 43305 465 43350 585
rect 43470 465 43515 585
rect 43635 465 43690 585
rect 43810 465 43855 585
rect 43975 465 44020 585
rect 44140 465 44185 585
rect 44305 465 44360 585
rect 44480 465 44525 585
rect 44645 465 44690 585
rect 44810 465 44855 585
rect 44975 465 45030 585
rect 45150 465 45195 585
rect 45315 465 45360 585
rect 45480 465 45525 585
rect 45645 465 45700 585
rect 45820 465 45865 585
rect 45985 465 46030 585
rect 46150 465 46195 585
rect 46315 465 46370 585
rect 46490 465 46535 585
rect 46655 465 46700 585
rect 46820 465 46865 585
rect 46985 465 47040 585
rect 47160 465 47205 585
rect 47325 465 47370 585
rect 47490 465 47535 585
rect 47655 465 47665 585
rect 42165 420 47665 465
rect 42165 300 42175 420
rect 42295 300 42350 420
rect 42470 300 42515 420
rect 42635 300 42680 420
rect 42800 300 42845 420
rect 42965 300 43020 420
rect 43140 300 43185 420
rect 43305 300 43350 420
rect 43470 300 43515 420
rect 43635 300 43690 420
rect 43810 300 43855 420
rect 43975 300 44020 420
rect 44140 300 44185 420
rect 44305 300 44360 420
rect 44480 300 44525 420
rect 44645 300 44690 420
rect 44810 300 44855 420
rect 44975 300 45030 420
rect 45150 300 45195 420
rect 45315 300 45360 420
rect 45480 300 45525 420
rect 45645 300 45700 420
rect 45820 300 45865 420
rect 45985 300 46030 420
rect 46150 300 46195 420
rect 46315 300 46370 420
rect 46490 300 46535 420
rect 46655 300 46700 420
rect 46820 300 46865 420
rect 46985 300 47040 420
rect 47160 300 47205 420
rect 47325 300 47370 420
rect 47490 300 47535 420
rect 47655 300 47665 420
rect 42165 255 47665 300
rect 42165 135 42175 255
rect 42295 135 42350 255
rect 42470 135 42515 255
rect 42635 135 42680 255
rect 42800 135 42845 255
rect 42965 135 43020 255
rect 43140 135 43185 255
rect 43305 135 43350 255
rect 43470 135 43515 255
rect 43635 135 43690 255
rect 43810 135 43855 255
rect 43975 135 44020 255
rect 44140 135 44185 255
rect 44305 135 44360 255
rect 44480 135 44525 255
rect 44645 135 44690 255
rect 44810 135 44855 255
rect 44975 135 45030 255
rect 45150 135 45195 255
rect 45315 135 45360 255
rect 45480 135 45525 255
rect 45645 135 45700 255
rect 45820 135 45865 255
rect 45985 135 46030 255
rect 46150 135 46195 255
rect 46315 135 46370 255
rect 46490 135 46535 255
rect 46655 135 46700 255
rect 46820 135 46865 255
rect 46985 135 47040 255
rect 47160 135 47205 255
rect 47325 135 47370 255
rect 47490 135 47535 255
rect 47655 135 47665 255
rect 42165 80 47665 135
rect 42165 -40 42175 80
rect 42295 -40 42350 80
rect 42470 -40 42515 80
rect 42635 -40 42680 80
rect 42800 -40 42845 80
rect 42965 -40 43020 80
rect 43140 -40 43185 80
rect 43305 -40 43350 80
rect 43470 -40 43515 80
rect 43635 -40 43690 80
rect 43810 -40 43855 80
rect 43975 -40 44020 80
rect 44140 -40 44185 80
rect 44305 -40 44360 80
rect 44480 -40 44525 80
rect 44645 -40 44690 80
rect 44810 -40 44855 80
rect 44975 -40 45030 80
rect 45150 -40 45195 80
rect 45315 -40 45360 80
rect 45480 -40 45525 80
rect 45645 -40 45700 80
rect 45820 -40 45865 80
rect 45985 -40 46030 80
rect 46150 -40 46195 80
rect 46315 -40 46370 80
rect 46490 -40 46535 80
rect 46655 -40 46700 80
rect 46820 -40 46865 80
rect 46985 -40 47040 80
rect 47160 -40 47205 80
rect 47325 -40 47370 80
rect 47490 -40 47535 80
rect 47655 -40 47665 80
rect 42165 -85 47665 -40
rect 42165 -205 42175 -85
rect 42295 -205 42350 -85
rect 42470 -205 42515 -85
rect 42635 -205 42680 -85
rect 42800 -205 42845 -85
rect 42965 -205 43020 -85
rect 43140 -205 43185 -85
rect 43305 -205 43350 -85
rect 43470 -205 43515 -85
rect 43635 -205 43690 -85
rect 43810 -205 43855 -85
rect 43975 -205 44020 -85
rect 44140 -205 44185 -85
rect 44305 -205 44360 -85
rect 44480 -205 44525 -85
rect 44645 -205 44690 -85
rect 44810 -205 44855 -85
rect 44975 -205 45030 -85
rect 45150 -205 45195 -85
rect 45315 -205 45360 -85
rect 45480 -205 45525 -85
rect 45645 -205 45700 -85
rect 45820 -205 45865 -85
rect 45985 -205 46030 -85
rect 46150 -205 46195 -85
rect 46315 -205 46370 -85
rect 46490 -205 46535 -85
rect 46655 -205 46700 -85
rect 46820 -205 46865 -85
rect 46985 -205 47040 -85
rect 47160 -205 47205 -85
rect 47325 -205 47370 -85
rect 47490 -205 47535 -85
rect 47655 -205 47665 -85
rect 42165 -250 47665 -205
rect 42165 -370 42175 -250
rect 42295 -370 42350 -250
rect 42470 -370 42515 -250
rect 42635 -370 42680 -250
rect 42800 -370 42845 -250
rect 42965 -370 43020 -250
rect 43140 -370 43185 -250
rect 43305 -370 43350 -250
rect 43470 -370 43515 -250
rect 43635 -370 43690 -250
rect 43810 -370 43855 -250
rect 43975 -370 44020 -250
rect 44140 -370 44185 -250
rect 44305 -370 44360 -250
rect 44480 -370 44525 -250
rect 44645 -370 44690 -250
rect 44810 -370 44855 -250
rect 44975 -370 45030 -250
rect 45150 -370 45195 -250
rect 45315 -370 45360 -250
rect 45480 -370 45525 -250
rect 45645 -370 45700 -250
rect 45820 -370 45865 -250
rect 45985 -370 46030 -250
rect 46150 -370 46195 -250
rect 46315 -370 46370 -250
rect 46490 -370 46535 -250
rect 46655 -370 46700 -250
rect 46820 -370 46865 -250
rect 46985 -370 47040 -250
rect 47160 -370 47205 -250
rect 47325 -370 47370 -250
rect 47490 -370 47535 -250
rect 47655 -370 47665 -250
rect 42165 -415 47665 -370
rect 42165 -535 42175 -415
rect 42295 -535 42350 -415
rect 42470 -535 42515 -415
rect 42635 -535 42680 -415
rect 42800 -535 42845 -415
rect 42965 -535 43020 -415
rect 43140 -535 43185 -415
rect 43305 -535 43350 -415
rect 43470 -535 43515 -415
rect 43635 -535 43690 -415
rect 43810 -535 43855 -415
rect 43975 -535 44020 -415
rect 44140 -535 44185 -415
rect 44305 -535 44360 -415
rect 44480 -535 44525 -415
rect 44645 -535 44690 -415
rect 44810 -535 44855 -415
rect 44975 -535 45030 -415
rect 45150 -535 45195 -415
rect 45315 -535 45360 -415
rect 45480 -535 45525 -415
rect 45645 -535 45700 -415
rect 45820 -535 45865 -415
rect 45985 -535 46030 -415
rect 46150 -535 46195 -415
rect 46315 -535 46370 -415
rect 46490 -535 46535 -415
rect 46655 -535 46700 -415
rect 46820 -535 46865 -415
rect 46985 -535 47040 -415
rect 47160 -535 47205 -415
rect 47325 -535 47370 -415
rect 47490 -535 47535 -415
rect 47655 -535 47665 -415
rect 42165 -590 47665 -535
rect 42165 -710 42175 -590
rect 42295 -710 42350 -590
rect 42470 -710 42515 -590
rect 42635 -710 42680 -590
rect 42800 -710 42845 -590
rect 42965 -710 43020 -590
rect 43140 -710 43185 -590
rect 43305 -710 43350 -590
rect 43470 -710 43515 -590
rect 43635 -710 43690 -590
rect 43810 -710 43855 -590
rect 43975 -710 44020 -590
rect 44140 -710 44185 -590
rect 44305 -710 44360 -590
rect 44480 -710 44525 -590
rect 44645 -710 44690 -590
rect 44810 -710 44855 -590
rect 44975 -710 45030 -590
rect 45150 -710 45195 -590
rect 45315 -710 45360 -590
rect 45480 -710 45525 -590
rect 45645 -710 45700 -590
rect 45820 -710 45865 -590
rect 45985 -710 46030 -590
rect 46150 -710 46195 -590
rect 46315 -710 46370 -590
rect 46490 -710 46535 -590
rect 46655 -710 46700 -590
rect 46820 -710 46865 -590
rect 46985 -710 47040 -590
rect 47160 -710 47205 -590
rect 47325 -710 47370 -590
rect 47490 -710 47535 -590
rect 47655 -710 47665 -590
rect 42165 -755 47665 -710
rect 42165 -875 42175 -755
rect 42295 -875 42350 -755
rect 42470 -875 42515 -755
rect 42635 -875 42680 -755
rect 42800 -875 42845 -755
rect 42965 -875 43020 -755
rect 43140 -875 43185 -755
rect 43305 -875 43350 -755
rect 43470 -875 43515 -755
rect 43635 -875 43690 -755
rect 43810 -875 43855 -755
rect 43975 -875 44020 -755
rect 44140 -875 44185 -755
rect 44305 -875 44360 -755
rect 44480 -875 44525 -755
rect 44645 -875 44690 -755
rect 44810 -875 44855 -755
rect 44975 -875 45030 -755
rect 45150 -875 45195 -755
rect 45315 -875 45360 -755
rect 45480 -875 45525 -755
rect 45645 -875 45700 -755
rect 45820 -875 45865 -755
rect 45985 -875 46030 -755
rect 46150 -875 46195 -755
rect 46315 -875 46370 -755
rect 46490 -875 46535 -755
rect 46655 -875 46700 -755
rect 46820 -875 46865 -755
rect 46985 -875 47040 -755
rect 47160 -875 47205 -755
rect 47325 -875 47370 -755
rect 47490 -875 47535 -755
rect 47655 -875 47665 -755
rect 42165 -920 47665 -875
rect 42165 -1040 42175 -920
rect 42295 -1040 42350 -920
rect 42470 -1040 42515 -920
rect 42635 -1040 42680 -920
rect 42800 -1040 42845 -920
rect 42965 -1040 43020 -920
rect 43140 -1040 43185 -920
rect 43305 -1040 43350 -920
rect 43470 -1040 43515 -920
rect 43635 -1040 43690 -920
rect 43810 -1040 43855 -920
rect 43975 -1040 44020 -920
rect 44140 -1040 44185 -920
rect 44305 -1040 44360 -920
rect 44480 -1040 44525 -920
rect 44645 -1040 44690 -920
rect 44810 -1040 44855 -920
rect 44975 -1040 45030 -920
rect 45150 -1040 45195 -920
rect 45315 -1040 45360 -920
rect 45480 -1040 45525 -920
rect 45645 -1040 45700 -920
rect 45820 -1040 45865 -920
rect 45985 -1040 46030 -920
rect 46150 -1040 46195 -920
rect 46315 -1040 46370 -920
rect 46490 -1040 46535 -920
rect 46655 -1040 46700 -920
rect 46820 -1040 46865 -920
rect 46985 -1040 47040 -920
rect 47160 -1040 47205 -920
rect 47325 -1040 47370 -920
rect 47490 -1040 47535 -920
rect 47655 -1040 47665 -920
rect 42165 -1085 47665 -1040
rect 42165 -1205 42175 -1085
rect 42295 -1205 42350 -1085
rect 42470 -1205 42515 -1085
rect 42635 -1205 42680 -1085
rect 42800 -1205 42845 -1085
rect 42965 -1205 43020 -1085
rect 43140 -1205 43185 -1085
rect 43305 -1205 43350 -1085
rect 43470 -1205 43515 -1085
rect 43635 -1205 43690 -1085
rect 43810 -1205 43855 -1085
rect 43975 -1205 44020 -1085
rect 44140 -1205 44185 -1085
rect 44305 -1205 44360 -1085
rect 44480 -1205 44525 -1085
rect 44645 -1205 44690 -1085
rect 44810 -1205 44855 -1085
rect 44975 -1205 45030 -1085
rect 45150 -1205 45195 -1085
rect 45315 -1205 45360 -1085
rect 45480 -1205 45525 -1085
rect 45645 -1205 45700 -1085
rect 45820 -1205 45865 -1085
rect 45985 -1205 46030 -1085
rect 46150 -1205 46195 -1085
rect 46315 -1205 46370 -1085
rect 46490 -1205 46535 -1085
rect 46655 -1205 46700 -1085
rect 46820 -1205 46865 -1085
rect 46985 -1205 47040 -1085
rect 47160 -1205 47205 -1085
rect 47325 -1205 47370 -1085
rect 47490 -1205 47535 -1085
rect 47655 -1205 47665 -1085
rect 42165 -1260 47665 -1205
rect 42165 -1380 42175 -1260
rect 42295 -1380 42350 -1260
rect 42470 -1380 42515 -1260
rect 42635 -1380 42680 -1260
rect 42800 -1380 42845 -1260
rect 42965 -1380 43020 -1260
rect 43140 -1380 43185 -1260
rect 43305 -1380 43350 -1260
rect 43470 -1380 43515 -1260
rect 43635 -1380 43690 -1260
rect 43810 -1380 43855 -1260
rect 43975 -1380 44020 -1260
rect 44140 -1380 44185 -1260
rect 44305 -1380 44360 -1260
rect 44480 -1380 44525 -1260
rect 44645 -1380 44690 -1260
rect 44810 -1380 44855 -1260
rect 44975 -1380 45030 -1260
rect 45150 -1380 45195 -1260
rect 45315 -1380 45360 -1260
rect 45480 -1380 45525 -1260
rect 45645 -1380 45700 -1260
rect 45820 -1380 45865 -1260
rect 45985 -1380 46030 -1260
rect 46150 -1380 46195 -1260
rect 46315 -1380 46370 -1260
rect 46490 -1380 46535 -1260
rect 46655 -1380 46700 -1260
rect 46820 -1380 46865 -1260
rect 46985 -1380 47040 -1260
rect 47160 -1380 47205 -1260
rect 47325 -1380 47370 -1260
rect 47490 -1380 47535 -1260
rect 47655 -1380 47665 -1260
rect 42165 -1425 47665 -1380
rect 42165 -1545 42175 -1425
rect 42295 -1545 42350 -1425
rect 42470 -1545 42515 -1425
rect 42635 -1545 42680 -1425
rect 42800 -1545 42845 -1425
rect 42965 -1545 43020 -1425
rect 43140 -1545 43185 -1425
rect 43305 -1545 43350 -1425
rect 43470 -1545 43515 -1425
rect 43635 -1545 43690 -1425
rect 43810 -1545 43855 -1425
rect 43975 -1545 44020 -1425
rect 44140 -1545 44185 -1425
rect 44305 -1545 44360 -1425
rect 44480 -1545 44525 -1425
rect 44645 -1545 44690 -1425
rect 44810 -1545 44855 -1425
rect 44975 -1545 45030 -1425
rect 45150 -1545 45195 -1425
rect 45315 -1545 45360 -1425
rect 45480 -1545 45525 -1425
rect 45645 -1545 45700 -1425
rect 45820 -1545 45865 -1425
rect 45985 -1545 46030 -1425
rect 46150 -1545 46195 -1425
rect 46315 -1545 46370 -1425
rect 46490 -1545 46535 -1425
rect 46655 -1545 46700 -1425
rect 46820 -1545 46865 -1425
rect 46985 -1545 47040 -1425
rect 47160 -1545 47205 -1425
rect 47325 -1545 47370 -1425
rect 47490 -1545 47535 -1425
rect 47655 -1545 47665 -1425
rect 42165 -1590 47665 -1545
rect 42165 -1710 42175 -1590
rect 42295 -1710 42350 -1590
rect 42470 -1710 42515 -1590
rect 42635 -1710 42680 -1590
rect 42800 -1710 42845 -1590
rect 42965 -1710 43020 -1590
rect 43140 -1710 43185 -1590
rect 43305 -1710 43350 -1590
rect 43470 -1710 43515 -1590
rect 43635 -1710 43690 -1590
rect 43810 -1710 43855 -1590
rect 43975 -1710 44020 -1590
rect 44140 -1710 44185 -1590
rect 44305 -1710 44360 -1590
rect 44480 -1710 44525 -1590
rect 44645 -1710 44690 -1590
rect 44810 -1710 44855 -1590
rect 44975 -1710 45030 -1590
rect 45150 -1710 45195 -1590
rect 45315 -1710 45360 -1590
rect 45480 -1710 45525 -1590
rect 45645 -1710 45700 -1590
rect 45820 -1710 45865 -1590
rect 45985 -1710 46030 -1590
rect 46150 -1710 46195 -1590
rect 46315 -1710 46370 -1590
rect 46490 -1710 46535 -1590
rect 46655 -1710 46700 -1590
rect 46820 -1710 46865 -1590
rect 46985 -1710 47040 -1590
rect 47160 -1710 47205 -1590
rect 47325 -1710 47370 -1590
rect 47490 -1710 47535 -1590
rect 47655 -1710 47665 -1590
rect 42165 -1755 47665 -1710
rect 42165 -1875 42175 -1755
rect 42295 -1875 42350 -1755
rect 42470 -1875 42515 -1755
rect 42635 -1875 42680 -1755
rect 42800 -1875 42845 -1755
rect 42965 -1875 43020 -1755
rect 43140 -1875 43185 -1755
rect 43305 -1875 43350 -1755
rect 43470 -1875 43515 -1755
rect 43635 -1875 43690 -1755
rect 43810 -1875 43855 -1755
rect 43975 -1875 44020 -1755
rect 44140 -1875 44185 -1755
rect 44305 -1875 44360 -1755
rect 44480 -1875 44525 -1755
rect 44645 -1875 44690 -1755
rect 44810 -1875 44855 -1755
rect 44975 -1875 45030 -1755
rect 45150 -1875 45195 -1755
rect 45315 -1875 45360 -1755
rect 45480 -1875 45525 -1755
rect 45645 -1875 45700 -1755
rect 45820 -1875 45865 -1755
rect 45985 -1875 46030 -1755
rect 46150 -1875 46195 -1755
rect 46315 -1875 46370 -1755
rect 46490 -1875 46535 -1755
rect 46655 -1875 46700 -1755
rect 46820 -1875 46865 -1755
rect 46985 -1875 47040 -1755
rect 47160 -1875 47205 -1755
rect 47325 -1875 47370 -1755
rect 47490 -1875 47535 -1755
rect 47655 -1875 47665 -1755
rect 42165 -1930 47665 -1875
rect 42165 -2050 42175 -1930
rect 42295 -2050 42350 -1930
rect 42470 -2050 42515 -1930
rect 42635 -2050 42680 -1930
rect 42800 -2050 42845 -1930
rect 42965 -2050 43020 -1930
rect 43140 -2050 43185 -1930
rect 43305 -2050 43350 -1930
rect 43470 -2050 43515 -1930
rect 43635 -2050 43690 -1930
rect 43810 -2050 43855 -1930
rect 43975 -2050 44020 -1930
rect 44140 -2050 44185 -1930
rect 44305 -2050 44360 -1930
rect 44480 -2050 44525 -1930
rect 44645 -2050 44690 -1930
rect 44810 -2050 44855 -1930
rect 44975 -2050 45030 -1930
rect 45150 -2050 45195 -1930
rect 45315 -2050 45360 -1930
rect 45480 -2050 45525 -1930
rect 45645 -2050 45700 -1930
rect 45820 -2050 45865 -1930
rect 45985 -2050 46030 -1930
rect 46150 -2050 46195 -1930
rect 46315 -2050 46370 -1930
rect 46490 -2050 46535 -1930
rect 46655 -2050 46700 -1930
rect 46820 -2050 46865 -1930
rect 46985 -2050 47040 -1930
rect 47160 -2050 47205 -1930
rect 47325 -2050 47370 -1930
rect 47490 -2050 47535 -1930
rect 47655 -2050 47665 -1930
rect 42165 -2095 47665 -2050
rect 42165 -2215 42175 -2095
rect 42295 -2215 42350 -2095
rect 42470 -2215 42515 -2095
rect 42635 -2215 42680 -2095
rect 42800 -2215 42845 -2095
rect 42965 -2215 43020 -2095
rect 43140 -2215 43185 -2095
rect 43305 -2215 43350 -2095
rect 43470 -2215 43515 -2095
rect 43635 -2215 43690 -2095
rect 43810 -2215 43855 -2095
rect 43975 -2215 44020 -2095
rect 44140 -2215 44185 -2095
rect 44305 -2215 44360 -2095
rect 44480 -2215 44525 -2095
rect 44645 -2215 44690 -2095
rect 44810 -2215 44855 -2095
rect 44975 -2215 45030 -2095
rect 45150 -2215 45195 -2095
rect 45315 -2215 45360 -2095
rect 45480 -2215 45525 -2095
rect 45645 -2215 45700 -2095
rect 45820 -2215 45865 -2095
rect 45985 -2215 46030 -2095
rect 46150 -2215 46195 -2095
rect 46315 -2215 46370 -2095
rect 46490 -2215 46535 -2095
rect 46655 -2215 46700 -2095
rect 46820 -2215 46865 -2095
rect 46985 -2215 47040 -2095
rect 47160 -2215 47205 -2095
rect 47325 -2215 47370 -2095
rect 47490 -2215 47535 -2095
rect 47655 -2215 47665 -2095
rect 42165 -2260 47665 -2215
rect 42165 -2380 42175 -2260
rect 42295 -2380 42350 -2260
rect 42470 -2380 42515 -2260
rect 42635 -2380 42680 -2260
rect 42800 -2380 42845 -2260
rect 42965 -2380 43020 -2260
rect 43140 -2380 43185 -2260
rect 43305 -2380 43350 -2260
rect 43470 -2380 43515 -2260
rect 43635 -2380 43690 -2260
rect 43810 -2380 43855 -2260
rect 43975 -2380 44020 -2260
rect 44140 -2380 44185 -2260
rect 44305 -2380 44360 -2260
rect 44480 -2380 44525 -2260
rect 44645 -2380 44690 -2260
rect 44810 -2380 44855 -2260
rect 44975 -2380 45030 -2260
rect 45150 -2380 45195 -2260
rect 45315 -2380 45360 -2260
rect 45480 -2380 45525 -2260
rect 45645 -2380 45700 -2260
rect 45820 -2380 45865 -2260
rect 45985 -2380 46030 -2260
rect 46150 -2380 46195 -2260
rect 46315 -2380 46370 -2260
rect 46490 -2380 46535 -2260
rect 46655 -2380 46700 -2260
rect 46820 -2380 46865 -2260
rect 46985 -2380 47040 -2260
rect 47160 -2380 47205 -2260
rect 47325 -2380 47370 -2260
rect 47490 -2380 47535 -2260
rect 47655 -2380 47665 -2260
rect 42165 -2425 47665 -2380
rect 42165 -2545 42175 -2425
rect 42295 -2545 42350 -2425
rect 42470 -2545 42515 -2425
rect 42635 -2545 42680 -2425
rect 42800 -2545 42845 -2425
rect 42965 -2545 43020 -2425
rect 43140 -2545 43185 -2425
rect 43305 -2545 43350 -2425
rect 43470 -2545 43515 -2425
rect 43635 -2545 43690 -2425
rect 43810 -2545 43855 -2425
rect 43975 -2545 44020 -2425
rect 44140 -2545 44185 -2425
rect 44305 -2545 44360 -2425
rect 44480 -2545 44525 -2425
rect 44645 -2545 44690 -2425
rect 44810 -2545 44855 -2425
rect 44975 -2545 45030 -2425
rect 45150 -2545 45195 -2425
rect 45315 -2545 45360 -2425
rect 45480 -2545 45525 -2425
rect 45645 -2545 45700 -2425
rect 45820 -2545 45865 -2425
rect 45985 -2545 46030 -2425
rect 46150 -2545 46195 -2425
rect 46315 -2545 46370 -2425
rect 46490 -2545 46535 -2425
rect 46655 -2545 46700 -2425
rect 46820 -2545 46865 -2425
rect 46985 -2545 47040 -2425
rect 47160 -2545 47205 -2425
rect 47325 -2545 47370 -2425
rect 47490 -2545 47535 -2425
rect 47655 -2545 47665 -2425
rect 42165 -2600 47665 -2545
rect 42165 -2720 42175 -2600
rect 42295 -2720 42350 -2600
rect 42470 -2720 42515 -2600
rect 42635 -2720 42680 -2600
rect 42800 -2720 42845 -2600
rect 42965 -2720 43020 -2600
rect 43140 -2720 43185 -2600
rect 43305 -2720 43350 -2600
rect 43470 -2720 43515 -2600
rect 43635 -2720 43690 -2600
rect 43810 -2720 43855 -2600
rect 43975 -2720 44020 -2600
rect 44140 -2720 44185 -2600
rect 44305 -2720 44360 -2600
rect 44480 -2720 44525 -2600
rect 44645 -2720 44690 -2600
rect 44810 -2720 44855 -2600
rect 44975 -2720 45030 -2600
rect 45150 -2720 45195 -2600
rect 45315 -2720 45360 -2600
rect 45480 -2720 45525 -2600
rect 45645 -2720 45700 -2600
rect 45820 -2720 45865 -2600
rect 45985 -2720 46030 -2600
rect 46150 -2720 46195 -2600
rect 46315 -2720 46370 -2600
rect 46490 -2720 46535 -2600
rect 46655 -2720 46700 -2600
rect 46820 -2720 46865 -2600
rect 46985 -2720 47040 -2600
rect 47160 -2720 47205 -2600
rect 47325 -2720 47370 -2600
rect 47490 -2720 47535 -2600
rect 47655 -2720 47665 -2600
rect 42165 -2765 47665 -2720
rect 42165 -2885 42175 -2765
rect 42295 -2885 42350 -2765
rect 42470 -2885 42515 -2765
rect 42635 -2885 42680 -2765
rect 42800 -2885 42845 -2765
rect 42965 -2885 43020 -2765
rect 43140 -2885 43185 -2765
rect 43305 -2885 43350 -2765
rect 43470 -2885 43515 -2765
rect 43635 -2885 43690 -2765
rect 43810 -2885 43855 -2765
rect 43975 -2885 44020 -2765
rect 44140 -2885 44185 -2765
rect 44305 -2885 44360 -2765
rect 44480 -2885 44525 -2765
rect 44645 -2885 44690 -2765
rect 44810 -2885 44855 -2765
rect 44975 -2885 45030 -2765
rect 45150 -2885 45195 -2765
rect 45315 -2885 45360 -2765
rect 45480 -2885 45525 -2765
rect 45645 -2885 45700 -2765
rect 45820 -2885 45865 -2765
rect 45985 -2885 46030 -2765
rect 46150 -2885 46195 -2765
rect 46315 -2885 46370 -2765
rect 46490 -2885 46535 -2765
rect 46655 -2885 46700 -2765
rect 46820 -2885 46865 -2765
rect 46985 -2885 47040 -2765
rect 47160 -2885 47205 -2765
rect 47325 -2885 47370 -2765
rect 47490 -2885 47535 -2765
rect 47655 -2885 47665 -2765
rect 42165 -2930 47665 -2885
rect 42165 -3050 42175 -2930
rect 42295 -3050 42350 -2930
rect 42470 -3050 42515 -2930
rect 42635 -3050 42680 -2930
rect 42800 -3050 42845 -2930
rect 42965 -3050 43020 -2930
rect 43140 -3050 43185 -2930
rect 43305 -3050 43350 -2930
rect 43470 -3050 43515 -2930
rect 43635 -3050 43690 -2930
rect 43810 -3050 43855 -2930
rect 43975 -3050 44020 -2930
rect 44140 -3050 44185 -2930
rect 44305 -3050 44360 -2930
rect 44480 -3050 44525 -2930
rect 44645 -3050 44690 -2930
rect 44810 -3050 44855 -2930
rect 44975 -3050 45030 -2930
rect 45150 -3050 45195 -2930
rect 45315 -3050 45360 -2930
rect 45480 -3050 45525 -2930
rect 45645 -3050 45700 -2930
rect 45820 -3050 45865 -2930
rect 45985 -3050 46030 -2930
rect 46150 -3050 46195 -2930
rect 46315 -3050 46370 -2930
rect 46490 -3050 46535 -2930
rect 46655 -3050 46700 -2930
rect 46820 -3050 46865 -2930
rect 46985 -3050 47040 -2930
rect 47160 -3050 47205 -2930
rect 47325 -3050 47370 -2930
rect 47490 -3050 47535 -2930
rect 47655 -3050 47665 -2930
rect 42165 -3095 47665 -3050
rect 42165 -3215 42175 -3095
rect 42295 -3215 42350 -3095
rect 42470 -3215 42515 -3095
rect 42635 -3215 42680 -3095
rect 42800 -3215 42845 -3095
rect 42965 -3215 43020 -3095
rect 43140 -3215 43185 -3095
rect 43305 -3215 43350 -3095
rect 43470 -3215 43515 -3095
rect 43635 -3215 43690 -3095
rect 43810 -3215 43855 -3095
rect 43975 -3215 44020 -3095
rect 44140 -3215 44185 -3095
rect 44305 -3215 44360 -3095
rect 44480 -3215 44525 -3095
rect 44645 -3215 44690 -3095
rect 44810 -3215 44855 -3095
rect 44975 -3215 45030 -3095
rect 45150 -3215 45195 -3095
rect 45315 -3215 45360 -3095
rect 45480 -3215 45525 -3095
rect 45645 -3215 45700 -3095
rect 45820 -3215 45865 -3095
rect 45985 -3215 46030 -3095
rect 46150 -3215 46195 -3095
rect 46315 -3215 46370 -3095
rect 46490 -3215 46535 -3095
rect 46655 -3215 46700 -3095
rect 46820 -3215 46865 -3095
rect 46985 -3215 47040 -3095
rect 47160 -3215 47205 -3095
rect 47325 -3215 47370 -3095
rect 47490 -3215 47535 -3095
rect 47655 -3215 47665 -3095
rect 42165 -3270 47665 -3215
rect 42165 -3390 42175 -3270
rect 42295 -3390 42350 -3270
rect 42470 -3390 42515 -3270
rect 42635 -3390 42680 -3270
rect 42800 -3390 42845 -3270
rect 42965 -3390 43020 -3270
rect 43140 -3390 43185 -3270
rect 43305 -3390 43350 -3270
rect 43470 -3390 43515 -3270
rect 43635 -3390 43690 -3270
rect 43810 -3390 43855 -3270
rect 43975 -3390 44020 -3270
rect 44140 -3390 44185 -3270
rect 44305 -3390 44360 -3270
rect 44480 -3390 44525 -3270
rect 44645 -3390 44690 -3270
rect 44810 -3390 44855 -3270
rect 44975 -3390 45030 -3270
rect 45150 -3390 45195 -3270
rect 45315 -3390 45360 -3270
rect 45480 -3390 45525 -3270
rect 45645 -3390 45700 -3270
rect 45820 -3390 45865 -3270
rect 45985 -3390 46030 -3270
rect 46150 -3390 46195 -3270
rect 46315 -3390 46370 -3270
rect 46490 -3390 46535 -3270
rect 46655 -3390 46700 -3270
rect 46820 -3390 46865 -3270
rect 46985 -3390 47040 -3270
rect 47160 -3390 47205 -3270
rect 47325 -3390 47370 -3270
rect 47490 -3390 47535 -3270
rect 47655 -3390 47665 -3270
rect 42165 -3435 47665 -3390
rect 42165 -3555 42175 -3435
rect 42295 -3555 42350 -3435
rect 42470 -3555 42515 -3435
rect 42635 -3555 42680 -3435
rect 42800 -3555 42845 -3435
rect 42965 -3555 43020 -3435
rect 43140 -3555 43185 -3435
rect 43305 -3555 43350 -3435
rect 43470 -3555 43515 -3435
rect 43635 -3555 43690 -3435
rect 43810 -3555 43855 -3435
rect 43975 -3555 44020 -3435
rect 44140 -3555 44185 -3435
rect 44305 -3555 44360 -3435
rect 44480 -3555 44525 -3435
rect 44645 -3555 44690 -3435
rect 44810 -3555 44855 -3435
rect 44975 -3555 45030 -3435
rect 45150 -3555 45195 -3435
rect 45315 -3555 45360 -3435
rect 45480 -3555 45525 -3435
rect 45645 -3555 45700 -3435
rect 45820 -3555 45865 -3435
rect 45985 -3555 46030 -3435
rect 46150 -3555 46195 -3435
rect 46315 -3555 46370 -3435
rect 46490 -3555 46535 -3435
rect 46655 -3555 46700 -3435
rect 46820 -3555 46865 -3435
rect 46985 -3555 47040 -3435
rect 47160 -3555 47205 -3435
rect 47325 -3555 47370 -3435
rect 47490 -3555 47535 -3435
rect 47655 -3555 47665 -3435
rect 42165 -3600 47665 -3555
rect 42165 -3720 42175 -3600
rect 42295 -3720 42350 -3600
rect 42470 -3720 42515 -3600
rect 42635 -3720 42680 -3600
rect 42800 -3720 42845 -3600
rect 42965 -3720 43020 -3600
rect 43140 -3720 43185 -3600
rect 43305 -3720 43350 -3600
rect 43470 -3720 43515 -3600
rect 43635 -3720 43690 -3600
rect 43810 -3720 43855 -3600
rect 43975 -3720 44020 -3600
rect 44140 -3720 44185 -3600
rect 44305 -3720 44360 -3600
rect 44480 -3720 44525 -3600
rect 44645 -3720 44690 -3600
rect 44810 -3720 44855 -3600
rect 44975 -3720 45030 -3600
rect 45150 -3720 45195 -3600
rect 45315 -3720 45360 -3600
rect 45480 -3720 45525 -3600
rect 45645 -3720 45700 -3600
rect 45820 -3720 45865 -3600
rect 45985 -3720 46030 -3600
rect 46150 -3720 46195 -3600
rect 46315 -3720 46370 -3600
rect 46490 -3720 46535 -3600
rect 46655 -3720 46700 -3600
rect 46820 -3720 46865 -3600
rect 46985 -3720 47040 -3600
rect 47160 -3720 47205 -3600
rect 47325 -3720 47370 -3600
rect 47490 -3720 47535 -3600
rect 47655 -3720 47665 -3600
rect 42165 -3765 47665 -3720
rect 42165 -3885 42175 -3765
rect 42295 -3885 42350 -3765
rect 42470 -3885 42515 -3765
rect 42635 -3885 42680 -3765
rect 42800 -3885 42845 -3765
rect 42965 -3885 43020 -3765
rect 43140 -3885 43185 -3765
rect 43305 -3885 43350 -3765
rect 43470 -3885 43515 -3765
rect 43635 -3885 43690 -3765
rect 43810 -3885 43855 -3765
rect 43975 -3885 44020 -3765
rect 44140 -3885 44185 -3765
rect 44305 -3885 44360 -3765
rect 44480 -3885 44525 -3765
rect 44645 -3885 44690 -3765
rect 44810 -3885 44855 -3765
rect 44975 -3885 45030 -3765
rect 45150 -3885 45195 -3765
rect 45315 -3885 45360 -3765
rect 45480 -3885 45525 -3765
rect 45645 -3885 45700 -3765
rect 45820 -3885 45865 -3765
rect 45985 -3885 46030 -3765
rect 46150 -3885 46195 -3765
rect 46315 -3885 46370 -3765
rect 46490 -3885 46535 -3765
rect 46655 -3885 46700 -3765
rect 46820 -3885 46865 -3765
rect 46985 -3885 47040 -3765
rect 47160 -3885 47205 -3765
rect 47325 -3885 47370 -3765
rect 47490 -3885 47535 -3765
rect 47655 -3885 47665 -3765
rect 42165 -3940 47665 -3885
rect 42165 -4060 42175 -3940
rect 42295 -4060 42350 -3940
rect 42470 -4060 42515 -3940
rect 42635 -4060 42680 -3940
rect 42800 -4060 42845 -3940
rect 42965 -4060 43020 -3940
rect 43140 -4060 43185 -3940
rect 43305 -4060 43350 -3940
rect 43470 -4060 43515 -3940
rect 43635 -4060 43690 -3940
rect 43810 -4060 43855 -3940
rect 43975 -4060 44020 -3940
rect 44140 -4060 44185 -3940
rect 44305 -4060 44360 -3940
rect 44480 -4060 44525 -3940
rect 44645 -4060 44690 -3940
rect 44810 -4060 44855 -3940
rect 44975 -4060 45030 -3940
rect 45150 -4060 45195 -3940
rect 45315 -4060 45360 -3940
rect 45480 -4060 45525 -3940
rect 45645 -4060 45700 -3940
rect 45820 -4060 45865 -3940
rect 45985 -4060 46030 -3940
rect 46150 -4060 46195 -3940
rect 46315 -4060 46370 -3940
rect 46490 -4060 46535 -3940
rect 46655 -4060 46700 -3940
rect 46820 -4060 46865 -3940
rect 46985 -4060 47040 -3940
rect 47160 -4060 47205 -3940
rect 47325 -4060 47370 -3940
rect 47490 -4060 47535 -3940
rect 47655 -4060 47665 -3940
rect 42165 -4070 47665 -4060
rect 47855 1420 53355 1430
rect 47855 1300 47865 1420
rect 47985 1300 48040 1420
rect 48160 1300 48205 1420
rect 48325 1300 48370 1420
rect 48490 1300 48535 1420
rect 48655 1300 48710 1420
rect 48830 1300 48875 1420
rect 48995 1300 49040 1420
rect 49160 1300 49205 1420
rect 49325 1300 49380 1420
rect 49500 1300 49545 1420
rect 49665 1300 49710 1420
rect 49830 1300 49875 1420
rect 49995 1300 50050 1420
rect 50170 1300 50215 1420
rect 50335 1300 50380 1420
rect 50500 1300 50545 1420
rect 50665 1300 50720 1420
rect 50840 1300 50885 1420
rect 51005 1300 51050 1420
rect 51170 1300 51215 1420
rect 51335 1300 51390 1420
rect 51510 1300 51555 1420
rect 51675 1300 51720 1420
rect 51840 1300 51885 1420
rect 52005 1300 52060 1420
rect 52180 1300 52225 1420
rect 52345 1300 52390 1420
rect 52510 1300 52555 1420
rect 52675 1300 52730 1420
rect 52850 1300 52895 1420
rect 53015 1300 53060 1420
rect 53180 1300 53225 1420
rect 53345 1300 53355 1420
rect 47855 1255 53355 1300
rect 47855 1135 47865 1255
rect 47985 1135 48040 1255
rect 48160 1135 48205 1255
rect 48325 1135 48370 1255
rect 48490 1135 48535 1255
rect 48655 1135 48710 1255
rect 48830 1135 48875 1255
rect 48995 1135 49040 1255
rect 49160 1135 49205 1255
rect 49325 1135 49380 1255
rect 49500 1135 49545 1255
rect 49665 1135 49710 1255
rect 49830 1135 49875 1255
rect 49995 1135 50050 1255
rect 50170 1135 50215 1255
rect 50335 1135 50380 1255
rect 50500 1135 50545 1255
rect 50665 1135 50720 1255
rect 50840 1135 50885 1255
rect 51005 1135 51050 1255
rect 51170 1135 51215 1255
rect 51335 1135 51390 1255
rect 51510 1135 51555 1255
rect 51675 1135 51720 1255
rect 51840 1135 51885 1255
rect 52005 1135 52060 1255
rect 52180 1135 52225 1255
rect 52345 1135 52390 1255
rect 52510 1135 52555 1255
rect 52675 1135 52730 1255
rect 52850 1135 52895 1255
rect 53015 1135 53060 1255
rect 53180 1135 53225 1255
rect 53345 1135 53355 1255
rect 47855 1090 53355 1135
rect 47855 970 47865 1090
rect 47985 970 48040 1090
rect 48160 970 48205 1090
rect 48325 970 48370 1090
rect 48490 970 48535 1090
rect 48655 970 48710 1090
rect 48830 970 48875 1090
rect 48995 970 49040 1090
rect 49160 970 49205 1090
rect 49325 970 49380 1090
rect 49500 970 49545 1090
rect 49665 970 49710 1090
rect 49830 970 49875 1090
rect 49995 970 50050 1090
rect 50170 970 50215 1090
rect 50335 970 50380 1090
rect 50500 970 50545 1090
rect 50665 970 50720 1090
rect 50840 970 50885 1090
rect 51005 970 51050 1090
rect 51170 970 51215 1090
rect 51335 970 51390 1090
rect 51510 970 51555 1090
rect 51675 970 51720 1090
rect 51840 970 51885 1090
rect 52005 970 52060 1090
rect 52180 970 52225 1090
rect 52345 970 52390 1090
rect 52510 970 52555 1090
rect 52675 970 52730 1090
rect 52850 970 52895 1090
rect 53015 970 53060 1090
rect 53180 970 53225 1090
rect 53345 970 53355 1090
rect 47855 925 53355 970
rect 47855 805 47865 925
rect 47985 805 48040 925
rect 48160 805 48205 925
rect 48325 805 48370 925
rect 48490 805 48535 925
rect 48655 805 48710 925
rect 48830 805 48875 925
rect 48995 805 49040 925
rect 49160 805 49205 925
rect 49325 805 49380 925
rect 49500 805 49545 925
rect 49665 805 49710 925
rect 49830 805 49875 925
rect 49995 805 50050 925
rect 50170 805 50215 925
rect 50335 805 50380 925
rect 50500 805 50545 925
rect 50665 805 50720 925
rect 50840 805 50885 925
rect 51005 805 51050 925
rect 51170 805 51215 925
rect 51335 805 51390 925
rect 51510 805 51555 925
rect 51675 805 51720 925
rect 51840 805 51885 925
rect 52005 805 52060 925
rect 52180 805 52225 925
rect 52345 805 52390 925
rect 52510 805 52555 925
rect 52675 805 52730 925
rect 52850 805 52895 925
rect 53015 805 53060 925
rect 53180 805 53225 925
rect 53345 805 53355 925
rect 47855 750 53355 805
rect 47855 630 47865 750
rect 47985 630 48040 750
rect 48160 630 48205 750
rect 48325 630 48370 750
rect 48490 630 48535 750
rect 48655 630 48710 750
rect 48830 630 48875 750
rect 48995 630 49040 750
rect 49160 630 49205 750
rect 49325 630 49380 750
rect 49500 630 49545 750
rect 49665 630 49710 750
rect 49830 630 49875 750
rect 49995 630 50050 750
rect 50170 630 50215 750
rect 50335 630 50380 750
rect 50500 630 50545 750
rect 50665 630 50720 750
rect 50840 630 50885 750
rect 51005 630 51050 750
rect 51170 630 51215 750
rect 51335 630 51390 750
rect 51510 630 51555 750
rect 51675 630 51720 750
rect 51840 630 51885 750
rect 52005 630 52060 750
rect 52180 630 52225 750
rect 52345 630 52390 750
rect 52510 630 52555 750
rect 52675 630 52730 750
rect 52850 630 52895 750
rect 53015 630 53060 750
rect 53180 630 53225 750
rect 53345 630 53355 750
rect 47855 585 53355 630
rect 47855 465 47865 585
rect 47985 465 48040 585
rect 48160 465 48205 585
rect 48325 465 48370 585
rect 48490 465 48535 585
rect 48655 465 48710 585
rect 48830 465 48875 585
rect 48995 465 49040 585
rect 49160 465 49205 585
rect 49325 465 49380 585
rect 49500 465 49545 585
rect 49665 465 49710 585
rect 49830 465 49875 585
rect 49995 465 50050 585
rect 50170 465 50215 585
rect 50335 465 50380 585
rect 50500 465 50545 585
rect 50665 465 50720 585
rect 50840 465 50885 585
rect 51005 465 51050 585
rect 51170 465 51215 585
rect 51335 465 51390 585
rect 51510 465 51555 585
rect 51675 465 51720 585
rect 51840 465 51885 585
rect 52005 465 52060 585
rect 52180 465 52225 585
rect 52345 465 52390 585
rect 52510 465 52555 585
rect 52675 465 52730 585
rect 52850 465 52895 585
rect 53015 465 53060 585
rect 53180 465 53225 585
rect 53345 465 53355 585
rect 47855 420 53355 465
rect 47855 300 47865 420
rect 47985 300 48040 420
rect 48160 300 48205 420
rect 48325 300 48370 420
rect 48490 300 48535 420
rect 48655 300 48710 420
rect 48830 300 48875 420
rect 48995 300 49040 420
rect 49160 300 49205 420
rect 49325 300 49380 420
rect 49500 300 49545 420
rect 49665 300 49710 420
rect 49830 300 49875 420
rect 49995 300 50050 420
rect 50170 300 50215 420
rect 50335 300 50380 420
rect 50500 300 50545 420
rect 50665 300 50720 420
rect 50840 300 50885 420
rect 51005 300 51050 420
rect 51170 300 51215 420
rect 51335 300 51390 420
rect 51510 300 51555 420
rect 51675 300 51720 420
rect 51840 300 51885 420
rect 52005 300 52060 420
rect 52180 300 52225 420
rect 52345 300 52390 420
rect 52510 300 52555 420
rect 52675 300 52730 420
rect 52850 300 52895 420
rect 53015 300 53060 420
rect 53180 300 53225 420
rect 53345 300 53355 420
rect 47855 255 53355 300
rect 47855 135 47865 255
rect 47985 135 48040 255
rect 48160 135 48205 255
rect 48325 135 48370 255
rect 48490 135 48535 255
rect 48655 135 48710 255
rect 48830 135 48875 255
rect 48995 135 49040 255
rect 49160 135 49205 255
rect 49325 135 49380 255
rect 49500 135 49545 255
rect 49665 135 49710 255
rect 49830 135 49875 255
rect 49995 135 50050 255
rect 50170 135 50215 255
rect 50335 135 50380 255
rect 50500 135 50545 255
rect 50665 135 50720 255
rect 50840 135 50885 255
rect 51005 135 51050 255
rect 51170 135 51215 255
rect 51335 135 51390 255
rect 51510 135 51555 255
rect 51675 135 51720 255
rect 51840 135 51885 255
rect 52005 135 52060 255
rect 52180 135 52225 255
rect 52345 135 52390 255
rect 52510 135 52555 255
rect 52675 135 52730 255
rect 52850 135 52895 255
rect 53015 135 53060 255
rect 53180 135 53225 255
rect 53345 135 53355 255
rect 47855 80 53355 135
rect 47855 -40 47865 80
rect 47985 -40 48040 80
rect 48160 -40 48205 80
rect 48325 -40 48370 80
rect 48490 -40 48535 80
rect 48655 -40 48710 80
rect 48830 -40 48875 80
rect 48995 -40 49040 80
rect 49160 -40 49205 80
rect 49325 -40 49380 80
rect 49500 -40 49545 80
rect 49665 -40 49710 80
rect 49830 -40 49875 80
rect 49995 -40 50050 80
rect 50170 -40 50215 80
rect 50335 -40 50380 80
rect 50500 -40 50545 80
rect 50665 -40 50720 80
rect 50840 -40 50885 80
rect 51005 -40 51050 80
rect 51170 -40 51215 80
rect 51335 -40 51390 80
rect 51510 -40 51555 80
rect 51675 -40 51720 80
rect 51840 -40 51885 80
rect 52005 -40 52060 80
rect 52180 -40 52225 80
rect 52345 -40 52390 80
rect 52510 -40 52555 80
rect 52675 -40 52730 80
rect 52850 -40 52895 80
rect 53015 -40 53060 80
rect 53180 -40 53225 80
rect 53345 -40 53355 80
rect 47855 -85 53355 -40
rect 47855 -205 47865 -85
rect 47985 -205 48040 -85
rect 48160 -205 48205 -85
rect 48325 -205 48370 -85
rect 48490 -205 48535 -85
rect 48655 -205 48710 -85
rect 48830 -205 48875 -85
rect 48995 -205 49040 -85
rect 49160 -205 49205 -85
rect 49325 -205 49380 -85
rect 49500 -205 49545 -85
rect 49665 -205 49710 -85
rect 49830 -205 49875 -85
rect 49995 -205 50050 -85
rect 50170 -205 50215 -85
rect 50335 -205 50380 -85
rect 50500 -205 50545 -85
rect 50665 -205 50720 -85
rect 50840 -205 50885 -85
rect 51005 -205 51050 -85
rect 51170 -205 51215 -85
rect 51335 -205 51390 -85
rect 51510 -205 51555 -85
rect 51675 -205 51720 -85
rect 51840 -205 51885 -85
rect 52005 -205 52060 -85
rect 52180 -205 52225 -85
rect 52345 -205 52390 -85
rect 52510 -205 52555 -85
rect 52675 -205 52730 -85
rect 52850 -205 52895 -85
rect 53015 -205 53060 -85
rect 53180 -205 53225 -85
rect 53345 -205 53355 -85
rect 47855 -250 53355 -205
rect 47855 -370 47865 -250
rect 47985 -370 48040 -250
rect 48160 -370 48205 -250
rect 48325 -370 48370 -250
rect 48490 -370 48535 -250
rect 48655 -370 48710 -250
rect 48830 -370 48875 -250
rect 48995 -370 49040 -250
rect 49160 -370 49205 -250
rect 49325 -370 49380 -250
rect 49500 -370 49545 -250
rect 49665 -370 49710 -250
rect 49830 -370 49875 -250
rect 49995 -370 50050 -250
rect 50170 -370 50215 -250
rect 50335 -370 50380 -250
rect 50500 -370 50545 -250
rect 50665 -370 50720 -250
rect 50840 -370 50885 -250
rect 51005 -370 51050 -250
rect 51170 -370 51215 -250
rect 51335 -370 51390 -250
rect 51510 -370 51555 -250
rect 51675 -370 51720 -250
rect 51840 -370 51885 -250
rect 52005 -370 52060 -250
rect 52180 -370 52225 -250
rect 52345 -370 52390 -250
rect 52510 -370 52555 -250
rect 52675 -370 52730 -250
rect 52850 -370 52895 -250
rect 53015 -370 53060 -250
rect 53180 -370 53225 -250
rect 53345 -370 53355 -250
rect 47855 -415 53355 -370
rect 47855 -535 47865 -415
rect 47985 -535 48040 -415
rect 48160 -535 48205 -415
rect 48325 -535 48370 -415
rect 48490 -535 48535 -415
rect 48655 -535 48710 -415
rect 48830 -535 48875 -415
rect 48995 -535 49040 -415
rect 49160 -535 49205 -415
rect 49325 -535 49380 -415
rect 49500 -535 49545 -415
rect 49665 -535 49710 -415
rect 49830 -535 49875 -415
rect 49995 -535 50050 -415
rect 50170 -535 50215 -415
rect 50335 -535 50380 -415
rect 50500 -535 50545 -415
rect 50665 -535 50720 -415
rect 50840 -535 50885 -415
rect 51005 -535 51050 -415
rect 51170 -535 51215 -415
rect 51335 -535 51390 -415
rect 51510 -535 51555 -415
rect 51675 -535 51720 -415
rect 51840 -535 51885 -415
rect 52005 -535 52060 -415
rect 52180 -535 52225 -415
rect 52345 -535 52390 -415
rect 52510 -535 52555 -415
rect 52675 -535 52730 -415
rect 52850 -535 52895 -415
rect 53015 -535 53060 -415
rect 53180 -535 53225 -415
rect 53345 -535 53355 -415
rect 47855 -590 53355 -535
rect 47855 -710 47865 -590
rect 47985 -710 48040 -590
rect 48160 -710 48205 -590
rect 48325 -710 48370 -590
rect 48490 -710 48535 -590
rect 48655 -710 48710 -590
rect 48830 -710 48875 -590
rect 48995 -710 49040 -590
rect 49160 -710 49205 -590
rect 49325 -710 49380 -590
rect 49500 -710 49545 -590
rect 49665 -710 49710 -590
rect 49830 -710 49875 -590
rect 49995 -710 50050 -590
rect 50170 -710 50215 -590
rect 50335 -710 50380 -590
rect 50500 -710 50545 -590
rect 50665 -710 50720 -590
rect 50840 -710 50885 -590
rect 51005 -710 51050 -590
rect 51170 -710 51215 -590
rect 51335 -710 51390 -590
rect 51510 -710 51555 -590
rect 51675 -710 51720 -590
rect 51840 -710 51885 -590
rect 52005 -710 52060 -590
rect 52180 -710 52225 -590
rect 52345 -710 52390 -590
rect 52510 -710 52555 -590
rect 52675 -710 52730 -590
rect 52850 -710 52895 -590
rect 53015 -710 53060 -590
rect 53180 -710 53225 -590
rect 53345 -710 53355 -590
rect 47855 -755 53355 -710
rect 47855 -875 47865 -755
rect 47985 -875 48040 -755
rect 48160 -875 48205 -755
rect 48325 -875 48370 -755
rect 48490 -875 48535 -755
rect 48655 -875 48710 -755
rect 48830 -875 48875 -755
rect 48995 -875 49040 -755
rect 49160 -875 49205 -755
rect 49325 -875 49380 -755
rect 49500 -875 49545 -755
rect 49665 -875 49710 -755
rect 49830 -875 49875 -755
rect 49995 -875 50050 -755
rect 50170 -875 50215 -755
rect 50335 -875 50380 -755
rect 50500 -875 50545 -755
rect 50665 -875 50720 -755
rect 50840 -875 50885 -755
rect 51005 -875 51050 -755
rect 51170 -875 51215 -755
rect 51335 -875 51390 -755
rect 51510 -875 51555 -755
rect 51675 -875 51720 -755
rect 51840 -875 51885 -755
rect 52005 -875 52060 -755
rect 52180 -875 52225 -755
rect 52345 -875 52390 -755
rect 52510 -875 52555 -755
rect 52675 -875 52730 -755
rect 52850 -875 52895 -755
rect 53015 -875 53060 -755
rect 53180 -875 53225 -755
rect 53345 -875 53355 -755
rect 47855 -920 53355 -875
rect 47855 -1040 47865 -920
rect 47985 -1040 48040 -920
rect 48160 -1040 48205 -920
rect 48325 -1040 48370 -920
rect 48490 -1040 48535 -920
rect 48655 -1040 48710 -920
rect 48830 -1040 48875 -920
rect 48995 -1040 49040 -920
rect 49160 -1040 49205 -920
rect 49325 -1040 49380 -920
rect 49500 -1040 49545 -920
rect 49665 -1040 49710 -920
rect 49830 -1040 49875 -920
rect 49995 -1040 50050 -920
rect 50170 -1040 50215 -920
rect 50335 -1040 50380 -920
rect 50500 -1040 50545 -920
rect 50665 -1040 50720 -920
rect 50840 -1040 50885 -920
rect 51005 -1040 51050 -920
rect 51170 -1040 51215 -920
rect 51335 -1040 51390 -920
rect 51510 -1040 51555 -920
rect 51675 -1040 51720 -920
rect 51840 -1040 51885 -920
rect 52005 -1040 52060 -920
rect 52180 -1040 52225 -920
rect 52345 -1040 52390 -920
rect 52510 -1040 52555 -920
rect 52675 -1040 52730 -920
rect 52850 -1040 52895 -920
rect 53015 -1040 53060 -920
rect 53180 -1040 53225 -920
rect 53345 -1040 53355 -920
rect 47855 -1085 53355 -1040
rect 47855 -1205 47865 -1085
rect 47985 -1205 48040 -1085
rect 48160 -1205 48205 -1085
rect 48325 -1205 48370 -1085
rect 48490 -1205 48535 -1085
rect 48655 -1205 48710 -1085
rect 48830 -1205 48875 -1085
rect 48995 -1205 49040 -1085
rect 49160 -1205 49205 -1085
rect 49325 -1205 49380 -1085
rect 49500 -1205 49545 -1085
rect 49665 -1205 49710 -1085
rect 49830 -1205 49875 -1085
rect 49995 -1205 50050 -1085
rect 50170 -1205 50215 -1085
rect 50335 -1205 50380 -1085
rect 50500 -1205 50545 -1085
rect 50665 -1205 50720 -1085
rect 50840 -1205 50885 -1085
rect 51005 -1205 51050 -1085
rect 51170 -1205 51215 -1085
rect 51335 -1205 51390 -1085
rect 51510 -1205 51555 -1085
rect 51675 -1205 51720 -1085
rect 51840 -1205 51885 -1085
rect 52005 -1205 52060 -1085
rect 52180 -1205 52225 -1085
rect 52345 -1205 52390 -1085
rect 52510 -1205 52555 -1085
rect 52675 -1205 52730 -1085
rect 52850 -1205 52895 -1085
rect 53015 -1205 53060 -1085
rect 53180 -1205 53225 -1085
rect 53345 -1205 53355 -1085
rect 47855 -1260 53355 -1205
rect 47855 -1380 47865 -1260
rect 47985 -1380 48040 -1260
rect 48160 -1380 48205 -1260
rect 48325 -1380 48370 -1260
rect 48490 -1380 48535 -1260
rect 48655 -1380 48710 -1260
rect 48830 -1380 48875 -1260
rect 48995 -1380 49040 -1260
rect 49160 -1380 49205 -1260
rect 49325 -1380 49380 -1260
rect 49500 -1380 49545 -1260
rect 49665 -1380 49710 -1260
rect 49830 -1380 49875 -1260
rect 49995 -1380 50050 -1260
rect 50170 -1380 50215 -1260
rect 50335 -1380 50380 -1260
rect 50500 -1380 50545 -1260
rect 50665 -1380 50720 -1260
rect 50840 -1380 50885 -1260
rect 51005 -1380 51050 -1260
rect 51170 -1380 51215 -1260
rect 51335 -1380 51390 -1260
rect 51510 -1380 51555 -1260
rect 51675 -1380 51720 -1260
rect 51840 -1380 51885 -1260
rect 52005 -1380 52060 -1260
rect 52180 -1380 52225 -1260
rect 52345 -1380 52390 -1260
rect 52510 -1380 52555 -1260
rect 52675 -1380 52730 -1260
rect 52850 -1380 52895 -1260
rect 53015 -1380 53060 -1260
rect 53180 -1380 53225 -1260
rect 53345 -1380 53355 -1260
rect 47855 -1425 53355 -1380
rect 47855 -1545 47865 -1425
rect 47985 -1545 48040 -1425
rect 48160 -1545 48205 -1425
rect 48325 -1545 48370 -1425
rect 48490 -1545 48535 -1425
rect 48655 -1545 48710 -1425
rect 48830 -1545 48875 -1425
rect 48995 -1545 49040 -1425
rect 49160 -1545 49205 -1425
rect 49325 -1545 49380 -1425
rect 49500 -1545 49545 -1425
rect 49665 -1545 49710 -1425
rect 49830 -1545 49875 -1425
rect 49995 -1545 50050 -1425
rect 50170 -1545 50215 -1425
rect 50335 -1545 50380 -1425
rect 50500 -1545 50545 -1425
rect 50665 -1545 50720 -1425
rect 50840 -1545 50885 -1425
rect 51005 -1545 51050 -1425
rect 51170 -1545 51215 -1425
rect 51335 -1545 51390 -1425
rect 51510 -1545 51555 -1425
rect 51675 -1545 51720 -1425
rect 51840 -1545 51885 -1425
rect 52005 -1545 52060 -1425
rect 52180 -1545 52225 -1425
rect 52345 -1545 52390 -1425
rect 52510 -1545 52555 -1425
rect 52675 -1545 52730 -1425
rect 52850 -1545 52895 -1425
rect 53015 -1545 53060 -1425
rect 53180 -1545 53225 -1425
rect 53345 -1545 53355 -1425
rect 47855 -1590 53355 -1545
rect 47855 -1710 47865 -1590
rect 47985 -1710 48040 -1590
rect 48160 -1710 48205 -1590
rect 48325 -1710 48370 -1590
rect 48490 -1710 48535 -1590
rect 48655 -1710 48710 -1590
rect 48830 -1710 48875 -1590
rect 48995 -1710 49040 -1590
rect 49160 -1710 49205 -1590
rect 49325 -1710 49380 -1590
rect 49500 -1710 49545 -1590
rect 49665 -1710 49710 -1590
rect 49830 -1710 49875 -1590
rect 49995 -1710 50050 -1590
rect 50170 -1710 50215 -1590
rect 50335 -1710 50380 -1590
rect 50500 -1710 50545 -1590
rect 50665 -1710 50720 -1590
rect 50840 -1710 50885 -1590
rect 51005 -1710 51050 -1590
rect 51170 -1710 51215 -1590
rect 51335 -1710 51390 -1590
rect 51510 -1710 51555 -1590
rect 51675 -1710 51720 -1590
rect 51840 -1710 51885 -1590
rect 52005 -1710 52060 -1590
rect 52180 -1710 52225 -1590
rect 52345 -1710 52390 -1590
rect 52510 -1710 52555 -1590
rect 52675 -1710 52730 -1590
rect 52850 -1710 52895 -1590
rect 53015 -1710 53060 -1590
rect 53180 -1710 53225 -1590
rect 53345 -1710 53355 -1590
rect 47855 -1755 53355 -1710
rect 47855 -1875 47865 -1755
rect 47985 -1875 48040 -1755
rect 48160 -1875 48205 -1755
rect 48325 -1875 48370 -1755
rect 48490 -1875 48535 -1755
rect 48655 -1875 48710 -1755
rect 48830 -1875 48875 -1755
rect 48995 -1875 49040 -1755
rect 49160 -1875 49205 -1755
rect 49325 -1875 49380 -1755
rect 49500 -1875 49545 -1755
rect 49665 -1875 49710 -1755
rect 49830 -1875 49875 -1755
rect 49995 -1875 50050 -1755
rect 50170 -1875 50215 -1755
rect 50335 -1875 50380 -1755
rect 50500 -1875 50545 -1755
rect 50665 -1875 50720 -1755
rect 50840 -1875 50885 -1755
rect 51005 -1875 51050 -1755
rect 51170 -1875 51215 -1755
rect 51335 -1875 51390 -1755
rect 51510 -1875 51555 -1755
rect 51675 -1875 51720 -1755
rect 51840 -1875 51885 -1755
rect 52005 -1875 52060 -1755
rect 52180 -1875 52225 -1755
rect 52345 -1875 52390 -1755
rect 52510 -1875 52555 -1755
rect 52675 -1875 52730 -1755
rect 52850 -1875 52895 -1755
rect 53015 -1875 53060 -1755
rect 53180 -1875 53225 -1755
rect 53345 -1875 53355 -1755
rect 47855 -1930 53355 -1875
rect 47855 -2050 47865 -1930
rect 47985 -2050 48040 -1930
rect 48160 -2050 48205 -1930
rect 48325 -2050 48370 -1930
rect 48490 -2050 48535 -1930
rect 48655 -2050 48710 -1930
rect 48830 -2050 48875 -1930
rect 48995 -2050 49040 -1930
rect 49160 -2050 49205 -1930
rect 49325 -2050 49380 -1930
rect 49500 -2050 49545 -1930
rect 49665 -2050 49710 -1930
rect 49830 -2050 49875 -1930
rect 49995 -2050 50050 -1930
rect 50170 -2050 50215 -1930
rect 50335 -2050 50380 -1930
rect 50500 -2050 50545 -1930
rect 50665 -2050 50720 -1930
rect 50840 -2050 50885 -1930
rect 51005 -2050 51050 -1930
rect 51170 -2050 51215 -1930
rect 51335 -2050 51390 -1930
rect 51510 -2050 51555 -1930
rect 51675 -2050 51720 -1930
rect 51840 -2050 51885 -1930
rect 52005 -2050 52060 -1930
rect 52180 -2050 52225 -1930
rect 52345 -2050 52390 -1930
rect 52510 -2050 52555 -1930
rect 52675 -2050 52730 -1930
rect 52850 -2050 52895 -1930
rect 53015 -2050 53060 -1930
rect 53180 -2050 53225 -1930
rect 53345 -2050 53355 -1930
rect 47855 -2095 53355 -2050
rect 47855 -2215 47865 -2095
rect 47985 -2215 48040 -2095
rect 48160 -2215 48205 -2095
rect 48325 -2215 48370 -2095
rect 48490 -2215 48535 -2095
rect 48655 -2215 48710 -2095
rect 48830 -2215 48875 -2095
rect 48995 -2215 49040 -2095
rect 49160 -2215 49205 -2095
rect 49325 -2215 49380 -2095
rect 49500 -2215 49545 -2095
rect 49665 -2215 49710 -2095
rect 49830 -2215 49875 -2095
rect 49995 -2215 50050 -2095
rect 50170 -2215 50215 -2095
rect 50335 -2215 50380 -2095
rect 50500 -2215 50545 -2095
rect 50665 -2215 50720 -2095
rect 50840 -2215 50885 -2095
rect 51005 -2215 51050 -2095
rect 51170 -2215 51215 -2095
rect 51335 -2215 51390 -2095
rect 51510 -2215 51555 -2095
rect 51675 -2215 51720 -2095
rect 51840 -2215 51885 -2095
rect 52005 -2215 52060 -2095
rect 52180 -2215 52225 -2095
rect 52345 -2215 52390 -2095
rect 52510 -2215 52555 -2095
rect 52675 -2215 52730 -2095
rect 52850 -2215 52895 -2095
rect 53015 -2215 53060 -2095
rect 53180 -2215 53225 -2095
rect 53345 -2215 53355 -2095
rect 47855 -2260 53355 -2215
rect 47855 -2380 47865 -2260
rect 47985 -2380 48040 -2260
rect 48160 -2380 48205 -2260
rect 48325 -2380 48370 -2260
rect 48490 -2380 48535 -2260
rect 48655 -2380 48710 -2260
rect 48830 -2380 48875 -2260
rect 48995 -2380 49040 -2260
rect 49160 -2380 49205 -2260
rect 49325 -2380 49380 -2260
rect 49500 -2380 49545 -2260
rect 49665 -2380 49710 -2260
rect 49830 -2380 49875 -2260
rect 49995 -2380 50050 -2260
rect 50170 -2380 50215 -2260
rect 50335 -2380 50380 -2260
rect 50500 -2380 50545 -2260
rect 50665 -2380 50720 -2260
rect 50840 -2380 50885 -2260
rect 51005 -2380 51050 -2260
rect 51170 -2380 51215 -2260
rect 51335 -2380 51390 -2260
rect 51510 -2380 51555 -2260
rect 51675 -2380 51720 -2260
rect 51840 -2380 51885 -2260
rect 52005 -2380 52060 -2260
rect 52180 -2380 52225 -2260
rect 52345 -2380 52390 -2260
rect 52510 -2380 52555 -2260
rect 52675 -2380 52730 -2260
rect 52850 -2380 52895 -2260
rect 53015 -2380 53060 -2260
rect 53180 -2380 53225 -2260
rect 53345 -2380 53355 -2260
rect 47855 -2425 53355 -2380
rect 47855 -2545 47865 -2425
rect 47985 -2545 48040 -2425
rect 48160 -2545 48205 -2425
rect 48325 -2545 48370 -2425
rect 48490 -2545 48535 -2425
rect 48655 -2545 48710 -2425
rect 48830 -2545 48875 -2425
rect 48995 -2545 49040 -2425
rect 49160 -2545 49205 -2425
rect 49325 -2545 49380 -2425
rect 49500 -2545 49545 -2425
rect 49665 -2545 49710 -2425
rect 49830 -2545 49875 -2425
rect 49995 -2545 50050 -2425
rect 50170 -2545 50215 -2425
rect 50335 -2545 50380 -2425
rect 50500 -2545 50545 -2425
rect 50665 -2545 50720 -2425
rect 50840 -2545 50885 -2425
rect 51005 -2545 51050 -2425
rect 51170 -2545 51215 -2425
rect 51335 -2545 51390 -2425
rect 51510 -2545 51555 -2425
rect 51675 -2545 51720 -2425
rect 51840 -2545 51885 -2425
rect 52005 -2545 52060 -2425
rect 52180 -2545 52225 -2425
rect 52345 -2545 52390 -2425
rect 52510 -2545 52555 -2425
rect 52675 -2545 52730 -2425
rect 52850 -2545 52895 -2425
rect 53015 -2545 53060 -2425
rect 53180 -2545 53225 -2425
rect 53345 -2545 53355 -2425
rect 47855 -2600 53355 -2545
rect 47855 -2720 47865 -2600
rect 47985 -2720 48040 -2600
rect 48160 -2720 48205 -2600
rect 48325 -2720 48370 -2600
rect 48490 -2720 48535 -2600
rect 48655 -2720 48710 -2600
rect 48830 -2720 48875 -2600
rect 48995 -2720 49040 -2600
rect 49160 -2720 49205 -2600
rect 49325 -2720 49380 -2600
rect 49500 -2720 49545 -2600
rect 49665 -2720 49710 -2600
rect 49830 -2720 49875 -2600
rect 49995 -2720 50050 -2600
rect 50170 -2720 50215 -2600
rect 50335 -2720 50380 -2600
rect 50500 -2720 50545 -2600
rect 50665 -2720 50720 -2600
rect 50840 -2720 50885 -2600
rect 51005 -2720 51050 -2600
rect 51170 -2720 51215 -2600
rect 51335 -2720 51390 -2600
rect 51510 -2720 51555 -2600
rect 51675 -2720 51720 -2600
rect 51840 -2720 51885 -2600
rect 52005 -2720 52060 -2600
rect 52180 -2720 52225 -2600
rect 52345 -2720 52390 -2600
rect 52510 -2720 52555 -2600
rect 52675 -2720 52730 -2600
rect 52850 -2720 52895 -2600
rect 53015 -2720 53060 -2600
rect 53180 -2720 53225 -2600
rect 53345 -2720 53355 -2600
rect 47855 -2765 53355 -2720
rect 47855 -2885 47865 -2765
rect 47985 -2885 48040 -2765
rect 48160 -2885 48205 -2765
rect 48325 -2885 48370 -2765
rect 48490 -2885 48535 -2765
rect 48655 -2885 48710 -2765
rect 48830 -2885 48875 -2765
rect 48995 -2885 49040 -2765
rect 49160 -2885 49205 -2765
rect 49325 -2885 49380 -2765
rect 49500 -2885 49545 -2765
rect 49665 -2885 49710 -2765
rect 49830 -2885 49875 -2765
rect 49995 -2885 50050 -2765
rect 50170 -2885 50215 -2765
rect 50335 -2885 50380 -2765
rect 50500 -2885 50545 -2765
rect 50665 -2885 50720 -2765
rect 50840 -2885 50885 -2765
rect 51005 -2885 51050 -2765
rect 51170 -2885 51215 -2765
rect 51335 -2885 51390 -2765
rect 51510 -2885 51555 -2765
rect 51675 -2885 51720 -2765
rect 51840 -2885 51885 -2765
rect 52005 -2885 52060 -2765
rect 52180 -2885 52225 -2765
rect 52345 -2885 52390 -2765
rect 52510 -2885 52555 -2765
rect 52675 -2885 52730 -2765
rect 52850 -2885 52895 -2765
rect 53015 -2885 53060 -2765
rect 53180 -2885 53225 -2765
rect 53345 -2885 53355 -2765
rect 47855 -2930 53355 -2885
rect 47855 -3050 47865 -2930
rect 47985 -3050 48040 -2930
rect 48160 -3050 48205 -2930
rect 48325 -3050 48370 -2930
rect 48490 -3050 48535 -2930
rect 48655 -3050 48710 -2930
rect 48830 -3050 48875 -2930
rect 48995 -3050 49040 -2930
rect 49160 -3050 49205 -2930
rect 49325 -3050 49380 -2930
rect 49500 -3050 49545 -2930
rect 49665 -3050 49710 -2930
rect 49830 -3050 49875 -2930
rect 49995 -3050 50050 -2930
rect 50170 -3050 50215 -2930
rect 50335 -3050 50380 -2930
rect 50500 -3050 50545 -2930
rect 50665 -3050 50720 -2930
rect 50840 -3050 50885 -2930
rect 51005 -3050 51050 -2930
rect 51170 -3050 51215 -2930
rect 51335 -3050 51390 -2930
rect 51510 -3050 51555 -2930
rect 51675 -3050 51720 -2930
rect 51840 -3050 51885 -2930
rect 52005 -3050 52060 -2930
rect 52180 -3050 52225 -2930
rect 52345 -3050 52390 -2930
rect 52510 -3050 52555 -2930
rect 52675 -3050 52730 -2930
rect 52850 -3050 52895 -2930
rect 53015 -3050 53060 -2930
rect 53180 -3050 53225 -2930
rect 53345 -3050 53355 -2930
rect 47855 -3095 53355 -3050
rect 47855 -3215 47865 -3095
rect 47985 -3215 48040 -3095
rect 48160 -3215 48205 -3095
rect 48325 -3215 48370 -3095
rect 48490 -3215 48535 -3095
rect 48655 -3215 48710 -3095
rect 48830 -3215 48875 -3095
rect 48995 -3215 49040 -3095
rect 49160 -3215 49205 -3095
rect 49325 -3215 49380 -3095
rect 49500 -3215 49545 -3095
rect 49665 -3215 49710 -3095
rect 49830 -3215 49875 -3095
rect 49995 -3215 50050 -3095
rect 50170 -3215 50215 -3095
rect 50335 -3215 50380 -3095
rect 50500 -3215 50545 -3095
rect 50665 -3215 50720 -3095
rect 50840 -3215 50885 -3095
rect 51005 -3215 51050 -3095
rect 51170 -3215 51215 -3095
rect 51335 -3215 51390 -3095
rect 51510 -3215 51555 -3095
rect 51675 -3215 51720 -3095
rect 51840 -3215 51885 -3095
rect 52005 -3215 52060 -3095
rect 52180 -3215 52225 -3095
rect 52345 -3215 52390 -3095
rect 52510 -3215 52555 -3095
rect 52675 -3215 52730 -3095
rect 52850 -3215 52895 -3095
rect 53015 -3215 53060 -3095
rect 53180 -3215 53225 -3095
rect 53345 -3215 53355 -3095
rect 47855 -3270 53355 -3215
rect 47855 -3390 47865 -3270
rect 47985 -3390 48040 -3270
rect 48160 -3390 48205 -3270
rect 48325 -3390 48370 -3270
rect 48490 -3390 48535 -3270
rect 48655 -3390 48710 -3270
rect 48830 -3390 48875 -3270
rect 48995 -3390 49040 -3270
rect 49160 -3390 49205 -3270
rect 49325 -3390 49380 -3270
rect 49500 -3390 49545 -3270
rect 49665 -3390 49710 -3270
rect 49830 -3390 49875 -3270
rect 49995 -3390 50050 -3270
rect 50170 -3390 50215 -3270
rect 50335 -3390 50380 -3270
rect 50500 -3390 50545 -3270
rect 50665 -3390 50720 -3270
rect 50840 -3390 50885 -3270
rect 51005 -3390 51050 -3270
rect 51170 -3390 51215 -3270
rect 51335 -3390 51390 -3270
rect 51510 -3390 51555 -3270
rect 51675 -3390 51720 -3270
rect 51840 -3390 51885 -3270
rect 52005 -3390 52060 -3270
rect 52180 -3390 52225 -3270
rect 52345 -3390 52390 -3270
rect 52510 -3390 52555 -3270
rect 52675 -3390 52730 -3270
rect 52850 -3390 52895 -3270
rect 53015 -3390 53060 -3270
rect 53180 -3390 53225 -3270
rect 53345 -3390 53355 -3270
rect 47855 -3435 53355 -3390
rect 47855 -3555 47865 -3435
rect 47985 -3555 48040 -3435
rect 48160 -3555 48205 -3435
rect 48325 -3555 48370 -3435
rect 48490 -3555 48535 -3435
rect 48655 -3555 48710 -3435
rect 48830 -3555 48875 -3435
rect 48995 -3555 49040 -3435
rect 49160 -3555 49205 -3435
rect 49325 -3555 49380 -3435
rect 49500 -3555 49545 -3435
rect 49665 -3555 49710 -3435
rect 49830 -3555 49875 -3435
rect 49995 -3555 50050 -3435
rect 50170 -3555 50215 -3435
rect 50335 -3555 50380 -3435
rect 50500 -3555 50545 -3435
rect 50665 -3555 50720 -3435
rect 50840 -3555 50885 -3435
rect 51005 -3555 51050 -3435
rect 51170 -3555 51215 -3435
rect 51335 -3555 51390 -3435
rect 51510 -3555 51555 -3435
rect 51675 -3555 51720 -3435
rect 51840 -3555 51885 -3435
rect 52005 -3555 52060 -3435
rect 52180 -3555 52225 -3435
rect 52345 -3555 52390 -3435
rect 52510 -3555 52555 -3435
rect 52675 -3555 52730 -3435
rect 52850 -3555 52895 -3435
rect 53015 -3555 53060 -3435
rect 53180 -3555 53225 -3435
rect 53345 -3555 53355 -3435
rect 47855 -3600 53355 -3555
rect 47855 -3720 47865 -3600
rect 47985 -3720 48040 -3600
rect 48160 -3720 48205 -3600
rect 48325 -3720 48370 -3600
rect 48490 -3720 48535 -3600
rect 48655 -3720 48710 -3600
rect 48830 -3720 48875 -3600
rect 48995 -3720 49040 -3600
rect 49160 -3720 49205 -3600
rect 49325 -3720 49380 -3600
rect 49500 -3720 49545 -3600
rect 49665 -3720 49710 -3600
rect 49830 -3720 49875 -3600
rect 49995 -3720 50050 -3600
rect 50170 -3720 50215 -3600
rect 50335 -3720 50380 -3600
rect 50500 -3720 50545 -3600
rect 50665 -3720 50720 -3600
rect 50840 -3720 50885 -3600
rect 51005 -3720 51050 -3600
rect 51170 -3720 51215 -3600
rect 51335 -3720 51390 -3600
rect 51510 -3720 51555 -3600
rect 51675 -3720 51720 -3600
rect 51840 -3720 51885 -3600
rect 52005 -3720 52060 -3600
rect 52180 -3720 52225 -3600
rect 52345 -3720 52390 -3600
rect 52510 -3720 52555 -3600
rect 52675 -3720 52730 -3600
rect 52850 -3720 52895 -3600
rect 53015 -3720 53060 -3600
rect 53180 -3720 53225 -3600
rect 53345 -3720 53355 -3600
rect 47855 -3765 53355 -3720
rect 47855 -3885 47865 -3765
rect 47985 -3885 48040 -3765
rect 48160 -3885 48205 -3765
rect 48325 -3885 48370 -3765
rect 48490 -3885 48535 -3765
rect 48655 -3885 48710 -3765
rect 48830 -3885 48875 -3765
rect 48995 -3885 49040 -3765
rect 49160 -3885 49205 -3765
rect 49325 -3885 49380 -3765
rect 49500 -3885 49545 -3765
rect 49665 -3885 49710 -3765
rect 49830 -3885 49875 -3765
rect 49995 -3885 50050 -3765
rect 50170 -3885 50215 -3765
rect 50335 -3885 50380 -3765
rect 50500 -3885 50545 -3765
rect 50665 -3885 50720 -3765
rect 50840 -3885 50885 -3765
rect 51005 -3885 51050 -3765
rect 51170 -3885 51215 -3765
rect 51335 -3885 51390 -3765
rect 51510 -3885 51555 -3765
rect 51675 -3885 51720 -3765
rect 51840 -3885 51885 -3765
rect 52005 -3885 52060 -3765
rect 52180 -3885 52225 -3765
rect 52345 -3885 52390 -3765
rect 52510 -3885 52555 -3765
rect 52675 -3885 52730 -3765
rect 52850 -3885 52895 -3765
rect 53015 -3885 53060 -3765
rect 53180 -3885 53225 -3765
rect 53345 -3885 53355 -3765
rect 47855 -3940 53355 -3885
rect 47855 -4060 47865 -3940
rect 47985 -4060 48040 -3940
rect 48160 -4060 48205 -3940
rect 48325 -4060 48370 -3940
rect 48490 -4060 48535 -3940
rect 48655 -4060 48710 -3940
rect 48830 -4060 48875 -3940
rect 48995 -4060 49040 -3940
rect 49160 -4060 49205 -3940
rect 49325 -4060 49380 -3940
rect 49500 -4060 49545 -3940
rect 49665 -4060 49710 -3940
rect 49830 -4060 49875 -3940
rect 49995 -4060 50050 -3940
rect 50170 -4060 50215 -3940
rect 50335 -4060 50380 -3940
rect 50500 -4060 50545 -3940
rect 50665 -4060 50720 -3940
rect 50840 -4060 50885 -3940
rect 51005 -4060 51050 -3940
rect 51170 -4060 51215 -3940
rect 51335 -4060 51390 -3940
rect 51510 -4060 51555 -3940
rect 51675 -4060 51720 -3940
rect 51840 -4060 51885 -3940
rect 52005 -4060 52060 -3940
rect 52180 -4060 52225 -3940
rect 52345 -4060 52390 -3940
rect 52510 -4060 52555 -3940
rect 52675 -4060 52730 -3940
rect 52850 -4060 52895 -3940
rect 53015 -4060 53060 -3940
rect 53180 -4060 53225 -3940
rect 53345 -4060 53355 -3940
rect 47855 -4070 53355 -4060
rect 30785 -4270 36285 -4260
rect 30785 -4390 30795 -4270
rect 30915 -4390 30960 -4270
rect 31080 -4390 31125 -4270
rect 31245 -4390 31290 -4270
rect 31410 -4390 31465 -4270
rect 31585 -4390 31630 -4270
rect 31750 -4390 31795 -4270
rect 31915 -4390 31960 -4270
rect 32080 -4390 32135 -4270
rect 32255 -4390 32300 -4270
rect 32420 -4390 32465 -4270
rect 32585 -4390 32630 -4270
rect 32750 -4390 32805 -4270
rect 32925 -4390 32970 -4270
rect 33090 -4390 33135 -4270
rect 33255 -4390 33300 -4270
rect 33420 -4390 33475 -4270
rect 33595 -4390 33640 -4270
rect 33760 -4390 33805 -4270
rect 33925 -4390 33970 -4270
rect 34090 -4390 34145 -4270
rect 34265 -4390 34310 -4270
rect 34430 -4390 34475 -4270
rect 34595 -4390 34640 -4270
rect 34760 -4390 34815 -4270
rect 34935 -4390 34980 -4270
rect 35100 -4390 35145 -4270
rect 35265 -4390 35310 -4270
rect 35430 -4390 35485 -4270
rect 35605 -4390 35650 -4270
rect 35770 -4390 35815 -4270
rect 35935 -4390 35980 -4270
rect 36100 -4390 36155 -4270
rect 36275 -4390 36285 -4270
rect 30785 -4445 36285 -4390
rect 30785 -4565 30795 -4445
rect 30915 -4565 30960 -4445
rect 31080 -4565 31125 -4445
rect 31245 -4565 31290 -4445
rect 31410 -4565 31465 -4445
rect 31585 -4565 31630 -4445
rect 31750 -4565 31795 -4445
rect 31915 -4565 31960 -4445
rect 32080 -4565 32135 -4445
rect 32255 -4565 32300 -4445
rect 32420 -4565 32465 -4445
rect 32585 -4565 32630 -4445
rect 32750 -4565 32805 -4445
rect 32925 -4565 32970 -4445
rect 33090 -4565 33135 -4445
rect 33255 -4565 33300 -4445
rect 33420 -4565 33475 -4445
rect 33595 -4565 33640 -4445
rect 33760 -4565 33805 -4445
rect 33925 -4565 33970 -4445
rect 34090 -4565 34145 -4445
rect 34265 -4565 34310 -4445
rect 34430 -4565 34475 -4445
rect 34595 -4565 34640 -4445
rect 34760 -4565 34815 -4445
rect 34935 -4565 34980 -4445
rect 35100 -4565 35145 -4445
rect 35265 -4565 35310 -4445
rect 35430 -4565 35485 -4445
rect 35605 -4565 35650 -4445
rect 35770 -4565 35815 -4445
rect 35935 -4565 35980 -4445
rect 36100 -4565 36155 -4445
rect 36275 -4565 36285 -4445
rect 30785 -4610 36285 -4565
rect 30785 -4730 30795 -4610
rect 30915 -4730 30960 -4610
rect 31080 -4730 31125 -4610
rect 31245 -4730 31290 -4610
rect 31410 -4730 31465 -4610
rect 31585 -4730 31630 -4610
rect 31750 -4730 31795 -4610
rect 31915 -4730 31960 -4610
rect 32080 -4730 32135 -4610
rect 32255 -4730 32300 -4610
rect 32420 -4730 32465 -4610
rect 32585 -4730 32630 -4610
rect 32750 -4730 32805 -4610
rect 32925 -4730 32970 -4610
rect 33090 -4730 33135 -4610
rect 33255 -4730 33300 -4610
rect 33420 -4730 33475 -4610
rect 33595 -4730 33640 -4610
rect 33760 -4730 33805 -4610
rect 33925 -4730 33970 -4610
rect 34090 -4730 34145 -4610
rect 34265 -4730 34310 -4610
rect 34430 -4730 34475 -4610
rect 34595 -4730 34640 -4610
rect 34760 -4730 34815 -4610
rect 34935 -4730 34980 -4610
rect 35100 -4730 35145 -4610
rect 35265 -4730 35310 -4610
rect 35430 -4730 35485 -4610
rect 35605 -4730 35650 -4610
rect 35770 -4730 35815 -4610
rect 35935 -4730 35980 -4610
rect 36100 -4730 36155 -4610
rect 36275 -4730 36285 -4610
rect 30785 -4775 36285 -4730
rect 30785 -4895 30795 -4775
rect 30915 -4895 30960 -4775
rect 31080 -4895 31125 -4775
rect 31245 -4895 31290 -4775
rect 31410 -4895 31465 -4775
rect 31585 -4895 31630 -4775
rect 31750 -4895 31795 -4775
rect 31915 -4895 31960 -4775
rect 32080 -4895 32135 -4775
rect 32255 -4895 32300 -4775
rect 32420 -4895 32465 -4775
rect 32585 -4895 32630 -4775
rect 32750 -4895 32805 -4775
rect 32925 -4895 32970 -4775
rect 33090 -4895 33135 -4775
rect 33255 -4895 33300 -4775
rect 33420 -4895 33475 -4775
rect 33595 -4895 33640 -4775
rect 33760 -4895 33805 -4775
rect 33925 -4895 33970 -4775
rect 34090 -4895 34145 -4775
rect 34265 -4895 34310 -4775
rect 34430 -4895 34475 -4775
rect 34595 -4895 34640 -4775
rect 34760 -4895 34815 -4775
rect 34935 -4895 34980 -4775
rect 35100 -4895 35145 -4775
rect 35265 -4895 35310 -4775
rect 35430 -4895 35485 -4775
rect 35605 -4895 35650 -4775
rect 35770 -4895 35815 -4775
rect 35935 -4895 35980 -4775
rect 36100 -4895 36155 -4775
rect 36275 -4895 36285 -4775
rect 30785 -4940 36285 -4895
rect 30785 -5060 30795 -4940
rect 30915 -5060 30960 -4940
rect 31080 -5060 31125 -4940
rect 31245 -5060 31290 -4940
rect 31410 -5060 31465 -4940
rect 31585 -5060 31630 -4940
rect 31750 -5060 31795 -4940
rect 31915 -5060 31960 -4940
rect 32080 -5060 32135 -4940
rect 32255 -5060 32300 -4940
rect 32420 -5060 32465 -4940
rect 32585 -5060 32630 -4940
rect 32750 -5060 32805 -4940
rect 32925 -5060 32970 -4940
rect 33090 -5060 33135 -4940
rect 33255 -5060 33300 -4940
rect 33420 -5060 33475 -4940
rect 33595 -5060 33640 -4940
rect 33760 -5060 33805 -4940
rect 33925 -5060 33970 -4940
rect 34090 -5060 34145 -4940
rect 34265 -5060 34310 -4940
rect 34430 -5060 34475 -4940
rect 34595 -5060 34640 -4940
rect 34760 -5060 34815 -4940
rect 34935 -5060 34980 -4940
rect 35100 -5060 35145 -4940
rect 35265 -5060 35310 -4940
rect 35430 -5060 35485 -4940
rect 35605 -5060 35650 -4940
rect 35770 -5060 35815 -4940
rect 35935 -5060 35980 -4940
rect 36100 -5060 36155 -4940
rect 36275 -5060 36285 -4940
rect 30785 -5115 36285 -5060
rect 30785 -5235 30795 -5115
rect 30915 -5235 30960 -5115
rect 31080 -5235 31125 -5115
rect 31245 -5235 31290 -5115
rect 31410 -5235 31465 -5115
rect 31585 -5235 31630 -5115
rect 31750 -5235 31795 -5115
rect 31915 -5235 31960 -5115
rect 32080 -5235 32135 -5115
rect 32255 -5235 32300 -5115
rect 32420 -5235 32465 -5115
rect 32585 -5235 32630 -5115
rect 32750 -5235 32805 -5115
rect 32925 -5235 32970 -5115
rect 33090 -5235 33135 -5115
rect 33255 -5235 33300 -5115
rect 33420 -5235 33475 -5115
rect 33595 -5235 33640 -5115
rect 33760 -5235 33805 -5115
rect 33925 -5235 33970 -5115
rect 34090 -5235 34145 -5115
rect 34265 -5235 34310 -5115
rect 34430 -5235 34475 -5115
rect 34595 -5235 34640 -5115
rect 34760 -5235 34815 -5115
rect 34935 -5235 34980 -5115
rect 35100 -5235 35145 -5115
rect 35265 -5235 35310 -5115
rect 35430 -5235 35485 -5115
rect 35605 -5235 35650 -5115
rect 35770 -5235 35815 -5115
rect 35935 -5235 35980 -5115
rect 36100 -5235 36155 -5115
rect 36275 -5235 36285 -5115
rect 30785 -5280 36285 -5235
rect 30785 -5400 30795 -5280
rect 30915 -5400 30960 -5280
rect 31080 -5400 31125 -5280
rect 31245 -5400 31290 -5280
rect 31410 -5400 31465 -5280
rect 31585 -5400 31630 -5280
rect 31750 -5400 31795 -5280
rect 31915 -5400 31960 -5280
rect 32080 -5400 32135 -5280
rect 32255 -5400 32300 -5280
rect 32420 -5400 32465 -5280
rect 32585 -5400 32630 -5280
rect 32750 -5400 32805 -5280
rect 32925 -5400 32970 -5280
rect 33090 -5400 33135 -5280
rect 33255 -5400 33300 -5280
rect 33420 -5400 33475 -5280
rect 33595 -5400 33640 -5280
rect 33760 -5400 33805 -5280
rect 33925 -5400 33970 -5280
rect 34090 -5400 34145 -5280
rect 34265 -5400 34310 -5280
rect 34430 -5400 34475 -5280
rect 34595 -5400 34640 -5280
rect 34760 -5400 34815 -5280
rect 34935 -5400 34980 -5280
rect 35100 -5400 35145 -5280
rect 35265 -5400 35310 -5280
rect 35430 -5400 35485 -5280
rect 35605 -5400 35650 -5280
rect 35770 -5400 35815 -5280
rect 35935 -5400 35980 -5280
rect 36100 -5400 36155 -5280
rect 36275 -5400 36285 -5280
rect 30785 -5445 36285 -5400
rect 30785 -5565 30795 -5445
rect 30915 -5565 30960 -5445
rect 31080 -5565 31125 -5445
rect 31245 -5565 31290 -5445
rect 31410 -5565 31465 -5445
rect 31585 -5565 31630 -5445
rect 31750 -5565 31795 -5445
rect 31915 -5565 31960 -5445
rect 32080 -5565 32135 -5445
rect 32255 -5565 32300 -5445
rect 32420 -5565 32465 -5445
rect 32585 -5565 32630 -5445
rect 32750 -5565 32805 -5445
rect 32925 -5565 32970 -5445
rect 33090 -5565 33135 -5445
rect 33255 -5565 33300 -5445
rect 33420 -5565 33475 -5445
rect 33595 -5565 33640 -5445
rect 33760 -5565 33805 -5445
rect 33925 -5565 33970 -5445
rect 34090 -5565 34145 -5445
rect 34265 -5565 34310 -5445
rect 34430 -5565 34475 -5445
rect 34595 -5565 34640 -5445
rect 34760 -5565 34815 -5445
rect 34935 -5565 34980 -5445
rect 35100 -5565 35145 -5445
rect 35265 -5565 35310 -5445
rect 35430 -5565 35485 -5445
rect 35605 -5565 35650 -5445
rect 35770 -5565 35815 -5445
rect 35935 -5565 35980 -5445
rect 36100 -5565 36155 -5445
rect 36275 -5565 36285 -5445
rect 30785 -5610 36285 -5565
rect 30785 -5730 30795 -5610
rect 30915 -5730 30960 -5610
rect 31080 -5730 31125 -5610
rect 31245 -5730 31290 -5610
rect 31410 -5730 31465 -5610
rect 31585 -5730 31630 -5610
rect 31750 -5730 31795 -5610
rect 31915 -5730 31960 -5610
rect 32080 -5730 32135 -5610
rect 32255 -5730 32300 -5610
rect 32420 -5730 32465 -5610
rect 32585 -5730 32630 -5610
rect 32750 -5730 32805 -5610
rect 32925 -5730 32970 -5610
rect 33090 -5730 33135 -5610
rect 33255 -5730 33300 -5610
rect 33420 -5730 33475 -5610
rect 33595 -5730 33640 -5610
rect 33760 -5730 33805 -5610
rect 33925 -5730 33970 -5610
rect 34090 -5730 34145 -5610
rect 34265 -5730 34310 -5610
rect 34430 -5730 34475 -5610
rect 34595 -5730 34640 -5610
rect 34760 -5730 34815 -5610
rect 34935 -5730 34980 -5610
rect 35100 -5730 35145 -5610
rect 35265 -5730 35310 -5610
rect 35430 -5730 35485 -5610
rect 35605 -5730 35650 -5610
rect 35770 -5730 35815 -5610
rect 35935 -5730 35980 -5610
rect 36100 -5730 36155 -5610
rect 36275 -5730 36285 -5610
rect 30785 -5785 36285 -5730
rect 30785 -5905 30795 -5785
rect 30915 -5905 30960 -5785
rect 31080 -5905 31125 -5785
rect 31245 -5905 31290 -5785
rect 31410 -5905 31465 -5785
rect 31585 -5905 31630 -5785
rect 31750 -5905 31795 -5785
rect 31915 -5905 31960 -5785
rect 32080 -5905 32135 -5785
rect 32255 -5905 32300 -5785
rect 32420 -5905 32465 -5785
rect 32585 -5905 32630 -5785
rect 32750 -5905 32805 -5785
rect 32925 -5905 32970 -5785
rect 33090 -5905 33135 -5785
rect 33255 -5905 33300 -5785
rect 33420 -5905 33475 -5785
rect 33595 -5905 33640 -5785
rect 33760 -5905 33805 -5785
rect 33925 -5905 33970 -5785
rect 34090 -5905 34145 -5785
rect 34265 -5905 34310 -5785
rect 34430 -5905 34475 -5785
rect 34595 -5905 34640 -5785
rect 34760 -5905 34815 -5785
rect 34935 -5905 34980 -5785
rect 35100 -5905 35145 -5785
rect 35265 -5905 35310 -5785
rect 35430 -5905 35485 -5785
rect 35605 -5905 35650 -5785
rect 35770 -5905 35815 -5785
rect 35935 -5905 35980 -5785
rect 36100 -5905 36155 -5785
rect 36275 -5905 36285 -5785
rect 30785 -5950 36285 -5905
rect 30785 -6070 30795 -5950
rect 30915 -6070 30960 -5950
rect 31080 -6070 31125 -5950
rect 31245 -6070 31290 -5950
rect 31410 -6070 31465 -5950
rect 31585 -6070 31630 -5950
rect 31750 -6070 31795 -5950
rect 31915 -6070 31960 -5950
rect 32080 -6070 32135 -5950
rect 32255 -6070 32300 -5950
rect 32420 -6070 32465 -5950
rect 32585 -6070 32630 -5950
rect 32750 -6070 32805 -5950
rect 32925 -6070 32970 -5950
rect 33090 -6070 33135 -5950
rect 33255 -6070 33300 -5950
rect 33420 -6070 33475 -5950
rect 33595 -6070 33640 -5950
rect 33760 -6070 33805 -5950
rect 33925 -6070 33970 -5950
rect 34090 -6070 34145 -5950
rect 34265 -6070 34310 -5950
rect 34430 -6070 34475 -5950
rect 34595 -6070 34640 -5950
rect 34760 -6070 34815 -5950
rect 34935 -6070 34980 -5950
rect 35100 -6070 35145 -5950
rect 35265 -6070 35310 -5950
rect 35430 -6070 35485 -5950
rect 35605 -6070 35650 -5950
rect 35770 -6070 35815 -5950
rect 35935 -6070 35980 -5950
rect 36100 -6070 36155 -5950
rect 36275 -6070 36285 -5950
rect 30785 -6115 36285 -6070
rect 30785 -6235 30795 -6115
rect 30915 -6235 30960 -6115
rect 31080 -6235 31125 -6115
rect 31245 -6235 31290 -6115
rect 31410 -6235 31465 -6115
rect 31585 -6235 31630 -6115
rect 31750 -6235 31795 -6115
rect 31915 -6235 31960 -6115
rect 32080 -6235 32135 -6115
rect 32255 -6235 32300 -6115
rect 32420 -6235 32465 -6115
rect 32585 -6235 32630 -6115
rect 32750 -6235 32805 -6115
rect 32925 -6235 32970 -6115
rect 33090 -6235 33135 -6115
rect 33255 -6235 33300 -6115
rect 33420 -6235 33475 -6115
rect 33595 -6235 33640 -6115
rect 33760 -6235 33805 -6115
rect 33925 -6235 33970 -6115
rect 34090 -6235 34145 -6115
rect 34265 -6235 34310 -6115
rect 34430 -6235 34475 -6115
rect 34595 -6235 34640 -6115
rect 34760 -6235 34815 -6115
rect 34935 -6235 34980 -6115
rect 35100 -6235 35145 -6115
rect 35265 -6235 35310 -6115
rect 35430 -6235 35485 -6115
rect 35605 -6235 35650 -6115
rect 35770 -6235 35815 -6115
rect 35935 -6235 35980 -6115
rect 36100 -6235 36155 -6115
rect 36275 -6235 36285 -6115
rect 30785 -6280 36285 -6235
rect 30785 -6400 30795 -6280
rect 30915 -6400 30960 -6280
rect 31080 -6400 31125 -6280
rect 31245 -6400 31290 -6280
rect 31410 -6400 31465 -6280
rect 31585 -6400 31630 -6280
rect 31750 -6400 31795 -6280
rect 31915 -6400 31960 -6280
rect 32080 -6400 32135 -6280
rect 32255 -6400 32300 -6280
rect 32420 -6400 32465 -6280
rect 32585 -6400 32630 -6280
rect 32750 -6400 32805 -6280
rect 32925 -6400 32970 -6280
rect 33090 -6400 33135 -6280
rect 33255 -6400 33300 -6280
rect 33420 -6400 33475 -6280
rect 33595 -6400 33640 -6280
rect 33760 -6400 33805 -6280
rect 33925 -6400 33970 -6280
rect 34090 -6400 34145 -6280
rect 34265 -6400 34310 -6280
rect 34430 -6400 34475 -6280
rect 34595 -6400 34640 -6280
rect 34760 -6400 34815 -6280
rect 34935 -6400 34980 -6280
rect 35100 -6400 35145 -6280
rect 35265 -6400 35310 -6280
rect 35430 -6400 35485 -6280
rect 35605 -6400 35650 -6280
rect 35770 -6400 35815 -6280
rect 35935 -6400 35980 -6280
rect 36100 -6400 36155 -6280
rect 36275 -6400 36285 -6280
rect 30785 -6455 36285 -6400
rect 30785 -6575 30795 -6455
rect 30915 -6575 30960 -6455
rect 31080 -6575 31125 -6455
rect 31245 -6575 31290 -6455
rect 31410 -6575 31465 -6455
rect 31585 -6575 31630 -6455
rect 31750 -6575 31795 -6455
rect 31915 -6575 31960 -6455
rect 32080 -6575 32135 -6455
rect 32255 -6575 32300 -6455
rect 32420 -6575 32465 -6455
rect 32585 -6575 32630 -6455
rect 32750 -6575 32805 -6455
rect 32925 -6575 32970 -6455
rect 33090 -6575 33135 -6455
rect 33255 -6575 33300 -6455
rect 33420 -6575 33475 -6455
rect 33595 -6575 33640 -6455
rect 33760 -6575 33805 -6455
rect 33925 -6575 33970 -6455
rect 34090 -6575 34145 -6455
rect 34265 -6575 34310 -6455
rect 34430 -6575 34475 -6455
rect 34595 -6575 34640 -6455
rect 34760 -6575 34815 -6455
rect 34935 -6575 34980 -6455
rect 35100 -6575 35145 -6455
rect 35265 -6575 35310 -6455
rect 35430 -6575 35485 -6455
rect 35605 -6575 35650 -6455
rect 35770 -6575 35815 -6455
rect 35935 -6575 35980 -6455
rect 36100 -6575 36155 -6455
rect 36275 -6575 36285 -6455
rect 30785 -6620 36285 -6575
rect 30785 -6740 30795 -6620
rect 30915 -6740 30960 -6620
rect 31080 -6740 31125 -6620
rect 31245 -6740 31290 -6620
rect 31410 -6740 31465 -6620
rect 31585 -6740 31630 -6620
rect 31750 -6740 31795 -6620
rect 31915 -6740 31960 -6620
rect 32080 -6740 32135 -6620
rect 32255 -6740 32300 -6620
rect 32420 -6740 32465 -6620
rect 32585 -6740 32630 -6620
rect 32750 -6740 32805 -6620
rect 32925 -6740 32970 -6620
rect 33090 -6740 33135 -6620
rect 33255 -6740 33300 -6620
rect 33420 -6740 33475 -6620
rect 33595 -6740 33640 -6620
rect 33760 -6740 33805 -6620
rect 33925 -6740 33970 -6620
rect 34090 -6740 34145 -6620
rect 34265 -6740 34310 -6620
rect 34430 -6740 34475 -6620
rect 34595 -6740 34640 -6620
rect 34760 -6740 34815 -6620
rect 34935 -6740 34980 -6620
rect 35100 -6740 35145 -6620
rect 35265 -6740 35310 -6620
rect 35430 -6740 35485 -6620
rect 35605 -6740 35650 -6620
rect 35770 -6740 35815 -6620
rect 35935 -6740 35980 -6620
rect 36100 -6740 36155 -6620
rect 36275 -6740 36285 -6620
rect 30785 -6785 36285 -6740
rect 30785 -6905 30795 -6785
rect 30915 -6905 30960 -6785
rect 31080 -6905 31125 -6785
rect 31245 -6905 31290 -6785
rect 31410 -6905 31465 -6785
rect 31585 -6905 31630 -6785
rect 31750 -6905 31795 -6785
rect 31915 -6905 31960 -6785
rect 32080 -6905 32135 -6785
rect 32255 -6905 32300 -6785
rect 32420 -6905 32465 -6785
rect 32585 -6905 32630 -6785
rect 32750 -6905 32805 -6785
rect 32925 -6905 32970 -6785
rect 33090 -6905 33135 -6785
rect 33255 -6905 33300 -6785
rect 33420 -6905 33475 -6785
rect 33595 -6905 33640 -6785
rect 33760 -6905 33805 -6785
rect 33925 -6905 33970 -6785
rect 34090 -6905 34145 -6785
rect 34265 -6905 34310 -6785
rect 34430 -6905 34475 -6785
rect 34595 -6905 34640 -6785
rect 34760 -6905 34815 -6785
rect 34935 -6905 34980 -6785
rect 35100 -6905 35145 -6785
rect 35265 -6905 35310 -6785
rect 35430 -6905 35485 -6785
rect 35605 -6905 35650 -6785
rect 35770 -6905 35815 -6785
rect 35935 -6905 35980 -6785
rect 36100 -6905 36155 -6785
rect 36275 -6905 36285 -6785
rect 30785 -6950 36285 -6905
rect 30785 -7070 30795 -6950
rect 30915 -7070 30960 -6950
rect 31080 -7070 31125 -6950
rect 31245 -7070 31290 -6950
rect 31410 -7070 31465 -6950
rect 31585 -7070 31630 -6950
rect 31750 -7070 31795 -6950
rect 31915 -7070 31960 -6950
rect 32080 -7070 32135 -6950
rect 32255 -7070 32300 -6950
rect 32420 -7070 32465 -6950
rect 32585 -7070 32630 -6950
rect 32750 -7070 32805 -6950
rect 32925 -7070 32970 -6950
rect 33090 -7070 33135 -6950
rect 33255 -7070 33300 -6950
rect 33420 -7070 33475 -6950
rect 33595 -7070 33640 -6950
rect 33760 -7070 33805 -6950
rect 33925 -7070 33970 -6950
rect 34090 -7070 34145 -6950
rect 34265 -7070 34310 -6950
rect 34430 -7070 34475 -6950
rect 34595 -7070 34640 -6950
rect 34760 -7070 34815 -6950
rect 34935 -7070 34980 -6950
rect 35100 -7070 35145 -6950
rect 35265 -7070 35310 -6950
rect 35430 -7070 35485 -6950
rect 35605 -7070 35650 -6950
rect 35770 -7070 35815 -6950
rect 35935 -7070 35980 -6950
rect 36100 -7070 36155 -6950
rect 36275 -7070 36285 -6950
rect 30785 -7125 36285 -7070
rect 30785 -7245 30795 -7125
rect 30915 -7245 30960 -7125
rect 31080 -7245 31125 -7125
rect 31245 -7245 31290 -7125
rect 31410 -7245 31465 -7125
rect 31585 -7245 31630 -7125
rect 31750 -7245 31795 -7125
rect 31915 -7245 31960 -7125
rect 32080 -7245 32135 -7125
rect 32255 -7245 32300 -7125
rect 32420 -7245 32465 -7125
rect 32585 -7245 32630 -7125
rect 32750 -7245 32805 -7125
rect 32925 -7245 32970 -7125
rect 33090 -7245 33135 -7125
rect 33255 -7245 33300 -7125
rect 33420 -7245 33475 -7125
rect 33595 -7245 33640 -7125
rect 33760 -7245 33805 -7125
rect 33925 -7245 33970 -7125
rect 34090 -7245 34145 -7125
rect 34265 -7245 34310 -7125
rect 34430 -7245 34475 -7125
rect 34595 -7245 34640 -7125
rect 34760 -7245 34815 -7125
rect 34935 -7245 34980 -7125
rect 35100 -7245 35145 -7125
rect 35265 -7245 35310 -7125
rect 35430 -7245 35485 -7125
rect 35605 -7245 35650 -7125
rect 35770 -7245 35815 -7125
rect 35935 -7245 35980 -7125
rect 36100 -7245 36155 -7125
rect 36275 -7245 36285 -7125
rect 30785 -7290 36285 -7245
rect 30785 -7410 30795 -7290
rect 30915 -7410 30960 -7290
rect 31080 -7410 31125 -7290
rect 31245 -7410 31290 -7290
rect 31410 -7410 31465 -7290
rect 31585 -7410 31630 -7290
rect 31750 -7410 31795 -7290
rect 31915 -7410 31960 -7290
rect 32080 -7410 32135 -7290
rect 32255 -7410 32300 -7290
rect 32420 -7410 32465 -7290
rect 32585 -7410 32630 -7290
rect 32750 -7410 32805 -7290
rect 32925 -7410 32970 -7290
rect 33090 -7410 33135 -7290
rect 33255 -7410 33300 -7290
rect 33420 -7410 33475 -7290
rect 33595 -7410 33640 -7290
rect 33760 -7410 33805 -7290
rect 33925 -7410 33970 -7290
rect 34090 -7410 34145 -7290
rect 34265 -7410 34310 -7290
rect 34430 -7410 34475 -7290
rect 34595 -7410 34640 -7290
rect 34760 -7410 34815 -7290
rect 34935 -7410 34980 -7290
rect 35100 -7410 35145 -7290
rect 35265 -7410 35310 -7290
rect 35430 -7410 35485 -7290
rect 35605 -7410 35650 -7290
rect 35770 -7410 35815 -7290
rect 35935 -7410 35980 -7290
rect 36100 -7410 36155 -7290
rect 36275 -7410 36285 -7290
rect 30785 -7455 36285 -7410
rect 30785 -7575 30795 -7455
rect 30915 -7575 30960 -7455
rect 31080 -7575 31125 -7455
rect 31245 -7575 31290 -7455
rect 31410 -7575 31465 -7455
rect 31585 -7575 31630 -7455
rect 31750 -7575 31795 -7455
rect 31915 -7575 31960 -7455
rect 32080 -7575 32135 -7455
rect 32255 -7575 32300 -7455
rect 32420 -7575 32465 -7455
rect 32585 -7575 32630 -7455
rect 32750 -7575 32805 -7455
rect 32925 -7575 32970 -7455
rect 33090 -7575 33135 -7455
rect 33255 -7575 33300 -7455
rect 33420 -7575 33475 -7455
rect 33595 -7575 33640 -7455
rect 33760 -7575 33805 -7455
rect 33925 -7575 33970 -7455
rect 34090 -7575 34145 -7455
rect 34265 -7575 34310 -7455
rect 34430 -7575 34475 -7455
rect 34595 -7575 34640 -7455
rect 34760 -7575 34815 -7455
rect 34935 -7575 34980 -7455
rect 35100 -7575 35145 -7455
rect 35265 -7575 35310 -7455
rect 35430 -7575 35485 -7455
rect 35605 -7575 35650 -7455
rect 35770 -7575 35815 -7455
rect 35935 -7575 35980 -7455
rect 36100 -7575 36155 -7455
rect 36275 -7575 36285 -7455
rect 30785 -7620 36285 -7575
rect 30785 -7740 30795 -7620
rect 30915 -7740 30960 -7620
rect 31080 -7740 31125 -7620
rect 31245 -7740 31290 -7620
rect 31410 -7740 31465 -7620
rect 31585 -7740 31630 -7620
rect 31750 -7740 31795 -7620
rect 31915 -7740 31960 -7620
rect 32080 -7740 32135 -7620
rect 32255 -7740 32300 -7620
rect 32420 -7740 32465 -7620
rect 32585 -7740 32630 -7620
rect 32750 -7740 32805 -7620
rect 32925 -7740 32970 -7620
rect 33090 -7740 33135 -7620
rect 33255 -7740 33300 -7620
rect 33420 -7740 33475 -7620
rect 33595 -7740 33640 -7620
rect 33760 -7740 33805 -7620
rect 33925 -7740 33970 -7620
rect 34090 -7740 34145 -7620
rect 34265 -7740 34310 -7620
rect 34430 -7740 34475 -7620
rect 34595 -7740 34640 -7620
rect 34760 -7740 34815 -7620
rect 34935 -7740 34980 -7620
rect 35100 -7740 35145 -7620
rect 35265 -7740 35310 -7620
rect 35430 -7740 35485 -7620
rect 35605 -7740 35650 -7620
rect 35770 -7740 35815 -7620
rect 35935 -7740 35980 -7620
rect 36100 -7740 36155 -7620
rect 36275 -7740 36285 -7620
rect 30785 -7795 36285 -7740
rect 30785 -7915 30795 -7795
rect 30915 -7915 30960 -7795
rect 31080 -7915 31125 -7795
rect 31245 -7915 31290 -7795
rect 31410 -7915 31465 -7795
rect 31585 -7915 31630 -7795
rect 31750 -7915 31795 -7795
rect 31915 -7915 31960 -7795
rect 32080 -7915 32135 -7795
rect 32255 -7915 32300 -7795
rect 32420 -7915 32465 -7795
rect 32585 -7915 32630 -7795
rect 32750 -7915 32805 -7795
rect 32925 -7915 32970 -7795
rect 33090 -7915 33135 -7795
rect 33255 -7915 33300 -7795
rect 33420 -7915 33475 -7795
rect 33595 -7915 33640 -7795
rect 33760 -7915 33805 -7795
rect 33925 -7915 33970 -7795
rect 34090 -7915 34145 -7795
rect 34265 -7915 34310 -7795
rect 34430 -7915 34475 -7795
rect 34595 -7915 34640 -7795
rect 34760 -7915 34815 -7795
rect 34935 -7915 34980 -7795
rect 35100 -7915 35145 -7795
rect 35265 -7915 35310 -7795
rect 35430 -7915 35485 -7795
rect 35605 -7915 35650 -7795
rect 35770 -7915 35815 -7795
rect 35935 -7915 35980 -7795
rect 36100 -7915 36155 -7795
rect 36275 -7915 36285 -7795
rect 30785 -7960 36285 -7915
rect 30785 -8080 30795 -7960
rect 30915 -8080 30960 -7960
rect 31080 -8080 31125 -7960
rect 31245 -8080 31290 -7960
rect 31410 -8080 31465 -7960
rect 31585 -8080 31630 -7960
rect 31750 -8080 31795 -7960
rect 31915 -8080 31960 -7960
rect 32080 -8080 32135 -7960
rect 32255 -8080 32300 -7960
rect 32420 -8080 32465 -7960
rect 32585 -8080 32630 -7960
rect 32750 -8080 32805 -7960
rect 32925 -8080 32970 -7960
rect 33090 -8080 33135 -7960
rect 33255 -8080 33300 -7960
rect 33420 -8080 33475 -7960
rect 33595 -8080 33640 -7960
rect 33760 -8080 33805 -7960
rect 33925 -8080 33970 -7960
rect 34090 -8080 34145 -7960
rect 34265 -8080 34310 -7960
rect 34430 -8080 34475 -7960
rect 34595 -8080 34640 -7960
rect 34760 -8080 34815 -7960
rect 34935 -8080 34980 -7960
rect 35100 -8080 35145 -7960
rect 35265 -8080 35310 -7960
rect 35430 -8080 35485 -7960
rect 35605 -8080 35650 -7960
rect 35770 -8080 35815 -7960
rect 35935 -8080 35980 -7960
rect 36100 -8080 36155 -7960
rect 36275 -8080 36285 -7960
rect 30785 -8125 36285 -8080
rect 30785 -8245 30795 -8125
rect 30915 -8245 30960 -8125
rect 31080 -8245 31125 -8125
rect 31245 -8245 31290 -8125
rect 31410 -8245 31465 -8125
rect 31585 -8245 31630 -8125
rect 31750 -8245 31795 -8125
rect 31915 -8245 31960 -8125
rect 32080 -8245 32135 -8125
rect 32255 -8245 32300 -8125
rect 32420 -8245 32465 -8125
rect 32585 -8245 32630 -8125
rect 32750 -8245 32805 -8125
rect 32925 -8245 32970 -8125
rect 33090 -8245 33135 -8125
rect 33255 -8245 33300 -8125
rect 33420 -8245 33475 -8125
rect 33595 -8245 33640 -8125
rect 33760 -8245 33805 -8125
rect 33925 -8245 33970 -8125
rect 34090 -8245 34145 -8125
rect 34265 -8245 34310 -8125
rect 34430 -8245 34475 -8125
rect 34595 -8245 34640 -8125
rect 34760 -8245 34815 -8125
rect 34935 -8245 34980 -8125
rect 35100 -8245 35145 -8125
rect 35265 -8245 35310 -8125
rect 35430 -8245 35485 -8125
rect 35605 -8245 35650 -8125
rect 35770 -8245 35815 -8125
rect 35935 -8245 35980 -8125
rect 36100 -8245 36155 -8125
rect 36275 -8245 36285 -8125
rect 30785 -8290 36285 -8245
rect 30785 -8410 30795 -8290
rect 30915 -8410 30960 -8290
rect 31080 -8410 31125 -8290
rect 31245 -8410 31290 -8290
rect 31410 -8410 31465 -8290
rect 31585 -8410 31630 -8290
rect 31750 -8410 31795 -8290
rect 31915 -8410 31960 -8290
rect 32080 -8410 32135 -8290
rect 32255 -8410 32300 -8290
rect 32420 -8410 32465 -8290
rect 32585 -8410 32630 -8290
rect 32750 -8410 32805 -8290
rect 32925 -8410 32970 -8290
rect 33090 -8410 33135 -8290
rect 33255 -8410 33300 -8290
rect 33420 -8410 33475 -8290
rect 33595 -8410 33640 -8290
rect 33760 -8410 33805 -8290
rect 33925 -8410 33970 -8290
rect 34090 -8410 34145 -8290
rect 34265 -8410 34310 -8290
rect 34430 -8410 34475 -8290
rect 34595 -8410 34640 -8290
rect 34760 -8410 34815 -8290
rect 34935 -8410 34980 -8290
rect 35100 -8410 35145 -8290
rect 35265 -8410 35310 -8290
rect 35430 -8410 35485 -8290
rect 35605 -8410 35650 -8290
rect 35770 -8410 35815 -8290
rect 35935 -8410 35980 -8290
rect 36100 -8410 36155 -8290
rect 36275 -8410 36285 -8290
rect 30785 -8465 36285 -8410
rect 30785 -8585 30795 -8465
rect 30915 -8585 30960 -8465
rect 31080 -8585 31125 -8465
rect 31245 -8585 31290 -8465
rect 31410 -8585 31465 -8465
rect 31585 -8585 31630 -8465
rect 31750 -8585 31795 -8465
rect 31915 -8585 31960 -8465
rect 32080 -8585 32135 -8465
rect 32255 -8585 32300 -8465
rect 32420 -8585 32465 -8465
rect 32585 -8585 32630 -8465
rect 32750 -8585 32805 -8465
rect 32925 -8585 32970 -8465
rect 33090 -8585 33135 -8465
rect 33255 -8585 33300 -8465
rect 33420 -8585 33475 -8465
rect 33595 -8585 33640 -8465
rect 33760 -8585 33805 -8465
rect 33925 -8585 33970 -8465
rect 34090 -8585 34145 -8465
rect 34265 -8585 34310 -8465
rect 34430 -8585 34475 -8465
rect 34595 -8585 34640 -8465
rect 34760 -8585 34815 -8465
rect 34935 -8585 34980 -8465
rect 35100 -8585 35145 -8465
rect 35265 -8585 35310 -8465
rect 35430 -8585 35485 -8465
rect 35605 -8585 35650 -8465
rect 35770 -8585 35815 -8465
rect 35935 -8585 35980 -8465
rect 36100 -8585 36155 -8465
rect 36275 -8585 36285 -8465
rect 30785 -8630 36285 -8585
rect 30785 -8750 30795 -8630
rect 30915 -8750 30960 -8630
rect 31080 -8750 31125 -8630
rect 31245 -8750 31290 -8630
rect 31410 -8750 31465 -8630
rect 31585 -8750 31630 -8630
rect 31750 -8750 31795 -8630
rect 31915 -8750 31960 -8630
rect 32080 -8750 32135 -8630
rect 32255 -8750 32300 -8630
rect 32420 -8750 32465 -8630
rect 32585 -8750 32630 -8630
rect 32750 -8750 32805 -8630
rect 32925 -8750 32970 -8630
rect 33090 -8750 33135 -8630
rect 33255 -8750 33300 -8630
rect 33420 -8750 33475 -8630
rect 33595 -8750 33640 -8630
rect 33760 -8750 33805 -8630
rect 33925 -8750 33970 -8630
rect 34090 -8750 34145 -8630
rect 34265 -8750 34310 -8630
rect 34430 -8750 34475 -8630
rect 34595 -8750 34640 -8630
rect 34760 -8750 34815 -8630
rect 34935 -8750 34980 -8630
rect 35100 -8750 35145 -8630
rect 35265 -8750 35310 -8630
rect 35430 -8750 35485 -8630
rect 35605 -8750 35650 -8630
rect 35770 -8750 35815 -8630
rect 35935 -8750 35980 -8630
rect 36100 -8750 36155 -8630
rect 36275 -8750 36285 -8630
rect 30785 -8795 36285 -8750
rect 30785 -8915 30795 -8795
rect 30915 -8915 30960 -8795
rect 31080 -8915 31125 -8795
rect 31245 -8915 31290 -8795
rect 31410 -8915 31465 -8795
rect 31585 -8915 31630 -8795
rect 31750 -8915 31795 -8795
rect 31915 -8915 31960 -8795
rect 32080 -8915 32135 -8795
rect 32255 -8915 32300 -8795
rect 32420 -8915 32465 -8795
rect 32585 -8915 32630 -8795
rect 32750 -8915 32805 -8795
rect 32925 -8915 32970 -8795
rect 33090 -8915 33135 -8795
rect 33255 -8915 33300 -8795
rect 33420 -8915 33475 -8795
rect 33595 -8915 33640 -8795
rect 33760 -8915 33805 -8795
rect 33925 -8915 33970 -8795
rect 34090 -8915 34145 -8795
rect 34265 -8915 34310 -8795
rect 34430 -8915 34475 -8795
rect 34595 -8915 34640 -8795
rect 34760 -8915 34815 -8795
rect 34935 -8915 34980 -8795
rect 35100 -8915 35145 -8795
rect 35265 -8915 35310 -8795
rect 35430 -8915 35485 -8795
rect 35605 -8915 35650 -8795
rect 35770 -8915 35815 -8795
rect 35935 -8915 35980 -8795
rect 36100 -8915 36155 -8795
rect 36275 -8915 36285 -8795
rect 30785 -8960 36285 -8915
rect 30785 -9080 30795 -8960
rect 30915 -9080 30960 -8960
rect 31080 -9080 31125 -8960
rect 31245 -9080 31290 -8960
rect 31410 -9080 31465 -8960
rect 31585 -9080 31630 -8960
rect 31750 -9080 31795 -8960
rect 31915 -9080 31960 -8960
rect 32080 -9080 32135 -8960
rect 32255 -9080 32300 -8960
rect 32420 -9080 32465 -8960
rect 32585 -9080 32630 -8960
rect 32750 -9080 32805 -8960
rect 32925 -9080 32970 -8960
rect 33090 -9080 33135 -8960
rect 33255 -9080 33300 -8960
rect 33420 -9080 33475 -8960
rect 33595 -9080 33640 -8960
rect 33760 -9080 33805 -8960
rect 33925 -9080 33970 -8960
rect 34090 -9080 34145 -8960
rect 34265 -9080 34310 -8960
rect 34430 -9080 34475 -8960
rect 34595 -9080 34640 -8960
rect 34760 -9080 34815 -8960
rect 34935 -9080 34980 -8960
rect 35100 -9080 35145 -8960
rect 35265 -9080 35310 -8960
rect 35430 -9080 35485 -8960
rect 35605 -9080 35650 -8960
rect 35770 -9080 35815 -8960
rect 35935 -9080 35980 -8960
rect 36100 -9080 36155 -8960
rect 36275 -9080 36285 -8960
rect 30785 -9135 36285 -9080
rect 30785 -9255 30795 -9135
rect 30915 -9255 30960 -9135
rect 31080 -9255 31125 -9135
rect 31245 -9255 31290 -9135
rect 31410 -9255 31465 -9135
rect 31585 -9255 31630 -9135
rect 31750 -9255 31795 -9135
rect 31915 -9255 31960 -9135
rect 32080 -9255 32135 -9135
rect 32255 -9255 32300 -9135
rect 32420 -9255 32465 -9135
rect 32585 -9255 32630 -9135
rect 32750 -9255 32805 -9135
rect 32925 -9255 32970 -9135
rect 33090 -9255 33135 -9135
rect 33255 -9255 33300 -9135
rect 33420 -9255 33475 -9135
rect 33595 -9255 33640 -9135
rect 33760 -9255 33805 -9135
rect 33925 -9255 33970 -9135
rect 34090 -9255 34145 -9135
rect 34265 -9255 34310 -9135
rect 34430 -9255 34475 -9135
rect 34595 -9255 34640 -9135
rect 34760 -9255 34815 -9135
rect 34935 -9255 34980 -9135
rect 35100 -9255 35145 -9135
rect 35265 -9255 35310 -9135
rect 35430 -9255 35485 -9135
rect 35605 -9255 35650 -9135
rect 35770 -9255 35815 -9135
rect 35935 -9255 35980 -9135
rect 36100 -9255 36155 -9135
rect 36275 -9255 36285 -9135
rect 30785 -9300 36285 -9255
rect 30785 -9420 30795 -9300
rect 30915 -9420 30960 -9300
rect 31080 -9420 31125 -9300
rect 31245 -9420 31290 -9300
rect 31410 -9420 31465 -9300
rect 31585 -9420 31630 -9300
rect 31750 -9420 31795 -9300
rect 31915 -9420 31960 -9300
rect 32080 -9420 32135 -9300
rect 32255 -9420 32300 -9300
rect 32420 -9420 32465 -9300
rect 32585 -9420 32630 -9300
rect 32750 -9420 32805 -9300
rect 32925 -9420 32970 -9300
rect 33090 -9420 33135 -9300
rect 33255 -9420 33300 -9300
rect 33420 -9420 33475 -9300
rect 33595 -9420 33640 -9300
rect 33760 -9420 33805 -9300
rect 33925 -9420 33970 -9300
rect 34090 -9420 34145 -9300
rect 34265 -9420 34310 -9300
rect 34430 -9420 34475 -9300
rect 34595 -9420 34640 -9300
rect 34760 -9420 34815 -9300
rect 34935 -9420 34980 -9300
rect 35100 -9420 35145 -9300
rect 35265 -9420 35310 -9300
rect 35430 -9420 35485 -9300
rect 35605 -9420 35650 -9300
rect 35770 -9420 35815 -9300
rect 35935 -9420 35980 -9300
rect 36100 -9420 36155 -9300
rect 36275 -9420 36285 -9300
rect 30785 -9465 36285 -9420
rect 30785 -9585 30795 -9465
rect 30915 -9585 30960 -9465
rect 31080 -9585 31125 -9465
rect 31245 -9585 31290 -9465
rect 31410 -9585 31465 -9465
rect 31585 -9585 31630 -9465
rect 31750 -9585 31795 -9465
rect 31915 -9585 31960 -9465
rect 32080 -9585 32135 -9465
rect 32255 -9585 32300 -9465
rect 32420 -9585 32465 -9465
rect 32585 -9585 32630 -9465
rect 32750 -9585 32805 -9465
rect 32925 -9585 32970 -9465
rect 33090 -9585 33135 -9465
rect 33255 -9585 33300 -9465
rect 33420 -9585 33475 -9465
rect 33595 -9585 33640 -9465
rect 33760 -9585 33805 -9465
rect 33925 -9585 33970 -9465
rect 34090 -9585 34145 -9465
rect 34265 -9585 34310 -9465
rect 34430 -9585 34475 -9465
rect 34595 -9585 34640 -9465
rect 34760 -9585 34815 -9465
rect 34935 -9585 34980 -9465
rect 35100 -9585 35145 -9465
rect 35265 -9585 35310 -9465
rect 35430 -9585 35485 -9465
rect 35605 -9585 35650 -9465
rect 35770 -9585 35815 -9465
rect 35935 -9585 35980 -9465
rect 36100 -9585 36155 -9465
rect 36275 -9585 36285 -9465
rect 30785 -9630 36285 -9585
rect 30785 -9750 30795 -9630
rect 30915 -9750 30960 -9630
rect 31080 -9750 31125 -9630
rect 31245 -9750 31290 -9630
rect 31410 -9750 31465 -9630
rect 31585 -9750 31630 -9630
rect 31750 -9750 31795 -9630
rect 31915 -9750 31960 -9630
rect 32080 -9750 32135 -9630
rect 32255 -9750 32300 -9630
rect 32420 -9750 32465 -9630
rect 32585 -9750 32630 -9630
rect 32750 -9750 32805 -9630
rect 32925 -9750 32970 -9630
rect 33090 -9750 33135 -9630
rect 33255 -9750 33300 -9630
rect 33420 -9750 33475 -9630
rect 33595 -9750 33640 -9630
rect 33760 -9750 33805 -9630
rect 33925 -9750 33970 -9630
rect 34090 -9750 34145 -9630
rect 34265 -9750 34310 -9630
rect 34430 -9750 34475 -9630
rect 34595 -9750 34640 -9630
rect 34760 -9750 34815 -9630
rect 34935 -9750 34980 -9630
rect 35100 -9750 35145 -9630
rect 35265 -9750 35310 -9630
rect 35430 -9750 35485 -9630
rect 35605 -9750 35650 -9630
rect 35770 -9750 35815 -9630
rect 35935 -9750 35980 -9630
rect 36100 -9750 36155 -9630
rect 36275 -9750 36285 -9630
rect 30785 -9760 36285 -9750
rect 36475 -4270 41975 -4260
rect 36475 -4390 36485 -4270
rect 36605 -4390 36650 -4270
rect 36770 -4390 36815 -4270
rect 36935 -4390 36980 -4270
rect 37100 -4390 37155 -4270
rect 37275 -4390 37320 -4270
rect 37440 -4390 37485 -4270
rect 37605 -4390 37650 -4270
rect 37770 -4390 37825 -4270
rect 37945 -4390 37990 -4270
rect 38110 -4390 38155 -4270
rect 38275 -4390 38320 -4270
rect 38440 -4390 38495 -4270
rect 38615 -4390 38660 -4270
rect 38780 -4390 38825 -4270
rect 38945 -4390 38990 -4270
rect 39110 -4390 39165 -4270
rect 39285 -4390 39330 -4270
rect 39450 -4390 39495 -4270
rect 39615 -4390 39660 -4270
rect 39780 -4390 39835 -4270
rect 39955 -4390 40000 -4270
rect 40120 -4390 40165 -4270
rect 40285 -4390 40330 -4270
rect 40450 -4390 40505 -4270
rect 40625 -4390 40670 -4270
rect 40790 -4390 40835 -4270
rect 40955 -4390 41000 -4270
rect 41120 -4390 41175 -4270
rect 41295 -4390 41340 -4270
rect 41460 -4390 41505 -4270
rect 41625 -4390 41670 -4270
rect 41790 -4390 41845 -4270
rect 41965 -4390 41975 -4270
rect 36475 -4445 41975 -4390
rect 36475 -4565 36485 -4445
rect 36605 -4565 36650 -4445
rect 36770 -4565 36815 -4445
rect 36935 -4565 36980 -4445
rect 37100 -4565 37155 -4445
rect 37275 -4565 37320 -4445
rect 37440 -4565 37485 -4445
rect 37605 -4565 37650 -4445
rect 37770 -4565 37825 -4445
rect 37945 -4565 37990 -4445
rect 38110 -4565 38155 -4445
rect 38275 -4565 38320 -4445
rect 38440 -4565 38495 -4445
rect 38615 -4565 38660 -4445
rect 38780 -4565 38825 -4445
rect 38945 -4565 38990 -4445
rect 39110 -4565 39165 -4445
rect 39285 -4565 39330 -4445
rect 39450 -4565 39495 -4445
rect 39615 -4565 39660 -4445
rect 39780 -4565 39835 -4445
rect 39955 -4565 40000 -4445
rect 40120 -4565 40165 -4445
rect 40285 -4565 40330 -4445
rect 40450 -4565 40505 -4445
rect 40625 -4565 40670 -4445
rect 40790 -4565 40835 -4445
rect 40955 -4565 41000 -4445
rect 41120 -4565 41175 -4445
rect 41295 -4565 41340 -4445
rect 41460 -4565 41505 -4445
rect 41625 -4565 41670 -4445
rect 41790 -4565 41845 -4445
rect 41965 -4565 41975 -4445
rect 36475 -4610 41975 -4565
rect 36475 -4730 36485 -4610
rect 36605 -4730 36650 -4610
rect 36770 -4730 36815 -4610
rect 36935 -4730 36980 -4610
rect 37100 -4730 37155 -4610
rect 37275 -4730 37320 -4610
rect 37440 -4730 37485 -4610
rect 37605 -4730 37650 -4610
rect 37770 -4730 37825 -4610
rect 37945 -4730 37990 -4610
rect 38110 -4730 38155 -4610
rect 38275 -4730 38320 -4610
rect 38440 -4730 38495 -4610
rect 38615 -4730 38660 -4610
rect 38780 -4730 38825 -4610
rect 38945 -4730 38990 -4610
rect 39110 -4730 39165 -4610
rect 39285 -4730 39330 -4610
rect 39450 -4730 39495 -4610
rect 39615 -4730 39660 -4610
rect 39780 -4730 39835 -4610
rect 39955 -4730 40000 -4610
rect 40120 -4730 40165 -4610
rect 40285 -4730 40330 -4610
rect 40450 -4730 40505 -4610
rect 40625 -4730 40670 -4610
rect 40790 -4730 40835 -4610
rect 40955 -4730 41000 -4610
rect 41120 -4730 41175 -4610
rect 41295 -4730 41340 -4610
rect 41460 -4730 41505 -4610
rect 41625 -4730 41670 -4610
rect 41790 -4730 41845 -4610
rect 41965 -4730 41975 -4610
rect 36475 -4775 41975 -4730
rect 36475 -4895 36485 -4775
rect 36605 -4895 36650 -4775
rect 36770 -4895 36815 -4775
rect 36935 -4895 36980 -4775
rect 37100 -4895 37155 -4775
rect 37275 -4895 37320 -4775
rect 37440 -4895 37485 -4775
rect 37605 -4895 37650 -4775
rect 37770 -4895 37825 -4775
rect 37945 -4895 37990 -4775
rect 38110 -4895 38155 -4775
rect 38275 -4895 38320 -4775
rect 38440 -4895 38495 -4775
rect 38615 -4895 38660 -4775
rect 38780 -4895 38825 -4775
rect 38945 -4895 38990 -4775
rect 39110 -4895 39165 -4775
rect 39285 -4895 39330 -4775
rect 39450 -4895 39495 -4775
rect 39615 -4895 39660 -4775
rect 39780 -4895 39835 -4775
rect 39955 -4895 40000 -4775
rect 40120 -4895 40165 -4775
rect 40285 -4895 40330 -4775
rect 40450 -4895 40505 -4775
rect 40625 -4895 40670 -4775
rect 40790 -4895 40835 -4775
rect 40955 -4895 41000 -4775
rect 41120 -4895 41175 -4775
rect 41295 -4895 41340 -4775
rect 41460 -4895 41505 -4775
rect 41625 -4895 41670 -4775
rect 41790 -4895 41845 -4775
rect 41965 -4895 41975 -4775
rect 36475 -4940 41975 -4895
rect 36475 -5060 36485 -4940
rect 36605 -5060 36650 -4940
rect 36770 -5060 36815 -4940
rect 36935 -5060 36980 -4940
rect 37100 -5060 37155 -4940
rect 37275 -5060 37320 -4940
rect 37440 -5060 37485 -4940
rect 37605 -5060 37650 -4940
rect 37770 -5060 37825 -4940
rect 37945 -5060 37990 -4940
rect 38110 -5060 38155 -4940
rect 38275 -5060 38320 -4940
rect 38440 -5060 38495 -4940
rect 38615 -5060 38660 -4940
rect 38780 -5060 38825 -4940
rect 38945 -5060 38990 -4940
rect 39110 -5060 39165 -4940
rect 39285 -5060 39330 -4940
rect 39450 -5060 39495 -4940
rect 39615 -5060 39660 -4940
rect 39780 -5060 39835 -4940
rect 39955 -5060 40000 -4940
rect 40120 -5060 40165 -4940
rect 40285 -5060 40330 -4940
rect 40450 -5060 40505 -4940
rect 40625 -5060 40670 -4940
rect 40790 -5060 40835 -4940
rect 40955 -5060 41000 -4940
rect 41120 -5060 41175 -4940
rect 41295 -5060 41340 -4940
rect 41460 -5060 41505 -4940
rect 41625 -5060 41670 -4940
rect 41790 -5060 41845 -4940
rect 41965 -5060 41975 -4940
rect 36475 -5115 41975 -5060
rect 36475 -5235 36485 -5115
rect 36605 -5235 36650 -5115
rect 36770 -5235 36815 -5115
rect 36935 -5235 36980 -5115
rect 37100 -5235 37155 -5115
rect 37275 -5235 37320 -5115
rect 37440 -5235 37485 -5115
rect 37605 -5235 37650 -5115
rect 37770 -5235 37825 -5115
rect 37945 -5235 37990 -5115
rect 38110 -5235 38155 -5115
rect 38275 -5235 38320 -5115
rect 38440 -5235 38495 -5115
rect 38615 -5235 38660 -5115
rect 38780 -5235 38825 -5115
rect 38945 -5235 38990 -5115
rect 39110 -5235 39165 -5115
rect 39285 -5235 39330 -5115
rect 39450 -5235 39495 -5115
rect 39615 -5235 39660 -5115
rect 39780 -5235 39835 -5115
rect 39955 -5235 40000 -5115
rect 40120 -5235 40165 -5115
rect 40285 -5235 40330 -5115
rect 40450 -5235 40505 -5115
rect 40625 -5235 40670 -5115
rect 40790 -5235 40835 -5115
rect 40955 -5235 41000 -5115
rect 41120 -5235 41175 -5115
rect 41295 -5235 41340 -5115
rect 41460 -5235 41505 -5115
rect 41625 -5235 41670 -5115
rect 41790 -5235 41845 -5115
rect 41965 -5235 41975 -5115
rect 36475 -5280 41975 -5235
rect 36475 -5400 36485 -5280
rect 36605 -5400 36650 -5280
rect 36770 -5400 36815 -5280
rect 36935 -5400 36980 -5280
rect 37100 -5400 37155 -5280
rect 37275 -5400 37320 -5280
rect 37440 -5400 37485 -5280
rect 37605 -5400 37650 -5280
rect 37770 -5400 37825 -5280
rect 37945 -5400 37990 -5280
rect 38110 -5400 38155 -5280
rect 38275 -5400 38320 -5280
rect 38440 -5400 38495 -5280
rect 38615 -5400 38660 -5280
rect 38780 -5400 38825 -5280
rect 38945 -5400 38990 -5280
rect 39110 -5400 39165 -5280
rect 39285 -5400 39330 -5280
rect 39450 -5400 39495 -5280
rect 39615 -5400 39660 -5280
rect 39780 -5400 39835 -5280
rect 39955 -5400 40000 -5280
rect 40120 -5400 40165 -5280
rect 40285 -5400 40330 -5280
rect 40450 -5400 40505 -5280
rect 40625 -5400 40670 -5280
rect 40790 -5400 40835 -5280
rect 40955 -5400 41000 -5280
rect 41120 -5400 41175 -5280
rect 41295 -5400 41340 -5280
rect 41460 -5400 41505 -5280
rect 41625 -5400 41670 -5280
rect 41790 -5400 41845 -5280
rect 41965 -5400 41975 -5280
rect 36475 -5445 41975 -5400
rect 36475 -5565 36485 -5445
rect 36605 -5565 36650 -5445
rect 36770 -5565 36815 -5445
rect 36935 -5565 36980 -5445
rect 37100 -5565 37155 -5445
rect 37275 -5565 37320 -5445
rect 37440 -5565 37485 -5445
rect 37605 -5565 37650 -5445
rect 37770 -5565 37825 -5445
rect 37945 -5565 37990 -5445
rect 38110 -5565 38155 -5445
rect 38275 -5565 38320 -5445
rect 38440 -5565 38495 -5445
rect 38615 -5565 38660 -5445
rect 38780 -5565 38825 -5445
rect 38945 -5565 38990 -5445
rect 39110 -5565 39165 -5445
rect 39285 -5565 39330 -5445
rect 39450 -5565 39495 -5445
rect 39615 -5565 39660 -5445
rect 39780 -5565 39835 -5445
rect 39955 -5565 40000 -5445
rect 40120 -5565 40165 -5445
rect 40285 -5565 40330 -5445
rect 40450 -5565 40505 -5445
rect 40625 -5565 40670 -5445
rect 40790 -5565 40835 -5445
rect 40955 -5565 41000 -5445
rect 41120 -5565 41175 -5445
rect 41295 -5565 41340 -5445
rect 41460 -5565 41505 -5445
rect 41625 -5565 41670 -5445
rect 41790 -5565 41845 -5445
rect 41965 -5565 41975 -5445
rect 36475 -5610 41975 -5565
rect 36475 -5730 36485 -5610
rect 36605 -5730 36650 -5610
rect 36770 -5730 36815 -5610
rect 36935 -5730 36980 -5610
rect 37100 -5730 37155 -5610
rect 37275 -5730 37320 -5610
rect 37440 -5730 37485 -5610
rect 37605 -5730 37650 -5610
rect 37770 -5730 37825 -5610
rect 37945 -5730 37990 -5610
rect 38110 -5730 38155 -5610
rect 38275 -5730 38320 -5610
rect 38440 -5730 38495 -5610
rect 38615 -5730 38660 -5610
rect 38780 -5730 38825 -5610
rect 38945 -5730 38990 -5610
rect 39110 -5730 39165 -5610
rect 39285 -5730 39330 -5610
rect 39450 -5730 39495 -5610
rect 39615 -5730 39660 -5610
rect 39780 -5730 39835 -5610
rect 39955 -5730 40000 -5610
rect 40120 -5730 40165 -5610
rect 40285 -5730 40330 -5610
rect 40450 -5730 40505 -5610
rect 40625 -5730 40670 -5610
rect 40790 -5730 40835 -5610
rect 40955 -5730 41000 -5610
rect 41120 -5730 41175 -5610
rect 41295 -5730 41340 -5610
rect 41460 -5730 41505 -5610
rect 41625 -5730 41670 -5610
rect 41790 -5730 41845 -5610
rect 41965 -5730 41975 -5610
rect 36475 -5785 41975 -5730
rect 36475 -5905 36485 -5785
rect 36605 -5905 36650 -5785
rect 36770 -5905 36815 -5785
rect 36935 -5905 36980 -5785
rect 37100 -5905 37155 -5785
rect 37275 -5905 37320 -5785
rect 37440 -5905 37485 -5785
rect 37605 -5905 37650 -5785
rect 37770 -5905 37825 -5785
rect 37945 -5905 37990 -5785
rect 38110 -5905 38155 -5785
rect 38275 -5905 38320 -5785
rect 38440 -5905 38495 -5785
rect 38615 -5905 38660 -5785
rect 38780 -5905 38825 -5785
rect 38945 -5905 38990 -5785
rect 39110 -5905 39165 -5785
rect 39285 -5905 39330 -5785
rect 39450 -5905 39495 -5785
rect 39615 -5905 39660 -5785
rect 39780 -5905 39835 -5785
rect 39955 -5905 40000 -5785
rect 40120 -5905 40165 -5785
rect 40285 -5905 40330 -5785
rect 40450 -5905 40505 -5785
rect 40625 -5905 40670 -5785
rect 40790 -5905 40835 -5785
rect 40955 -5905 41000 -5785
rect 41120 -5905 41175 -5785
rect 41295 -5905 41340 -5785
rect 41460 -5905 41505 -5785
rect 41625 -5905 41670 -5785
rect 41790 -5905 41845 -5785
rect 41965 -5905 41975 -5785
rect 36475 -5950 41975 -5905
rect 36475 -6070 36485 -5950
rect 36605 -6070 36650 -5950
rect 36770 -6070 36815 -5950
rect 36935 -6070 36980 -5950
rect 37100 -6070 37155 -5950
rect 37275 -6070 37320 -5950
rect 37440 -6070 37485 -5950
rect 37605 -6070 37650 -5950
rect 37770 -6070 37825 -5950
rect 37945 -6070 37990 -5950
rect 38110 -6070 38155 -5950
rect 38275 -6070 38320 -5950
rect 38440 -6070 38495 -5950
rect 38615 -6070 38660 -5950
rect 38780 -6070 38825 -5950
rect 38945 -6070 38990 -5950
rect 39110 -6070 39165 -5950
rect 39285 -6070 39330 -5950
rect 39450 -6070 39495 -5950
rect 39615 -6070 39660 -5950
rect 39780 -6070 39835 -5950
rect 39955 -6070 40000 -5950
rect 40120 -6070 40165 -5950
rect 40285 -6070 40330 -5950
rect 40450 -6070 40505 -5950
rect 40625 -6070 40670 -5950
rect 40790 -6070 40835 -5950
rect 40955 -6070 41000 -5950
rect 41120 -6070 41175 -5950
rect 41295 -6070 41340 -5950
rect 41460 -6070 41505 -5950
rect 41625 -6070 41670 -5950
rect 41790 -6070 41845 -5950
rect 41965 -6070 41975 -5950
rect 36475 -6115 41975 -6070
rect 36475 -6235 36485 -6115
rect 36605 -6235 36650 -6115
rect 36770 -6235 36815 -6115
rect 36935 -6235 36980 -6115
rect 37100 -6235 37155 -6115
rect 37275 -6235 37320 -6115
rect 37440 -6235 37485 -6115
rect 37605 -6235 37650 -6115
rect 37770 -6235 37825 -6115
rect 37945 -6235 37990 -6115
rect 38110 -6235 38155 -6115
rect 38275 -6235 38320 -6115
rect 38440 -6235 38495 -6115
rect 38615 -6235 38660 -6115
rect 38780 -6235 38825 -6115
rect 38945 -6235 38990 -6115
rect 39110 -6235 39165 -6115
rect 39285 -6235 39330 -6115
rect 39450 -6235 39495 -6115
rect 39615 -6235 39660 -6115
rect 39780 -6235 39835 -6115
rect 39955 -6235 40000 -6115
rect 40120 -6235 40165 -6115
rect 40285 -6235 40330 -6115
rect 40450 -6235 40505 -6115
rect 40625 -6235 40670 -6115
rect 40790 -6235 40835 -6115
rect 40955 -6235 41000 -6115
rect 41120 -6235 41175 -6115
rect 41295 -6235 41340 -6115
rect 41460 -6235 41505 -6115
rect 41625 -6235 41670 -6115
rect 41790 -6235 41845 -6115
rect 41965 -6235 41975 -6115
rect 36475 -6280 41975 -6235
rect 36475 -6400 36485 -6280
rect 36605 -6400 36650 -6280
rect 36770 -6400 36815 -6280
rect 36935 -6400 36980 -6280
rect 37100 -6400 37155 -6280
rect 37275 -6400 37320 -6280
rect 37440 -6400 37485 -6280
rect 37605 -6400 37650 -6280
rect 37770 -6400 37825 -6280
rect 37945 -6400 37990 -6280
rect 38110 -6400 38155 -6280
rect 38275 -6400 38320 -6280
rect 38440 -6400 38495 -6280
rect 38615 -6400 38660 -6280
rect 38780 -6400 38825 -6280
rect 38945 -6400 38990 -6280
rect 39110 -6400 39165 -6280
rect 39285 -6400 39330 -6280
rect 39450 -6400 39495 -6280
rect 39615 -6400 39660 -6280
rect 39780 -6400 39835 -6280
rect 39955 -6400 40000 -6280
rect 40120 -6400 40165 -6280
rect 40285 -6400 40330 -6280
rect 40450 -6400 40505 -6280
rect 40625 -6400 40670 -6280
rect 40790 -6400 40835 -6280
rect 40955 -6400 41000 -6280
rect 41120 -6400 41175 -6280
rect 41295 -6400 41340 -6280
rect 41460 -6400 41505 -6280
rect 41625 -6400 41670 -6280
rect 41790 -6400 41845 -6280
rect 41965 -6400 41975 -6280
rect 36475 -6455 41975 -6400
rect 36475 -6575 36485 -6455
rect 36605 -6575 36650 -6455
rect 36770 -6575 36815 -6455
rect 36935 -6575 36980 -6455
rect 37100 -6575 37155 -6455
rect 37275 -6575 37320 -6455
rect 37440 -6575 37485 -6455
rect 37605 -6575 37650 -6455
rect 37770 -6575 37825 -6455
rect 37945 -6575 37990 -6455
rect 38110 -6575 38155 -6455
rect 38275 -6575 38320 -6455
rect 38440 -6575 38495 -6455
rect 38615 -6575 38660 -6455
rect 38780 -6575 38825 -6455
rect 38945 -6575 38990 -6455
rect 39110 -6575 39165 -6455
rect 39285 -6575 39330 -6455
rect 39450 -6575 39495 -6455
rect 39615 -6575 39660 -6455
rect 39780 -6575 39835 -6455
rect 39955 -6575 40000 -6455
rect 40120 -6575 40165 -6455
rect 40285 -6575 40330 -6455
rect 40450 -6575 40505 -6455
rect 40625 -6575 40670 -6455
rect 40790 -6575 40835 -6455
rect 40955 -6575 41000 -6455
rect 41120 -6575 41175 -6455
rect 41295 -6575 41340 -6455
rect 41460 -6575 41505 -6455
rect 41625 -6575 41670 -6455
rect 41790 -6575 41845 -6455
rect 41965 -6575 41975 -6455
rect 36475 -6620 41975 -6575
rect 36475 -6740 36485 -6620
rect 36605 -6740 36650 -6620
rect 36770 -6740 36815 -6620
rect 36935 -6740 36980 -6620
rect 37100 -6740 37155 -6620
rect 37275 -6740 37320 -6620
rect 37440 -6740 37485 -6620
rect 37605 -6740 37650 -6620
rect 37770 -6740 37825 -6620
rect 37945 -6740 37990 -6620
rect 38110 -6740 38155 -6620
rect 38275 -6740 38320 -6620
rect 38440 -6740 38495 -6620
rect 38615 -6740 38660 -6620
rect 38780 -6740 38825 -6620
rect 38945 -6740 38990 -6620
rect 39110 -6740 39165 -6620
rect 39285 -6740 39330 -6620
rect 39450 -6740 39495 -6620
rect 39615 -6740 39660 -6620
rect 39780 -6740 39835 -6620
rect 39955 -6740 40000 -6620
rect 40120 -6740 40165 -6620
rect 40285 -6740 40330 -6620
rect 40450 -6740 40505 -6620
rect 40625 -6740 40670 -6620
rect 40790 -6740 40835 -6620
rect 40955 -6740 41000 -6620
rect 41120 -6740 41175 -6620
rect 41295 -6740 41340 -6620
rect 41460 -6740 41505 -6620
rect 41625 -6740 41670 -6620
rect 41790 -6740 41845 -6620
rect 41965 -6740 41975 -6620
rect 36475 -6785 41975 -6740
rect 36475 -6905 36485 -6785
rect 36605 -6905 36650 -6785
rect 36770 -6905 36815 -6785
rect 36935 -6905 36980 -6785
rect 37100 -6905 37155 -6785
rect 37275 -6905 37320 -6785
rect 37440 -6905 37485 -6785
rect 37605 -6905 37650 -6785
rect 37770 -6905 37825 -6785
rect 37945 -6905 37990 -6785
rect 38110 -6905 38155 -6785
rect 38275 -6905 38320 -6785
rect 38440 -6905 38495 -6785
rect 38615 -6905 38660 -6785
rect 38780 -6905 38825 -6785
rect 38945 -6905 38990 -6785
rect 39110 -6905 39165 -6785
rect 39285 -6905 39330 -6785
rect 39450 -6905 39495 -6785
rect 39615 -6905 39660 -6785
rect 39780 -6905 39835 -6785
rect 39955 -6905 40000 -6785
rect 40120 -6905 40165 -6785
rect 40285 -6905 40330 -6785
rect 40450 -6905 40505 -6785
rect 40625 -6905 40670 -6785
rect 40790 -6905 40835 -6785
rect 40955 -6905 41000 -6785
rect 41120 -6905 41175 -6785
rect 41295 -6905 41340 -6785
rect 41460 -6905 41505 -6785
rect 41625 -6905 41670 -6785
rect 41790 -6905 41845 -6785
rect 41965 -6905 41975 -6785
rect 36475 -6950 41975 -6905
rect 36475 -7070 36485 -6950
rect 36605 -7070 36650 -6950
rect 36770 -7070 36815 -6950
rect 36935 -7070 36980 -6950
rect 37100 -7070 37155 -6950
rect 37275 -7070 37320 -6950
rect 37440 -7070 37485 -6950
rect 37605 -7070 37650 -6950
rect 37770 -7070 37825 -6950
rect 37945 -7070 37990 -6950
rect 38110 -7070 38155 -6950
rect 38275 -7070 38320 -6950
rect 38440 -7070 38495 -6950
rect 38615 -7070 38660 -6950
rect 38780 -7070 38825 -6950
rect 38945 -7070 38990 -6950
rect 39110 -7070 39165 -6950
rect 39285 -7070 39330 -6950
rect 39450 -7070 39495 -6950
rect 39615 -7070 39660 -6950
rect 39780 -7070 39835 -6950
rect 39955 -7070 40000 -6950
rect 40120 -7070 40165 -6950
rect 40285 -7070 40330 -6950
rect 40450 -7070 40505 -6950
rect 40625 -7070 40670 -6950
rect 40790 -7070 40835 -6950
rect 40955 -7070 41000 -6950
rect 41120 -7070 41175 -6950
rect 41295 -7070 41340 -6950
rect 41460 -7070 41505 -6950
rect 41625 -7070 41670 -6950
rect 41790 -7070 41845 -6950
rect 41965 -7070 41975 -6950
rect 36475 -7125 41975 -7070
rect 36475 -7245 36485 -7125
rect 36605 -7245 36650 -7125
rect 36770 -7245 36815 -7125
rect 36935 -7245 36980 -7125
rect 37100 -7245 37155 -7125
rect 37275 -7245 37320 -7125
rect 37440 -7245 37485 -7125
rect 37605 -7245 37650 -7125
rect 37770 -7245 37825 -7125
rect 37945 -7245 37990 -7125
rect 38110 -7245 38155 -7125
rect 38275 -7245 38320 -7125
rect 38440 -7245 38495 -7125
rect 38615 -7245 38660 -7125
rect 38780 -7245 38825 -7125
rect 38945 -7245 38990 -7125
rect 39110 -7245 39165 -7125
rect 39285 -7245 39330 -7125
rect 39450 -7245 39495 -7125
rect 39615 -7245 39660 -7125
rect 39780 -7245 39835 -7125
rect 39955 -7245 40000 -7125
rect 40120 -7245 40165 -7125
rect 40285 -7245 40330 -7125
rect 40450 -7245 40505 -7125
rect 40625 -7245 40670 -7125
rect 40790 -7245 40835 -7125
rect 40955 -7245 41000 -7125
rect 41120 -7245 41175 -7125
rect 41295 -7245 41340 -7125
rect 41460 -7245 41505 -7125
rect 41625 -7245 41670 -7125
rect 41790 -7245 41845 -7125
rect 41965 -7245 41975 -7125
rect 36475 -7290 41975 -7245
rect 36475 -7410 36485 -7290
rect 36605 -7410 36650 -7290
rect 36770 -7410 36815 -7290
rect 36935 -7410 36980 -7290
rect 37100 -7410 37155 -7290
rect 37275 -7410 37320 -7290
rect 37440 -7410 37485 -7290
rect 37605 -7410 37650 -7290
rect 37770 -7410 37825 -7290
rect 37945 -7410 37990 -7290
rect 38110 -7410 38155 -7290
rect 38275 -7410 38320 -7290
rect 38440 -7410 38495 -7290
rect 38615 -7410 38660 -7290
rect 38780 -7410 38825 -7290
rect 38945 -7410 38990 -7290
rect 39110 -7410 39165 -7290
rect 39285 -7410 39330 -7290
rect 39450 -7410 39495 -7290
rect 39615 -7410 39660 -7290
rect 39780 -7410 39835 -7290
rect 39955 -7410 40000 -7290
rect 40120 -7410 40165 -7290
rect 40285 -7410 40330 -7290
rect 40450 -7410 40505 -7290
rect 40625 -7410 40670 -7290
rect 40790 -7410 40835 -7290
rect 40955 -7410 41000 -7290
rect 41120 -7410 41175 -7290
rect 41295 -7410 41340 -7290
rect 41460 -7410 41505 -7290
rect 41625 -7410 41670 -7290
rect 41790 -7410 41845 -7290
rect 41965 -7410 41975 -7290
rect 36475 -7455 41975 -7410
rect 36475 -7575 36485 -7455
rect 36605 -7575 36650 -7455
rect 36770 -7575 36815 -7455
rect 36935 -7575 36980 -7455
rect 37100 -7575 37155 -7455
rect 37275 -7575 37320 -7455
rect 37440 -7575 37485 -7455
rect 37605 -7575 37650 -7455
rect 37770 -7575 37825 -7455
rect 37945 -7575 37990 -7455
rect 38110 -7575 38155 -7455
rect 38275 -7575 38320 -7455
rect 38440 -7575 38495 -7455
rect 38615 -7575 38660 -7455
rect 38780 -7575 38825 -7455
rect 38945 -7575 38990 -7455
rect 39110 -7575 39165 -7455
rect 39285 -7575 39330 -7455
rect 39450 -7575 39495 -7455
rect 39615 -7575 39660 -7455
rect 39780 -7575 39835 -7455
rect 39955 -7575 40000 -7455
rect 40120 -7575 40165 -7455
rect 40285 -7575 40330 -7455
rect 40450 -7575 40505 -7455
rect 40625 -7575 40670 -7455
rect 40790 -7575 40835 -7455
rect 40955 -7575 41000 -7455
rect 41120 -7575 41175 -7455
rect 41295 -7575 41340 -7455
rect 41460 -7575 41505 -7455
rect 41625 -7575 41670 -7455
rect 41790 -7575 41845 -7455
rect 41965 -7575 41975 -7455
rect 36475 -7620 41975 -7575
rect 36475 -7740 36485 -7620
rect 36605 -7740 36650 -7620
rect 36770 -7740 36815 -7620
rect 36935 -7740 36980 -7620
rect 37100 -7740 37155 -7620
rect 37275 -7740 37320 -7620
rect 37440 -7740 37485 -7620
rect 37605 -7740 37650 -7620
rect 37770 -7740 37825 -7620
rect 37945 -7740 37990 -7620
rect 38110 -7740 38155 -7620
rect 38275 -7740 38320 -7620
rect 38440 -7740 38495 -7620
rect 38615 -7740 38660 -7620
rect 38780 -7740 38825 -7620
rect 38945 -7740 38990 -7620
rect 39110 -7740 39165 -7620
rect 39285 -7740 39330 -7620
rect 39450 -7740 39495 -7620
rect 39615 -7740 39660 -7620
rect 39780 -7740 39835 -7620
rect 39955 -7740 40000 -7620
rect 40120 -7740 40165 -7620
rect 40285 -7740 40330 -7620
rect 40450 -7740 40505 -7620
rect 40625 -7740 40670 -7620
rect 40790 -7740 40835 -7620
rect 40955 -7740 41000 -7620
rect 41120 -7740 41175 -7620
rect 41295 -7740 41340 -7620
rect 41460 -7740 41505 -7620
rect 41625 -7740 41670 -7620
rect 41790 -7740 41845 -7620
rect 41965 -7740 41975 -7620
rect 36475 -7795 41975 -7740
rect 36475 -7915 36485 -7795
rect 36605 -7915 36650 -7795
rect 36770 -7915 36815 -7795
rect 36935 -7915 36980 -7795
rect 37100 -7915 37155 -7795
rect 37275 -7915 37320 -7795
rect 37440 -7915 37485 -7795
rect 37605 -7915 37650 -7795
rect 37770 -7915 37825 -7795
rect 37945 -7915 37990 -7795
rect 38110 -7915 38155 -7795
rect 38275 -7915 38320 -7795
rect 38440 -7915 38495 -7795
rect 38615 -7915 38660 -7795
rect 38780 -7915 38825 -7795
rect 38945 -7915 38990 -7795
rect 39110 -7915 39165 -7795
rect 39285 -7915 39330 -7795
rect 39450 -7915 39495 -7795
rect 39615 -7915 39660 -7795
rect 39780 -7915 39835 -7795
rect 39955 -7915 40000 -7795
rect 40120 -7915 40165 -7795
rect 40285 -7915 40330 -7795
rect 40450 -7915 40505 -7795
rect 40625 -7915 40670 -7795
rect 40790 -7915 40835 -7795
rect 40955 -7915 41000 -7795
rect 41120 -7915 41175 -7795
rect 41295 -7915 41340 -7795
rect 41460 -7915 41505 -7795
rect 41625 -7915 41670 -7795
rect 41790 -7915 41845 -7795
rect 41965 -7915 41975 -7795
rect 36475 -7960 41975 -7915
rect 36475 -8080 36485 -7960
rect 36605 -8080 36650 -7960
rect 36770 -8080 36815 -7960
rect 36935 -8080 36980 -7960
rect 37100 -8080 37155 -7960
rect 37275 -8080 37320 -7960
rect 37440 -8080 37485 -7960
rect 37605 -8080 37650 -7960
rect 37770 -8080 37825 -7960
rect 37945 -8080 37990 -7960
rect 38110 -8080 38155 -7960
rect 38275 -8080 38320 -7960
rect 38440 -8080 38495 -7960
rect 38615 -8080 38660 -7960
rect 38780 -8080 38825 -7960
rect 38945 -8080 38990 -7960
rect 39110 -8080 39165 -7960
rect 39285 -8080 39330 -7960
rect 39450 -8080 39495 -7960
rect 39615 -8080 39660 -7960
rect 39780 -8080 39835 -7960
rect 39955 -8080 40000 -7960
rect 40120 -8080 40165 -7960
rect 40285 -8080 40330 -7960
rect 40450 -8080 40505 -7960
rect 40625 -8080 40670 -7960
rect 40790 -8080 40835 -7960
rect 40955 -8080 41000 -7960
rect 41120 -8080 41175 -7960
rect 41295 -8080 41340 -7960
rect 41460 -8080 41505 -7960
rect 41625 -8080 41670 -7960
rect 41790 -8080 41845 -7960
rect 41965 -8080 41975 -7960
rect 36475 -8125 41975 -8080
rect 36475 -8245 36485 -8125
rect 36605 -8245 36650 -8125
rect 36770 -8245 36815 -8125
rect 36935 -8245 36980 -8125
rect 37100 -8245 37155 -8125
rect 37275 -8245 37320 -8125
rect 37440 -8245 37485 -8125
rect 37605 -8245 37650 -8125
rect 37770 -8245 37825 -8125
rect 37945 -8245 37990 -8125
rect 38110 -8245 38155 -8125
rect 38275 -8245 38320 -8125
rect 38440 -8245 38495 -8125
rect 38615 -8245 38660 -8125
rect 38780 -8245 38825 -8125
rect 38945 -8245 38990 -8125
rect 39110 -8245 39165 -8125
rect 39285 -8245 39330 -8125
rect 39450 -8245 39495 -8125
rect 39615 -8245 39660 -8125
rect 39780 -8245 39835 -8125
rect 39955 -8245 40000 -8125
rect 40120 -8245 40165 -8125
rect 40285 -8245 40330 -8125
rect 40450 -8245 40505 -8125
rect 40625 -8245 40670 -8125
rect 40790 -8245 40835 -8125
rect 40955 -8245 41000 -8125
rect 41120 -8245 41175 -8125
rect 41295 -8245 41340 -8125
rect 41460 -8245 41505 -8125
rect 41625 -8245 41670 -8125
rect 41790 -8245 41845 -8125
rect 41965 -8245 41975 -8125
rect 36475 -8290 41975 -8245
rect 36475 -8410 36485 -8290
rect 36605 -8410 36650 -8290
rect 36770 -8410 36815 -8290
rect 36935 -8410 36980 -8290
rect 37100 -8410 37155 -8290
rect 37275 -8410 37320 -8290
rect 37440 -8410 37485 -8290
rect 37605 -8410 37650 -8290
rect 37770 -8410 37825 -8290
rect 37945 -8410 37990 -8290
rect 38110 -8410 38155 -8290
rect 38275 -8410 38320 -8290
rect 38440 -8410 38495 -8290
rect 38615 -8410 38660 -8290
rect 38780 -8410 38825 -8290
rect 38945 -8410 38990 -8290
rect 39110 -8410 39165 -8290
rect 39285 -8410 39330 -8290
rect 39450 -8410 39495 -8290
rect 39615 -8410 39660 -8290
rect 39780 -8410 39835 -8290
rect 39955 -8410 40000 -8290
rect 40120 -8410 40165 -8290
rect 40285 -8410 40330 -8290
rect 40450 -8410 40505 -8290
rect 40625 -8410 40670 -8290
rect 40790 -8410 40835 -8290
rect 40955 -8410 41000 -8290
rect 41120 -8410 41175 -8290
rect 41295 -8410 41340 -8290
rect 41460 -8410 41505 -8290
rect 41625 -8410 41670 -8290
rect 41790 -8410 41845 -8290
rect 41965 -8410 41975 -8290
rect 36475 -8465 41975 -8410
rect 36475 -8585 36485 -8465
rect 36605 -8585 36650 -8465
rect 36770 -8585 36815 -8465
rect 36935 -8585 36980 -8465
rect 37100 -8585 37155 -8465
rect 37275 -8585 37320 -8465
rect 37440 -8585 37485 -8465
rect 37605 -8585 37650 -8465
rect 37770 -8585 37825 -8465
rect 37945 -8585 37990 -8465
rect 38110 -8585 38155 -8465
rect 38275 -8585 38320 -8465
rect 38440 -8585 38495 -8465
rect 38615 -8585 38660 -8465
rect 38780 -8585 38825 -8465
rect 38945 -8585 38990 -8465
rect 39110 -8585 39165 -8465
rect 39285 -8585 39330 -8465
rect 39450 -8585 39495 -8465
rect 39615 -8585 39660 -8465
rect 39780 -8585 39835 -8465
rect 39955 -8585 40000 -8465
rect 40120 -8585 40165 -8465
rect 40285 -8585 40330 -8465
rect 40450 -8585 40505 -8465
rect 40625 -8585 40670 -8465
rect 40790 -8585 40835 -8465
rect 40955 -8585 41000 -8465
rect 41120 -8585 41175 -8465
rect 41295 -8585 41340 -8465
rect 41460 -8585 41505 -8465
rect 41625 -8585 41670 -8465
rect 41790 -8585 41845 -8465
rect 41965 -8585 41975 -8465
rect 36475 -8630 41975 -8585
rect 36475 -8750 36485 -8630
rect 36605 -8750 36650 -8630
rect 36770 -8750 36815 -8630
rect 36935 -8750 36980 -8630
rect 37100 -8750 37155 -8630
rect 37275 -8750 37320 -8630
rect 37440 -8750 37485 -8630
rect 37605 -8750 37650 -8630
rect 37770 -8750 37825 -8630
rect 37945 -8750 37990 -8630
rect 38110 -8750 38155 -8630
rect 38275 -8750 38320 -8630
rect 38440 -8750 38495 -8630
rect 38615 -8750 38660 -8630
rect 38780 -8750 38825 -8630
rect 38945 -8750 38990 -8630
rect 39110 -8750 39165 -8630
rect 39285 -8750 39330 -8630
rect 39450 -8750 39495 -8630
rect 39615 -8750 39660 -8630
rect 39780 -8750 39835 -8630
rect 39955 -8750 40000 -8630
rect 40120 -8750 40165 -8630
rect 40285 -8750 40330 -8630
rect 40450 -8750 40505 -8630
rect 40625 -8750 40670 -8630
rect 40790 -8750 40835 -8630
rect 40955 -8750 41000 -8630
rect 41120 -8750 41175 -8630
rect 41295 -8750 41340 -8630
rect 41460 -8750 41505 -8630
rect 41625 -8750 41670 -8630
rect 41790 -8750 41845 -8630
rect 41965 -8750 41975 -8630
rect 36475 -8795 41975 -8750
rect 36475 -8915 36485 -8795
rect 36605 -8915 36650 -8795
rect 36770 -8915 36815 -8795
rect 36935 -8915 36980 -8795
rect 37100 -8915 37155 -8795
rect 37275 -8915 37320 -8795
rect 37440 -8915 37485 -8795
rect 37605 -8915 37650 -8795
rect 37770 -8915 37825 -8795
rect 37945 -8915 37990 -8795
rect 38110 -8915 38155 -8795
rect 38275 -8915 38320 -8795
rect 38440 -8915 38495 -8795
rect 38615 -8915 38660 -8795
rect 38780 -8915 38825 -8795
rect 38945 -8915 38990 -8795
rect 39110 -8915 39165 -8795
rect 39285 -8915 39330 -8795
rect 39450 -8915 39495 -8795
rect 39615 -8915 39660 -8795
rect 39780 -8915 39835 -8795
rect 39955 -8915 40000 -8795
rect 40120 -8915 40165 -8795
rect 40285 -8915 40330 -8795
rect 40450 -8915 40505 -8795
rect 40625 -8915 40670 -8795
rect 40790 -8915 40835 -8795
rect 40955 -8915 41000 -8795
rect 41120 -8915 41175 -8795
rect 41295 -8915 41340 -8795
rect 41460 -8915 41505 -8795
rect 41625 -8915 41670 -8795
rect 41790 -8915 41845 -8795
rect 41965 -8915 41975 -8795
rect 36475 -8960 41975 -8915
rect 36475 -9080 36485 -8960
rect 36605 -9080 36650 -8960
rect 36770 -9080 36815 -8960
rect 36935 -9080 36980 -8960
rect 37100 -9080 37155 -8960
rect 37275 -9080 37320 -8960
rect 37440 -9080 37485 -8960
rect 37605 -9080 37650 -8960
rect 37770 -9080 37825 -8960
rect 37945 -9080 37990 -8960
rect 38110 -9080 38155 -8960
rect 38275 -9080 38320 -8960
rect 38440 -9080 38495 -8960
rect 38615 -9080 38660 -8960
rect 38780 -9080 38825 -8960
rect 38945 -9080 38990 -8960
rect 39110 -9080 39165 -8960
rect 39285 -9080 39330 -8960
rect 39450 -9080 39495 -8960
rect 39615 -9080 39660 -8960
rect 39780 -9080 39835 -8960
rect 39955 -9080 40000 -8960
rect 40120 -9080 40165 -8960
rect 40285 -9080 40330 -8960
rect 40450 -9080 40505 -8960
rect 40625 -9080 40670 -8960
rect 40790 -9080 40835 -8960
rect 40955 -9080 41000 -8960
rect 41120 -9080 41175 -8960
rect 41295 -9080 41340 -8960
rect 41460 -9080 41505 -8960
rect 41625 -9080 41670 -8960
rect 41790 -9080 41845 -8960
rect 41965 -9080 41975 -8960
rect 36475 -9135 41975 -9080
rect 36475 -9255 36485 -9135
rect 36605 -9255 36650 -9135
rect 36770 -9255 36815 -9135
rect 36935 -9255 36980 -9135
rect 37100 -9255 37155 -9135
rect 37275 -9255 37320 -9135
rect 37440 -9255 37485 -9135
rect 37605 -9255 37650 -9135
rect 37770 -9255 37825 -9135
rect 37945 -9255 37990 -9135
rect 38110 -9255 38155 -9135
rect 38275 -9255 38320 -9135
rect 38440 -9255 38495 -9135
rect 38615 -9255 38660 -9135
rect 38780 -9255 38825 -9135
rect 38945 -9255 38990 -9135
rect 39110 -9255 39165 -9135
rect 39285 -9255 39330 -9135
rect 39450 -9255 39495 -9135
rect 39615 -9255 39660 -9135
rect 39780 -9255 39835 -9135
rect 39955 -9255 40000 -9135
rect 40120 -9255 40165 -9135
rect 40285 -9255 40330 -9135
rect 40450 -9255 40505 -9135
rect 40625 -9255 40670 -9135
rect 40790 -9255 40835 -9135
rect 40955 -9255 41000 -9135
rect 41120 -9255 41175 -9135
rect 41295 -9255 41340 -9135
rect 41460 -9255 41505 -9135
rect 41625 -9255 41670 -9135
rect 41790 -9255 41845 -9135
rect 41965 -9255 41975 -9135
rect 36475 -9300 41975 -9255
rect 36475 -9420 36485 -9300
rect 36605 -9420 36650 -9300
rect 36770 -9420 36815 -9300
rect 36935 -9420 36980 -9300
rect 37100 -9420 37155 -9300
rect 37275 -9420 37320 -9300
rect 37440 -9420 37485 -9300
rect 37605 -9420 37650 -9300
rect 37770 -9420 37825 -9300
rect 37945 -9420 37990 -9300
rect 38110 -9420 38155 -9300
rect 38275 -9420 38320 -9300
rect 38440 -9420 38495 -9300
rect 38615 -9420 38660 -9300
rect 38780 -9420 38825 -9300
rect 38945 -9420 38990 -9300
rect 39110 -9420 39165 -9300
rect 39285 -9420 39330 -9300
rect 39450 -9420 39495 -9300
rect 39615 -9420 39660 -9300
rect 39780 -9420 39835 -9300
rect 39955 -9420 40000 -9300
rect 40120 -9420 40165 -9300
rect 40285 -9420 40330 -9300
rect 40450 -9420 40505 -9300
rect 40625 -9420 40670 -9300
rect 40790 -9420 40835 -9300
rect 40955 -9420 41000 -9300
rect 41120 -9420 41175 -9300
rect 41295 -9420 41340 -9300
rect 41460 -9420 41505 -9300
rect 41625 -9420 41670 -9300
rect 41790 -9420 41845 -9300
rect 41965 -9420 41975 -9300
rect 36475 -9465 41975 -9420
rect 36475 -9585 36485 -9465
rect 36605 -9585 36650 -9465
rect 36770 -9585 36815 -9465
rect 36935 -9585 36980 -9465
rect 37100 -9585 37155 -9465
rect 37275 -9585 37320 -9465
rect 37440 -9585 37485 -9465
rect 37605 -9585 37650 -9465
rect 37770 -9585 37825 -9465
rect 37945 -9585 37990 -9465
rect 38110 -9585 38155 -9465
rect 38275 -9585 38320 -9465
rect 38440 -9585 38495 -9465
rect 38615 -9585 38660 -9465
rect 38780 -9585 38825 -9465
rect 38945 -9585 38990 -9465
rect 39110 -9585 39165 -9465
rect 39285 -9585 39330 -9465
rect 39450 -9585 39495 -9465
rect 39615 -9585 39660 -9465
rect 39780 -9585 39835 -9465
rect 39955 -9585 40000 -9465
rect 40120 -9585 40165 -9465
rect 40285 -9585 40330 -9465
rect 40450 -9585 40505 -9465
rect 40625 -9585 40670 -9465
rect 40790 -9585 40835 -9465
rect 40955 -9585 41000 -9465
rect 41120 -9585 41175 -9465
rect 41295 -9585 41340 -9465
rect 41460 -9585 41505 -9465
rect 41625 -9585 41670 -9465
rect 41790 -9585 41845 -9465
rect 41965 -9585 41975 -9465
rect 36475 -9630 41975 -9585
rect 36475 -9750 36485 -9630
rect 36605 -9750 36650 -9630
rect 36770 -9750 36815 -9630
rect 36935 -9750 36980 -9630
rect 37100 -9750 37155 -9630
rect 37275 -9750 37320 -9630
rect 37440 -9750 37485 -9630
rect 37605 -9750 37650 -9630
rect 37770 -9750 37825 -9630
rect 37945 -9750 37990 -9630
rect 38110 -9750 38155 -9630
rect 38275 -9750 38320 -9630
rect 38440 -9750 38495 -9630
rect 38615 -9750 38660 -9630
rect 38780 -9750 38825 -9630
rect 38945 -9750 38990 -9630
rect 39110 -9750 39165 -9630
rect 39285 -9750 39330 -9630
rect 39450 -9750 39495 -9630
rect 39615 -9750 39660 -9630
rect 39780 -9750 39835 -9630
rect 39955 -9750 40000 -9630
rect 40120 -9750 40165 -9630
rect 40285 -9750 40330 -9630
rect 40450 -9750 40505 -9630
rect 40625 -9750 40670 -9630
rect 40790 -9750 40835 -9630
rect 40955 -9750 41000 -9630
rect 41120 -9750 41175 -9630
rect 41295 -9750 41340 -9630
rect 41460 -9750 41505 -9630
rect 41625 -9750 41670 -9630
rect 41790 -9750 41845 -9630
rect 41965 -9750 41975 -9630
rect 36475 -9760 41975 -9750
rect 42165 -4270 47665 -4260
rect 42165 -4390 42175 -4270
rect 42295 -4390 42340 -4270
rect 42460 -4390 42505 -4270
rect 42625 -4390 42670 -4270
rect 42790 -4390 42845 -4270
rect 42965 -4390 43010 -4270
rect 43130 -4390 43175 -4270
rect 43295 -4390 43340 -4270
rect 43460 -4390 43515 -4270
rect 43635 -4390 43680 -4270
rect 43800 -4390 43845 -4270
rect 43965 -4390 44010 -4270
rect 44130 -4390 44185 -4270
rect 44305 -4390 44350 -4270
rect 44470 -4390 44515 -4270
rect 44635 -4390 44680 -4270
rect 44800 -4390 44855 -4270
rect 44975 -4390 45020 -4270
rect 45140 -4390 45185 -4270
rect 45305 -4390 45350 -4270
rect 45470 -4390 45525 -4270
rect 45645 -4390 45690 -4270
rect 45810 -4390 45855 -4270
rect 45975 -4390 46020 -4270
rect 46140 -4390 46195 -4270
rect 46315 -4390 46360 -4270
rect 46480 -4390 46525 -4270
rect 46645 -4390 46690 -4270
rect 46810 -4390 46865 -4270
rect 46985 -4390 47030 -4270
rect 47150 -4390 47195 -4270
rect 47315 -4390 47360 -4270
rect 47480 -4390 47535 -4270
rect 47655 -4390 47665 -4270
rect 42165 -4445 47665 -4390
rect 42165 -4565 42175 -4445
rect 42295 -4565 42340 -4445
rect 42460 -4565 42505 -4445
rect 42625 -4565 42670 -4445
rect 42790 -4565 42845 -4445
rect 42965 -4565 43010 -4445
rect 43130 -4565 43175 -4445
rect 43295 -4565 43340 -4445
rect 43460 -4565 43515 -4445
rect 43635 -4565 43680 -4445
rect 43800 -4565 43845 -4445
rect 43965 -4565 44010 -4445
rect 44130 -4565 44185 -4445
rect 44305 -4565 44350 -4445
rect 44470 -4565 44515 -4445
rect 44635 -4565 44680 -4445
rect 44800 -4565 44855 -4445
rect 44975 -4565 45020 -4445
rect 45140 -4565 45185 -4445
rect 45305 -4565 45350 -4445
rect 45470 -4565 45525 -4445
rect 45645 -4565 45690 -4445
rect 45810 -4565 45855 -4445
rect 45975 -4565 46020 -4445
rect 46140 -4565 46195 -4445
rect 46315 -4565 46360 -4445
rect 46480 -4565 46525 -4445
rect 46645 -4565 46690 -4445
rect 46810 -4565 46865 -4445
rect 46985 -4565 47030 -4445
rect 47150 -4565 47195 -4445
rect 47315 -4565 47360 -4445
rect 47480 -4565 47535 -4445
rect 47655 -4565 47665 -4445
rect 42165 -4610 47665 -4565
rect 42165 -4730 42175 -4610
rect 42295 -4730 42340 -4610
rect 42460 -4730 42505 -4610
rect 42625 -4730 42670 -4610
rect 42790 -4730 42845 -4610
rect 42965 -4730 43010 -4610
rect 43130 -4730 43175 -4610
rect 43295 -4730 43340 -4610
rect 43460 -4730 43515 -4610
rect 43635 -4730 43680 -4610
rect 43800 -4730 43845 -4610
rect 43965 -4730 44010 -4610
rect 44130 -4730 44185 -4610
rect 44305 -4730 44350 -4610
rect 44470 -4730 44515 -4610
rect 44635 -4730 44680 -4610
rect 44800 -4730 44855 -4610
rect 44975 -4730 45020 -4610
rect 45140 -4730 45185 -4610
rect 45305 -4730 45350 -4610
rect 45470 -4730 45525 -4610
rect 45645 -4730 45690 -4610
rect 45810 -4730 45855 -4610
rect 45975 -4730 46020 -4610
rect 46140 -4730 46195 -4610
rect 46315 -4730 46360 -4610
rect 46480 -4730 46525 -4610
rect 46645 -4730 46690 -4610
rect 46810 -4730 46865 -4610
rect 46985 -4730 47030 -4610
rect 47150 -4730 47195 -4610
rect 47315 -4730 47360 -4610
rect 47480 -4730 47535 -4610
rect 47655 -4730 47665 -4610
rect 42165 -4775 47665 -4730
rect 42165 -4895 42175 -4775
rect 42295 -4895 42340 -4775
rect 42460 -4895 42505 -4775
rect 42625 -4895 42670 -4775
rect 42790 -4895 42845 -4775
rect 42965 -4895 43010 -4775
rect 43130 -4895 43175 -4775
rect 43295 -4895 43340 -4775
rect 43460 -4895 43515 -4775
rect 43635 -4895 43680 -4775
rect 43800 -4895 43845 -4775
rect 43965 -4895 44010 -4775
rect 44130 -4895 44185 -4775
rect 44305 -4895 44350 -4775
rect 44470 -4895 44515 -4775
rect 44635 -4895 44680 -4775
rect 44800 -4895 44855 -4775
rect 44975 -4895 45020 -4775
rect 45140 -4895 45185 -4775
rect 45305 -4895 45350 -4775
rect 45470 -4895 45525 -4775
rect 45645 -4895 45690 -4775
rect 45810 -4895 45855 -4775
rect 45975 -4895 46020 -4775
rect 46140 -4895 46195 -4775
rect 46315 -4895 46360 -4775
rect 46480 -4895 46525 -4775
rect 46645 -4895 46690 -4775
rect 46810 -4895 46865 -4775
rect 46985 -4895 47030 -4775
rect 47150 -4895 47195 -4775
rect 47315 -4895 47360 -4775
rect 47480 -4895 47535 -4775
rect 47655 -4895 47665 -4775
rect 42165 -4940 47665 -4895
rect 42165 -5060 42175 -4940
rect 42295 -5060 42340 -4940
rect 42460 -5060 42505 -4940
rect 42625 -5060 42670 -4940
rect 42790 -5060 42845 -4940
rect 42965 -5060 43010 -4940
rect 43130 -5060 43175 -4940
rect 43295 -5060 43340 -4940
rect 43460 -5060 43515 -4940
rect 43635 -5060 43680 -4940
rect 43800 -5060 43845 -4940
rect 43965 -5060 44010 -4940
rect 44130 -5060 44185 -4940
rect 44305 -5060 44350 -4940
rect 44470 -5060 44515 -4940
rect 44635 -5060 44680 -4940
rect 44800 -5060 44855 -4940
rect 44975 -5060 45020 -4940
rect 45140 -5060 45185 -4940
rect 45305 -5060 45350 -4940
rect 45470 -5060 45525 -4940
rect 45645 -5060 45690 -4940
rect 45810 -5060 45855 -4940
rect 45975 -5060 46020 -4940
rect 46140 -5060 46195 -4940
rect 46315 -5060 46360 -4940
rect 46480 -5060 46525 -4940
rect 46645 -5060 46690 -4940
rect 46810 -5060 46865 -4940
rect 46985 -5060 47030 -4940
rect 47150 -5060 47195 -4940
rect 47315 -5060 47360 -4940
rect 47480 -5060 47535 -4940
rect 47655 -5060 47665 -4940
rect 42165 -5115 47665 -5060
rect 42165 -5235 42175 -5115
rect 42295 -5235 42340 -5115
rect 42460 -5235 42505 -5115
rect 42625 -5235 42670 -5115
rect 42790 -5235 42845 -5115
rect 42965 -5235 43010 -5115
rect 43130 -5235 43175 -5115
rect 43295 -5235 43340 -5115
rect 43460 -5235 43515 -5115
rect 43635 -5235 43680 -5115
rect 43800 -5235 43845 -5115
rect 43965 -5235 44010 -5115
rect 44130 -5235 44185 -5115
rect 44305 -5235 44350 -5115
rect 44470 -5235 44515 -5115
rect 44635 -5235 44680 -5115
rect 44800 -5235 44855 -5115
rect 44975 -5235 45020 -5115
rect 45140 -5235 45185 -5115
rect 45305 -5235 45350 -5115
rect 45470 -5235 45525 -5115
rect 45645 -5235 45690 -5115
rect 45810 -5235 45855 -5115
rect 45975 -5235 46020 -5115
rect 46140 -5235 46195 -5115
rect 46315 -5235 46360 -5115
rect 46480 -5235 46525 -5115
rect 46645 -5235 46690 -5115
rect 46810 -5235 46865 -5115
rect 46985 -5235 47030 -5115
rect 47150 -5235 47195 -5115
rect 47315 -5235 47360 -5115
rect 47480 -5235 47535 -5115
rect 47655 -5235 47665 -5115
rect 42165 -5280 47665 -5235
rect 42165 -5400 42175 -5280
rect 42295 -5400 42340 -5280
rect 42460 -5400 42505 -5280
rect 42625 -5400 42670 -5280
rect 42790 -5400 42845 -5280
rect 42965 -5400 43010 -5280
rect 43130 -5400 43175 -5280
rect 43295 -5400 43340 -5280
rect 43460 -5400 43515 -5280
rect 43635 -5400 43680 -5280
rect 43800 -5400 43845 -5280
rect 43965 -5400 44010 -5280
rect 44130 -5400 44185 -5280
rect 44305 -5400 44350 -5280
rect 44470 -5400 44515 -5280
rect 44635 -5400 44680 -5280
rect 44800 -5400 44855 -5280
rect 44975 -5400 45020 -5280
rect 45140 -5400 45185 -5280
rect 45305 -5400 45350 -5280
rect 45470 -5400 45525 -5280
rect 45645 -5400 45690 -5280
rect 45810 -5400 45855 -5280
rect 45975 -5400 46020 -5280
rect 46140 -5400 46195 -5280
rect 46315 -5400 46360 -5280
rect 46480 -5400 46525 -5280
rect 46645 -5400 46690 -5280
rect 46810 -5400 46865 -5280
rect 46985 -5400 47030 -5280
rect 47150 -5400 47195 -5280
rect 47315 -5400 47360 -5280
rect 47480 -5400 47535 -5280
rect 47655 -5400 47665 -5280
rect 42165 -5445 47665 -5400
rect 42165 -5565 42175 -5445
rect 42295 -5565 42340 -5445
rect 42460 -5565 42505 -5445
rect 42625 -5565 42670 -5445
rect 42790 -5565 42845 -5445
rect 42965 -5565 43010 -5445
rect 43130 -5565 43175 -5445
rect 43295 -5565 43340 -5445
rect 43460 -5565 43515 -5445
rect 43635 -5565 43680 -5445
rect 43800 -5565 43845 -5445
rect 43965 -5565 44010 -5445
rect 44130 -5565 44185 -5445
rect 44305 -5565 44350 -5445
rect 44470 -5565 44515 -5445
rect 44635 -5565 44680 -5445
rect 44800 -5565 44855 -5445
rect 44975 -5565 45020 -5445
rect 45140 -5565 45185 -5445
rect 45305 -5565 45350 -5445
rect 45470 -5565 45525 -5445
rect 45645 -5565 45690 -5445
rect 45810 -5565 45855 -5445
rect 45975 -5565 46020 -5445
rect 46140 -5565 46195 -5445
rect 46315 -5565 46360 -5445
rect 46480 -5565 46525 -5445
rect 46645 -5565 46690 -5445
rect 46810 -5565 46865 -5445
rect 46985 -5565 47030 -5445
rect 47150 -5565 47195 -5445
rect 47315 -5565 47360 -5445
rect 47480 -5565 47535 -5445
rect 47655 -5565 47665 -5445
rect 42165 -5610 47665 -5565
rect 42165 -5730 42175 -5610
rect 42295 -5730 42340 -5610
rect 42460 -5730 42505 -5610
rect 42625 -5730 42670 -5610
rect 42790 -5730 42845 -5610
rect 42965 -5730 43010 -5610
rect 43130 -5730 43175 -5610
rect 43295 -5730 43340 -5610
rect 43460 -5730 43515 -5610
rect 43635 -5730 43680 -5610
rect 43800 -5730 43845 -5610
rect 43965 -5730 44010 -5610
rect 44130 -5730 44185 -5610
rect 44305 -5730 44350 -5610
rect 44470 -5730 44515 -5610
rect 44635 -5730 44680 -5610
rect 44800 -5730 44855 -5610
rect 44975 -5730 45020 -5610
rect 45140 -5730 45185 -5610
rect 45305 -5730 45350 -5610
rect 45470 -5730 45525 -5610
rect 45645 -5730 45690 -5610
rect 45810 -5730 45855 -5610
rect 45975 -5730 46020 -5610
rect 46140 -5730 46195 -5610
rect 46315 -5730 46360 -5610
rect 46480 -5730 46525 -5610
rect 46645 -5730 46690 -5610
rect 46810 -5730 46865 -5610
rect 46985 -5730 47030 -5610
rect 47150 -5730 47195 -5610
rect 47315 -5730 47360 -5610
rect 47480 -5730 47535 -5610
rect 47655 -5730 47665 -5610
rect 42165 -5785 47665 -5730
rect 42165 -5905 42175 -5785
rect 42295 -5905 42340 -5785
rect 42460 -5905 42505 -5785
rect 42625 -5905 42670 -5785
rect 42790 -5905 42845 -5785
rect 42965 -5905 43010 -5785
rect 43130 -5905 43175 -5785
rect 43295 -5905 43340 -5785
rect 43460 -5905 43515 -5785
rect 43635 -5905 43680 -5785
rect 43800 -5905 43845 -5785
rect 43965 -5905 44010 -5785
rect 44130 -5905 44185 -5785
rect 44305 -5905 44350 -5785
rect 44470 -5905 44515 -5785
rect 44635 -5905 44680 -5785
rect 44800 -5905 44855 -5785
rect 44975 -5905 45020 -5785
rect 45140 -5905 45185 -5785
rect 45305 -5905 45350 -5785
rect 45470 -5905 45525 -5785
rect 45645 -5905 45690 -5785
rect 45810 -5905 45855 -5785
rect 45975 -5905 46020 -5785
rect 46140 -5905 46195 -5785
rect 46315 -5905 46360 -5785
rect 46480 -5905 46525 -5785
rect 46645 -5905 46690 -5785
rect 46810 -5905 46865 -5785
rect 46985 -5905 47030 -5785
rect 47150 -5905 47195 -5785
rect 47315 -5905 47360 -5785
rect 47480 -5905 47535 -5785
rect 47655 -5905 47665 -5785
rect 42165 -5950 47665 -5905
rect 42165 -6070 42175 -5950
rect 42295 -6070 42340 -5950
rect 42460 -6070 42505 -5950
rect 42625 -6070 42670 -5950
rect 42790 -6070 42845 -5950
rect 42965 -6070 43010 -5950
rect 43130 -6070 43175 -5950
rect 43295 -6070 43340 -5950
rect 43460 -6070 43515 -5950
rect 43635 -6070 43680 -5950
rect 43800 -6070 43845 -5950
rect 43965 -6070 44010 -5950
rect 44130 -6070 44185 -5950
rect 44305 -6070 44350 -5950
rect 44470 -6070 44515 -5950
rect 44635 -6070 44680 -5950
rect 44800 -6070 44855 -5950
rect 44975 -6070 45020 -5950
rect 45140 -6070 45185 -5950
rect 45305 -6070 45350 -5950
rect 45470 -6070 45525 -5950
rect 45645 -6070 45690 -5950
rect 45810 -6070 45855 -5950
rect 45975 -6070 46020 -5950
rect 46140 -6070 46195 -5950
rect 46315 -6070 46360 -5950
rect 46480 -6070 46525 -5950
rect 46645 -6070 46690 -5950
rect 46810 -6070 46865 -5950
rect 46985 -6070 47030 -5950
rect 47150 -6070 47195 -5950
rect 47315 -6070 47360 -5950
rect 47480 -6070 47535 -5950
rect 47655 -6070 47665 -5950
rect 42165 -6115 47665 -6070
rect 42165 -6235 42175 -6115
rect 42295 -6235 42340 -6115
rect 42460 -6235 42505 -6115
rect 42625 -6235 42670 -6115
rect 42790 -6235 42845 -6115
rect 42965 -6235 43010 -6115
rect 43130 -6235 43175 -6115
rect 43295 -6235 43340 -6115
rect 43460 -6235 43515 -6115
rect 43635 -6235 43680 -6115
rect 43800 -6235 43845 -6115
rect 43965 -6235 44010 -6115
rect 44130 -6235 44185 -6115
rect 44305 -6235 44350 -6115
rect 44470 -6235 44515 -6115
rect 44635 -6235 44680 -6115
rect 44800 -6235 44855 -6115
rect 44975 -6235 45020 -6115
rect 45140 -6235 45185 -6115
rect 45305 -6235 45350 -6115
rect 45470 -6235 45525 -6115
rect 45645 -6235 45690 -6115
rect 45810 -6235 45855 -6115
rect 45975 -6235 46020 -6115
rect 46140 -6235 46195 -6115
rect 46315 -6235 46360 -6115
rect 46480 -6235 46525 -6115
rect 46645 -6235 46690 -6115
rect 46810 -6235 46865 -6115
rect 46985 -6235 47030 -6115
rect 47150 -6235 47195 -6115
rect 47315 -6235 47360 -6115
rect 47480 -6235 47535 -6115
rect 47655 -6235 47665 -6115
rect 42165 -6280 47665 -6235
rect 42165 -6400 42175 -6280
rect 42295 -6400 42340 -6280
rect 42460 -6400 42505 -6280
rect 42625 -6400 42670 -6280
rect 42790 -6400 42845 -6280
rect 42965 -6400 43010 -6280
rect 43130 -6400 43175 -6280
rect 43295 -6400 43340 -6280
rect 43460 -6400 43515 -6280
rect 43635 -6400 43680 -6280
rect 43800 -6400 43845 -6280
rect 43965 -6400 44010 -6280
rect 44130 -6400 44185 -6280
rect 44305 -6400 44350 -6280
rect 44470 -6400 44515 -6280
rect 44635 -6400 44680 -6280
rect 44800 -6400 44855 -6280
rect 44975 -6400 45020 -6280
rect 45140 -6400 45185 -6280
rect 45305 -6400 45350 -6280
rect 45470 -6400 45525 -6280
rect 45645 -6400 45690 -6280
rect 45810 -6400 45855 -6280
rect 45975 -6400 46020 -6280
rect 46140 -6400 46195 -6280
rect 46315 -6400 46360 -6280
rect 46480 -6400 46525 -6280
rect 46645 -6400 46690 -6280
rect 46810 -6400 46865 -6280
rect 46985 -6400 47030 -6280
rect 47150 -6400 47195 -6280
rect 47315 -6400 47360 -6280
rect 47480 -6400 47535 -6280
rect 47655 -6400 47665 -6280
rect 42165 -6455 47665 -6400
rect 42165 -6575 42175 -6455
rect 42295 -6575 42340 -6455
rect 42460 -6575 42505 -6455
rect 42625 -6575 42670 -6455
rect 42790 -6575 42845 -6455
rect 42965 -6575 43010 -6455
rect 43130 -6575 43175 -6455
rect 43295 -6575 43340 -6455
rect 43460 -6575 43515 -6455
rect 43635 -6575 43680 -6455
rect 43800 -6575 43845 -6455
rect 43965 -6575 44010 -6455
rect 44130 -6575 44185 -6455
rect 44305 -6575 44350 -6455
rect 44470 -6575 44515 -6455
rect 44635 -6575 44680 -6455
rect 44800 -6575 44855 -6455
rect 44975 -6575 45020 -6455
rect 45140 -6575 45185 -6455
rect 45305 -6575 45350 -6455
rect 45470 -6575 45525 -6455
rect 45645 -6575 45690 -6455
rect 45810 -6575 45855 -6455
rect 45975 -6575 46020 -6455
rect 46140 -6575 46195 -6455
rect 46315 -6575 46360 -6455
rect 46480 -6575 46525 -6455
rect 46645 -6575 46690 -6455
rect 46810 -6575 46865 -6455
rect 46985 -6575 47030 -6455
rect 47150 -6575 47195 -6455
rect 47315 -6575 47360 -6455
rect 47480 -6575 47535 -6455
rect 47655 -6575 47665 -6455
rect 42165 -6620 47665 -6575
rect 42165 -6740 42175 -6620
rect 42295 -6740 42340 -6620
rect 42460 -6740 42505 -6620
rect 42625 -6740 42670 -6620
rect 42790 -6740 42845 -6620
rect 42965 -6740 43010 -6620
rect 43130 -6740 43175 -6620
rect 43295 -6740 43340 -6620
rect 43460 -6740 43515 -6620
rect 43635 -6740 43680 -6620
rect 43800 -6740 43845 -6620
rect 43965 -6740 44010 -6620
rect 44130 -6740 44185 -6620
rect 44305 -6740 44350 -6620
rect 44470 -6740 44515 -6620
rect 44635 -6740 44680 -6620
rect 44800 -6740 44855 -6620
rect 44975 -6740 45020 -6620
rect 45140 -6740 45185 -6620
rect 45305 -6740 45350 -6620
rect 45470 -6740 45525 -6620
rect 45645 -6740 45690 -6620
rect 45810 -6740 45855 -6620
rect 45975 -6740 46020 -6620
rect 46140 -6740 46195 -6620
rect 46315 -6740 46360 -6620
rect 46480 -6740 46525 -6620
rect 46645 -6740 46690 -6620
rect 46810 -6740 46865 -6620
rect 46985 -6740 47030 -6620
rect 47150 -6740 47195 -6620
rect 47315 -6740 47360 -6620
rect 47480 -6740 47535 -6620
rect 47655 -6740 47665 -6620
rect 42165 -6785 47665 -6740
rect 42165 -6905 42175 -6785
rect 42295 -6905 42340 -6785
rect 42460 -6905 42505 -6785
rect 42625 -6905 42670 -6785
rect 42790 -6905 42845 -6785
rect 42965 -6905 43010 -6785
rect 43130 -6905 43175 -6785
rect 43295 -6905 43340 -6785
rect 43460 -6905 43515 -6785
rect 43635 -6905 43680 -6785
rect 43800 -6905 43845 -6785
rect 43965 -6905 44010 -6785
rect 44130 -6905 44185 -6785
rect 44305 -6905 44350 -6785
rect 44470 -6905 44515 -6785
rect 44635 -6905 44680 -6785
rect 44800 -6905 44855 -6785
rect 44975 -6905 45020 -6785
rect 45140 -6905 45185 -6785
rect 45305 -6905 45350 -6785
rect 45470 -6905 45525 -6785
rect 45645 -6905 45690 -6785
rect 45810 -6905 45855 -6785
rect 45975 -6905 46020 -6785
rect 46140 -6905 46195 -6785
rect 46315 -6905 46360 -6785
rect 46480 -6905 46525 -6785
rect 46645 -6905 46690 -6785
rect 46810 -6905 46865 -6785
rect 46985 -6905 47030 -6785
rect 47150 -6905 47195 -6785
rect 47315 -6905 47360 -6785
rect 47480 -6905 47535 -6785
rect 47655 -6905 47665 -6785
rect 42165 -6950 47665 -6905
rect 42165 -7070 42175 -6950
rect 42295 -7070 42340 -6950
rect 42460 -7070 42505 -6950
rect 42625 -7070 42670 -6950
rect 42790 -7070 42845 -6950
rect 42965 -7070 43010 -6950
rect 43130 -7070 43175 -6950
rect 43295 -7070 43340 -6950
rect 43460 -7070 43515 -6950
rect 43635 -7070 43680 -6950
rect 43800 -7070 43845 -6950
rect 43965 -7070 44010 -6950
rect 44130 -7070 44185 -6950
rect 44305 -7070 44350 -6950
rect 44470 -7070 44515 -6950
rect 44635 -7070 44680 -6950
rect 44800 -7070 44855 -6950
rect 44975 -7070 45020 -6950
rect 45140 -7070 45185 -6950
rect 45305 -7070 45350 -6950
rect 45470 -7070 45525 -6950
rect 45645 -7070 45690 -6950
rect 45810 -7070 45855 -6950
rect 45975 -7070 46020 -6950
rect 46140 -7070 46195 -6950
rect 46315 -7070 46360 -6950
rect 46480 -7070 46525 -6950
rect 46645 -7070 46690 -6950
rect 46810 -7070 46865 -6950
rect 46985 -7070 47030 -6950
rect 47150 -7070 47195 -6950
rect 47315 -7070 47360 -6950
rect 47480 -7070 47535 -6950
rect 47655 -7070 47665 -6950
rect 42165 -7125 47665 -7070
rect 42165 -7245 42175 -7125
rect 42295 -7245 42340 -7125
rect 42460 -7245 42505 -7125
rect 42625 -7245 42670 -7125
rect 42790 -7245 42845 -7125
rect 42965 -7245 43010 -7125
rect 43130 -7245 43175 -7125
rect 43295 -7245 43340 -7125
rect 43460 -7245 43515 -7125
rect 43635 -7245 43680 -7125
rect 43800 -7245 43845 -7125
rect 43965 -7245 44010 -7125
rect 44130 -7245 44185 -7125
rect 44305 -7245 44350 -7125
rect 44470 -7245 44515 -7125
rect 44635 -7245 44680 -7125
rect 44800 -7245 44855 -7125
rect 44975 -7245 45020 -7125
rect 45140 -7245 45185 -7125
rect 45305 -7245 45350 -7125
rect 45470 -7245 45525 -7125
rect 45645 -7245 45690 -7125
rect 45810 -7245 45855 -7125
rect 45975 -7245 46020 -7125
rect 46140 -7245 46195 -7125
rect 46315 -7245 46360 -7125
rect 46480 -7245 46525 -7125
rect 46645 -7245 46690 -7125
rect 46810 -7245 46865 -7125
rect 46985 -7245 47030 -7125
rect 47150 -7245 47195 -7125
rect 47315 -7245 47360 -7125
rect 47480 -7245 47535 -7125
rect 47655 -7245 47665 -7125
rect 42165 -7290 47665 -7245
rect 42165 -7410 42175 -7290
rect 42295 -7410 42340 -7290
rect 42460 -7410 42505 -7290
rect 42625 -7410 42670 -7290
rect 42790 -7410 42845 -7290
rect 42965 -7410 43010 -7290
rect 43130 -7410 43175 -7290
rect 43295 -7410 43340 -7290
rect 43460 -7410 43515 -7290
rect 43635 -7410 43680 -7290
rect 43800 -7410 43845 -7290
rect 43965 -7410 44010 -7290
rect 44130 -7410 44185 -7290
rect 44305 -7410 44350 -7290
rect 44470 -7410 44515 -7290
rect 44635 -7410 44680 -7290
rect 44800 -7410 44855 -7290
rect 44975 -7410 45020 -7290
rect 45140 -7410 45185 -7290
rect 45305 -7410 45350 -7290
rect 45470 -7410 45525 -7290
rect 45645 -7410 45690 -7290
rect 45810 -7410 45855 -7290
rect 45975 -7410 46020 -7290
rect 46140 -7410 46195 -7290
rect 46315 -7410 46360 -7290
rect 46480 -7410 46525 -7290
rect 46645 -7410 46690 -7290
rect 46810 -7410 46865 -7290
rect 46985 -7410 47030 -7290
rect 47150 -7410 47195 -7290
rect 47315 -7410 47360 -7290
rect 47480 -7410 47535 -7290
rect 47655 -7410 47665 -7290
rect 42165 -7455 47665 -7410
rect 42165 -7575 42175 -7455
rect 42295 -7575 42340 -7455
rect 42460 -7575 42505 -7455
rect 42625 -7575 42670 -7455
rect 42790 -7575 42845 -7455
rect 42965 -7575 43010 -7455
rect 43130 -7575 43175 -7455
rect 43295 -7575 43340 -7455
rect 43460 -7575 43515 -7455
rect 43635 -7575 43680 -7455
rect 43800 -7575 43845 -7455
rect 43965 -7575 44010 -7455
rect 44130 -7575 44185 -7455
rect 44305 -7575 44350 -7455
rect 44470 -7575 44515 -7455
rect 44635 -7575 44680 -7455
rect 44800 -7575 44855 -7455
rect 44975 -7575 45020 -7455
rect 45140 -7575 45185 -7455
rect 45305 -7575 45350 -7455
rect 45470 -7575 45525 -7455
rect 45645 -7575 45690 -7455
rect 45810 -7575 45855 -7455
rect 45975 -7575 46020 -7455
rect 46140 -7575 46195 -7455
rect 46315 -7575 46360 -7455
rect 46480 -7575 46525 -7455
rect 46645 -7575 46690 -7455
rect 46810 -7575 46865 -7455
rect 46985 -7575 47030 -7455
rect 47150 -7575 47195 -7455
rect 47315 -7575 47360 -7455
rect 47480 -7575 47535 -7455
rect 47655 -7575 47665 -7455
rect 42165 -7620 47665 -7575
rect 42165 -7740 42175 -7620
rect 42295 -7740 42340 -7620
rect 42460 -7740 42505 -7620
rect 42625 -7740 42670 -7620
rect 42790 -7740 42845 -7620
rect 42965 -7740 43010 -7620
rect 43130 -7740 43175 -7620
rect 43295 -7740 43340 -7620
rect 43460 -7740 43515 -7620
rect 43635 -7740 43680 -7620
rect 43800 -7740 43845 -7620
rect 43965 -7740 44010 -7620
rect 44130 -7740 44185 -7620
rect 44305 -7740 44350 -7620
rect 44470 -7740 44515 -7620
rect 44635 -7740 44680 -7620
rect 44800 -7740 44855 -7620
rect 44975 -7740 45020 -7620
rect 45140 -7740 45185 -7620
rect 45305 -7740 45350 -7620
rect 45470 -7740 45525 -7620
rect 45645 -7740 45690 -7620
rect 45810 -7740 45855 -7620
rect 45975 -7740 46020 -7620
rect 46140 -7740 46195 -7620
rect 46315 -7740 46360 -7620
rect 46480 -7740 46525 -7620
rect 46645 -7740 46690 -7620
rect 46810 -7740 46865 -7620
rect 46985 -7740 47030 -7620
rect 47150 -7740 47195 -7620
rect 47315 -7740 47360 -7620
rect 47480 -7740 47535 -7620
rect 47655 -7740 47665 -7620
rect 42165 -7795 47665 -7740
rect 42165 -7915 42175 -7795
rect 42295 -7915 42340 -7795
rect 42460 -7915 42505 -7795
rect 42625 -7915 42670 -7795
rect 42790 -7915 42845 -7795
rect 42965 -7915 43010 -7795
rect 43130 -7915 43175 -7795
rect 43295 -7915 43340 -7795
rect 43460 -7915 43515 -7795
rect 43635 -7915 43680 -7795
rect 43800 -7915 43845 -7795
rect 43965 -7915 44010 -7795
rect 44130 -7915 44185 -7795
rect 44305 -7915 44350 -7795
rect 44470 -7915 44515 -7795
rect 44635 -7915 44680 -7795
rect 44800 -7915 44855 -7795
rect 44975 -7915 45020 -7795
rect 45140 -7915 45185 -7795
rect 45305 -7915 45350 -7795
rect 45470 -7915 45525 -7795
rect 45645 -7915 45690 -7795
rect 45810 -7915 45855 -7795
rect 45975 -7915 46020 -7795
rect 46140 -7915 46195 -7795
rect 46315 -7915 46360 -7795
rect 46480 -7915 46525 -7795
rect 46645 -7915 46690 -7795
rect 46810 -7915 46865 -7795
rect 46985 -7915 47030 -7795
rect 47150 -7915 47195 -7795
rect 47315 -7915 47360 -7795
rect 47480 -7915 47535 -7795
rect 47655 -7915 47665 -7795
rect 42165 -7960 47665 -7915
rect 42165 -8080 42175 -7960
rect 42295 -8080 42340 -7960
rect 42460 -8080 42505 -7960
rect 42625 -8080 42670 -7960
rect 42790 -8080 42845 -7960
rect 42965 -8080 43010 -7960
rect 43130 -8080 43175 -7960
rect 43295 -8080 43340 -7960
rect 43460 -8080 43515 -7960
rect 43635 -8080 43680 -7960
rect 43800 -8080 43845 -7960
rect 43965 -8080 44010 -7960
rect 44130 -8080 44185 -7960
rect 44305 -8080 44350 -7960
rect 44470 -8080 44515 -7960
rect 44635 -8080 44680 -7960
rect 44800 -8080 44855 -7960
rect 44975 -8080 45020 -7960
rect 45140 -8080 45185 -7960
rect 45305 -8080 45350 -7960
rect 45470 -8080 45525 -7960
rect 45645 -8080 45690 -7960
rect 45810 -8080 45855 -7960
rect 45975 -8080 46020 -7960
rect 46140 -8080 46195 -7960
rect 46315 -8080 46360 -7960
rect 46480 -8080 46525 -7960
rect 46645 -8080 46690 -7960
rect 46810 -8080 46865 -7960
rect 46985 -8080 47030 -7960
rect 47150 -8080 47195 -7960
rect 47315 -8080 47360 -7960
rect 47480 -8080 47535 -7960
rect 47655 -8080 47665 -7960
rect 42165 -8125 47665 -8080
rect 42165 -8245 42175 -8125
rect 42295 -8245 42340 -8125
rect 42460 -8245 42505 -8125
rect 42625 -8245 42670 -8125
rect 42790 -8245 42845 -8125
rect 42965 -8245 43010 -8125
rect 43130 -8245 43175 -8125
rect 43295 -8245 43340 -8125
rect 43460 -8245 43515 -8125
rect 43635 -8245 43680 -8125
rect 43800 -8245 43845 -8125
rect 43965 -8245 44010 -8125
rect 44130 -8245 44185 -8125
rect 44305 -8245 44350 -8125
rect 44470 -8245 44515 -8125
rect 44635 -8245 44680 -8125
rect 44800 -8245 44855 -8125
rect 44975 -8245 45020 -8125
rect 45140 -8245 45185 -8125
rect 45305 -8245 45350 -8125
rect 45470 -8245 45525 -8125
rect 45645 -8245 45690 -8125
rect 45810 -8245 45855 -8125
rect 45975 -8245 46020 -8125
rect 46140 -8245 46195 -8125
rect 46315 -8245 46360 -8125
rect 46480 -8245 46525 -8125
rect 46645 -8245 46690 -8125
rect 46810 -8245 46865 -8125
rect 46985 -8245 47030 -8125
rect 47150 -8245 47195 -8125
rect 47315 -8245 47360 -8125
rect 47480 -8245 47535 -8125
rect 47655 -8245 47665 -8125
rect 42165 -8290 47665 -8245
rect 42165 -8410 42175 -8290
rect 42295 -8410 42340 -8290
rect 42460 -8410 42505 -8290
rect 42625 -8410 42670 -8290
rect 42790 -8410 42845 -8290
rect 42965 -8410 43010 -8290
rect 43130 -8410 43175 -8290
rect 43295 -8410 43340 -8290
rect 43460 -8410 43515 -8290
rect 43635 -8410 43680 -8290
rect 43800 -8410 43845 -8290
rect 43965 -8410 44010 -8290
rect 44130 -8410 44185 -8290
rect 44305 -8410 44350 -8290
rect 44470 -8410 44515 -8290
rect 44635 -8410 44680 -8290
rect 44800 -8410 44855 -8290
rect 44975 -8410 45020 -8290
rect 45140 -8410 45185 -8290
rect 45305 -8410 45350 -8290
rect 45470 -8410 45525 -8290
rect 45645 -8410 45690 -8290
rect 45810 -8410 45855 -8290
rect 45975 -8410 46020 -8290
rect 46140 -8410 46195 -8290
rect 46315 -8410 46360 -8290
rect 46480 -8410 46525 -8290
rect 46645 -8410 46690 -8290
rect 46810 -8410 46865 -8290
rect 46985 -8410 47030 -8290
rect 47150 -8410 47195 -8290
rect 47315 -8410 47360 -8290
rect 47480 -8410 47535 -8290
rect 47655 -8410 47665 -8290
rect 42165 -8465 47665 -8410
rect 42165 -8585 42175 -8465
rect 42295 -8585 42340 -8465
rect 42460 -8585 42505 -8465
rect 42625 -8585 42670 -8465
rect 42790 -8585 42845 -8465
rect 42965 -8585 43010 -8465
rect 43130 -8585 43175 -8465
rect 43295 -8585 43340 -8465
rect 43460 -8585 43515 -8465
rect 43635 -8585 43680 -8465
rect 43800 -8585 43845 -8465
rect 43965 -8585 44010 -8465
rect 44130 -8585 44185 -8465
rect 44305 -8585 44350 -8465
rect 44470 -8585 44515 -8465
rect 44635 -8585 44680 -8465
rect 44800 -8585 44855 -8465
rect 44975 -8585 45020 -8465
rect 45140 -8585 45185 -8465
rect 45305 -8585 45350 -8465
rect 45470 -8585 45525 -8465
rect 45645 -8585 45690 -8465
rect 45810 -8585 45855 -8465
rect 45975 -8585 46020 -8465
rect 46140 -8585 46195 -8465
rect 46315 -8585 46360 -8465
rect 46480 -8585 46525 -8465
rect 46645 -8585 46690 -8465
rect 46810 -8585 46865 -8465
rect 46985 -8585 47030 -8465
rect 47150 -8585 47195 -8465
rect 47315 -8585 47360 -8465
rect 47480 -8585 47535 -8465
rect 47655 -8585 47665 -8465
rect 42165 -8630 47665 -8585
rect 42165 -8750 42175 -8630
rect 42295 -8750 42340 -8630
rect 42460 -8750 42505 -8630
rect 42625 -8750 42670 -8630
rect 42790 -8750 42845 -8630
rect 42965 -8750 43010 -8630
rect 43130 -8750 43175 -8630
rect 43295 -8750 43340 -8630
rect 43460 -8750 43515 -8630
rect 43635 -8750 43680 -8630
rect 43800 -8750 43845 -8630
rect 43965 -8750 44010 -8630
rect 44130 -8750 44185 -8630
rect 44305 -8750 44350 -8630
rect 44470 -8750 44515 -8630
rect 44635 -8750 44680 -8630
rect 44800 -8750 44855 -8630
rect 44975 -8750 45020 -8630
rect 45140 -8750 45185 -8630
rect 45305 -8750 45350 -8630
rect 45470 -8750 45525 -8630
rect 45645 -8750 45690 -8630
rect 45810 -8750 45855 -8630
rect 45975 -8750 46020 -8630
rect 46140 -8750 46195 -8630
rect 46315 -8750 46360 -8630
rect 46480 -8750 46525 -8630
rect 46645 -8750 46690 -8630
rect 46810 -8750 46865 -8630
rect 46985 -8750 47030 -8630
rect 47150 -8750 47195 -8630
rect 47315 -8750 47360 -8630
rect 47480 -8750 47535 -8630
rect 47655 -8750 47665 -8630
rect 42165 -8795 47665 -8750
rect 42165 -8915 42175 -8795
rect 42295 -8915 42340 -8795
rect 42460 -8915 42505 -8795
rect 42625 -8915 42670 -8795
rect 42790 -8915 42845 -8795
rect 42965 -8915 43010 -8795
rect 43130 -8915 43175 -8795
rect 43295 -8915 43340 -8795
rect 43460 -8915 43515 -8795
rect 43635 -8915 43680 -8795
rect 43800 -8915 43845 -8795
rect 43965 -8915 44010 -8795
rect 44130 -8915 44185 -8795
rect 44305 -8915 44350 -8795
rect 44470 -8915 44515 -8795
rect 44635 -8915 44680 -8795
rect 44800 -8915 44855 -8795
rect 44975 -8915 45020 -8795
rect 45140 -8915 45185 -8795
rect 45305 -8915 45350 -8795
rect 45470 -8915 45525 -8795
rect 45645 -8915 45690 -8795
rect 45810 -8915 45855 -8795
rect 45975 -8915 46020 -8795
rect 46140 -8915 46195 -8795
rect 46315 -8915 46360 -8795
rect 46480 -8915 46525 -8795
rect 46645 -8915 46690 -8795
rect 46810 -8915 46865 -8795
rect 46985 -8915 47030 -8795
rect 47150 -8915 47195 -8795
rect 47315 -8915 47360 -8795
rect 47480 -8915 47535 -8795
rect 47655 -8915 47665 -8795
rect 42165 -8960 47665 -8915
rect 42165 -9080 42175 -8960
rect 42295 -9080 42340 -8960
rect 42460 -9080 42505 -8960
rect 42625 -9080 42670 -8960
rect 42790 -9080 42845 -8960
rect 42965 -9080 43010 -8960
rect 43130 -9080 43175 -8960
rect 43295 -9080 43340 -8960
rect 43460 -9080 43515 -8960
rect 43635 -9080 43680 -8960
rect 43800 -9080 43845 -8960
rect 43965 -9080 44010 -8960
rect 44130 -9080 44185 -8960
rect 44305 -9080 44350 -8960
rect 44470 -9080 44515 -8960
rect 44635 -9080 44680 -8960
rect 44800 -9080 44855 -8960
rect 44975 -9080 45020 -8960
rect 45140 -9080 45185 -8960
rect 45305 -9080 45350 -8960
rect 45470 -9080 45525 -8960
rect 45645 -9080 45690 -8960
rect 45810 -9080 45855 -8960
rect 45975 -9080 46020 -8960
rect 46140 -9080 46195 -8960
rect 46315 -9080 46360 -8960
rect 46480 -9080 46525 -8960
rect 46645 -9080 46690 -8960
rect 46810 -9080 46865 -8960
rect 46985 -9080 47030 -8960
rect 47150 -9080 47195 -8960
rect 47315 -9080 47360 -8960
rect 47480 -9080 47535 -8960
rect 47655 -9080 47665 -8960
rect 42165 -9135 47665 -9080
rect 42165 -9255 42175 -9135
rect 42295 -9255 42340 -9135
rect 42460 -9255 42505 -9135
rect 42625 -9255 42670 -9135
rect 42790 -9255 42845 -9135
rect 42965 -9255 43010 -9135
rect 43130 -9255 43175 -9135
rect 43295 -9255 43340 -9135
rect 43460 -9255 43515 -9135
rect 43635 -9255 43680 -9135
rect 43800 -9255 43845 -9135
rect 43965 -9255 44010 -9135
rect 44130 -9255 44185 -9135
rect 44305 -9255 44350 -9135
rect 44470 -9255 44515 -9135
rect 44635 -9255 44680 -9135
rect 44800 -9255 44855 -9135
rect 44975 -9255 45020 -9135
rect 45140 -9255 45185 -9135
rect 45305 -9255 45350 -9135
rect 45470 -9255 45525 -9135
rect 45645 -9255 45690 -9135
rect 45810 -9255 45855 -9135
rect 45975 -9255 46020 -9135
rect 46140 -9255 46195 -9135
rect 46315 -9255 46360 -9135
rect 46480 -9255 46525 -9135
rect 46645 -9255 46690 -9135
rect 46810 -9255 46865 -9135
rect 46985 -9255 47030 -9135
rect 47150 -9255 47195 -9135
rect 47315 -9255 47360 -9135
rect 47480 -9255 47535 -9135
rect 47655 -9255 47665 -9135
rect 42165 -9300 47665 -9255
rect 42165 -9420 42175 -9300
rect 42295 -9420 42340 -9300
rect 42460 -9420 42505 -9300
rect 42625 -9420 42670 -9300
rect 42790 -9420 42845 -9300
rect 42965 -9420 43010 -9300
rect 43130 -9420 43175 -9300
rect 43295 -9420 43340 -9300
rect 43460 -9420 43515 -9300
rect 43635 -9420 43680 -9300
rect 43800 -9420 43845 -9300
rect 43965 -9420 44010 -9300
rect 44130 -9420 44185 -9300
rect 44305 -9420 44350 -9300
rect 44470 -9420 44515 -9300
rect 44635 -9420 44680 -9300
rect 44800 -9420 44855 -9300
rect 44975 -9420 45020 -9300
rect 45140 -9420 45185 -9300
rect 45305 -9420 45350 -9300
rect 45470 -9420 45525 -9300
rect 45645 -9420 45690 -9300
rect 45810 -9420 45855 -9300
rect 45975 -9420 46020 -9300
rect 46140 -9420 46195 -9300
rect 46315 -9420 46360 -9300
rect 46480 -9420 46525 -9300
rect 46645 -9420 46690 -9300
rect 46810 -9420 46865 -9300
rect 46985 -9420 47030 -9300
rect 47150 -9420 47195 -9300
rect 47315 -9420 47360 -9300
rect 47480 -9420 47535 -9300
rect 47655 -9420 47665 -9300
rect 42165 -9465 47665 -9420
rect 42165 -9585 42175 -9465
rect 42295 -9585 42340 -9465
rect 42460 -9585 42505 -9465
rect 42625 -9585 42670 -9465
rect 42790 -9585 42845 -9465
rect 42965 -9585 43010 -9465
rect 43130 -9585 43175 -9465
rect 43295 -9585 43340 -9465
rect 43460 -9585 43515 -9465
rect 43635 -9585 43680 -9465
rect 43800 -9585 43845 -9465
rect 43965 -9585 44010 -9465
rect 44130 -9585 44185 -9465
rect 44305 -9585 44350 -9465
rect 44470 -9585 44515 -9465
rect 44635 -9585 44680 -9465
rect 44800 -9585 44855 -9465
rect 44975 -9585 45020 -9465
rect 45140 -9585 45185 -9465
rect 45305 -9585 45350 -9465
rect 45470 -9585 45525 -9465
rect 45645 -9585 45690 -9465
rect 45810 -9585 45855 -9465
rect 45975 -9585 46020 -9465
rect 46140 -9585 46195 -9465
rect 46315 -9585 46360 -9465
rect 46480 -9585 46525 -9465
rect 46645 -9585 46690 -9465
rect 46810 -9585 46865 -9465
rect 46985 -9585 47030 -9465
rect 47150 -9585 47195 -9465
rect 47315 -9585 47360 -9465
rect 47480 -9585 47535 -9465
rect 47655 -9585 47665 -9465
rect 42165 -9630 47665 -9585
rect 42165 -9750 42175 -9630
rect 42295 -9750 42340 -9630
rect 42460 -9750 42505 -9630
rect 42625 -9750 42670 -9630
rect 42790 -9750 42845 -9630
rect 42965 -9750 43010 -9630
rect 43130 -9750 43175 -9630
rect 43295 -9750 43340 -9630
rect 43460 -9750 43515 -9630
rect 43635 -9750 43680 -9630
rect 43800 -9750 43845 -9630
rect 43965 -9750 44010 -9630
rect 44130 -9750 44185 -9630
rect 44305 -9750 44350 -9630
rect 44470 -9750 44515 -9630
rect 44635 -9750 44680 -9630
rect 44800 -9750 44855 -9630
rect 44975 -9750 45020 -9630
rect 45140 -9750 45185 -9630
rect 45305 -9750 45350 -9630
rect 45470 -9750 45525 -9630
rect 45645 -9750 45690 -9630
rect 45810 -9750 45855 -9630
rect 45975 -9750 46020 -9630
rect 46140 -9750 46195 -9630
rect 46315 -9750 46360 -9630
rect 46480 -9750 46525 -9630
rect 46645 -9750 46690 -9630
rect 46810 -9750 46865 -9630
rect 46985 -9750 47030 -9630
rect 47150 -9750 47195 -9630
rect 47315 -9750 47360 -9630
rect 47480 -9750 47535 -9630
rect 47655 -9750 47665 -9630
rect 42165 -9760 47665 -9750
rect 47855 -4270 53355 -4260
rect 47855 -4390 47865 -4270
rect 47985 -4390 48030 -4270
rect 48150 -4390 48195 -4270
rect 48315 -4390 48360 -4270
rect 48480 -4390 48535 -4270
rect 48655 -4390 48700 -4270
rect 48820 -4390 48865 -4270
rect 48985 -4390 49030 -4270
rect 49150 -4390 49205 -4270
rect 49325 -4390 49370 -4270
rect 49490 -4390 49535 -4270
rect 49655 -4390 49700 -4270
rect 49820 -4390 49875 -4270
rect 49995 -4390 50040 -4270
rect 50160 -4390 50205 -4270
rect 50325 -4390 50370 -4270
rect 50490 -4390 50545 -4270
rect 50665 -4390 50710 -4270
rect 50830 -4390 50875 -4270
rect 50995 -4390 51040 -4270
rect 51160 -4390 51215 -4270
rect 51335 -4390 51380 -4270
rect 51500 -4390 51545 -4270
rect 51665 -4390 51710 -4270
rect 51830 -4390 51885 -4270
rect 52005 -4390 52050 -4270
rect 52170 -4390 52215 -4270
rect 52335 -4390 52380 -4270
rect 52500 -4390 52555 -4270
rect 52675 -4390 52720 -4270
rect 52840 -4390 52885 -4270
rect 53005 -4390 53050 -4270
rect 53170 -4390 53225 -4270
rect 53345 -4390 53355 -4270
rect 47855 -4445 53355 -4390
rect 47855 -4565 47865 -4445
rect 47985 -4565 48030 -4445
rect 48150 -4565 48195 -4445
rect 48315 -4565 48360 -4445
rect 48480 -4565 48535 -4445
rect 48655 -4565 48700 -4445
rect 48820 -4565 48865 -4445
rect 48985 -4565 49030 -4445
rect 49150 -4565 49205 -4445
rect 49325 -4565 49370 -4445
rect 49490 -4565 49535 -4445
rect 49655 -4565 49700 -4445
rect 49820 -4565 49875 -4445
rect 49995 -4565 50040 -4445
rect 50160 -4565 50205 -4445
rect 50325 -4565 50370 -4445
rect 50490 -4565 50545 -4445
rect 50665 -4565 50710 -4445
rect 50830 -4565 50875 -4445
rect 50995 -4565 51040 -4445
rect 51160 -4565 51215 -4445
rect 51335 -4565 51380 -4445
rect 51500 -4565 51545 -4445
rect 51665 -4565 51710 -4445
rect 51830 -4565 51885 -4445
rect 52005 -4565 52050 -4445
rect 52170 -4565 52215 -4445
rect 52335 -4565 52380 -4445
rect 52500 -4565 52555 -4445
rect 52675 -4565 52720 -4445
rect 52840 -4565 52885 -4445
rect 53005 -4565 53050 -4445
rect 53170 -4565 53225 -4445
rect 53345 -4565 53355 -4445
rect 47855 -4610 53355 -4565
rect 47855 -4730 47865 -4610
rect 47985 -4730 48030 -4610
rect 48150 -4730 48195 -4610
rect 48315 -4730 48360 -4610
rect 48480 -4730 48535 -4610
rect 48655 -4730 48700 -4610
rect 48820 -4730 48865 -4610
rect 48985 -4730 49030 -4610
rect 49150 -4730 49205 -4610
rect 49325 -4730 49370 -4610
rect 49490 -4730 49535 -4610
rect 49655 -4730 49700 -4610
rect 49820 -4730 49875 -4610
rect 49995 -4730 50040 -4610
rect 50160 -4730 50205 -4610
rect 50325 -4730 50370 -4610
rect 50490 -4730 50545 -4610
rect 50665 -4730 50710 -4610
rect 50830 -4730 50875 -4610
rect 50995 -4730 51040 -4610
rect 51160 -4730 51215 -4610
rect 51335 -4730 51380 -4610
rect 51500 -4730 51545 -4610
rect 51665 -4730 51710 -4610
rect 51830 -4730 51885 -4610
rect 52005 -4730 52050 -4610
rect 52170 -4730 52215 -4610
rect 52335 -4730 52380 -4610
rect 52500 -4730 52555 -4610
rect 52675 -4730 52720 -4610
rect 52840 -4730 52885 -4610
rect 53005 -4730 53050 -4610
rect 53170 -4730 53225 -4610
rect 53345 -4730 53355 -4610
rect 47855 -4775 53355 -4730
rect 47855 -4895 47865 -4775
rect 47985 -4895 48030 -4775
rect 48150 -4895 48195 -4775
rect 48315 -4895 48360 -4775
rect 48480 -4895 48535 -4775
rect 48655 -4895 48700 -4775
rect 48820 -4895 48865 -4775
rect 48985 -4895 49030 -4775
rect 49150 -4895 49205 -4775
rect 49325 -4895 49370 -4775
rect 49490 -4895 49535 -4775
rect 49655 -4895 49700 -4775
rect 49820 -4895 49875 -4775
rect 49995 -4895 50040 -4775
rect 50160 -4895 50205 -4775
rect 50325 -4895 50370 -4775
rect 50490 -4895 50545 -4775
rect 50665 -4895 50710 -4775
rect 50830 -4895 50875 -4775
rect 50995 -4895 51040 -4775
rect 51160 -4895 51215 -4775
rect 51335 -4895 51380 -4775
rect 51500 -4895 51545 -4775
rect 51665 -4895 51710 -4775
rect 51830 -4895 51885 -4775
rect 52005 -4895 52050 -4775
rect 52170 -4895 52215 -4775
rect 52335 -4895 52380 -4775
rect 52500 -4895 52555 -4775
rect 52675 -4895 52720 -4775
rect 52840 -4895 52885 -4775
rect 53005 -4895 53050 -4775
rect 53170 -4895 53225 -4775
rect 53345 -4895 53355 -4775
rect 47855 -4940 53355 -4895
rect 47855 -5060 47865 -4940
rect 47985 -5060 48030 -4940
rect 48150 -5060 48195 -4940
rect 48315 -5060 48360 -4940
rect 48480 -5060 48535 -4940
rect 48655 -5060 48700 -4940
rect 48820 -5060 48865 -4940
rect 48985 -5060 49030 -4940
rect 49150 -5060 49205 -4940
rect 49325 -5060 49370 -4940
rect 49490 -5060 49535 -4940
rect 49655 -5060 49700 -4940
rect 49820 -5060 49875 -4940
rect 49995 -5060 50040 -4940
rect 50160 -5060 50205 -4940
rect 50325 -5060 50370 -4940
rect 50490 -5060 50545 -4940
rect 50665 -5060 50710 -4940
rect 50830 -5060 50875 -4940
rect 50995 -5060 51040 -4940
rect 51160 -5060 51215 -4940
rect 51335 -5060 51380 -4940
rect 51500 -5060 51545 -4940
rect 51665 -5060 51710 -4940
rect 51830 -5060 51885 -4940
rect 52005 -5060 52050 -4940
rect 52170 -5060 52215 -4940
rect 52335 -5060 52380 -4940
rect 52500 -5060 52555 -4940
rect 52675 -5060 52720 -4940
rect 52840 -5060 52885 -4940
rect 53005 -5060 53050 -4940
rect 53170 -5060 53225 -4940
rect 53345 -5060 53355 -4940
rect 47855 -5115 53355 -5060
rect 47855 -5235 47865 -5115
rect 47985 -5235 48030 -5115
rect 48150 -5235 48195 -5115
rect 48315 -5235 48360 -5115
rect 48480 -5235 48535 -5115
rect 48655 -5235 48700 -5115
rect 48820 -5235 48865 -5115
rect 48985 -5235 49030 -5115
rect 49150 -5235 49205 -5115
rect 49325 -5235 49370 -5115
rect 49490 -5235 49535 -5115
rect 49655 -5235 49700 -5115
rect 49820 -5235 49875 -5115
rect 49995 -5235 50040 -5115
rect 50160 -5235 50205 -5115
rect 50325 -5235 50370 -5115
rect 50490 -5235 50545 -5115
rect 50665 -5235 50710 -5115
rect 50830 -5235 50875 -5115
rect 50995 -5235 51040 -5115
rect 51160 -5235 51215 -5115
rect 51335 -5235 51380 -5115
rect 51500 -5235 51545 -5115
rect 51665 -5235 51710 -5115
rect 51830 -5235 51885 -5115
rect 52005 -5235 52050 -5115
rect 52170 -5235 52215 -5115
rect 52335 -5235 52380 -5115
rect 52500 -5235 52555 -5115
rect 52675 -5235 52720 -5115
rect 52840 -5235 52885 -5115
rect 53005 -5235 53050 -5115
rect 53170 -5235 53225 -5115
rect 53345 -5235 53355 -5115
rect 47855 -5280 53355 -5235
rect 47855 -5400 47865 -5280
rect 47985 -5400 48030 -5280
rect 48150 -5400 48195 -5280
rect 48315 -5400 48360 -5280
rect 48480 -5400 48535 -5280
rect 48655 -5400 48700 -5280
rect 48820 -5400 48865 -5280
rect 48985 -5400 49030 -5280
rect 49150 -5400 49205 -5280
rect 49325 -5400 49370 -5280
rect 49490 -5400 49535 -5280
rect 49655 -5400 49700 -5280
rect 49820 -5400 49875 -5280
rect 49995 -5400 50040 -5280
rect 50160 -5400 50205 -5280
rect 50325 -5400 50370 -5280
rect 50490 -5400 50545 -5280
rect 50665 -5400 50710 -5280
rect 50830 -5400 50875 -5280
rect 50995 -5400 51040 -5280
rect 51160 -5400 51215 -5280
rect 51335 -5400 51380 -5280
rect 51500 -5400 51545 -5280
rect 51665 -5400 51710 -5280
rect 51830 -5400 51885 -5280
rect 52005 -5400 52050 -5280
rect 52170 -5400 52215 -5280
rect 52335 -5400 52380 -5280
rect 52500 -5400 52555 -5280
rect 52675 -5400 52720 -5280
rect 52840 -5400 52885 -5280
rect 53005 -5400 53050 -5280
rect 53170 -5400 53225 -5280
rect 53345 -5400 53355 -5280
rect 47855 -5445 53355 -5400
rect 47855 -5565 47865 -5445
rect 47985 -5565 48030 -5445
rect 48150 -5565 48195 -5445
rect 48315 -5565 48360 -5445
rect 48480 -5565 48535 -5445
rect 48655 -5565 48700 -5445
rect 48820 -5565 48865 -5445
rect 48985 -5565 49030 -5445
rect 49150 -5565 49205 -5445
rect 49325 -5565 49370 -5445
rect 49490 -5565 49535 -5445
rect 49655 -5565 49700 -5445
rect 49820 -5565 49875 -5445
rect 49995 -5565 50040 -5445
rect 50160 -5565 50205 -5445
rect 50325 -5565 50370 -5445
rect 50490 -5565 50545 -5445
rect 50665 -5565 50710 -5445
rect 50830 -5565 50875 -5445
rect 50995 -5565 51040 -5445
rect 51160 -5565 51215 -5445
rect 51335 -5565 51380 -5445
rect 51500 -5565 51545 -5445
rect 51665 -5565 51710 -5445
rect 51830 -5565 51885 -5445
rect 52005 -5565 52050 -5445
rect 52170 -5565 52215 -5445
rect 52335 -5565 52380 -5445
rect 52500 -5565 52555 -5445
rect 52675 -5565 52720 -5445
rect 52840 -5565 52885 -5445
rect 53005 -5565 53050 -5445
rect 53170 -5565 53225 -5445
rect 53345 -5565 53355 -5445
rect 47855 -5610 53355 -5565
rect 47855 -5730 47865 -5610
rect 47985 -5730 48030 -5610
rect 48150 -5730 48195 -5610
rect 48315 -5730 48360 -5610
rect 48480 -5730 48535 -5610
rect 48655 -5730 48700 -5610
rect 48820 -5730 48865 -5610
rect 48985 -5730 49030 -5610
rect 49150 -5730 49205 -5610
rect 49325 -5730 49370 -5610
rect 49490 -5730 49535 -5610
rect 49655 -5730 49700 -5610
rect 49820 -5730 49875 -5610
rect 49995 -5730 50040 -5610
rect 50160 -5730 50205 -5610
rect 50325 -5730 50370 -5610
rect 50490 -5730 50545 -5610
rect 50665 -5730 50710 -5610
rect 50830 -5730 50875 -5610
rect 50995 -5730 51040 -5610
rect 51160 -5730 51215 -5610
rect 51335 -5730 51380 -5610
rect 51500 -5730 51545 -5610
rect 51665 -5730 51710 -5610
rect 51830 -5730 51885 -5610
rect 52005 -5730 52050 -5610
rect 52170 -5730 52215 -5610
rect 52335 -5730 52380 -5610
rect 52500 -5730 52555 -5610
rect 52675 -5730 52720 -5610
rect 52840 -5730 52885 -5610
rect 53005 -5730 53050 -5610
rect 53170 -5730 53225 -5610
rect 53345 -5730 53355 -5610
rect 47855 -5785 53355 -5730
rect 47855 -5905 47865 -5785
rect 47985 -5905 48030 -5785
rect 48150 -5905 48195 -5785
rect 48315 -5905 48360 -5785
rect 48480 -5905 48535 -5785
rect 48655 -5905 48700 -5785
rect 48820 -5905 48865 -5785
rect 48985 -5905 49030 -5785
rect 49150 -5905 49205 -5785
rect 49325 -5905 49370 -5785
rect 49490 -5905 49535 -5785
rect 49655 -5905 49700 -5785
rect 49820 -5905 49875 -5785
rect 49995 -5905 50040 -5785
rect 50160 -5905 50205 -5785
rect 50325 -5905 50370 -5785
rect 50490 -5905 50545 -5785
rect 50665 -5905 50710 -5785
rect 50830 -5905 50875 -5785
rect 50995 -5905 51040 -5785
rect 51160 -5905 51215 -5785
rect 51335 -5905 51380 -5785
rect 51500 -5905 51545 -5785
rect 51665 -5905 51710 -5785
rect 51830 -5905 51885 -5785
rect 52005 -5905 52050 -5785
rect 52170 -5905 52215 -5785
rect 52335 -5905 52380 -5785
rect 52500 -5905 52555 -5785
rect 52675 -5905 52720 -5785
rect 52840 -5905 52885 -5785
rect 53005 -5905 53050 -5785
rect 53170 -5905 53225 -5785
rect 53345 -5905 53355 -5785
rect 47855 -5950 53355 -5905
rect 47855 -6070 47865 -5950
rect 47985 -6070 48030 -5950
rect 48150 -6070 48195 -5950
rect 48315 -6070 48360 -5950
rect 48480 -6070 48535 -5950
rect 48655 -6070 48700 -5950
rect 48820 -6070 48865 -5950
rect 48985 -6070 49030 -5950
rect 49150 -6070 49205 -5950
rect 49325 -6070 49370 -5950
rect 49490 -6070 49535 -5950
rect 49655 -6070 49700 -5950
rect 49820 -6070 49875 -5950
rect 49995 -6070 50040 -5950
rect 50160 -6070 50205 -5950
rect 50325 -6070 50370 -5950
rect 50490 -6070 50545 -5950
rect 50665 -6070 50710 -5950
rect 50830 -6070 50875 -5950
rect 50995 -6070 51040 -5950
rect 51160 -6070 51215 -5950
rect 51335 -6070 51380 -5950
rect 51500 -6070 51545 -5950
rect 51665 -6070 51710 -5950
rect 51830 -6070 51885 -5950
rect 52005 -6070 52050 -5950
rect 52170 -6070 52215 -5950
rect 52335 -6070 52380 -5950
rect 52500 -6070 52555 -5950
rect 52675 -6070 52720 -5950
rect 52840 -6070 52885 -5950
rect 53005 -6070 53050 -5950
rect 53170 -6070 53225 -5950
rect 53345 -6070 53355 -5950
rect 47855 -6115 53355 -6070
rect 47855 -6235 47865 -6115
rect 47985 -6235 48030 -6115
rect 48150 -6235 48195 -6115
rect 48315 -6235 48360 -6115
rect 48480 -6235 48535 -6115
rect 48655 -6235 48700 -6115
rect 48820 -6235 48865 -6115
rect 48985 -6235 49030 -6115
rect 49150 -6235 49205 -6115
rect 49325 -6235 49370 -6115
rect 49490 -6235 49535 -6115
rect 49655 -6235 49700 -6115
rect 49820 -6235 49875 -6115
rect 49995 -6235 50040 -6115
rect 50160 -6235 50205 -6115
rect 50325 -6235 50370 -6115
rect 50490 -6235 50545 -6115
rect 50665 -6235 50710 -6115
rect 50830 -6235 50875 -6115
rect 50995 -6235 51040 -6115
rect 51160 -6235 51215 -6115
rect 51335 -6235 51380 -6115
rect 51500 -6235 51545 -6115
rect 51665 -6235 51710 -6115
rect 51830 -6235 51885 -6115
rect 52005 -6235 52050 -6115
rect 52170 -6235 52215 -6115
rect 52335 -6235 52380 -6115
rect 52500 -6235 52555 -6115
rect 52675 -6235 52720 -6115
rect 52840 -6235 52885 -6115
rect 53005 -6235 53050 -6115
rect 53170 -6235 53225 -6115
rect 53345 -6235 53355 -6115
rect 47855 -6280 53355 -6235
rect 47855 -6400 47865 -6280
rect 47985 -6400 48030 -6280
rect 48150 -6400 48195 -6280
rect 48315 -6400 48360 -6280
rect 48480 -6400 48535 -6280
rect 48655 -6400 48700 -6280
rect 48820 -6400 48865 -6280
rect 48985 -6400 49030 -6280
rect 49150 -6400 49205 -6280
rect 49325 -6400 49370 -6280
rect 49490 -6400 49535 -6280
rect 49655 -6400 49700 -6280
rect 49820 -6400 49875 -6280
rect 49995 -6400 50040 -6280
rect 50160 -6400 50205 -6280
rect 50325 -6400 50370 -6280
rect 50490 -6400 50545 -6280
rect 50665 -6400 50710 -6280
rect 50830 -6400 50875 -6280
rect 50995 -6400 51040 -6280
rect 51160 -6400 51215 -6280
rect 51335 -6400 51380 -6280
rect 51500 -6400 51545 -6280
rect 51665 -6400 51710 -6280
rect 51830 -6400 51885 -6280
rect 52005 -6400 52050 -6280
rect 52170 -6400 52215 -6280
rect 52335 -6400 52380 -6280
rect 52500 -6400 52555 -6280
rect 52675 -6400 52720 -6280
rect 52840 -6400 52885 -6280
rect 53005 -6400 53050 -6280
rect 53170 -6400 53225 -6280
rect 53345 -6400 53355 -6280
rect 47855 -6455 53355 -6400
rect 47855 -6575 47865 -6455
rect 47985 -6575 48030 -6455
rect 48150 -6575 48195 -6455
rect 48315 -6575 48360 -6455
rect 48480 -6575 48535 -6455
rect 48655 -6575 48700 -6455
rect 48820 -6575 48865 -6455
rect 48985 -6575 49030 -6455
rect 49150 -6575 49205 -6455
rect 49325 -6575 49370 -6455
rect 49490 -6575 49535 -6455
rect 49655 -6575 49700 -6455
rect 49820 -6575 49875 -6455
rect 49995 -6575 50040 -6455
rect 50160 -6575 50205 -6455
rect 50325 -6575 50370 -6455
rect 50490 -6575 50545 -6455
rect 50665 -6575 50710 -6455
rect 50830 -6575 50875 -6455
rect 50995 -6575 51040 -6455
rect 51160 -6575 51215 -6455
rect 51335 -6575 51380 -6455
rect 51500 -6575 51545 -6455
rect 51665 -6575 51710 -6455
rect 51830 -6575 51885 -6455
rect 52005 -6575 52050 -6455
rect 52170 -6575 52215 -6455
rect 52335 -6575 52380 -6455
rect 52500 -6575 52555 -6455
rect 52675 -6575 52720 -6455
rect 52840 -6575 52885 -6455
rect 53005 -6575 53050 -6455
rect 53170 -6575 53225 -6455
rect 53345 -6575 53355 -6455
rect 47855 -6620 53355 -6575
rect 47855 -6740 47865 -6620
rect 47985 -6740 48030 -6620
rect 48150 -6740 48195 -6620
rect 48315 -6740 48360 -6620
rect 48480 -6740 48535 -6620
rect 48655 -6740 48700 -6620
rect 48820 -6740 48865 -6620
rect 48985 -6740 49030 -6620
rect 49150 -6740 49205 -6620
rect 49325 -6740 49370 -6620
rect 49490 -6740 49535 -6620
rect 49655 -6740 49700 -6620
rect 49820 -6740 49875 -6620
rect 49995 -6740 50040 -6620
rect 50160 -6740 50205 -6620
rect 50325 -6740 50370 -6620
rect 50490 -6740 50545 -6620
rect 50665 -6740 50710 -6620
rect 50830 -6740 50875 -6620
rect 50995 -6740 51040 -6620
rect 51160 -6740 51215 -6620
rect 51335 -6740 51380 -6620
rect 51500 -6740 51545 -6620
rect 51665 -6740 51710 -6620
rect 51830 -6740 51885 -6620
rect 52005 -6740 52050 -6620
rect 52170 -6740 52215 -6620
rect 52335 -6740 52380 -6620
rect 52500 -6740 52555 -6620
rect 52675 -6740 52720 -6620
rect 52840 -6740 52885 -6620
rect 53005 -6740 53050 -6620
rect 53170 -6740 53225 -6620
rect 53345 -6740 53355 -6620
rect 47855 -6785 53355 -6740
rect 47855 -6905 47865 -6785
rect 47985 -6905 48030 -6785
rect 48150 -6905 48195 -6785
rect 48315 -6905 48360 -6785
rect 48480 -6905 48535 -6785
rect 48655 -6905 48700 -6785
rect 48820 -6905 48865 -6785
rect 48985 -6905 49030 -6785
rect 49150 -6905 49205 -6785
rect 49325 -6905 49370 -6785
rect 49490 -6905 49535 -6785
rect 49655 -6905 49700 -6785
rect 49820 -6905 49875 -6785
rect 49995 -6905 50040 -6785
rect 50160 -6905 50205 -6785
rect 50325 -6905 50370 -6785
rect 50490 -6905 50545 -6785
rect 50665 -6905 50710 -6785
rect 50830 -6905 50875 -6785
rect 50995 -6905 51040 -6785
rect 51160 -6905 51215 -6785
rect 51335 -6905 51380 -6785
rect 51500 -6905 51545 -6785
rect 51665 -6905 51710 -6785
rect 51830 -6905 51885 -6785
rect 52005 -6905 52050 -6785
rect 52170 -6905 52215 -6785
rect 52335 -6905 52380 -6785
rect 52500 -6905 52555 -6785
rect 52675 -6905 52720 -6785
rect 52840 -6905 52885 -6785
rect 53005 -6905 53050 -6785
rect 53170 -6905 53225 -6785
rect 53345 -6905 53355 -6785
rect 47855 -6950 53355 -6905
rect 47855 -7070 47865 -6950
rect 47985 -7070 48030 -6950
rect 48150 -7070 48195 -6950
rect 48315 -7070 48360 -6950
rect 48480 -7070 48535 -6950
rect 48655 -7070 48700 -6950
rect 48820 -7070 48865 -6950
rect 48985 -7070 49030 -6950
rect 49150 -7070 49205 -6950
rect 49325 -7070 49370 -6950
rect 49490 -7070 49535 -6950
rect 49655 -7070 49700 -6950
rect 49820 -7070 49875 -6950
rect 49995 -7070 50040 -6950
rect 50160 -7070 50205 -6950
rect 50325 -7070 50370 -6950
rect 50490 -7070 50545 -6950
rect 50665 -7070 50710 -6950
rect 50830 -7070 50875 -6950
rect 50995 -7070 51040 -6950
rect 51160 -7070 51215 -6950
rect 51335 -7070 51380 -6950
rect 51500 -7070 51545 -6950
rect 51665 -7070 51710 -6950
rect 51830 -7070 51885 -6950
rect 52005 -7070 52050 -6950
rect 52170 -7070 52215 -6950
rect 52335 -7070 52380 -6950
rect 52500 -7070 52555 -6950
rect 52675 -7070 52720 -6950
rect 52840 -7070 52885 -6950
rect 53005 -7070 53050 -6950
rect 53170 -7070 53225 -6950
rect 53345 -7070 53355 -6950
rect 47855 -7125 53355 -7070
rect 47855 -7245 47865 -7125
rect 47985 -7245 48030 -7125
rect 48150 -7245 48195 -7125
rect 48315 -7245 48360 -7125
rect 48480 -7245 48535 -7125
rect 48655 -7245 48700 -7125
rect 48820 -7245 48865 -7125
rect 48985 -7245 49030 -7125
rect 49150 -7245 49205 -7125
rect 49325 -7245 49370 -7125
rect 49490 -7245 49535 -7125
rect 49655 -7245 49700 -7125
rect 49820 -7245 49875 -7125
rect 49995 -7245 50040 -7125
rect 50160 -7245 50205 -7125
rect 50325 -7245 50370 -7125
rect 50490 -7245 50545 -7125
rect 50665 -7245 50710 -7125
rect 50830 -7245 50875 -7125
rect 50995 -7245 51040 -7125
rect 51160 -7245 51215 -7125
rect 51335 -7245 51380 -7125
rect 51500 -7245 51545 -7125
rect 51665 -7245 51710 -7125
rect 51830 -7245 51885 -7125
rect 52005 -7245 52050 -7125
rect 52170 -7245 52215 -7125
rect 52335 -7245 52380 -7125
rect 52500 -7245 52555 -7125
rect 52675 -7245 52720 -7125
rect 52840 -7245 52885 -7125
rect 53005 -7245 53050 -7125
rect 53170 -7245 53225 -7125
rect 53345 -7245 53355 -7125
rect 47855 -7290 53355 -7245
rect 47855 -7410 47865 -7290
rect 47985 -7410 48030 -7290
rect 48150 -7410 48195 -7290
rect 48315 -7410 48360 -7290
rect 48480 -7410 48535 -7290
rect 48655 -7410 48700 -7290
rect 48820 -7410 48865 -7290
rect 48985 -7410 49030 -7290
rect 49150 -7410 49205 -7290
rect 49325 -7410 49370 -7290
rect 49490 -7410 49535 -7290
rect 49655 -7410 49700 -7290
rect 49820 -7410 49875 -7290
rect 49995 -7410 50040 -7290
rect 50160 -7410 50205 -7290
rect 50325 -7410 50370 -7290
rect 50490 -7410 50545 -7290
rect 50665 -7410 50710 -7290
rect 50830 -7410 50875 -7290
rect 50995 -7410 51040 -7290
rect 51160 -7410 51215 -7290
rect 51335 -7410 51380 -7290
rect 51500 -7410 51545 -7290
rect 51665 -7410 51710 -7290
rect 51830 -7410 51885 -7290
rect 52005 -7410 52050 -7290
rect 52170 -7410 52215 -7290
rect 52335 -7410 52380 -7290
rect 52500 -7410 52555 -7290
rect 52675 -7410 52720 -7290
rect 52840 -7410 52885 -7290
rect 53005 -7410 53050 -7290
rect 53170 -7410 53225 -7290
rect 53345 -7410 53355 -7290
rect 47855 -7455 53355 -7410
rect 47855 -7575 47865 -7455
rect 47985 -7575 48030 -7455
rect 48150 -7575 48195 -7455
rect 48315 -7575 48360 -7455
rect 48480 -7575 48535 -7455
rect 48655 -7575 48700 -7455
rect 48820 -7575 48865 -7455
rect 48985 -7575 49030 -7455
rect 49150 -7575 49205 -7455
rect 49325 -7575 49370 -7455
rect 49490 -7575 49535 -7455
rect 49655 -7575 49700 -7455
rect 49820 -7575 49875 -7455
rect 49995 -7575 50040 -7455
rect 50160 -7575 50205 -7455
rect 50325 -7575 50370 -7455
rect 50490 -7575 50545 -7455
rect 50665 -7575 50710 -7455
rect 50830 -7575 50875 -7455
rect 50995 -7575 51040 -7455
rect 51160 -7575 51215 -7455
rect 51335 -7575 51380 -7455
rect 51500 -7575 51545 -7455
rect 51665 -7575 51710 -7455
rect 51830 -7575 51885 -7455
rect 52005 -7575 52050 -7455
rect 52170 -7575 52215 -7455
rect 52335 -7575 52380 -7455
rect 52500 -7575 52555 -7455
rect 52675 -7575 52720 -7455
rect 52840 -7575 52885 -7455
rect 53005 -7575 53050 -7455
rect 53170 -7575 53225 -7455
rect 53345 -7575 53355 -7455
rect 47855 -7620 53355 -7575
rect 47855 -7740 47865 -7620
rect 47985 -7740 48030 -7620
rect 48150 -7740 48195 -7620
rect 48315 -7740 48360 -7620
rect 48480 -7740 48535 -7620
rect 48655 -7740 48700 -7620
rect 48820 -7740 48865 -7620
rect 48985 -7740 49030 -7620
rect 49150 -7740 49205 -7620
rect 49325 -7740 49370 -7620
rect 49490 -7740 49535 -7620
rect 49655 -7740 49700 -7620
rect 49820 -7740 49875 -7620
rect 49995 -7740 50040 -7620
rect 50160 -7740 50205 -7620
rect 50325 -7740 50370 -7620
rect 50490 -7740 50545 -7620
rect 50665 -7740 50710 -7620
rect 50830 -7740 50875 -7620
rect 50995 -7740 51040 -7620
rect 51160 -7740 51215 -7620
rect 51335 -7740 51380 -7620
rect 51500 -7740 51545 -7620
rect 51665 -7740 51710 -7620
rect 51830 -7740 51885 -7620
rect 52005 -7740 52050 -7620
rect 52170 -7740 52215 -7620
rect 52335 -7740 52380 -7620
rect 52500 -7740 52555 -7620
rect 52675 -7740 52720 -7620
rect 52840 -7740 52885 -7620
rect 53005 -7740 53050 -7620
rect 53170 -7740 53225 -7620
rect 53345 -7740 53355 -7620
rect 47855 -7795 53355 -7740
rect 47855 -7915 47865 -7795
rect 47985 -7915 48030 -7795
rect 48150 -7915 48195 -7795
rect 48315 -7915 48360 -7795
rect 48480 -7915 48535 -7795
rect 48655 -7915 48700 -7795
rect 48820 -7915 48865 -7795
rect 48985 -7915 49030 -7795
rect 49150 -7915 49205 -7795
rect 49325 -7915 49370 -7795
rect 49490 -7915 49535 -7795
rect 49655 -7915 49700 -7795
rect 49820 -7915 49875 -7795
rect 49995 -7915 50040 -7795
rect 50160 -7915 50205 -7795
rect 50325 -7915 50370 -7795
rect 50490 -7915 50545 -7795
rect 50665 -7915 50710 -7795
rect 50830 -7915 50875 -7795
rect 50995 -7915 51040 -7795
rect 51160 -7915 51215 -7795
rect 51335 -7915 51380 -7795
rect 51500 -7915 51545 -7795
rect 51665 -7915 51710 -7795
rect 51830 -7915 51885 -7795
rect 52005 -7915 52050 -7795
rect 52170 -7915 52215 -7795
rect 52335 -7915 52380 -7795
rect 52500 -7915 52555 -7795
rect 52675 -7915 52720 -7795
rect 52840 -7915 52885 -7795
rect 53005 -7915 53050 -7795
rect 53170 -7915 53225 -7795
rect 53345 -7915 53355 -7795
rect 47855 -7960 53355 -7915
rect 47855 -8080 47865 -7960
rect 47985 -8080 48030 -7960
rect 48150 -8080 48195 -7960
rect 48315 -8080 48360 -7960
rect 48480 -8080 48535 -7960
rect 48655 -8080 48700 -7960
rect 48820 -8080 48865 -7960
rect 48985 -8080 49030 -7960
rect 49150 -8080 49205 -7960
rect 49325 -8080 49370 -7960
rect 49490 -8080 49535 -7960
rect 49655 -8080 49700 -7960
rect 49820 -8080 49875 -7960
rect 49995 -8080 50040 -7960
rect 50160 -8080 50205 -7960
rect 50325 -8080 50370 -7960
rect 50490 -8080 50545 -7960
rect 50665 -8080 50710 -7960
rect 50830 -8080 50875 -7960
rect 50995 -8080 51040 -7960
rect 51160 -8080 51215 -7960
rect 51335 -8080 51380 -7960
rect 51500 -8080 51545 -7960
rect 51665 -8080 51710 -7960
rect 51830 -8080 51885 -7960
rect 52005 -8080 52050 -7960
rect 52170 -8080 52215 -7960
rect 52335 -8080 52380 -7960
rect 52500 -8080 52555 -7960
rect 52675 -8080 52720 -7960
rect 52840 -8080 52885 -7960
rect 53005 -8080 53050 -7960
rect 53170 -8080 53225 -7960
rect 53345 -8080 53355 -7960
rect 47855 -8125 53355 -8080
rect 47855 -8245 47865 -8125
rect 47985 -8245 48030 -8125
rect 48150 -8245 48195 -8125
rect 48315 -8245 48360 -8125
rect 48480 -8245 48535 -8125
rect 48655 -8245 48700 -8125
rect 48820 -8245 48865 -8125
rect 48985 -8245 49030 -8125
rect 49150 -8245 49205 -8125
rect 49325 -8245 49370 -8125
rect 49490 -8245 49535 -8125
rect 49655 -8245 49700 -8125
rect 49820 -8245 49875 -8125
rect 49995 -8245 50040 -8125
rect 50160 -8245 50205 -8125
rect 50325 -8245 50370 -8125
rect 50490 -8245 50545 -8125
rect 50665 -8245 50710 -8125
rect 50830 -8245 50875 -8125
rect 50995 -8245 51040 -8125
rect 51160 -8245 51215 -8125
rect 51335 -8245 51380 -8125
rect 51500 -8245 51545 -8125
rect 51665 -8245 51710 -8125
rect 51830 -8245 51885 -8125
rect 52005 -8245 52050 -8125
rect 52170 -8245 52215 -8125
rect 52335 -8245 52380 -8125
rect 52500 -8245 52555 -8125
rect 52675 -8245 52720 -8125
rect 52840 -8245 52885 -8125
rect 53005 -8245 53050 -8125
rect 53170 -8245 53225 -8125
rect 53345 -8245 53355 -8125
rect 47855 -8290 53355 -8245
rect 47855 -8410 47865 -8290
rect 47985 -8410 48030 -8290
rect 48150 -8410 48195 -8290
rect 48315 -8410 48360 -8290
rect 48480 -8410 48535 -8290
rect 48655 -8410 48700 -8290
rect 48820 -8410 48865 -8290
rect 48985 -8410 49030 -8290
rect 49150 -8410 49205 -8290
rect 49325 -8410 49370 -8290
rect 49490 -8410 49535 -8290
rect 49655 -8410 49700 -8290
rect 49820 -8410 49875 -8290
rect 49995 -8410 50040 -8290
rect 50160 -8410 50205 -8290
rect 50325 -8410 50370 -8290
rect 50490 -8410 50545 -8290
rect 50665 -8410 50710 -8290
rect 50830 -8410 50875 -8290
rect 50995 -8410 51040 -8290
rect 51160 -8410 51215 -8290
rect 51335 -8410 51380 -8290
rect 51500 -8410 51545 -8290
rect 51665 -8410 51710 -8290
rect 51830 -8410 51885 -8290
rect 52005 -8410 52050 -8290
rect 52170 -8410 52215 -8290
rect 52335 -8410 52380 -8290
rect 52500 -8410 52555 -8290
rect 52675 -8410 52720 -8290
rect 52840 -8410 52885 -8290
rect 53005 -8410 53050 -8290
rect 53170 -8410 53225 -8290
rect 53345 -8410 53355 -8290
rect 47855 -8465 53355 -8410
rect 47855 -8585 47865 -8465
rect 47985 -8585 48030 -8465
rect 48150 -8585 48195 -8465
rect 48315 -8585 48360 -8465
rect 48480 -8585 48535 -8465
rect 48655 -8585 48700 -8465
rect 48820 -8585 48865 -8465
rect 48985 -8585 49030 -8465
rect 49150 -8585 49205 -8465
rect 49325 -8585 49370 -8465
rect 49490 -8585 49535 -8465
rect 49655 -8585 49700 -8465
rect 49820 -8585 49875 -8465
rect 49995 -8585 50040 -8465
rect 50160 -8585 50205 -8465
rect 50325 -8585 50370 -8465
rect 50490 -8585 50545 -8465
rect 50665 -8585 50710 -8465
rect 50830 -8585 50875 -8465
rect 50995 -8585 51040 -8465
rect 51160 -8585 51215 -8465
rect 51335 -8585 51380 -8465
rect 51500 -8585 51545 -8465
rect 51665 -8585 51710 -8465
rect 51830 -8585 51885 -8465
rect 52005 -8585 52050 -8465
rect 52170 -8585 52215 -8465
rect 52335 -8585 52380 -8465
rect 52500 -8585 52555 -8465
rect 52675 -8585 52720 -8465
rect 52840 -8585 52885 -8465
rect 53005 -8585 53050 -8465
rect 53170 -8585 53225 -8465
rect 53345 -8585 53355 -8465
rect 47855 -8630 53355 -8585
rect 47855 -8750 47865 -8630
rect 47985 -8750 48030 -8630
rect 48150 -8750 48195 -8630
rect 48315 -8750 48360 -8630
rect 48480 -8750 48535 -8630
rect 48655 -8750 48700 -8630
rect 48820 -8750 48865 -8630
rect 48985 -8750 49030 -8630
rect 49150 -8750 49205 -8630
rect 49325 -8750 49370 -8630
rect 49490 -8750 49535 -8630
rect 49655 -8750 49700 -8630
rect 49820 -8750 49875 -8630
rect 49995 -8750 50040 -8630
rect 50160 -8750 50205 -8630
rect 50325 -8750 50370 -8630
rect 50490 -8750 50545 -8630
rect 50665 -8750 50710 -8630
rect 50830 -8750 50875 -8630
rect 50995 -8750 51040 -8630
rect 51160 -8750 51215 -8630
rect 51335 -8750 51380 -8630
rect 51500 -8750 51545 -8630
rect 51665 -8750 51710 -8630
rect 51830 -8750 51885 -8630
rect 52005 -8750 52050 -8630
rect 52170 -8750 52215 -8630
rect 52335 -8750 52380 -8630
rect 52500 -8750 52555 -8630
rect 52675 -8750 52720 -8630
rect 52840 -8750 52885 -8630
rect 53005 -8750 53050 -8630
rect 53170 -8750 53225 -8630
rect 53345 -8750 53355 -8630
rect 47855 -8795 53355 -8750
rect 47855 -8915 47865 -8795
rect 47985 -8915 48030 -8795
rect 48150 -8915 48195 -8795
rect 48315 -8915 48360 -8795
rect 48480 -8915 48535 -8795
rect 48655 -8915 48700 -8795
rect 48820 -8915 48865 -8795
rect 48985 -8915 49030 -8795
rect 49150 -8915 49205 -8795
rect 49325 -8915 49370 -8795
rect 49490 -8915 49535 -8795
rect 49655 -8915 49700 -8795
rect 49820 -8915 49875 -8795
rect 49995 -8915 50040 -8795
rect 50160 -8915 50205 -8795
rect 50325 -8915 50370 -8795
rect 50490 -8915 50545 -8795
rect 50665 -8915 50710 -8795
rect 50830 -8915 50875 -8795
rect 50995 -8915 51040 -8795
rect 51160 -8915 51215 -8795
rect 51335 -8915 51380 -8795
rect 51500 -8915 51545 -8795
rect 51665 -8915 51710 -8795
rect 51830 -8915 51885 -8795
rect 52005 -8915 52050 -8795
rect 52170 -8915 52215 -8795
rect 52335 -8915 52380 -8795
rect 52500 -8915 52555 -8795
rect 52675 -8915 52720 -8795
rect 52840 -8915 52885 -8795
rect 53005 -8915 53050 -8795
rect 53170 -8915 53225 -8795
rect 53345 -8915 53355 -8795
rect 47855 -8960 53355 -8915
rect 47855 -9080 47865 -8960
rect 47985 -9080 48030 -8960
rect 48150 -9080 48195 -8960
rect 48315 -9080 48360 -8960
rect 48480 -9080 48535 -8960
rect 48655 -9080 48700 -8960
rect 48820 -9080 48865 -8960
rect 48985 -9080 49030 -8960
rect 49150 -9080 49205 -8960
rect 49325 -9080 49370 -8960
rect 49490 -9080 49535 -8960
rect 49655 -9080 49700 -8960
rect 49820 -9080 49875 -8960
rect 49995 -9080 50040 -8960
rect 50160 -9080 50205 -8960
rect 50325 -9080 50370 -8960
rect 50490 -9080 50545 -8960
rect 50665 -9080 50710 -8960
rect 50830 -9080 50875 -8960
rect 50995 -9080 51040 -8960
rect 51160 -9080 51215 -8960
rect 51335 -9080 51380 -8960
rect 51500 -9080 51545 -8960
rect 51665 -9080 51710 -8960
rect 51830 -9080 51885 -8960
rect 52005 -9080 52050 -8960
rect 52170 -9080 52215 -8960
rect 52335 -9080 52380 -8960
rect 52500 -9080 52555 -8960
rect 52675 -9080 52720 -8960
rect 52840 -9080 52885 -8960
rect 53005 -9080 53050 -8960
rect 53170 -9080 53225 -8960
rect 53345 -9080 53355 -8960
rect 47855 -9135 53355 -9080
rect 47855 -9255 47865 -9135
rect 47985 -9255 48030 -9135
rect 48150 -9255 48195 -9135
rect 48315 -9255 48360 -9135
rect 48480 -9255 48535 -9135
rect 48655 -9255 48700 -9135
rect 48820 -9255 48865 -9135
rect 48985 -9255 49030 -9135
rect 49150 -9255 49205 -9135
rect 49325 -9255 49370 -9135
rect 49490 -9255 49535 -9135
rect 49655 -9255 49700 -9135
rect 49820 -9255 49875 -9135
rect 49995 -9255 50040 -9135
rect 50160 -9255 50205 -9135
rect 50325 -9255 50370 -9135
rect 50490 -9255 50545 -9135
rect 50665 -9255 50710 -9135
rect 50830 -9255 50875 -9135
rect 50995 -9255 51040 -9135
rect 51160 -9255 51215 -9135
rect 51335 -9255 51380 -9135
rect 51500 -9255 51545 -9135
rect 51665 -9255 51710 -9135
rect 51830 -9255 51885 -9135
rect 52005 -9255 52050 -9135
rect 52170 -9255 52215 -9135
rect 52335 -9255 52380 -9135
rect 52500 -9255 52555 -9135
rect 52675 -9255 52720 -9135
rect 52840 -9255 52885 -9135
rect 53005 -9255 53050 -9135
rect 53170 -9255 53225 -9135
rect 53345 -9255 53355 -9135
rect 47855 -9300 53355 -9255
rect 47855 -9420 47865 -9300
rect 47985 -9420 48030 -9300
rect 48150 -9420 48195 -9300
rect 48315 -9420 48360 -9300
rect 48480 -9420 48535 -9300
rect 48655 -9420 48700 -9300
rect 48820 -9420 48865 -9300
rect 48985 -9420 49030 -9300
rect 49150 -9420 49205 -9300
rect 49325 -9420 49370 -9300
rect 49490 -9420 49535 -9300
rect 49655 -9420 49700 -9300
rect 49820 -9420 49875 -9300
rect 49995 -9420 50040 -9300
rect 50160 -9420 50205 -9300
rect 50325 -9420 50370 -9300
rect 50490 -9420 50545 -9300
rect 50665 -9420 50710 -9300
rect 50830 -9420 50875 -9300
rect 50995 -9420 51040 -9300
rect 51160 -9420 51215 -9300
rect 51335 -9420 51380 -9300
rect 51500 -9420 51545 -9300
rect 51665 -9420 51710 -9300
rect 51830 -9420 51885 -9300
rect 52005 -9420 52050 -9300
rect 52170 -9420 52215 -9300
rect 52335 -9420 52380 -9300
rect 52500 -9420 52555 -9300
rect 52675 -9420 52720 -9300
rect 52840 -9420 52885 -9300
rect 53005 -9420 53050 -9300
rect 53170 -9420 53225 -9300
rect 53345 -9420 53355 -9300
rect 47855 -9465 53355 -9420
rect 47855 -9585 47865 -9465
rect 47985 -9585 48030 -9465
rect 48150 -9585 48195 -9465
rect 48315 -9585 48360 -9465
rect 48480 -9585 48535 -9465
rect 48655 -9585 48700 -9465
rect 48820 -9585 48865 -9465
rect 48985 -9585 49030 -9465
rect 49150 -9585 49205 -9465
rect 49325 -9585 49370 -9465
rect 49490 -9585 49535 -9465
rect 49655 -9585 49700 -9465
rect 49820 -9585 49875 -9465
rect 49995 -9585 50040 -9465
rect 50160 -9585 50205 -9465
rect 50325 -9585 50370 -9465
rect 50490 -9585 50545 -9465
rect 50665 -9585 50710 -9465
rect 50830 -9585 50875 -9465
rect 50995 -9585 51040 -9465
rect 51160 -9585 51215 -9465
rect 51335 -9585 51380 -9465
rect 51500 -9585 51545 -9465
rect 51665 -9585 51710 -9465
rect 51830 -9585 51885 -9465
rect 52005 -9585 52050 -9465
rect 52170 -9585 52215 -9465
rect 52335 -9585 52380 -9465
rect 52500 -9585 52555 -9465
rect 52675 -9585 52720 -9465
rect 52840 -9585 52885 -9465
rect 53005 -9585 53050 -9465
rect 53170 -9585 53225 -9465
rect 53345 -9585 53355 -9465
rect 47855 -9630 53355 -9585
rect 47855 -9750 47865 -9630
rect 47985 -9750 48030 -9630
rect 48150 -9750 48195 -9630
rect 48315 -9750 48360 -9630
rect 48480 -9750 48535 -9630
rect 48655 -9750 48700 -9630
rect 48820 -9750 48865 -9630
rect 48985 -9750 49030 -9630
rect 49150 -9750 49205 -9630
rect 49325 -9750 49370 -9630
rect 49490 -9750 49535 -9630
rect 49655 -9750 49700 -9630
rect 49820 -9750 49875 -9630
rect 49995 -9750 50040 -9630
rect 50160 -9750 50205 -9630
rect 50325 -9750 50370 -9630
rect 50490 -9750 50545 -9630
rect 50665 -9750 50710 -9630
rect 50830 -9750 50875 -9630
rect 50995 -9750 51040 -9630
rect 51160 -9750 51215 -9630
rect 51335 -9750 51380 -9630
rect 51500 -9750 51545 -9630
rect 51665 -9750 51710 -9630
rect 51830 -9750 51885 -9630
rect 52005 -9750 52050 -9630
rect 52170 -9750 52215 -9630
rect 52335 -9750 52380 -9630
rect 52500 -9750 52555 -9630
rect 52675 -9750 52720 -9630
rect 52840 -9750 52885 -9630
rect 53005 -9750 53050 -9630
rect 53170 -9750 53225 -9630
rect 53345 -9750 53355 -9630
rect 47855 -9760 53355 -9750
rect 30785 -10050 36285 -10040
rect 30785 -10170 30795 -10050
rect 30915 -10170 30970 -10050
rect 31090 -10170 31135 -10050
rect 31255 -10170 31300 -10050
rect 31420 -10170 31465 -10050
rect 31585 -10170 31640 -10050
rect 31760 -10170 31805 -10050
rect 31925 -10170 31970 -10050
rect 32090 -10170 32135 -10050
rect 32255 -10170 32310 -10050
rect 32430 -10170 32475 -10050
rect 32595 -10170 32640 -10050
rect 32760 -10170 32805 -10050
rect 32925 -10170 32980 -10050
rect 33100 -10170 33145 -10050
rect 33265 -10170 33310 -10050
rect 33430 -10170 33475 -10050
rect 33595 -10170 33650 -10050
rect 33770 -10170 33815 -10050
rect 33935 -10170 33980 -10050
rect 34100 -10170 34145 -10050
rect 34265 -10170 34320 -10050
rect 34440 -10170 34485 -10050
rect 34605 -10170 34650 -10050
rect 34770 -10170 34815 -10050
rect 34935 -10170 34990 -10050
rect 35110 -10170 35155 -10050
rect 35275 -10170 35320 -10050
rect 35440 -10170 35485 -10050
rect 35605 -10170 35660 -10050
rect 35780 -10170 35825 -10050
rect 35945 -10170 35990 -10050
rect 36110 -10170 36155 -10050
rect 36275 -10170 36285 -10050
rect 30785 -10215 36285 -10170
rect 30785 -10335 30795 -10215
rect 30915 -10335 30970 -10215
rect 31090 -10335 31135 -10215
rect 31255 -10335 31300 -10215
rect 31420 -10335 31465 -10215
rect 31585 -10335 31640 -10215
rect 31760 -10335 31805 -10215
rect 31925 -10335 31970 -10215
rect 32090 -10335 32135 -10215
rect 32255 -10335 32310 -10215
rect 32430 -10335 32475 -10215
rect 32595 -10335 32640 -10215
rect 32760 -10335 32805 -10215
rect 32925 -10335 32980 -10215
rect 33100 -10335 33145 -10215
rect 33265 -10335 33310 -10215
rect 33430 -10335 33475 -10215
rect 33595 -10335 33650 -10215
rect 33770 -10335 33815 -10215
rect 33935 -10335 33980 -10215
rect 34100 -10335 34145 -10215
rect 34265 -10335 34320 -10215
rect 34440 -10335 34485 -10215
rect 34605 -10335 34650 -10215
rect 34770 -10335 34815 -10215
rect 34935 -10335 34990 -10215
rect 35110 -10335 35155 -10215
rect 35275 -10335 35320 -10215
rect 35440 -10335 35485 -10215
rect 35605 -10335 35660 -10215
rect 35780 -10335 35825 -10215
rect 35945 -10335 35990 -10215
rect 36110 -10335 36155 -10215
rect 36275 -10335 36285 -10215
rect 30785 -10380 36285 -10335
rect 30785 -10500 30795 -10380
rect 30915 -10500 30970 -10380
rect 31090 -10500 31135 -10380
rect 31255 -10500 31300 -10380
rect 31420 -10500 31465 -10380
rect 31585 -10500 31640 -10380
rect 31760 -10500 31805 -10380
rect 31925 -10500 31970 -10380
rect 32090 -10500 32135 -10380
rect 32255 -10500 32310 -10380
rect 32430 -10500 32475 -10380
rect 32595 -10500 32640 -10380
rect 32760 -10500 32805 -10380
rect 32925 -10500 32980 -10380
rect 33100 -10500 33145 -10380
rect 33265 -10500 33310 -10380
rect 33430 -10500 33475 -10380
rect 33595 -10500 33650 -10380
rect 33770 -10500 33815 -10380
rect 33935 -10500 33980 -10380
rect 34100 -10500 34145 -10380
rect 34265 -10500 34320 -10380
rect 34440 -10500 34485 -10380
rect 34605 -10500 34650 -10380
rect 34770 -10500 34815 -10380
rect 34935 -10500 34990 -10380
rect 35110 -10500 35155 -10380
rect 35275 -10500 35320 -10380
rect 35440 -10500 35485 -10380
rect 35605 -10500 35660 -10380
rect 35780 -10500 35825 -10380
rect 35945 -10500 35990 -10380
rect 36110 -10500 36155 -10380
rect 36275 -10500 36285 -10380
rect 30785 -10545 36285 -10500
rect 30785 -10665 30795 -10545
rect 30915 -10665 30970 -10545
rect 31090 -10665 31135 -10545
rect 31255 -10665 31300 -10545
rect 31420 -10665 31465 -10545
rect 31585 -10665 31640 -10545
rect 31760 -10665 31805 -10545
rect 31925 -10665 31970 -10545
rect 32090 -10665 32135 -10545
rect 32255 -10665 32310 -10545
rect 32430 -10665 32475 -10545
rect 32595 -10665 32640 -10545
rect 32760 -10665 32805 -10545
rect 32925 -10665 32980 -10545
rect 33100 -10665 33145 -10545
rect 33265 -10665 33310 -10545
rect 33430 -10665 33475 -10545
rect 33595 -10665 33650 -10545
rect 33770 -10665 33815 -10545
rect 33935 -10665 33980 -10545
rect 34100 -10665 34145 -10545
rect 34265 -10665 34320 -10545
rect 34440 -10665 34485 -10545
rect 34605 -10665 34650 -10545
rect 34770 -10665 34815 -10545
rect 34935 -10665 34990 -10545
rect 35110 -10665 35155 -10545
rect 35275 -10665 35320 -10545
rect 35440 -10665 35485 -10545
rect 35605 -10665 35660 -10545
rect 35780 -10665 35825 -10545
rect 35945 -10665 35990 -10545
rect 36110 -10665 36155 -10545
rect 36275 -10665 36285 -10545
rect 30785 -10720 36285 -10665
rect 30785 -10840 30795 -10720
rect 30915 -10840 30970 -10720
rect 31090 -10840 31135 -10720
rect 31255 -10840 31300 -10720
rect 31420 -10840 31465 -10720
rect 31585 -10840 31640 -10720
rect 31760 -10840 31805 -10720
rect 31925 -10840 31970 -10720
rect 32090 -10840 32135 -10720
rect 32255 -10840 32310 -10720
rect 32430 -10840 32475 -10720
rect 32595 -10840 32640 -10720
rect 32760 -10840 32805 -10720
rect 32925 -10840 32980 -10720
rect 33100 -10840 33145 -10720
rect 33265 -10840 33310 -10720
rect 33430 -10840 33475 -10720
rect 33595 -10840 33650 -10720
rect 33770 -10840 33815 -10720
rect 33935 -10840 33980 -10720
rect 34100 -10840 34145 -10720
rect 34265 -10840 34320 -10720
rect 34440 -10840 34485 -10720
rect 34605 -10840 34650 -10720
rect 34770 -10840 34815 -10720
rect 34935 -10840 34990 -10720
rect 35110 -10840 35155 -10720
rect 35275 -10840 35320 -10720
rect 35440 -10840 35485 -10720
rect 35605 -10840 35660 -10720
rect 35780 -10840 35825 -10720
rect 35945 -10840 35990 -10720
rect 36110 -10840 36155 -10720
rect 36275 -10840 36285 -10720
rect 30785 -10885 36285 -10840
rect 30785 -11005 30795 -10885
rect 30915 -11005 30970 -10885
rect 31090 -11005 31135 -10885
rect 31255 -11005 31300 -10885
rect 31420 -11005 31465 -10885
rect 31585 -11005 31640 -10885
rect 31760 -11005 31805 -10885
rect 31925 -11005 31970 -10885
rect 32090 -11005 32135 -10885
rect 32255 -11005 32310 -10885
rect 32430 -11005 32475 -10885
rect 32595 -11005 32640 -10885
rect 32760 -11005 32805 -10885
rect 32925 -11005 32980 -10885
rect 33100 -11005 33145 -10885
rect 33265 -11005 33310 -10885
rect 33430 -11005 33475 -10885
rect 33595 -11005 33650 -10885
rect 33770 -11005 33815 -10885
rect 33935 -11005 33980 -10885
rect 34100 -11005 34145 -10885
rect 34265 -11005 34320 -10885
rect 34440 -11005 34485 -10885
rect 34605 -11005 34650 -10885
rect 34770 -11005 34815 -10885
rect 34935 -11005 34990 -10885
rect 35110 -11005 35155 -10885
rect 35275 -11005 35320 -10885
rect 35440 -11005 35485 -10885
rect 35605 -11005 35660 -10885
rect 35780 -11005 35825 -10885
rect 35945 -11005 35990 -10885
rect 36110 -11005 36155 -10885
rect 36275 -11005 36285 -10885
rect 30785 -11050 36285 -11005
rect 30785 -11170 30795 -11050
rect 30915 -11170 30970 -11050
rect 31090 -11170 31135 -11050
rect 31255 -11170 31300 -11050
rect 31420 -11170 31465 -11050
rect 31585 -11170 31640 -11050
rect 31760 -11170 31805 -11050
rect 31925 -11170 31970 -11050
rect 32090 -11170 32135 -11050
rect 32255 -11170 32310 -11050
rect 32430 -11170 32475 -11050
rect 32595 -11170 32640 -11050
rect 32760 -11170 32805 -11050
rect 32925 -11170 32980 -11050
rect 33100 -11170 33145 -11050
rect 33265 -11170 33310 -11050
rect 33430 -11170 33475 -11050
rect 33595 -11170 33650 -11050
rect 33770 -11170 33815 -11050
rect 33935 -11170 33980 -11050
rect 34100 -11170 34145 -11050
rect 34265 -11170 34320 -11050
rect 34440 -11170 34485 -11050
rect 34605 -11170 34650 -11050
rect 34770 -11170 34815 -11050
rect 34935 -11170 34990 -11050
rect 35110 -11170 35155 -11050
rect 35275 -11170 35320 -11050
rect 35440 -11170 35485 -11050
rect 35605 -11170 35660 -11050
rect 35780 -11170 35825 -11050
rect 35945 -11170 35990 -11050
rect 36110 -11170 36155 -11050
rect 36275 -11170 36285 -11050
rect 30785 -11215 36285 -11170
rect 30785 -11335 30795 -11215
rect 30915 -11335 30970 -11215
rect 31090 -11335 31135 -11215
rect 31255 -11335 31300 -11215
rect 31420 -11335 31465 -11215
rect 31585 -11335 31640 -11215
rect 31760 -11335 31805 -11215
rect 31925 -11335 31970 -11215
rect 32090 -11335 32135 -11215
rect 32255 -11335 32310 -11215
rect 32430 -11335 32475 -11215
rect 32595 -11335 32640 -11215
rect 32760 -11335 32805 -11215
rect 32925 -11335 32980 -11215
rect 33100 -11335 33145 -11215
rect 33265 -11335 33310 -11215
rect 33430 -11335 33475 -11215
rect 33595 -11335 33650 -11215
rect 33770 -11335 33815 -11215
rect 33935 -11335 33980 -11215
rect 34100 -11335 34145 -11215
rect 34265 -11335 34320 -11215
rect 34440 -11335 34485 -11215
rect 34605 -11335 34650 -11215
rect 34770 -11335 34815 -11215
rect 34935 -11335 34990 -11215
rect 35110 -11335 35155 -11215
rect 35275 -11335 35320 -11215
rect 35440 -11335 35485 -11215
rect 35605 -11335 35660 -11215
rect 35780 -11335 35825 -11215
rect 35945 -11335 35990 -11215
rect 36110 -11335 36155 -11215
rect 36275 -11335 36285 -11215
rect 30785 -11390 36285 -11335
rect 30785 -11510 30795 -11390
rect 30915 -11510 30970 -11390
rect 31090 -11510 31135 -11390
rect 31255 -11510 31300 -11390
rect 31420 -11510 31465 -11390
rect 31585 -11510 31640 -11390
rect 31760 -11510 31805 -11390
rect 31925 -11510 31970 -11390
rect 32090 -11510 32135 -11390
rect 32255 -11510 32310 -11390
rect 32430 -11510 32475 -11390
rect 32595 -11510 32640 -11390
rect 32760 -11510 32805 -11390
rect 32925 -11510 32980 -11390
rect 33100 -11510 33145 -11390
rect 33265 -11510 33310 -11390
rect 33430 -11510 33475 -11390
rect 33595 -11510 33650 -11390
rect 33770 -11510 33815 -11390
rect 33935 -11510 33980 -11390
rect 34100 -11510 34145 -11390
rect 34265 -11510 34320 -11390
rect 34440 -11510 34485 -11390
rect 34605 -11510 34650 -11390
rect 34770 -11510 34815 -11390
rect 34935 -11510 34990 -11390
rect 35110 -11510 35155 -11390
rect 35275 -11510 35320 -11390
rect 35440 -11510 35485 -11390
rect 35605 -11510 35660 -11390
rect 35780 -11510 35825 -11390
rect 35945 -11510 35990 -11390
rect 36110 -11510 36155 -11390
rect 36275 -11510 36285 -11390
rect 30785 -11555 36285 -11510
rect 30785 -11675 30795 -11555
rect 30915 -11675 30970 -11555
rect 31090 -11675 31135 -11555
rect 31255 -11675 31300 -11555
rect 31420 -11675 31465 -11555
rect 31585 -11675 31640 -11555
rect 31760 -11675 31805 -11555
rect 31925 -11675 31970 -11555
rect 32090 -11675 32135 -11555
rect 32255 -11675 32310 -11555
rect 32430 -11675 32475 -11555
rect 32595 -11675 32640 -11555
rect 32760 -11675 32805 -11555
rect 32925 -11675 32980 -11555
rect 33100 -11675 33145 -11555
rect 33265 -11675 33310 -11555
rect 33430 -11675 33475 -11555
rect 33595 -11675 33650 -11555
rect 33770 -11675 33815 -11555
rect 33935 -11675 33980 -11555
rect 34100 -11675 34145 -11555
rect 34265 -11675 34320 -11555
rect 34440 -11675 34485 -11555
rect 34605 -11675 34650 -11555
rect 34770 -11675 34815 -11555
rect 34935 -11675 34990 -11555
rect 35110 -11675 35155 -11555
rect 35275 -11675 35320 -11555
rect 35440 -11675 35485 -11555
rect 35605 -11675 35660 -11555
rect 35780 -11675 35825 -11555
rect 35945 -11675 35990 -11555
rect 36110 -11675 36155 -11555
rect 36275 -11675 36285 -11555
rect 30785 -11720 36285 -11675
rect 30785 -11840 30795 -11720
rect 30915 -11840 30970 -11720
rect 31090 -11840 31135 -11720
rect 31255 -11840 31300 -11720
rect 31420 -11840 31465 -11720
rect 31585 -11840 31640 -11720
rect 31760 -11840 31805 -11720
rect 31925 -11840 31970 -11720
rect 32090 -11840 32135 -11720
rect 32255 -11840 32310 -11720
rect 32430 -11840 32475 -11720
rect 32595 -11840 32640 -11720
rect 32760 -11840 32805 -11720
rect 32925 -11840 32980 -11720
rect 33100 -11840 33145 -11720
rect 33265 -11840 33310 -11720
rect 33430 -11840 33475 -11720
rect 33595 -11840 33650 -11720
rect 33770 -11840 33815 -11720
rect 33935 -11840 33980 -11720
rect 34100 -11840 34145 -11720
rect 34265 -11840 34320 -11720
rect 34440 -11840 34485 -11720
rect 34605 -11840 34650 -11720
rect 34770 -11840 34815 -11720
rect 34935 -11840 34990 -11720
rect 35110 -11840 35155 -11720
rect 35275 -11840 35320 -11720
rect 35440 -11840 35485 -11720
rect 35605 -11840 35660 -11720
rect 35780 -11840 35825 -11720
rect 35945 -11840 35990 -11720
rect 36110 -11840 36155 -11720
rect 36275 -11840 36285 -11720
rect 30785 -11885 36285 -11840
rect 30785 -12005 30795 -11885
rect 30915 -12005 30970 -11885
rect 31090 -12005 31135 -11885
rect 31255 -12005 31300 -11885
rect 31420 -12005 31465 -11885
rect 31585 -12005 31640 -11885
rect 31760 -12005 31805 -11885
rect 31925 -12005 31970 -11885
rect 32090 -12005 32135 -11885
rect 32255 -12005 32310 -11885
rect 32430 -12005 32475 -11885
rect 32595 -12005 32640 -11885
rect 32760 -12005 32805 -11885
rect 32925 -12005 32980 -11885
rect 33100 -12005 33145 -11885
rect 33265 -12005 33310 -11885
rect 33430 -12005 33475 -11885
rect 33595 -12005 33650 -11885
rect 33770 -12005 33815 -11885
rect 33935 -12005 33980 -11885
rect 34100 -12005 34145 -11885
rect 34265 -12005 34320 -11885
rect 34440 -12005 34485 -11885
rect 34605 -12005 34650 -11885
rect 34770 -12005 34815 -11885
rect 34935 -12005 34990 -11885
rect 35110 -12005 35155 -11885
rect 35275 -12005 35320 -11885
rect 35440 -12005 35485 -11885
rect 35605 -12005 35660 -11885
rect 35780 -12005 35825 -11885
rect 35945 -12005 35990 -11885
rect 36110 -12005 36155 -11885
rect 36275 -12005 36285 -11885
rect 30785 -12060 36285 -12005
rect 30785 -12180 30795 -12060
rect 30915 -12180 30970 -12060
rect 31090 -12180 31135 -12060
rect 31255 -12180 31300 -12060
rect 31420 -12180 31465 -12060
rect 31585 -12180 31640 -12060
rect 31760 -12180 31805 -12060
rect 31925 -12180 31970 -12060
rect 32090 -12180 32135 -12060
rect 32255 -12180 32310 -12060
rect 32430 -12180 32475 -12060
rect 32595 -12180 32640 -12060
rect 32760 -12180 32805 -12060
rect 32925 -12180 32980 -12060
rect 33100 -12180 33145 -12060
rect 33265 -12180 33310 -12060
rect 33430 -12180 33475 -12060
rect 33595 -12180 33650 -12060
rect 33770 -12180 33815 -12060
rect 33935 -12180 33980 -12060
rect 34100 -12180 34145 -12060
rect 34265 -12180 34320 -12060
rect 34440 -12180 34485 -12060
rect 34605 -12180 34650 -12060
rect 34770 -12180 34815 -12060
rect 34935 -12180 34990 -12060
rect 35110 -12180 35155 -12060
rect 35275 -12180 35320 -12060
rect 35440 -12180 35485 -12060
rect 35605 -12180 35660 -12060
rect 35780 -12180 35825 -12060
rect 35945 -12180 35990 -12060
rect 36110 -12180 36155 -12060
rect 36275 -12180 36285 -12060
rect 30785 -12225 36285 -12180
rect 30785 -12345 30795 -12225
rect 30915 -12345 30970 -12225
rect 31090 -12345 31135 -12225
rect 31255 -12345 31300 -12225
rect 31420 -12345 31465 -12225
rect 31585 -12345 31640 -12225
rect 31760 -12345 31805 -12225
rect 31925 -12345 31970 -12225
rect 32090 -12345 32135 -12225
rect 32255 -12345 32310 -12225
rect 32430 -12345 32475 -12225
rect 32595 -12345 32640 -12225
rect 32760 -12345 32805 -12225
rect 32925 -12345 32980 -12225
rect 33100 -12345 33145 -12225
rect 33265 -12345 33310 -12225
rect 33430 -12345 33475 -12225
rect 33595 -12345 33650 -12225
rect 33770 -12345 33815 -12225
rect 33935 -12345 33980 -12225
rect 34100 -12345 34145 -12225
rect 34265 -12345 34320 -12225
rect 34440 -12345 34485 -12225
rect 34605 -12345 34650 -12225
rect 34770 -12345 34815 -12225
rect 34935 -12345 34990 -12225
rect 35110 -12345 35155 -12225
rect 35275 -12345 35320 -12225
rect 35440 -12345 35485 -12225
rect 35605 -12345 35660 -12225
rect 35780 -12345 35825 -12225
rect 35945 -12345 35990 -12225
rect 36110 -12345 36155 -12225
rect 36275 -12345 36285 -12225
rect 30785 -12390 36285 -12345
rect 30785 -12510 30795 -12390
rect 30915 -12510 30970 -12390
rect 31090 -12510 31135 -12390
rect 31255 -12510 31300 -12390
rect 31420 -12510 31465 -12390
rect 31585 -12510 31640 -12390
rect 31760 -12510 31805 -12390
rect 31925 -12510 31970 -12390
rect 32090 -12510 32135 -12390
rect 32255 -12510 32310 -12390
rect 32430 -12510 32475 -12390
rect 32595 -12510 32640 -12390
rect 32760 -12510 32805 -12390
rect 32925 -12510 32980 -12390
rect 33100 -12510 33145 -12390
rect 33265 -12510 33310 -12390
rect 33430 -12510 33475 -12390
rect 33595 -12510 33650 -12390
rect 33770 -12510 33815 -12390
rect 33935 -12510 33980 -12390
rect 34100 -12510 34145 -12390
rect 34265 -12510 34320 -12390
rect 34440 -12510 34485 -12390
rect 34605 -12510 34650 -12390
rect 34770 -12510 34815 -12390
rect 34935 -12510 34990 -12390
rect 35110 -12510 35155 -12390
rect 35275 -12510 35320 -12390
rect 35440 -12510 35485 -12390
rect 35605 -12510 35660 -12390
rect 35780 -12510 35825 -12390
rect 35945 -12510 35990 -12390
rect 36110 -12510 36155 -12390
rect 36275 -12510 36285 -12390
rect 30785 -12555 36285 -12510
rect 30785 -12675 30795 -12555
rect 30915 -12675 30970 -12555
rect 31090 -12675 31135 -12555
rect 31255 -12675 31300 -12555
rect 31420 -12675 31465 -12555
rect 31585 -12675 31640 -12555
rect 31760 -12675 31805 -12555
rect 31925 -12675 31970 -12555
rect 32090 -12675 32135 -12555
rect 32255 -12675 32310 -12555
rect 32430 -12675 32475 -12555
rect 32595 -12675 32640 -12555
rect 32760 -12675 32805 -12555
rect 32925 -12675 32980 -12555
rect 33100 -12675 33145 -12555
rect 33265 -12675 33310 -12555
rect 33430 -12675 33475 -12555
rect 33595 -12675 33650 -12555
rect 33770 -12675 33815 -12555
rect 33935 -12675 33980 -12555
rect 34100 -12675 34145 -12555
rect 34265 -12675 34320 -12555
rect 34440 -12675 34485 -12555
rect 34605 -12675 34650 -12555
rect 34770 -12675 34815 -12555
rect 34935 -12675 34990 -12555
rect 35110 -12675 35155 -12555
rect 35275 -12675 35320 -12555
rect 35440 -12675 35485 -12555
rect 35605 -12675 35660 -12555
rect 35780 -12675 35825 -12555
rect 35945 -12675 35990 -12555
rect 36110 -12675 36155 -12555
rect 36275 -12675 36285 -12555
rect 30785 -12730 36285 -12675
rect 30785 -12850 30795 -12730
rect 30915 -12850 30970 -12730
rect 31090 -12850 31135 -12730
rect 31255 -12850 31300 -12730
rect 31420 -12850 31465 -12730
rect 31585 -12850 31640 -12730
rect 31760 -12850 31805 -12730
rect 31925 -12850 31970 -12730
rect 32090 -12850 32135 -12730
rect 32255 -12850 32310 -12730
rect 32430 -12850 32475 -12730
rect 32595 -12850 32640 -12730
rect 32760 -12850 32805 -12730
rect 32925 -12850 32980 -12730
rect 33100 -12850 33145 -12730
rect 33265 -12850 33310 -12730
rect 33430 -12850 33475 -12730
rect 33595 -12850 33650 -12730
rect 33770 -12850 33815 -12730
rect 33935 -12850 33980 -12730
rect 34100 -12850 34145 -12730
rect 34265 -12850 34320 -12730
rect 34440 -12850 34485 -12730
rect 34605 -12850 34650 -12730
rect 34770 -12850 34815 -12730
rect 34935 -12850 34990 -12730
rect 35110 -12850 35155 -12730
rect 35275 -12850 35320 -12730
rect 35440 -12850 35485 -12730
rect 35605 -12850 35660 -12730
rect 35780 -12850 35825 -12730
rect 35945 -12850 35990 -12730
rect 36110 -12850 36155 -12730
rect 36275 -12850 36285 -12730
rect 30785 -12895 36285 -12850
rect 30785 -13015 30795 -12895
rect 30915 -13015 30970 -12895
rect 31090 -13015 31135 -12895
rect 31255 -13015 31300 -12895
rect 31420 -13015 31465 -12895
rect 31585 -13015 31640 -12895
rect 31760 -13015 31805 -12895
rect 31925 -13015 31970 -12895
rect 32090 -13015 32135 -12895
rect 32255 -13015 32310 -12895
rect 32430 -13015 32475 -12895
rect 32595 -13015 32640 -12895
rect 32760 -13015 32805 -12895
rect 32925 -13015 32980 -12895
rect 33100 -13015 33145 -12895
rect 33265 -13015 33310 -12895
rect 33430 -13015 33475 -12895
rect 33595 -13015 33650 -12895
rect 33770 -13015 33815 -12895
rect 33935 -13015 33980 -12895
rect 34100 -13015 34145 -12895
rect 34265 -13015 34320 -12895
rect 34440 -13015 34485 -12895
rect 34605 -13015 34650 -12895
rect 34770 -13015 34815 -12895
rect 34935 -13015 34990 -12895
rect 35110 -13015 35155 -12895
rect 35275 -13015 35320 -12895
rect 35440 -13015 35485 -12895
rect 35605 -13015 35660 -12895
rect 35780 -13015 35825 -12895
rect 35945 -13015 35990 -12895
rect 36110 -13015 36155 -12895
rect 36275 -13015 36285 -12895
rect 30785 -13060 36285 -13015
rect 30785 -13180 30795 -13060
rect 30915 -13180 30970 -13060
rect 31090 -13180 31135 -13060
rect 31255 -13180 31300 -13060
rect 31420 -13180 31465 -13060
rect 31585 -13180 31640 -13060
rect 31760 -13180 31805 -13060
rect 31925 -13180 31970 -13060
rect 32090 -13180 32135 -13060
rect 32255 -13180 32310 -13060
rect 32430 -13180 32475 -13060
rect 32595 -13180 32640 -13060
rect 32760 -13180 32805 -13060
rect 32925 -13180 32980 -13060
rect 33100 -13180 33145 -13060
rect 33265 -13180 33310 -13060
rect 33430 -13180 33475 -13060
rect 33595 -13180 33650 -13060
rect 33770 -13180 33815 -13060
rect 33935 -13180 33980 -13060
rect 34100 -13180 34145 -13060
rect 34265 -13180 34320 -13060
rect 34440 -13180 34485 -13060
rect 34605 -13180 34650 -13060
rect 34770 -13180 34815 -13060
rect 34935 -13180 34990 -13060
rect 35110 -13180 35155 -13060
rect 35275 -13180 35320 -13060
rect 35440 -13180 35485 -13060
rect 35605 -13180 35660 -13060
rect 35780 -13180 35825 -13060
rect 35945 -13180 35990 -13060
rect 36110 -13180 36155 -13060
rect 36275 -13180 36285 -13060
rect 30785 -13225 36285 -13180
rect 30785 -13345 30795 -13225
rect 30915 -13345 30970 -13225
rect 31090 -13345 31135 -13225
rect 31255 -13345 31300 -13225
rect 31420 -13345 31465 -13225
rect 31585 -13345 31640 -13225
rect 31760 -13345 31805 -13225
rect 31925 -13345 31970 -13225
rect 32090 -13345 32135 -13225
rect 32255 -13345 32310 -13225
rect 32430 -13345 32475 -13225
rect 32595 -13345 32640 -13225
rect 32760 -13345 32805 -13225
rect 32925 -13345 32980 -13225
rect 33100 -13345 33145 -13225
rect 33265 -13345 33310 -13225
rect 33430 -13345 33475 -13225
rect 33595 -13345 33650 -13225
rect 33770 -13345 33815 -13225
rect 33935 -13345 33980 -13225
rect 34100 -13345 34145 -13225
rect 34265 -13345 34320 -13225
rect 34440 -13345 34485 -13225
rect 34605 -13345 34650 -13225
rect 34770 -13345 34815 -13225
rect 34935 -13345 34990 -13225
rect 35110 -13345 35155 -13225
rect 35275 -13345 35320 -13225
rect 35440 -13345 35485 -13225
rect 35605 -13345 35660 -13225
rect 35780 -13345 35825 -13225
rect 35945 -13345 35990 -13225
rect 36110 -13345 36155 -13225
rect 36275 -13345 36285 -13225
rect 30785 -13400 36285 -13345
rect 30785 -13520 30795 -13400
rect 30915 -13520 30970 -13400
rect 31090 -13520 31135 -13400
rect 31255 -13520 31300 -13400
rect 31420 -13520 31465 -13400
rect 31585 -13520 31640 -13400
rect 31760 -13520 31805 -13400
rect 31925 -13520 31970 -13400
rect 32090 -13520 32135 -13400
rect 32255 -13520 32310 -13400
rect 32430 -13520 32475 -13400
rect 32595 -13520 32640 -13400
rect 32760 -13520 32805 -13400
rect 32925 -13520 32980 -13400
rect 33100 -13520 33145 -13400
rect 33265 -13520 33310 -13400
rect 33430 -13520 33475 -13400
rect 33595 -13520 33650 -13400
rect 33770 -13520 33815 -13400
rect 33935 -13520 33980 -13400
rect 34100 -13520 34145 -13400
rect 34265 -13520 34320 -13400
rect 34440 -13520 34485 -13400
rect 34605 -13520 34650 -13400
rect 34770 -13520 34815 -13400
rect 34935 -13520 34990 -13400
rect 35110 -13520 35155 -13400
rect 35275 -13520 35320 -13400
rect 35440 -13520 35485 -13400
rect 35605 -13520 35660 -13400
rect 35780 -13520 35825 -13400
rect 35945 -13520 35990 -13400
rect 36110 -13520 36155 -13400
rect 36275 -13520 36285 -13400
rect 30785 -13565 36285 -13520
rect 30785 -13685 30795 -13565
rect 30915 -13685 30970 -13565
rect 31090 -13685 31135 -13565
rect 31255 -13685 31300 -13565
rect 31420 -13685 31465 -13565
rect 31585 -13685 31640 -13565
rect 31760 -13685 31805 -13565
rect 31925 -13685 31970 -13565
rect 32090 -13685 32135 -13565
rect 32255 -13685 32310 -13565
rect 32430 -13685 32475 -13565
rect 32595 -13685 32640 -13565
rect 32760 -13685 32805 -13565
rect 32925 -13685 32980 -13565
rect 33100 -13685 33145 -13565
rect 33265 -13685 33310 -13565
rect 33430 -13685 33475 -13565
rect 33595 -13685 33650 -13565
rect 33770 -13685 33815 -13565
rect 33935 -13685 33980 -13565
rect 34100 -13685 34145 -13565
rect 34265 -13685 34320 -13565
rect 34440 -13685 34485 -13565
rect 34605 -13685 34650 -13565
rect 34770 -13685 34815 -13565
rect 34935 -13685 34990 -13565
rect 35110 -13685 35155 -13565
rect 35275 -13685 35320 -13565
rect 35440 -13685 35485 -13565
rect 35605 -13685 35660 -13565
rect 35780 -13685 35825 -13565
rect 35945 -13685 35990 -13565
rect 36110 -13685 36155 -13565
rect 36275 -13685 36285 -13565
rect 30785 -13730 36285 -13685
rect 30785 -13850 30795 -13730
rect 30915 -13850 30970 -13730
rect 31090 -13850 31135 -13730
rect 31255 -13850 31300 -13730
rect 31420 -13850 31465 -13730
rect 31585 -13850 31640 -13730
rect 31760 -13850 31805 -13730
rect 31925 -13850 31970 -13730
rect 32090 -13850 32135 -13730
rect 32255 -13850 32310 -13730
rect 32430 -13850 32475 -13730
rect 32595 -13850 32640 -13730
rect 32760 -13850 32805 -13730
rect 32925 -13850 32980 -13730
rect 33100 -13850 33145 -13730
rect 33265 -13850 33310 -13730
rect 33430 -13850 33475 -13730
rect 33595 -13850 33650 -13730
rect 33770 -13850 33815 -13730
rect 33935 -13850 33980 -13730
rect 34100 -13850 34145 -13730
rect 34265 -13850 34320 -13730
rect 34440 -13850 34485 -13730
rect 34605 -13850 34650 -13730
rect 34770 -13850 34815 -13730
rect 34935 -13850 34990 -13730
rect 35110 -13850 35155 -13730
rect 35275 -13850 35320 -13730
rect 35440 -13850 35485 -13730
rect 35605 -13850 35660 -13730
rect 35780 -13850 35825 -13730
rect 35945 -13850 35990 -13730
rect 36110 -13850 36155 -13730
rect 36275 -13850 36285 -13730
rect 30785 -13895 36285 -13850
rect 30785 -14015 30795 -13895
rect 30915 -14015 30970 -13895
rect 31090 -14015 31135 -13895
rect 31255 -14015 31300 -13895
rect 31420 -14015 31465 -13895
rect 31585 -14015 31640 -13895
rect 31760 -14015 31805 -13895
rect 31925 -14015 31970 -13895
rect 32090 -14015 32135 -13895
rect 32255 -14015 32310 -13895
rect 32430 -14015 32475 -13895
rect 32595 -14015 32640 -13895
rect 32760 -14015 32805 -13895
rect 32925 -14015 32980 -13895
rect 33100 -14015 33145 -13895
rect 33265 -14015 33310 -13895
rect 33430 -14015 33475 -13895
rect 33595 -14015 33650 -13895
rect 33770 -14015 33815 -13895
rect 33935 -14015 33980 -13895
rect 34100 -14015 34145 -13895
rect 34265 -14015 34320 -13895
rect 34440 -14015 34485 -13895
rect 34605 -14015 34650 -13895
rect 34770 -14015 34815 -13895
rect 34935 -14015 34990 -13895
rect 35110 -14015 35155 -13895
rect 35275 -14015 35320 -13895
rect 35440 -14015 35485 -13895
rect 35605 -14015 35660 -13895
rect 35780 -14015 35825 -13895
rect 35945 -14015 35990 -13895
rect 36110 -14015 36155 -13895
rect 36275 -14015 36285 -13895
rect 30785 -14070 36285 -14015
rect 30785 -14190 30795 -14070
rect 30915 -14190 30970 -14070
rect 31090 -14190 31135 -14070
rect 31255 -14190 31300 -14070
rect 31420 -14190 31465 -14070
rect 31585 -14190 31640 -14070
rect 31760 -14190 31805 -14070
rect 31925 -14190 31970 -14070
rect 32090 -14190 32135 -14070
rect 32255 -14190 32310 -14070
rect 32430 -14190 32475 -14070
rect 32595 -14190 32640 -14070
rect 32760 -14190 32805 -14070
rect 32925 -14190 32980 -14070
rect 33100 -14190 33145 -14070
rect 33265 -14190 33310 -14070
rect 33430 -14190 33475 -14070
rect 33595 -14190 33650 -14070
rect 33770 -14190 33815 -14070
rect 33935 -14190 33980 -14070
rect 34100 -14190 34145 -14070
rect 34265 -14190 34320 -14070
rect 34440 -14190 34485 -14070
rect 34605 -14190 34650 -14070
rect 34770 -14190 34815 -14070
rect 34935 -14190 34990 -14070
rect 35110 -14190 35155 -14070
rect 35275 -14190 35320 -14070
rect 35440 -14190 35485 -14070
rect 35605 -14190 35660 -14070
rect 35780 -14190 35825 -14070
rect 35945 -14190 35990 -14070
rect 36110 -14190 36155 -14070
rect 36275 -14190 36285 -14070
rect 30785 -14235 36285 -14190
rect 30785 -14355 30795 -14235
rect 30915 -14355 30970 -14235
rect 31090 -14355 31135 -14235
rect 31255 -14355 31300 -14235
rect 31420 -14355 31465 -14235
rect 31585 -14355 31640 -14235
rect 31760 -14355 31805 -14235
rect 31925 -14355 31970 -14235
rect 32090 -14355 32135 -14235
rect 32255 -14355 32310 -14235
rect 32430 -14355 32475 -14235
rect 32595 -14355 32640 -14235
rect 32760 -14355 32805 -14235
rect 32925 -14355 32980 -14235
rect 33100 -14355 33145 -14235
rect 33265 -14355 33310 -14235
rect 33430 -14355 33475 -14235
rect 33595 -14355 33650 -14235
rect 33770 -14355 33815 -14235
rect 33935 -14355 33980 -14235
rect 34100 -14355 34145 -14235
rect 34265 -14355 34320 -14235
rect 34440 -14355 34485 -14235
rect 34605 -14355 34650 -14235
rect 34770 -14355 34815 -14235
rect 34935 -14355 34990 -14235
rect 35110 -14355 35155 -14235
rect 35275 -14355 35320 -14235
rect 35440 -14355 35485 -14235
rect 35605 -14355 35660 -14235
rect 35780 -14355 35825 -14235
rect 35945 -14355 35990 -14235
rect 36110 -14355 36155 -14235
rect 36275 -14355 36285 -14235
rect 30785 -14400 36285 -14355
rect 30785 -14520 30795 -14400
rect 30915 -14520 30970 -14400
rect 31090 -14520 31135 -14400
rect 31255 -14520 31300 -14400
rect 31420 -14520 31465 -14400
rect 31585 -14520 31640 -14400
rect 31760 -14520 31805 -14400
rect 31925 -14520 31970 -14400
rect 32090 -14520 32135 -14400
rect 32255 -14520 32310 -14400
rect 32430 -14520 32475 -14400
rect 32595 -14520 32640 -14400
rect 32760 -14520 32805 -14400
rect 32925 -14520 32980 -14400
rect 33100 -14520 33145 -14400
rect 33265 -14520 33310 -14400
rect 33430 -14520 33475 -14400
rect 33595 -14520 33650 -14400
rect 33770 -14520 33815 -14400
rect 33935 -14520 33980 -14400
rect 34100 -14520 34145 -14400
rect 34265 -14520 34320 -14400
rect 34440 -14520 34485 -14400
rect 34605 -14520 34650 -14400
rect 34770 -14520 34815 -14400
rect 34935 -14520 34990 -14400
rect 35110 -14520 35155 -14400
rect 35275 -14520 35320 -14400
rect 35440 -14520 35485 -14400
rect 35605 -14520 35660 -14400
rect 35780 -14520 35825 -14400
rect 35945 -14520 35990 -14400
rect 36110 -14520 36155 -14400
rect 36275 -14520 36285 -14400
rect 30785 -14565 36285 -14520
rect 30785 -14685 30795 -14565
rect 30915 -14685 30970 -14565
rect 31090 -14685 31135 -14565
rect 31255 -14685 31300 -14565
rect 31420 -14685 31465 -14565
rect 31585 -14685 31640 -14565
rect 31760 -14685 31805 -14565
rect 31925 -14685 31970 -14565
rect 32090 -14685 32135 -14565
rect 32255 -14685 32310 -14565
rect 32430 -14685 32475 -14565
rect 32595 -14685 32640 -14565
rect 32760 -14685 32805 -14565
rect 32925 -14685 32980 -14565
rect 33100 -14685 33145 -14565
rect 33265 -14685 33310 -14565
rect 33430 -14685 33475 -14565
rect 33595 -14685 33650 -14565
rect 33770 -14685 33815 -14565
rect 33935 -14685 33980 -14565
rect 34100 -14685 34145 -14565
rect 34265 -14685 34320 -14565
rect 34440 -14685 34485 -14565
rect 34605 -14685 34650 -14565
rect 34770 -14685 34815 -14565
rect 34935 -14685 34990 -14565
rect 35110 -14685 35155 -14565
rect 35275 -14685 35320 -14565
rect 35440 -14685 35485 -14565
rect 35605 -14685 35660 -14565
rect 35780 -14685 35825 -14565
rect 35945 -14685 35990 -14565
rect 36110 -14685 36155 -14565
rect 36275 -14685 36285 -14565
rect 30785 -14740 36285 -14685
rect 30785 -14860 30795 -14740
rect 30915 -14860 30970 -14740
rect 31090 -14860 31135 -14740
rect 31255 -14860 31300 -14740
rect 31420 -14860 31465 -14740
rect 31585 -14860 31640 -14740
rect 31760 -14860 31805 -14740
rect 31925 -14860 31970 -14740
rect 32090 -14860 32135 -14740
rect 32255 -14860 32310 -14740
rect 32430 -14860 32475 -14740
rect 32595 -14860 32640 -14740
rect 32760 -14860 32805 -14740
rect 32925 -14860 32980 -14740
rect 33100 -14860 33145 -14740
rect 33265 -14860 33310 -14740
rect 33430 -14860 33475 -14740
rect 33595 -14860 33650 -14740
rect 33770 -14860 33815 -14740
rect 33935 -14860 33980 -14740
rect 34100 -14860 34145 -14740
rect 34265 -14860 34320 -14740
rect 34440 -14860 34485 -14740
rect 34605 -14860 34650 -14740
rect 34770 -14860 34815 -14740
rect 34935 -14860 34990 -14740
rect 35110 -14860 35155 -14740
rect 35275 -14860 35320 -14740
rect 35440 -14860 35485 -14740
rect 35605 -14860 35660 -14740
rect 35780 -14860 35825 -14740
rect 35945 -14860 35990 -14740
rect 36110 -14860 36155 -14740
rect 36275 -14860 36285 -14740
rect 30785 -14905 36285 -14860
rect 30785 -15025 30795 -14905
rect 30915 -15025 30970 -14905
rect 31090 -15025 31135 -14905
rect 31255 -15025 31300 -14905
rect 31420 -15025 31465 -14905
rect 31585 -15025 31640 -14905
rect 31760 -15025 31805 -14905
rect 31925 -15025 31970 -14905
rect 32090 -15025 32135 -14905
rect 32255 -15025 32310 -14905
rect 32430 -15025 32475 -14905
rect 32595 -15025 32640 -14905
rect 32760 -15025 32805 -14905
rect 32925 -15025 32980 -14905
rect 33100 -15025 33145 -14905
rect 33265 -15025 33310 -14905
rect 33430 -15025 33475 -14905
rect 33595 -15025 33650 -14905
rect 33770 -15025 33815 -14905
rect 33935 -15025 33980 -14905
rect 34100 -15025 34145 -14905
rect 34265 -15025 34320 -14905
rect 34440 -15025 34485 -14905
rect 34605 -15025 34650 -14905
rect 34770 -15025 34815 -14905
rect 34935 -15025 34990 -14905
rect 35110 -15025 35155 -14905
rect 35275 -15025 35320 -14905
rect 35440 -15025 35485 -14905
rect 35605 -15025 35660 -14905
rect 35780 -15025 35825 -14905
rect 35945 -15025 35990 -14905
rect 36110 -15025 36155 -14905
rect 36275 -15025 36285 -14905
rect 30785 -15070 36285 -15025
rect 30785 -15190 30795 -15070
rect 30915 -15190 30970 -15070
rect 31090 -15190 31135 -15070
rect 31255 -15190 31300 -15070
rect 31420 -15190 31465 -15070
rect 31585 -15190 31640 -15070
rect 31760 -15190 31805 -15070
rect 31925 -15190 31970 -15070
rect 32090 -15190 32135 -15070
rect 32255 -15190 32310 -15070
rect 32430 -15190 32475 -15070
rect 32595 -15190 32640 -15070
rect 32760 -15190 32805 -15070
rect 32925 -15190 32980 -15070
rect 33100 -15190 33145 -15070
rect 33265 -15190 33310 -15070
rect 33430 -15190 33475 -15070
rect 33595 -15190 33650 -15070
rect 33770 -15190 33815 -15070
rect 33935 -15190 33980 -15070
rect 34100 -15190 34145 -15070
rect 34265 -15190 34320 -15070
rect 34440 -15190 34485 -15070
rect 34605 -15190 34650 -15070
rect 34770 -15190 34815 -15070
rect 34935 -15190 34990 -15070
rect 35110 -15190 35155 -15070
rect 35275 -15190 35320 -15070
rect 35440 -15190 35485 -15070
rect 35605 -15190 35660 -15070
rect 35780 -15190 35825 -15070
rect 35945 -15190 35990 -15070
rect 36110 -15190 36155 -15070
rect 36275 -15190 36285 -15070
rect 30785 -15235 36285 -15190
rect 30785 -15355 30795 -15235
rect 30915 -15355 30970 -15235
rect 31090 -15355 31135 -15235
rect 31255 -15355 31300 -15235
rect 31420 -15355 31465 -15235
rect 31585 -15355 31640 -15235
rect 31760 -15355 31805 -15235
rect 31925 -15355 31970 -15235
rect 32090 -15355 32135 -15235
rect 32255 -15355 32310 -15235
rect 32430 -15355 32475 -15235
rect 32595 -15355 32640 -15235
rect 32760 -15355 32805 -15235
rect 32925 -15355 32980 -15235
rect 33100 -15355 33145 -15235
rect 33265 -15355 33310 -15235
rect 33430 -15355 33475 -15235
rect 33595 -15355 33650 -15235
rect 33770 -15355 33815 -15235
rect 33935 -15355 33980 -15235
rect 34100 -15355 34145 -15235
rect 34265 -15355 34320 -15235
rect 34440 -15355 34485 -15235
rect 34605 -15355 34650 -15235
rect 34770 -15355 34815 -15235
rect 34935 -15355 34990 -15235
rect 35110 -15355 35155 -15235
rect 35275 -15355 35320 -15235
rect 35440 -15355 35485 -15235
rect 35605 -15355 35660 -15235
rect 35780 -15355 35825 -15235
rect 35945 -15355 35990 -15235
rect 36110 -15355 36155 -15235
rect 36275 -15355 36285 -15235
rect 30785 -15410 36285 -15355
rect 30785 -15530 30795 -15410
rect 30915 -15530 30970 -15410
rect 31090 -15530 31135 -15410
rect 31255 -15530 31300 -15410
rect 31420 -15530 31465 -15410
rect 31585 -15530 31640 -15410
rect 31760 -15530 31805 -15410
rect 31925 -15530 31970 -15410
rect 32090 -15530 32135 -15410
rect 32255 -15530 32310 -15410
rect 32430 -15530 32475 -15410
rect 32595 -15530 32640 -15410
rect 32760 -15530 32805 -15410
rect 32925 -15530 32980 -15410
rect 33100 -15530 33145 -15410
rect 33265 -15530 33310 -15410
rect 33430 -15530 33475 -15410
rect 33595 -15530 33650 -15410
rect 33770 -15530 33815 -15410
rect 33935 -15530 33980 -15410
rect 34100 -15530 34145 -15410
rect 34265 -15530 34320 -15410
rect 34440 -15530 34485 -15410
rect 34605 -15530 34650 -15410
rect 34770 -15530 34815 -15410
rect 34935 -15530 34990 -15410
rect 35110 -15530 35155 -15410
rect 35275 -15530 35320 -15410
rect 35440 -15530 35485 -15410
rect 35605 -15530 35660 -15410
rect 35780 -15530 35825 -15410
rect 35945 -15530 35990 -15410
rect 36110 -15530 36155 -15410
rect 36275 -15530 36285 -15410
rect 30785 -15540 36285 -15530
rect 36475 -10050 41975 -10040
rect 36475 -10170 36485 -10050
rect 36605 -10170 36660 -10050
rect 36780 -10170 36825 -10050
rect 36945 -10170 36990 -10050
rect 37110 -10170 37155 -10050
rect 37275 -10170 37330 -10050
rect 37450 -10170 37495 -10050
rect 37615 -10170 37660 -10050
rect 37780 -10170 37825 -10050
rect 37945 -10170 38000 -10050
rect 38120 -10170 38165 -10050
rect 38285 -10170 38330 -10050
rect 38450 -10170 38495 -10050
rect 38615 -10170 38670 -10050
rect 38790 -10170 38835 -10050
rect 38955 -10170 39000 -10050
rect 39120 -10170 39165 -10050
rect 39285 -10170 39340 -10050
rect 39460 -10170 39505 -10050
rect 39625 -10170 39670 -10050
rect 39790 -10170 39835 -10050
rect 39955 -10170 40010 -10050
rect 40130 -10170 40175 -10050
rect 40295 -10170 40340 -10050
rect 40460 -10170 40505 -10050
rect 40625 -10170 40680 -10050
rect 40800 -10170 40845 -10050
rect 40965 -10170 41010 -10050
rect 41130 -10170 41175 -10050
rect 41295 -10170 41350 -10050
rect 41470 -10170 41515 -10050
rect 41635 -10170 41680 -10050
rect 41800 -10170 41845 -10050
rect 41965 -10170 41975 -10050
rect 36475 -10215 41975 -10170
rect 36475 -10335 36485 -10215
rect 36605 -10335 36660 -10215
rect 36780 -10335 36825 -10215
rect 36945 -10335 36990 -10215
rect 37110 -10335 37155 -10215
rect 37275 -10335 37330 -10215
rect 37450 -10335 37495 -10215
rect 37615 -10335 37660 -10215
rect 37780 -10335 37825 -10215
rect 37945 -10335 38000 -10215
rect 38120 -10335 38165 -10215
rect 38285 -10335 38330 -10215
rect 38450 -10335 38495 -10215
rect 38615 -10335 38670 -10215
rect 38790 -10335 38835 -10215
rect 38955 -10335 39000 -10215
rect 39120 -10335 39165 -10215
rect 39285 -10335 39340 -10215
rect 39460 -10335 39505 -10215
rect 39625 -10335 39670 -10215
rect 39790 -10335 39835 -10215
rect 39955 -10335 40010 -10215
rect 40130 -10335 40175 -10215
rect 40295 -10335 40340 -10215
rect 40460 -10335 40505 -10215
rect 40625 -10335 40680 -10215
rect 40800 -10335 40845 -10215
rect 40965 -10335 41010 -10215
rect 41130 -10335 41175 -10215
rect 41295 -10335 41350 -10215
rect 41470 -10335 41515 -10215
rect 41635 -10335 41680 -10215
rect 41800 -10335 41845 -10215
rect 41965 -10335 41975 -10215
rect 36475 -10380 41975 -10335
rect 36475 -10500 36485 -10380
rect 36605 -10500 36660 -10380
rect 36780 -10500 36825 -10380
rect 36945 -10500 36990 -10380
rect 37110 -10500 37155 -10380
rect 37275 -10500 37330 -10380
rect 37450 -10500 37495 -10380
rect 37615 -10500 37660 -10380
rect 37780 -10500 37825 -10380
rect 37945 -10500 38000 -10380
rect 38120 -10500 38165 -10380
rect 38285 -10500 38330 -10380
rect 38450 -10500 38495 -10380
rect 38615 -10500 38670 -10380
rect 38790 -10500 38835 -10380
rect 38955 -10500 39000 -10380
rect 39120 -10500 39165 -10380
rect 39285 -10500 39340 -10380
rect 39460 -10500 39505 -10380
rect 39625 -10500 39670 -10380
rect 39790 -10500 39835 -10380
rect 39955 -10500 40010 -10380
rect 40130 -10500 40175 -10380
rect 40295 -10500 40340 -10380
rect 40460 -10500 40505 -10380
rect 40625 -10500 40680 -10380
rect 40800 -10500 40845 -10380
rect 40965 -10500 41010 -10380
rect 41130 -10500 41175 -10380
rect 41295 -10500 41350 -10380
rect 41470 -10500 41515 -10380
rect 41635 -10500 41680 -10380
rect 41800 -10500 41845 -10380
rect 41965 -10500 41975 -10380
rect 36475 -10545 41975 -10500
rect 36475 -10665 36485 -10545
rect 36605 -10665 36660 -10545
rect 36780 -10665 36825 -10545
rect 36945 -10665 36990 -10545
rect 37110 -10665 37155 -10545
rect 37275 -10665 37330 -10545
rect 37450 -10665 37495 -10545
rect 37615 -10665 37660 -10545
rect 37780 -10665 37825 -10545
rect 37945 -10665 38000 -10545
rect 38120 -10665 38165 -10545
rect 38285 -10665 38330 -10545
rect 38450 -10665 38495 -10545
rect 38615 -10665 38670 -10545
rect 38790 -10665 38835 -10545
rect 38955 -10665 39000 -10545
rect 39120 -10665 39165 -10545
rect 39285 -10665 39340 -10545
rect 39460 -10665 39505 -10545
rect 39625 -10665 39670 -10545
rect 39790 -10665 39835 -10545
rect 39955 -10665 40010 -10545
rect 40130 -10665 40175 -10545
rect 40295 -10665 40340 -10545
rect 40460 -10665 40505 -10545
rect 40625 -10665 40680 -10545
rect 40800 -10665 40845 -10545
rect 40965 -10665 41010 -10545
rect 41130 -10665 41175 -10545
rect 41295 -10665 41350 -10545
rect 41470 -10665 41515 -10545
rect 41635 -10665 41680 -10545
rect 41800 -10665 41845 -10545
rect 41965 -10665 41975 -10545
rect 36475 -10720 41975 -10665
rect 36475 -10840 36485 -10720
rect 36605 -10840 36660 -10720
rect 36780 -10840 36825 -10720
rect 36945 -10840 36990 -10720
rect 37110 -10840 37155 -10720
rect 37275 -10840 37330 -10720
rect 37450 -10840 37495 -10720
rect 37615 -10840 37660 -10720
rect 37780 -10840 37825 -10720
rect 37945 -10840 38000 -10720
rect 38120 -10840 38165 -10720
rect 38285 -10840 38330 -10720
rect 38450 -10840 38495 -10720
rect 38615 -10840 38670 -10720
rect 38790 -10840 38835 -10720
rect 38955 -10840 39000 -10720
rect 39120 -10840 39165 -10720
rect 39285 -10840 39340 -10720
rect 39460 -10840 39505 -10720
rect 39625 -10840 39670 -10720
rect 39790 -10840 39835 -10720
rect 39955 -10840 40010 -10720
rect 40130 -10840 40175 -10720
rect 40295 -10840 40340 -10720
rect 40460 -10840 40505 -10720
rect 40625 -10840 40680 -10720
rect 40800 -10840 40845 -10720
rect 40965 -10840 41010 -10720
rect 41130 -10840 41175 -10720
rect 41295 -10840 41350 -10720
rect 41470 -10840 41515 -10720
rect 41635 -10840 41680 -10720
rect 41800 -10840 41845 -10720
rect 41965 -10840 41975 -10720
rect 36475 -10885 41975 -10840
rect 36475 -11005 36485 -10885
rect 36605 -11005 36660 -10885
rect 36780 -11005 36825 -10885
rect 36945 -11005 36990 -10885
rect 37110 -11005 37155 -10885
rect 37275 -11005 37330 -10885
rect 37450 -11005 37495 -10885
rect 37615 -11005 37660 -10885
rect 37780 -11005 37825 -10885
rect 37945 -11005 38000 -10885
rect 38120 -11005 38165 -10885
rect 38285 -11005 38330 -10885
rect 38450 -11005 38495 -10885
rect 38615 -11005 38670 -10885
rect 38790 -11005 38835 -10885
rect 38955 -11005 39000 -10885
rect 39120 -11005 39165 -10885
rect 39285 -11005 39340 -10885
rect 39460 -11005 39505 -10885
rect 39625 -11005 39670 -10885
rect 39790 -11005 39835 -10885
rect 39955 -11005 40010 -10885
rect 40130 -11005 40175 -10885
rect 40295 -11005 40340 -10885
rect 40460 -11005 40505 -10885
rect 40625 -11005 40680 -10885
rect 40800 -11005 40845 -10885
rect 40965 -11005 41010 -10885
rect 41130 -11005 41175 -10885
rect 41295 -11005 41350 -10885
rect 41470 -11005 41515 -10885
rect 41635 -11005 41680 -10885
rect 41800 -11005 41845 -10885
rect 41965 -11005 41975 -10885
rect 36475 -11050 41975 -11005
rect 36475 -11170 36485 -11050
rect 36605 -11170 36660 -11050
rect 36780 -11170 36825 -11050
rect 36945 -11170 36990 -11050
rect 37110 -11170 37155 -11050
rect 37275 -11170 37330 -11050
rect 37450 -11170 37495 -11050
rect 37615 -11170 37660 -11050
rect 37780 -11170 37825 -11050
rect 37945 -11170 38000 -11050
rect 38120 -11170 38165 -11050
rect 38285 -11170 38330 -11050
rect 38450 -11170 38495 -11050
rect 38615 -11170 38670 -11050
rect 38790 -11170 38835 -11050
rect 38955 -11170 39000 -11050
rect 39120 -11170 39165 -11050
rect 39285 -11170 39340 -11050
rect 39460 -11170 39505 -11050
rect 39625 -11170 39670 -11050
rect 39790 -11170 39835 -11050
rect 39955 -11170 40010 -11050
rect 40130 -11170 40175 -11050
rect 40295 -11170 40340 -11050
rect 40460 -11170 40505 -11050
rect 40625 -11170 40680 -11050
rect 40800 -11170 40845 -11050
rect 40965 -11170 41010 -11050
rect 41130 -11170 41175 -11050
rect 41295 -11170 41350 -11050
rect 41470 -11170 41515 -11050
rect 41635 -11170 41680 -11050
rect 41800 -11170 41845 -11050
rect 41965 -11170 41975 -11050
rect 36475 -11215 41975 -11170
rect 36475 -11335 36485 -11215
rect 36605 -11335 36660 -11215
rect 36780 -11335 36825 -11215
rect 36945 -11335 36990 -11215
rect 37110 -11335 37155 -11215
rect 37275 -11335 37330 -11215
rect 37450 -11335 37495 -11215
rect 37615 -11335 37660 -11215
rect 37780 -11335 37825 -11215
rect 37945 -11335 38000 -11215
rect 38120 -11335 38165 -11215
rect 38285 -11335 38330 -11215
rect 38450 -11335 38495 -11215
rect 38615 -11335 38670 -11215
rect 38790 -11335 38835 -11215
rect 38955 -11335 39000 -11215
rect 39120 -11335 39165 -11215
rect 39285 -11335 39340 -11215
rect 39460 -11335 39505 -11215
rect 39625 -11335 39670 -11215
rect 39790 -11335 39835 -11215
rect 39955 -11335 40010 -11215
rect 40130 -11335 40175 -11215
rect 40295 -11335 40340 -11215
rect 40460 -11335 40505 -11215
rect 40625 -11335 40680 -11215
rect 40800 -11335 40845 -11215
rect 40965 -11335 41010 -11215
rect 41130 -11335 41175 -11215
rect 41295 -11335 41350 -11215
rect 41470 -11335 41515 -11215
rect 41635 -11335 41680 -11215
rect 41800 -11335 41845 -11215
rect 41965 -11335 41975 -11215
rect 36475 -11390 41975 -11335
rect 36475 -11510 36485 -11390
rect 36605 -11510 36660 -11390
rect 36780 -11510 36825 -11390
rect 36945 -11510 36990 -11390
rect 37110 -11510 37155 -11390
rect 37275 -11510 37330 -11390
rect 37450 -11510 37495 -11390
rect 37615 -11510 37660 -11390
rect 37780 -11510 37825 -11390
rect 37945 -11510 38000 -11390
rect 38120 -11510 38165 -11390
rect 38285 -11510 38330 -11390
rect 38450 -11510 38495 -11390
rect 38615 -11510 38670 -11390
rect 38790 -11510 38835 -11390
rect 38955 -11510 39000 -11390
rect 39120 -11510 39165 -11390
rect 39285 -11510 39340 -11390
rect 39460 -11510 39505 -11390
rect 39625 -11510 39670 -11390
rect 39790 -11510 39835 -11390
rect 39955 -11510 40010 -11390
rect 40130 -11510 40175 -11390
rect 40295 -11510 40340 -11390
rect 40460 -11510 40505 -11390
rect 40625 -11510 40680 -11390
rect 40800 -11510 40845 -11390
rect 40965 -11510 41010 -11390
rect 41130 -11510 41175 -11390
rect 41295 -11510 41350 -11390
rect 41470 -11510 41515 -11390
rect 41635 -11510 41680 -11390
rect 41800 -11510 41845 -11390
rect 41965 -11510 41975 -11390
rect 36475 -11555 41975 -11510
rect 36475 -11675 36485 -11555
rect 36605 -11675 36660 -11555
rect 36780 -11675 36825 -11555
rect 36945 -11675 36990 -11555
rect 37110 -11675 37155 -11555
rect 37275 -11675 37330 -11555
rect 37450 -11675 37495 -11555
rect 37615 -11675 37660 -11555
rect 37780 -11675 37825 -11555
rect 37945 -11675 38000 -11555
rect 38120 -11675 38165 -11555
rect 38285 -11675 38330 -11555
rect 38450 -11675 38495 -11555
rect 38615 -11675 38670 -11555
rect 38790 -11675 38835 -11555
rect 38955 -11675 39000 -11555
rect 39120 -11675 39165 -11555
rect 39285 -11675 39340 -11555
rect 39460 -11675 39505 -11555
rect 39625 -11675 39670 -11555
rect 39790 -11675 39835 -11555
rect 39955 -11675 40010 -11555
rect 40130 -11675 40175 -11555
rect 40295 -11675 40340 -11555
rect 40460 -11675 40505 -11555
rect 40625 -11675 40680 -11555
rect 40800 -11675 40845 -11555
rect 40965 -11675 41010 -11555
rect 41130 -11675 41175 -11555
rect 41295 -11675 41350 -11555
rect 41470 -11675 41515 -11555
rect 41635 -11675 41680 -11555
rect 41800 -11675 41845 -11555
rect 41965 -11675 41975 -11555
rect 36475 -11720 41975 -11675
rect 36475 -11840 36485 -11720
rect 36605 -11840 36660 -11720
rect 36780 -11840 36825 -11720
rect 36945 -11840 36990 -11720
rect 37110 -11840 37155 -11720
rect 37275 -11840 37330 -11720
rect 37450 -11840 37495 -11720
rect 37615 -11840 37660 -11720
rect 37780 -11840 37825 -11720
rect 37945 -11840 38000 -11720
rect 38120 -11840 38165 -11720
rect 38285 -11840 38330 -11720
rect 38450 -11840 38495 -11720
rect 38615 -11840 38670 -11720
rect 38790 -11840 38835 -11720
rect 38955 -11840 39000 -11720
rect 39120 -11840 39165 -11720
rect 39285 -11840 39340 -11720
rect 39460 -11840 39505 -11720
rect 39625 -11840 39670 -11720
rect 39790 -11840 39835 -11720
rect 39955 -11840 40010 -11720
rect 40130 -11840 40175 -11720
rect 40295 -11840 40340 -11720
rect 40460 -11840 40505 -11720
rect 40625 -11840 40680 -11720
rect 40800 -11840 40845 -11720
rect 40965 -11840 41010 -11720
rect 41130 -11840 41175 -11720
rect 41295 -11840 41350 -11720
rect 41470 -11840 41515 -11720
rect 41635 -11840 41680 -11720
rect 41800 -11840 41845 -11720
rect 41965 -11840 41975 -11720
rect 36475 -11885 41975 -11840
rect 36475 -12005 36485 -11885
rect 36605 -12005 36660 -11885
rect 36780 -12005 36825 -11885
rect 36945 -12005 36990 -11885
rect 37110 -12005 37155 -11885
rect 37275 -12005 37330 -11885
rect 37450 -12005 37495 -11885
rect 37615 -12005 37660 -11885
rect 37780 -12005 37825 -11885
rect 37945 -12005 38000 -11885
rect 38120 -12005 38165 -11885
rect 38285 -12005 38330 -11885
rect 38450 -12005 38495 -11885
rect 38615 -12005 38670 -11885
rect 38790 -12005 38835 -11885
rect 38955 -12005 39000 -11885
rect 39120 -12005 39165 -11885
rect 39285 -12005 39340 -11885
rect 39460 -12005 39505 -11885
rect 39625 -12005 39670 -11885
rect 39790 -12005 39835 -11885
rect 39955 -12005 40010 -11885
rect 40130 -12005 40175 -11885
rect 40295 -12005 40340 -11885
rect 40460 -12005 40505 -11885
rect 40625 -12005 40680 -11885
rect 40800 -12005 40845 -11885
rect 40965 -12005 41010 -11885
rect 41130 -12005 41175 -11885
rect 41295 -12005 41350 -11885
rect 41470 -12005 41515 -11885
rect 41635 -12005 41680 -11885
rect 41800 -12005 41845 -11885
rect 41965 -12005 41975 -11885
rect 36475 -12060 41975 -12005
rect 36475 -12180 36485 -12060
rect 36605 -12180 36660 -12060
rect 36780 -12180 36825 -12060
rect 36945 -12180 36990 -12060
rect 37110 -12180 37155 -12060
rect 37275 -12180 37330 -12060
rect 37450 -12180 37495 -12060
rect 37615 -12180 37660 -12060
rect 37780 -12180 37825 -12060
rect 37945 -12180 38000 -12060
rect 38120 -12180 38165 -12060
rect 38285 -12180 38330 -12060
rect 38450 -12180 38495 -12060
rect 38615 -12180 38670 -12060
rect 38790 -12180 38835 -12060
rect 38955 -12180 39000 -12060
rect 39120 -12180 39165 -12060
rect 39285 -12180 39340 -12060
rect 39460 -12180 39505 -12060
rect 39625 -12180 39670 -12060
rect 39790 -12180 39835 -12060
rect 39955 -12180 40010 -12060
rect 40130 -12180 40175 -12060
rect 40295 -12180 40340 -12060
rect 40460 -12180 40505 -12060
rect 40625 -12180 40680 -12060
rect 40800 -12180 40845 -12060
rect 40965 -12180 41010 -12060
rect 41130 -12180 41175 -12060
rect 41295 -12180 41350 -12060
rect 41470 -12180 41515 -12060
rect 41635 -12180 41680 -12060
rect 41800 -12180 41845 -12060
rect 41965 -12180 41975 -12060
rect 36475 -12225 41975 -12180
rect 36475 -12345 36485 -12225
rect 36605 -12345 36660 -12225
rect 36780 -12345 36825 -12225
rect 36945 -12345 36990 -12225
rect 37110 -12345 37155 -12225
rect 37275 -12345 37330 -12225
rect 37450 -12345 37495 -12225
rect 37615 -12345 37660 -12225
rect 37780 -12345 37825 -12225
rect 37945 -12345 38000 -12225
rect 38120 -12345 38165 -12225
rect 38285 -12345 38330 -12225
rect 38450 -12345 38495 -12225
rect 38615 -12345 38670 -12225
rect 38790 -12345 38835 -12225
rect 38955 -12345 39000 -12225
rect 39120 -12345 39165 -12225
rect 39285 -12345 39340 -12225
rect 39460 -12345 39505 -12225
rect 39625 -12345 39670 -12225
rect 39790 -12345 39835 -12225
rect 39955 -12345 40010 -12225
rect 40130 -12345 40175 -12225
rect 40295 -12345 40340 -12225
rect 40460 -12345 40505 -12225
rect 40625 -12345 40680 -12225
rect 40800 -12345 40845 -12225
rect 40965 -12345 41010 -12225
rect 41130 -12345 41175 -12225
rect 41295 -12345 41350 -12225
rect 41470 -12345 41515 -12225
rect 41635 -12345 41680 -12225
rect 41800 -12345 41845 -12225
rect 41965 -12345 41975 -12225
rect 36475 -12390 41975 -12345
rect 36475 -12510 36485 -12390
rect 36605 -12510 36660 -12390
rect 36780 -12510 36825 -12390
rect 36945 -12510 36990 -12390
rect 37110 -12510 37155 -12390
rect 37275 -12510 37330 -12390
rect 37450 -12510 37495 -12390
rect 37615 -12510 37660 -12390
rect 37780 -12510 37825 -12390
rect 37945 -12510 38000 -12390
rect 38120 -12510 38165 -12390
rect 38285 -12510 38330 -12390
rect 38450 -12510 38495 -12390
rect 38615 -12510 38670 -12390
rect 38790 -12510 38835 -12390
rect 38955 -12510 39000 -12390
rect 39120 -12510 39165 -12390
rect 39285 -12510 39340 -12390
rect 39460 -12510 39505 -12390
rect 39625 -12510 39670 -12390
rect 39790 -12510 39835 -12390
rect 39955 -12510 40010 -12390
rect 40130 -12510 40175 -12390
rect 40295 -12510 40340 -12390
rect 40460 -12510 40505 -12390
rect 40625 -12510 40680 -12390
rect 40800 -12510 40845 -12390
rect 40965 -12510 41010 -12390
rect 41130 -12510 41175 -12390
rect 41295 -12510 41350 -12390
rect 41470 -12510 41515 -12390
rect 41635 -12510 41680 -12390
rect 41800 -12510 41845 -12390
rect 41965 -12510 41975 -12390
rect 36475 -12555 41975 -12510
rect 36475 -12675 36485 -12555
rect 36605 -12675 36660 -12555
rect 36780 -12675 36825 -12555
rect 36945 -12675 36990 -12555
rect 37110 -12675 37155 -12555
rect 37275 -12675 37330 -12555
rect 37450 -12675 37495 -12555
rect 37615 -12675 37660 -12555
rect 37780 -12675 37825 -12555
rect 37945 -12675 38000 -12555
rect 38120 -12675 38165 -12555
rect 38285 -12675 38330 -12555
rect 38450 -12675 38495 -12555
rect 38615 -12675 38670 -12555
rect 38790 -12675 38835 -12555
rect 38955 -12675 39000 -12555
rect 39120 -12675 39165 -12555
rect 39285 -12675 39340 -12555
rect 39460 -12675 39505 -12555
rect 39625 -12675 39670 -12555
rect 39790 -12675 39835 -12555
rect 39955 -12675 40010 -12555
rect 40130 -12675 40175 -12555
rect 40295 -12675 40340 -12555
rect 40460 -12675 40505 -12555
rect 40625 -12675 40680 -12555
rect 40800 -12675 40845 -12555
rect 40965 -12675 41010 -12555
rect 41130 -12675 41175 -12555
rect 41295 -12675 41350 -12555
rect 41470 -12675 41515 -12555
rect 41635 -12675 41680 -12555
rect 41800 -12675 41845 -12555
rect 41965 -12675 41975 -12555
rect 36475 -12730 41975 -12675
rect 36475 -12850 36485 -12730
rect 36605 -12850 36660 -12730
rect 36780 -12850 36825 -12730
rect 36945 -12850 36990 -12730
rect 37110 -12850 37155 -12730
rect 37275 -12850 37330 -12730
rect 37450 -12850 37495 -12730
rect 37615 -12850 37660 -12730
rect 37780 -12850 37825 -12730
rect 37945 -12850 38000 -12730
rect 38120 -12850 38165 -12730
rect 38285 -12850 38330 -12730
rect 38450 -12850 38495 -12730
rect 38615 -12850 38670 -12730
rect 38790 -12850 38835 -12730
rect 38955 -12850 39000 -12730
rect 39120 -12850 39165 -12730
rect 39285 -12850 39340 -12730
rect 39460 -12850 39505 -12730
rect 39625 -12850 39670 -12730
rect 39790 -12850 39835 -12730
rect 39955 -12850 40010 -12730
rect 40130 -12850 40175 -12730
rect 40295 -12850 40340 -12730
rect 40460 -12850 40505 -12730
rect 40625 -12850 40680 -12730
rect 40800 -12850 40845 -12730
rect 40965 -12850 41010 -12730
rect 41130 -12850 41175 -12730
rect 41295 -12850 41350 -12730
rect 41470 -12850 41515 -12730
rect 41635 -12850 41680 -12730
rect 41800 -12850 41845 -12730
rect 41965 -12850 41975 -12730
rect 36475 -12895 41975 -12850
rect 36475 -13015 36485 -12895
rect 36605 -13015 36660 -12895
rect 36780 -13015 36825 -12895
rect 36945 -13015 36990 -12895
rect 37110 -13015 37155 -12895
rect 37275 -13015 37330 -12895
rect 37450 -13015 37495 -12895
rect 37615 -13015 37660 -12895
rect 37780 -13015 37825 -12895
rect 37945 -13015 38000 -12895
rect 38120 -13015 38165 -12895
rect 38285 -13015 38330 -12895
rect 38450 -13015 38495 -12895
rect 38615 -13015 38670 -12895
rect 38790 -13015 38835 -12895
rect 38955 -13015 39000 -12895
rect 39120 -13015 39165 -12895
rect 39285 -13015 39340 -12895
rect 39460 -13015 39505 -12895
rect 39625 -13015 39670 -12895
rect 39790 -13015 39835 -12895
rect 39955 -13015 40010 -12895
rect 40130 -13015 40175 -12895
rect 40295 -13015 40340 -12895
rect 40460 -13015 40505 -12895
rect 40625 -13015 40680 -12895
rect 40800 -13015 40845 -12895
rect 40965 -13015 41010 -12895
rect 41130 -13015 41175 -12895
rect 41295 -13015 41350 -12895
rect 41470 -13015 41515 -12895
rect 41635 -13015 41680 -12895
rect 41800 -13015 41845 -12895
rect 41965 -13015 41975 -12895
rect 36475 -13060 41975 -13015
rect 36475 -13180 36485 -13060
rect 36605 -13180 36660 -13060
rect 36780 -13180 36825 -13060
rect 36945 -13180 36990 -13060
rect 37110 -13180 37155 -13060
rect 37275 -13180 37330 -13060
rect 37450 -13180 37495 -13060
rect 37615 -13180 37660 -13060
rect 37780 -13180 37825 -13060
rect 37945 -13180 38000 -13060
rect 38120 -13180 38165 -13060
rect 38285 -13180 38330 -13060
rect 38450 -13180 38495 -13060
rect 38615 -13180 38670 -13060
rect 38790 -13180 38835 -13060
rect 38955 -13180 39000 -13060
rect 39120 -13180 39165 -13060
rect 39285 -13180 39340 -13060
rect 39460 -13180 39505 -13060
rect 39625 -13180 39670 -13060
rect 39790 -13180 39835 -13060
rect 39955 -13180 40010 -13060
rect 40130 -13180 40175 -13060
rect 40295 -13180 40340 -13060
rect 40460 -13180 40505 -13060
rect 40625 -13180 40680 -13060
rect 40800 -13180 40845 -13060
rect 40965 -13180 41010 -13060
rect 41130 -13180 41175 -13060
rect 41295 -13180 41350 -13060
rect 41470 -13180 41515 -13060
rect 41635 -13180 41680 -13060
rect 41800 -13180 41845 -13060
rect 41965 -13180 41975 -13060
rect 36475 -13225 41975 -13180
rect 36475 -13345 36485 -13225
rect 36605 -13345 36660 -13225
rect 36780 -13345 36825 -13225
rect 36945 -13345 36990 -13225
rect 37110 -13345 37155 -13225
rect 37275 -13345 37330 -13225
rect 37450 -13345 37495 -13225
rect 37615 -13345 37660 -13225
rect 37780 -13345 37825 -13225
rect 37945 -13345 38000 -13225
rect 38120 -13345 38165 -13225
rect 38285 -13345 38330 -13225
rect 38450 -13345 38495 -13225
rect 38615 -13345 38670 -13225
rect 38790 -13345 38835 -13225
rect 38955 -13345 39000 -13225
rect 39120 -13345 39165 -13225
rect 39285 -13345 39340 -13225
rect 39460 -13345 39505 -13225
rect 39625 -13345 39670 -13225
rect 39790 -13345 39835 -13225
rect 39955 -13345 40010 -13225
rect 40130 -13345 40175 -13225
rect 40295 -13345 40340 -13225
rect 40460 -13345 40505 -13225
rect 40625 -13345 40680 -13225
rect 40800 -13345 40845 -13225
rect 40965 -13345 41010 -13225
rect 41130 -13345 41175 -13225
rect 41295 -13345 41350 -13225
rect 41470 -13345 41515 -13225
rect 41635 -13345 41680 -13225
rect 41800 -13345 41845 -13225
rect 41965 -13345 41975 -13225
rect 36475 -13400 41975 -13345
rect 36475 -13520 36485 -13400
rect 36605 -13520 36660 -13400
rect 36780 -13520 36825 -13400
rect 36945 -13520 36990 -13400
rect 37110 -13520 37155 -13400
rect 37275 -13520 37330 -13400
rect 37450 -13520 37495 -13400
rect 37615 -13520 37660 -13400
rect 37780 -13520 37825 -13400
rect 37945 -13520 38000 -13400
rect 38120 -13520 38165 -13400
rect 38285 -13520 38330 -13400
rect 38450 -13520 38495 -13400
rect 38615 -13520 38670 -13400
rect 38790 -13520 38835 -13400
rect 38955 -13520 39000 -13400
rect 39120 -13520 39165 -13400
rect 39285 -13520 39340 -13400
rect 39460 -13520 39505 -13400
rect 39625 -13520 39670 -13400
rect 39790 -13520 39835 -13400
rect 39955 -13520 40010 -13400
rect 40130 -13520 40175 -13400
rect 40295 -13520 40340 -13400
rect 40460 -13520 40505 -13400
rect 40625 -13520 40680 -13400
rect 40800 -13520 40845 -13400
rect 40965 -13520 41010 -13400
rect 41130 -13520 41175 -13400
rect 41295 -13520 41350 -13400
rect 41470 -13520 41515 -13400
rect 41635 -13520 41680 -13400
rect 41800 -13520 41845 -13400
rect 41965 -13520 41975 -13400
rect 36475 -13565 41975 -13520
rect 36475 -13685 36485 -13565
rect 36605 -13685 36660 -13565
rect 36780 -13685 36825 -13565
rect 36945 -13685 36990 -13565
rect 37110 -13685 37155 -13565
rect 37275 -13685 37330 -13565
rect 37450 -13685 37495 -13565
rect 37615 -13685 37660 -13565
rect 37780 -13685 37825 -13565
rect 37945 -13685 38000 -13565
rect 38120 -13685 38165 -13565
rect 38285 -13685 38330 -13565
rect 38450 -13685 38495 -13565
rect 38615 -13685 38670 -13565
rect 38790 -13685 38835 -13565
rect 38955 -13685 39000 -13565
rect 39120 -13685 39165 -13565
rect 39285 -13685 39340 -13565
rect 39460 -13685 39505 -13565
rect 39625 -13685 39670 -13565
rect 39790 -13685 39835 -13565
rect 39955 -13685 40010 -13565
rect 40130 -13685 40175 -13565
rect 40295 -13685 40340 -13565
rect 40460 -13685 40505 -13565
rect 40625 -13685 40680 -13565
rect 40800 -13685 40845 -13565
rect 40965 -13685 41010 -13565
rect 41130 -13685 41175 -13565
rect 41295 -13685 41350 -13565
rect 41470 -13685 41515 -13565
rect 41635 -13685 41680 -13565
rect 41800 -13685 41845 -13565
rect 41965 -13685 41975 -13565
rect 36475 -13730 41975 -13685
rect 36475 -13850 36485 -13730
rect 36605 -13850 36660 -13730
rect 36780 -13850 36825 -13730
rect 36945 -13850 36990 -13730
rect 37110 -13850 37155 -13730
rect 37275 -13850 37330 -13730
rect 37450 -13850 37495 -13730
rect 37615 -13850 37660 -13730
rect 37780 -13850 37825 -13730
rect 37945 -13850 38000 -13730
rect 38120 -13850 38165 -13730
rect 38285 -13850 38330 -13730
rect 38450 -13850 38495 -13730
rect 38615 -13850 38670 -13730
rect 38790 -13850 38835 -13730
rect 38955 -13850 39000 -13730
rect 39120 -13850 39165 -13730
rect 39285 -13850 39340 -13730
rect 39460 -13850 39505 -13730
rect 39625 -13850 39670 -13730
rect 39790 -13850 39835 -13730
rect 39955 -13850 40010 -13730
rect 40130 -13850 40175 -13730
rect 40295 -13850 40340 -13730
rect 40460 -13850 40505 -13730
rect 40625 -13850 40680 -13730
rect 40800 -13850 40845 -13730
rect 40965 -13850 41010 -13730
rect 41130 -13850 41175 -13730
rect 41295 -13850 41350 -13730
rect 41470 -13850 41515 -13730
rect 41635 -13850 41680 -13730
rect 41800 -13850 41845 -13730
rect 41965 -13850 41975 -13730
rect 36475 -13895 41975 -13850
rect 36475 -14015 36485 -13895
rect 36605 -14015 36660 -13895
rect 36780 -14015 36825 -13895
rect 36945 -14015 36990 -13895
rect 37110 -14015 37155 -13895
rect 37275 -14015 37330 -13895
rect 37450 -14015 37495 -13895
rect 37615 -14015 37660 -13895
rect 37780 -14015 37825 -13895
rect 37945 -14015 38000 -13895
rect 38120 -14015 38165 -13895
rect 38285 -14015 38330 -13895
rect 38450 -14015 38495 -13895
rect 38615 -14015 38670 -13895
rect 38790 -14015 38835 -13895
rect 38955 -14015 39000 -13895
rect 39120 -14015 39165 -13895
rect 39285 -14015 39340 -13895
rect 39460 -14015 39505 -13895
rect 39625 -14015 39670 -13895
rect 39790 -14015 39835 -13895
rect 39955 -14015 40010 -13895
rect 40130 -14015 40175 -13895
rect 40295 -14015 40340 -13895
rect 40460 -14015 40505 -13895
rect 40625 -14015 40680 -13895
rect 40800 -14015 40845 -13895
rect 40965 -14015 41010 -13895
rect 41130 -14015 41175 -13895
rect 41295 -14015 41350 -13895
rect 41470 -14015 41515 -13895
rect 41635 -14015 41680 -13895
rect 41800 -14015 41845 -13895
rect 41965 -14015 41975 -13895
rect 36475 -14070 41975 -14015
rect 36475 -14190 36485 -14070
rect 36605 -14190 36660 -14070
rect 36780 -14190 36825 -14070
rect 36945 -14190 36990 -14070
rect 37110 -14190 37155 -14070
rect 37275 -14190 37330 -14070
rect 37450 -14190 37495 -14070
rect 37615 -14190 37660 -14070
rect 37780 -14190 37825 -14070
rect 37945 -14190 38000 -14070
rect 38120 -14190 38165 -14070
rect 38285 -14190 38330 -14070
rect 38450 -14190 38495 -14070
rect 38615 -14190 38670 -14070
rect 38790 -14190 38835 -14070
rect 38955 -14190 39000 -14070
rect 39120 -14190 39165 -14070
rect 39285 -14190 39340 -14070
rect 39460 -14190 39505 -14070
rect 39625 -14190 39670 -14070
rect 39790 -14190 39835 -14070
rect 39955 -14190 40010 -14070
rect 40130 -14190 40175 -14070
rect 40295 -14190 40340 -14070
rect 40460 -14190 40505 -14070
rect 40625 -14190 40680 -14070
rect 40800 -14190 40845 -14070
rect 40965 -14190 41010 -14070
rect 41130 -14190 41175 -14070
rect 41295 -14190 41350 -14070
rect 41470 -14190 41515 -14070
rect 41635 -14190 41680 -14070
rect 41800 -14190 41845 -14070
rect 41965 -14190 41975 -14070
rect 36475 -14235 41975 -14190
rect 36475 -14355 36485 -14235
rect 36605 -14355 36660 -14235
rect 36780 -14355 36825 -14235
rect 36945 -14355 36990 -14235
rect 37110 -14355 37155 -14235
rect 37275 -14355 37330 -14235
rect 37450 -14355 37495 -14235
rect 37615 -14355 37660 -14235
rect 37780 -14355 37825 -14235
rect 37945 -14355 38000 -14235
rect 38120 -14355 38165 -14235
rect 38285 -14355 38330 -14235
rect 38450 -14355 38495 -14235
rect 38615 -14355 38670 -14235
rect 38790 -14355 38835 -14235
rect 38955 -14355 39000 -14235
rect 39120 -14355 39165 -14235
rect 39285 -14355 39340 -14235
rect 39460 -14355 39505 -14235
rect 39625 -14355 39670 -14235
rect 39790 -14355 39835 -14235
rect 39955 -14355 40010 -14235
rect 40130 -14355 40175 -14235
rect 40295 -14355 40340 -14235
rect 40460 -14355 40505 -14235
rect 40625 -14355 40680 -14235
rect 40800 -14355 40845 -14235
rect 40965 -14355 41010 -14235
rect 41130 -14355 41175 -14235
rect 41295 -14355 41350 -14235
rect 41470 -14355 41515 -14235
rect 41635 -14355 41680 -14235
rect 41800 -14355 41845 -14235
rect 41965 -14355 41975 -14235
rect 36475 -14400 41975 -14355
rect 36475 -14520 36485 -14400
rect 36605 -14520 36660 -14400
rect 36780 -14520 36825 -14400
rect 36945 -14520 36990 -14400
rect 37110 -14520 37155 -14400
rect 37275 -14520 37330 -14400
rect 37450 -14520 37495 -14400
rect 37615 -14520 37660 -14400
rect 37780 -14520 37825 -14400
rect 37945 -14520 38000 -14400
rect 38120 -14520 38165 -14400
rect 38285 -14520 38330 -14400
rect 38450 -14520 38495 -14400
rect 38615 -14520 38670 -14400
rect 38790 -14520 38835 -14400
rect 38955 -14520 39000 -14400
rect 39120 -14520 39165 -14400
rect 39285 -14520 39340 -14400
rect 39460 -14520 39505 -14400
rect 39625 -14520 39670 -14400
rect 39790 -14520 39835 -14400
rect 39955 -14520 40010 -14400
rect 40130 -14520 40175 -14400
rect 40295 -14520 40340 -14400
rect 40460 -14520 40505 -14400
rect 40625 -14520 40680 -14400
rect 40800 -14520 40845 -14400
rect 40965 -14520 41010 -14400
rect 41130 -14520 41175 -14400
rect 41295 -14520 41350 -14400
rect 41470 -14520 41515 -14400
rect 41635 -14520 41680 -14400
rect 41800 -14520 41845 -14400
rect 41965 -14520 41975 -14400
rect 36475 -14565 41975 -14520
rect 36475 -14685 36485 -14565
rect 36605 -14685 36660 -14565
rect 36780 -14685 36825 -14565
rect 36945 -14685 36990 -14565
rect 37110 -14685 37155 -14565
rect 37275 -14685 37330 -14565
rect 37450 -14685 37495 -14565
rect 37615 -14685 37660 -14565
rect 37780 -14685 37825 -14565
rect 37945 -14685 38000 -14565
rect 38120 -14685 38165 -14565
rect 38285 -14685 38330 -14565
rect 38450 -14685 38495 -14565
rect 38615 -14685 38670 -14565
rect 38790 -14685 38835 -14565
rect 38955 -14685 39000 -14565
rect 39120 -14685 39165 -14565
rect 39285 -14685 39340 -14565
rect 39460 -14685 39505 -14565
rect 39625 -14685 39670 -14565
rect 39790 -14685 39835 -14565
rect 39955 -14685 40010 -14565
rect 40130 -14685 40175 -14565
rect 40295 -14685 40340 -14565
rect 40460 -14685 40505 -14565
rect 40625 -14685 40680 -14565
rect 40800 -14685 40845 -14565
rect 40965 -14685 41010 -14565
rect 41130 -14685 41175 -14565
rect 41295 -14685 41350 -14565
rect 41470 -14685 41515 -14565
rect 41635 -14685 41680 -14565
rect 41800 -14685 41845 -14565
rect 41965 -14685 41975 -14565
rect 36475 -14740 41975 -14685
rect 36475 -14860 36485 -14740
rect 36605 -14860 36660 -14740
rect 36780 -14860 36825 -14740
rect 36945 -14860 36990 -14740
rect 37110 -14860 37155 -14740
rect 37275 -14860 37330 -14740
rect 37450 -14860 37495 -14740
rect 37615 -14860 37660 -14740
rect 37780 -14860 37825 -14740
rect 37945 -14860 38000 -14740
rect 38120 -14860 38165 -14740
rect 38285 -14860 38330 -14740
rect 38450 -14860 38495 -14740
rect 38615 -14860 38670 -14740
rect 38790 -14860 38835 -14740
rect 38955 -14860 39000 -14740
rect 39120 -14860 39165 -14740
rect 39285 -14860 39340 -14740
rect 39460 -14860 39505 -14740
rect 39625 -14860 39670 -14740
rect 39790 -14860 39835 -14740
rect 39955 -14860 40010 -14740
rect 40130 -14860 40175 -14740
rect 40295 -14860 40340 -14740
rect 40460 -14860 40505 -14740
rect 40625 -14860 40680 -14740
rect 40800 -14860 40845 -14740
rect 40965 -14860 41010 -14740
rect 41130 -14860 41175 -14740
rect 41295 -14860 41350 -14740
rect 41470 -14860 41515 -14740
rect 41635 -14860 41680 -14740
rect 41800 -14860 41845 -14740
rect 41965 -14860 41975 -14740
rect 36475 -14905 41975 -14860
rect 36475 -15025 36485 -14905
rect 36605 -15025 36660 -14905
rect 36780 -15025 36825 -14905
rect 36945 -15025 36990 -14905
rect 37110 -15025 37155 -14905
rect 37275 -15025 37330 -14905
rect 37450 -15025 37495 -14905
rect 37615 -15025 37660 -14905
rect 37780 -15025 37825 -14905
rect 37945 -15025 38000 -14905
rect 38120 -15025 38165 -14905
rect 38285 -15025 38330 -14905
rect 38450 -15025 38495 -14905
rect 38615 -15025 38670 -14905
rect 38790 -15025 38835 -14905
rect 38955 -15025 39000 -14905
rect 39120 -15025 39165 -14905
rect 39285 -15025 39340 -14905
rect 39460 -15025 39505 -14905
rect 39625 -15025 39670 -14905
rect 39790 -15025 39835 -14905
rect 39955 -15025 40010 -14905
rect 40130 -15025 40175 -14905
rect 40295 -15025 40340 -14905
rect 40460 -15025 40505 -14905
rect 40625 -15025 40680 -14905
rect 40800 -15025 40845 -14905
rect 40965 -15025 41010 -14905
rect 41130 -15025 41175 -14905
rect 41295 -15025 41350 -14905
rect 41470 -15025 41515 -14905
rect 41635 -15025 41680 -14905
rect 41800 -15025 41845 -14905
rect 41965 -15025 41975 -14905
rect 36475 -15070 41975 -15025
rect 36475 -15190 36485 -15070
rect 36605 -15190 36660 -15070
rect 36780 -15190 36825 -15070
rect 36945 -15190 36990 -15070
rect 37110 -15190 37155 -15070
rect 37275 -15190 37330 -15070
rect 37450 -15190 37495 -15070
rect 37615 -15190 37660 -15070
rect 37780 -15190 37825 -15070
rect 37945 -15190 38000 -15070
rect 38120 -15190 38165 -15070
rect 38285 -15190 38330 -15070
rect 38450 -15190 38495 -15070
rect 38615 -15190 38670 -15070
rect 38790 -15190 38835 -15070
rect 38955 -15190 39000 -15070
rect 39120 -15190 39165 -15070
rect 39285 -15190 39340 -15070
rect 39460 -15190 39505 -15070
rect 39625 -15190 39670 -15070
rect 39790 -15190 39835 -15070
rect 39955 -15190 40010 -15070
rect 40130 -15190 40175 -15070
rect 40295 -15190 40340 -15070
rect 40460 -15190 40505 -15070
rect 40625 -15190 40680 -15070
rect 40800 -15190 40845 -15070
rect 40965 -15190 41010 -15070
rect 41130 -15190 41175 -15070
rect 41295 -15190 41350 -15070
rect 41470 -15190 41515 -15070
rect 41635 -15190 41680 -15070
rect 41800 -15190 41845 -15070
rect 41965 -15190 41975 -15070
rect 36475 -15235 41975 -15190
rect 36475 -15355 36485 -15235
rect 36605 -15355 36660 -15235
rect 36780 -15355 36825 -15235
rect 36945 -15355 36990 -15235
rect 37110 -15355 37155 -15235
rect 37275 -15355 37330 -15235
rect 37450 -15355 37495 -15235
rect 37615 -15355 37660 -15235
rect 37780 -15355 37825 -15235
rect 37945 -15355 38000 -15235
rect 38120 -15355 38165 -15235
rect 38285 -15355 38330 -15235
rect 38450 -15355 38495 -15235
rect 38615 -15355 38670 -15235
rect 38790 -15355 38835 -15235
rect 38955 -15355 39000 -15235
rect 39120 -15355 39165 -15235
rect 39285 -15355 39340 -15235
rect 39460 -15355 39505 -15235
rect 39625 -15355 39670 -15235
rect 39790 -15355 39835 -15235
rect 39955 -15355 40010 -15235
rect 40130 -15355 40175 -15235
rect 40295 -15355 40340 -15235
rect 40460 -15355 40505 -15235
rect 40625 -15355 40680 -15235
rect 40800 -15355 40845 -15235
rect 40965 -15355 41010 -15235
rect 41130 -15355 41175 -15235
rect 41295 -15355 41350 -15235
rect 41470 -15355 41515 -15235
rect 41635 -15355 41680 -15235
rect 41800 -15355 41845 -15235
rect 41965 -15355 41975 -15235
rect 36475 -15410 41975 -15355
rect 36475 -15530 36485 -15410
rect 36605 -15530 36660 -15410
rect 36780 -15530 36825 -15410
rect 36945 -15530 36990 -15410
rect 37110 -15530 37155 -15410
rect 37275 -15530 37330 -15410
rect 37450 -15530 37495 -15410
rect 37615 -15530 37660 -15410
rect 37780 -15530 37825 -15410
rect 37945 -15530 38000 -15410
rect 38120 -15530 38165 -15410
rect 38285 -15530 38330 -15410
rect 38450 -15530 38495 -15410
rect 38615 -15530 38670 -15410
rect 38790 -15530 38835 -15410
rect 38955 -15530 39000 -15410
rect 39120 -15530 39165 -15410
rect 39285 -15530 39340 -15410
rect 39460 -15530 39505 -15410
rect 39625 -15530 39670 -15410
rect 39790 -15530 39835 -15410
rect 39955 -15530 40010 -15410
rect 40130 -15530 40175 -15410
rect 40295 -15530 40340 -15410
rect 40460 -15530 40505 -15410
rect 40625 -15530 40680 -15410
rect 40800 -15530 40845 -15410
rect 40965 -15530 41010 -15410
rect 41130 -15530 41175 -15410
rect 41295 -15530 41350 -15410
rect 41470 -15530 41515 -15410
rect 41635 -15530 41680 -15410
rect 41800 -15530 41845 -15410
rect 41965 -15530 41975 -15410
rect 36475 -15540 41975 -15530
rect 42165 -10050 47665 -10040
rect 42165 -10170 42175 -10050
rect 42295 -10170 42350 -10050
rect 42470 -10170 42515 -10050
rect 42635 -10170 42680 -10050
rect 42800 -10170 42845 -10050
rect 42965 -10170 43020 -10050
rect 43140 -10170 43185 -10050
rect 43305 -10170 43350 -10050
rect 43470 -10170 43515 -10050
rect 43635 -10170 43690 -10050
rect 43810 -10170 43855 -10050
rect 43975 -10170 44020 -10050
rect 44140 -10170 44185 -10050
rect 44305 -10170 44360 -10050
rect 44480 -10170 44525 -10050
rect 44645 -10170 44690 -10050
rect 44810 -10170 44855 -10050
rect 44975 -10170 45030 -10050
rect 45150 -10170 45195 -10050
rect 45315 -10170 45360 -10050
rect 45480 -10170 45525 -10050
rect 45645 -10170 45700 -10050
rect 45820 -10170 45865 -10050
rect 45985 -10170 46030 -10050
rect 46150 -10170 46195 -10050
rect 46315 -10170 46370 -10050
rect 46490 -10170 46535 -10050
rect 46655 -10170 46700 -10050
rect 46820 -10170 46865 -10050
rect 46985 -10170 47040 -10050
rect 47160 -10170 47205 -10050
rect 47325 -10170 47370 -10050
rect 47490 -10170 47535 -10050
rect 47655 -10170 47665 -10050
rect 42165 -10215 47665 -10170
rect 42165 -10335 42175 -10215
rect 42295 -10335 42350 -10215
rect 42470 -10335 42515 -10215
rect 42635 -10335 42680 -10215
rect 42800 -10335 42845 -10215
rect 42965 -10335 43020 -10215
rect 43140 -10335 43185 -10215
rect 43305 -10335 43350 -10215
rect 43470 -10335 43515 -10215
rect 43635 -10335 43690 -10215
rect 43810 -10335 43855 -10215
rect 43975 -10335 44020 -10215
rect 44140 -10335 44185 -10215
rect 44305 -10335 44360 -10215
rect 44480 -10335 44525 -10215
rect 44645 -10335 44690 -10215
rect 44810 -10335 44855 -10215
rect 44975 -10335 45030 -10215
rect 45150 -10335 45195 -10215
rect 45315 -10335 45360 -10215
rect 45480 -10335 45525 -10215
rect 45645 -10335 45700 -10215
rect 45820 -10335 45865 -10215
rect 45985 -10335 46030 -10215
rect 46150 -10335 46195 -10215
rect 46315 -10335 46370 -10215
rect 46490 -10335 46535 -10215
rect 46655 -10335 46700 -10215
rect 46820 -10335 46865 -10215
rect 46985 -10335 47040 -10215
rect 47160 -10335 47205 -10215
rect 47325 -10335 47370 -10215
rect 47490 -10335 47535 -10215
rect 47655 -10335 47665 -10215
rect 42165 -10380 47665 -10335
rect 42165 -10500 42175 -10380
rect 42295 -10500 42350 -10380
rect 42470 -10500 42515 -10380
rect 42635 -10500 42680 -10380
rect 42800 -10500 42845 -10380
rect 42965 -10500 43020 -10380
rect 43140 -10500 43185 -10380
rect 43305 -10500 43350 -10380
rect 43470 -10500 43515 -10380
rect 43635 -10500 43690 -10380
rect 43810 -10500 43855 -10380
rect 43975 -10500 44020 -10380
rect 44140 -10500 44185 -10380
rect 44305 -10500 44360 -10380
rect 44480 -10500 44525 -10380
rect 44645 -10500 44690 -10380
rect 44810 -10500 44855 -10380
rect 44975 -10500 45030 -10380
rect 45150 -10500 45195 -10380
rect 45315 -10500 45360 -10380
rect 45480 -10500 45525 -10380
rect 45645 -10500 45700 -10380
rect 45820 -10500 45865 -10380
rect 45985 -10500 46030 -10380
rect 46150 -10500 46195 -10380
rect 46315 -10500 46370 -10380
rect 46490 -10500 46535 -10380
rect 46655 -10500 46700 -10380
rect 46820 -10500 46865 -10380
rect 46985 -10500 47040 -10380
rect 47160 -10500 47205 -10380
rect 47325 -10500 47370 -10380
rect 47490 -10500 47535 -10380
rect 47655 -10500 47665 -10380
rect 42165 -10545 47665 -10500
rect 42165 -10665 42175 -10545
rect 42295 -10665 42350 -10545
rect 42470 -10665 42515 -10545
rect 42635 -10665 42680 -10545
rect 42800 -10665 42845 -10545
rect 42965 -10665 43020 -10545
rect 43140 -10665 43185 -10545
rect 43305 -10665 43350 -10545
rect 43470 -10665 43515 -10545
rect 43635 -10665 43690 -10545
rect 43810 -10665 43855 -10545
rect 43975 -10665 44020 -10545
rect 44140 -10665 44185 -10545
rect 44305 -10665 44360 -10545
rect 44480 -10665 44525 -10545
rect 44645 -10665 44690 -10545
rect 44810 -10665 44855 -10545
rect 44975 -10665 45030 -10545
rect 45150 -10665 45195 -10545
rect 45315 -10665 45360 -10545
rect 45480 -10665 45525 -10545
rect 45645 -10665 45700 -10545
rect 45820 -10665 45865 -10545
rect 45985 -10665 46030 -10545
rect 46150 -10665 46195 -10545
rect 46315 -10665 46370 -10545
rect 46490 -10665 46535 -10545
rect 46655 -10665 46700 -10545
rect 46820 -10665 46865 -10545
rect 46985 -10665 47040 -10545
rect 47160 -10665 47205 -10545
rect 47325 -10665 47370 -10545
rect 47490 -10665 47535 -10545
rect 47655 -10665 47665 -10545
rect 42165 -10720 47665 -10665
rect 42165 -10840 42175 -10720
rect 42295 -10840 42350 -10720
rect 42470 -10840 42515 -10720
rect 42635 -10840 42680 -10720
rect 42800 -10840 42845 -10720
rect 42965 -10840 43020 -10720
rect 43140 -10840 43185 -10720
rect 43305 -10840 43350 -10720
rect 43470 -10840 43515 -10720
rect 43635 -10840 43690 -10720
rect 43810 -10840 43855 -10720
rect 43975 -10840 44020 -10720
rect 44140 -10840 44185 -10720
rect 44305 -10840 44360 -10720
rect 44480 -10840 44525 -10720
rect 44645 -10840 44690 -10720
rect 44810 -10840 44855 -10720
rect 44975 -10840 45030 -10720
rect 45150 -10840 45195 -10720
rect 45315 -10840 45360 -10720
rect 45480 -10840 45525 -10720
rect 45645 -10840 45700 -10720
rect 45820 -10840 45865 -10720
rect 45985 -10840 46030 -10720
rect 46150 -10840 46195 -10720
rect 46315 -10840 46370 -10720
rect 46490 -10840 46535 -10720
rect 46655 -10840 46700 -10720
rect 46820 -10840 46865 -10720
rect 46985 -10840 47040 -10720
rect 47160 -10840 47205 -10720
rect 47325 -10840 47370 -10720
rect 47490 -10840 47535 -10720
rect 47655 -10840 47665 -10720
rect 42165 -10885 47665 -10840
rect 42165 -11005 42175 -10885
rect 42295 -11005 42350 -10885
rect 42470 -11005 42515 -10885
rect 42635 -11005 42680 -10885
rect 42800 -11005 42845 -10885
rect 42965 -11005 43020 -10885
rect 43140 -11005 43185 -10885
rect 43305 -11005 43350 -10885
rect 43470 -11005 43515 -10885
rect 43635 -11005 43690 -10885
rect 43810 -11005 43855 -10885
rect 43975 -11005 44020 -10885
rect 44140 -11005 44185 -10885
rect 44305 -11005 44360 -10885
rect 44480 -11005 44525 -10885
rect 44645 -11005 44690 -10885
rect 44810 -11005 44855 -10885
rect 44975 -11005 45030 -10885
rect 45150 -11005 45195 -10885
rect 45315 -11005 45360 -10885
rect 45480 -11005 45525 -10885
rect 45645 -11005 45700 -10885
rect 45820 -11005 45865 -10885
rect 45985 -11005 46030 -10885
rect 46150 -11005 46195 -10885
rect 46315 -11005 46370 -10885
rect 46490 -11005 46535 -10885
rect 46655 -11005 46700 -10885
rect 46820 -11005 46865 -10885
rect 46985 -11005 47040 -10885
rect 47160 -11005 47205 -10885
rect 47325 -11005 47370 -10885
rect 47490 -11005 47535 -10885
rect 47655 -11005 47665 -10885
rect 42165 -11050 47665 -11005
rect 42165 -11170 42175 -11050
rect 42295 -11170 42350 -11050
rect 42470 -11170 42515 -11050
rect 42635 -11170 42680 -11050
rect 42800 -11170 42845 -11050
rect 42965 -11170 43020 -11050
rect 43140 -11170 43185 -11050
rect 43305 -11170 43350 -11050
rect 43470 -11170 43515 -11050
rect 43635 -11170 43690 -11050
rect 43810 -11170 43855 -11050
rect 43975 -11170 44020 -11050
rect 44140 -11170 44185 -11050
rect 44305 -11170 44360 -11050
rect 44480 -11170 44525 -11050
rect 44645 -11170 44690 -11050
rect 44810 -11170 44855 -11050
rect 44975 -11170 45030 -11050
rect 45150 -11170 45195 -11050
rect 45315 -11170 45360 -11050
rect 45480 -11170 45525 -11050
rect 45645 -11170 45700 -11050
rect 45820 -11170 45865 -11050
rect 45985 -11170 46030 -11050
rect 46150 -11170 46195 -11050
rect 46315 -11170 46370 -11050
rect 46490 -11170 46535 -11050
rect 46655 -11170 46700 -11050
rect 46820 -11170 46865 -11050
rect 46985 -11170 47040 -11050
rect 47160 -11170 47205 -11050
rect 47325 -11170 47370 -11050
rect 47490 -11170 47535 -11050
rect 47655 -11170 47665 -11050
rect 42165 -11215 47665 -11170
rect 42165 -11335 42175 -11215
rect 42295 -11335 42350 -11215
rect 42470 -11335 42515 -11215
rect 42635 -11335 42680 -11215
rect 42800 -11335 42845 -11215
rect 42965 -11335 43020 -11215
rect 43140 -11335 43185 -11215
rect 43305 -11335 43350 -11215
rect 43470 -11335 43515 -11215
rect 43635 -11335 43690 -11215
rect 43810 -11335 43855 -11215
rect 43975 -11335 44020 -11215
rect 44140 -11335 44185 -11215
rect 44305 -11335 44360 -11215
rect 44480 -11335 44525 -11215
rect 44645 -11335 44690 -11215
rect 44810 -11335 44855 -11215
rect 44975 -11335 45030 -11215
rect 45150 -11335 45195 -11215
rect 45315 -11335 45360 -11215
rect 45480 -11335 45525 -11215
rect 45645 -11335 45700 -11215
rect 45820 -11335 45865 -11215
rect 45985 -11335 46030 -11215
rect 46150 -11335 46195 -11215
rect 46315 -11335 46370 -11215
rect 46490 -11335 46535 -11215
rect 46655 -11335 46700 -11215
rect 46820 -11335 46865 -11215
rect 46985 -11335 47040 -11215
rect 47160 -11335 47205 -11215
rect 47325 -11335 47370 -11215
rect 47490 -11335 47535 -11215
rect 47655 -11335 47665 -11215
rect 42165 -11390 47665 -11335
rect 42165 -11510 42175 -11390
rect 42295 -11510 42350 -11390
rect 42470 -11510 42515 -11390
rect 42635 -11510 42680 -11390
rect 42800 -11510 42845 -11390
rect 42965 -11510 43020 -11390
rect 43140 -11510 43185 -11390
rect 43305 -11510 43350 -11390
rect 43470 -11510 43515 -11390
rect 43635 -11510 43690 -11390
rect 43810 -11510 43855 -11390
rect 43975 -11510 44020 -11390
rect 44140 -11510 44185 -11390
rect 44305 -11510 44360 -11390
rect 44480 -11510 44525 -11390
rect 44645 -11510 44690 -11390
rect 44810 -11510 44855 -11390
rect 44975 -11510 45030 -11390
rect 45150 -11510 45195 -11390
rect 45315 -11510 45360 -11390
rect 45480 -11510 45525 -11390
rect 45645 -11510 45700 -11390
rect 45820 -11510 45865 -11390
rect 45985 -11510 46030 -11390
rect 46150 -11510 46195 -11390
rect 46315 -11510 46370 -11390
rect 46490 -11510 46535 -11390
rect 46655 -11510 46700 -11390
rect 46820 -11510 46865 -11390
rect 46985 -11510 47040 -11390
rect 47160 -11510 47205 -11390
rect 47325 -11510 47370 -11390
rect 47490 -11510 47535 -11390
rect 47655 -11510 47665 -11390
rect 42165 -11555 47665 -11510
rect 42165 -11675 42175 -11555
rect 42295 -11675 42350 -11555
rect 42470 -11675 42515 -11555
rect 42635 -11675 42680 -11555
rect 42800 -11675 42845 -11555
rect 42965 -11675 43020 -11555
rect 43140 -11675 43185 -11555
rect 43305 -11675 43350 -11555
rect 43470 -11675 43515 -11555
rect 43635 -11675 43690 -11555
rect 43810 -11675 43855 -11555
rect 43975 -11675 44020 -11555
rect 44140 -11675 44185 -11555
rect 44305 -11675 44360 -11555
rect 44480 -11675 44525 -11555
rect 44645 -11675 44690 -11555
rect 44810 -11675 44855 -11555
rect 44975 -11675 45030 -11555
rect 45150 -11675 45195 -11555
rect 45315 -11675 45360 -11555
rect 45480 -11675 45525 -11555
rect 45645 -11675 45700 -11555
rect 45820 -11675 45865 -11555
rect 45985 -11675 46030 -11555
rect 46150 -11675 46195 -11555
rect 46315 -11675 46370 -11555
rect 46490 -11675 46535 -11555
rect 46655 -11675 46700 -11555
rect 46820 -11675 46865 -11555
rect 46985 -11675 47040 -11555
rect 47160 -11675 47205 -11555
rect 47325 -11675 47370 -11555
rect 47490 -11675 47535 -11555
rect 47655 -11675 47665 -11555
rect 42165 -11720 47665 -11675
rect 42165 -11840 42175 -11720
rect 42295 -11840 42350 -11720
rect 42470 -11840 42515 -11720
rect 42635 -11840 42680 -11720
rect 42800 -11840 42845 -11720
rect 42965 -11840 43020 -11720
rect 43140 -11840 43185 -11720
rect 43305 -11840 43350 -11720
rect 43470 -11840 43515 -11720
rect 43635 -11840 43690 -11720
rect 43810 -11840 43855 -11720
rect 43975 -11840 44020 -11720
rect 44140 -11840 44185 -11720
rect 44305 -11840 44360 -11720
rect 44480 -11840 44525 -11720
rect 44645 -11840 44690 -11720
rect 44810 -11840 44855 -11720
rect 44975 -11840 45030 -11720
rect 45150 -11840 45195 -11720
rect 45315 -11840 45360 -11720
rect 45480 -11840 45525 -11720
rect 45645 -11840 45700 -11720
rect 45820 -11840 45865 -11720
rect 45985 -11840 46030 -11720
rect 46150 -11840 46195 -11720
rect 46315 -11840 46370 -11720
rect 46490 -11840 46535 -11720
rect 46655 -11840 46700 -11720
rect 46820 -11840 46865 -11720
rect 46985 -11840 47040 -11720
rect 47160 -11840 47205 -11720
rect 47325 -11840 47370 -11720
rect 47490 -11840 47535 -11720
rect 47655 -11840 47665 -11720
rect 42165 -11885 47665 -11840
rect 42165 -12005 42175 -11885
rect 42295 -12005 42350 -11885
rect 42470 -12005 42515 -11885
rect 42635 -12005 42680 -11885
rect 42800 -12005 42845 -11885
rect 42965 -12005 43020 -11885
rect 43140 -12005 43185 -11885
rect 43305 -12005 43350 -11885
rect 43470 -12005 43515 -11885
rect 43635 -12005 43690 -11885
rect 43810 -12005 43855 -11885
rect 43975 -12005 44020 -11885
rect 44140 -12005 44185 -11885
rect 44305 -12005 44360 -11885
rect 44480 -12005 44525 -11885
rect 44645 -12005 44690 -11885
rect 44810 -12005 44855 -11885
rect 44975 -12005 45030 -11885
rect 45150 -12005 45195 -11885
rect 45315 -12005 45360 -11885
rect 45480 -12005 45525 -11885
rect 45645 -12005 45700 -11885
rect 45820 -12005 45865 -11885
rect 45985 -12005 46030 -11885
rect 46150 -12005 46195 -11885
rect 46315 -12005 46370 -11885
rect 46490 -12005 46535 -11885
rect 46655 -12005 46700 -11885
rect 46820 -12005 46865 -11885
rect 46985 -12005 47040 -11885
rect 47160 -12005 47205 -11885
rect 47325 -12005 47370 -11885
rect 47490 -12005 47535 -11885
rect 47655 -12005 47665 -11885
rect 42165 -12060 47665 -12005
rect 42165 -12180 42175 -12060
rect 42295 -12180 42350 -12060
rect 42470 -12180 42515 -12060
rect 42635 -12180 42680 -12060
rect 42800 -12180 42845 -12060
rect 42965 -12180 43020 -12060
rect 43140 -12180 43185 -12060
rect 43305 -12180 43350 -12060
rect 43470 -12180 43515 -12060
rect 43635 -12180 43690 -12060
rect 43810 -12180 43855 -12060
rect 43975 -12180 44020 -12060
rect 44140 -12180 44185 -12060
rect 44305 -12180 44360 -12060
rect 44480 -12180 44525 -12060
rect 44645 -12180 44690 -12060
rect 44810 -12180 44855 -12060
rect 44975 -12180 45030 -12060
rect 45150 -12180 45195 -12060
rect 45315 -12180 45360 -12060
rect 45480 -12180 45525 -12060
rect 45645 -12180 45700 -12060
rect 45820 -12180 45865 -12060
rect 45985 -12180 46030 -12060
rect 46150 -12180 46195 -12060
rect 46315 -12180 46370 -12060
rect 46490 -12180 46535 -12060
rect 46655 -12180 46700 -12060
rect 46820 -12180 46865 -12060
rect 46985 -12180 47040 -12060
rect 47160 -12180 47205 -12060
rect 47325 -12180 47370 -12060
rect 47490 -12180 47535 -12060
rect 47655 -12180 47665 -12060
rect 42165 -12225 47665 -12180
rect 42165 -12345 42175 -12225
rect 42295 -12345 42350 -12225
rect 42470 -12345 42515 -12225
rect 42635 -12345 42680 -12225
rect 42800 -12345 42845 -12225
rect 42965 -12345 43020 -12225
rect 43140 -12345 43185 -12225
rect 43305 -12345 43350 -12225
rect 43470 -12345 43515 -12225
rect 43635 -12345 43690 -12225
rect 43810 -12345 43855 -12225
rect 43975 -12345 44020 -12225
rect 44140 -12345 44185 -12225
rect 44305 -12345 44360 -12225
rect 44480 -12345 44525 -12225
rect 44645 -12345 44690 -12225
rect 44810 -12345 44855 -12225
rect 44975 -12345 45030 -12225
rect 45150 -12345 45195 -12225
rect 45315 -12345 45360 -12225
rect 45480 -12345 45525 -12225
rect 45645 -12345 45700 -12225
rect 45820 -12345 45865 -12225
rect 45985 -12345 46030 -12225
rect 46150 -12345 46195 -12225
rect 46315 -12345 46370 -12225
rect 46490 -12345 46535 -12225
rect 46655 -12345 46700 -12225
rect 46820 -12345 46865 -12225
rect 46985 -12345 47040 -12225
rect 47160 -12345 47205 -12225
rect 47325 -12345 47370 -12225
rect 47490 -12345 47535 -12225
rect 47655 -12345 47665 -12225
rect 42165 -12390 47665 -12345
rect 42165 -12510 42175 -12390
rect 42295 -12510 42350 -12390
rect 42470 -12510 42515 -12390
rect 42635 -12510 42680 -12390
rect 42800 -12510 42845 -12390
rect 42965 -12510 43020 -12390
rect 43140 -12510 43185 -12390
rect 43305 -12510 43350 -12390
rect 43470 -12510 43515 -12390
rect 43635 -12510 43690 -12390
rect 43810 -12510 43855 -12390
rect 43975 -12510 44020 -12390
rect 44140 -12510 44185 -12390
rect 44305 -12510 44360 -12390
rect 44480 -12510 44525 -12390
rect 44645 -12510 44690 -12390
rect 44810 -12510 44855 -12390
rect 44975 -12510 45030 -12390
rect 45150 -12510 45195 -12390
rect 45315 -12510 45360 -12390
rect 45480 -12510 45525 -12390
rect 45645 -12510 45700 -12390
rect 45820 -12510 45865 -12390
rect 45985 -12510 46030 -12390
rect 46150 -12510 46195 -12390
rect 46315 -12510 46370 -12390
rect 46490 -12510 46535 -12390
rect 46655 -12510 46700 -12390
rect 46820 -12510 46865 -12390
rect 46985 -12510 47040 -12390
rect 47160 -12510 47205 -12390
rect 47325 -12510 47370 -12390
rect 47490 -12510 47535 -12390
rect 47655 -12510 47665 -12390
rect 42165 -12555 47665 -12510
rect 42165 -12675 42175 -12555
rect 42295 -12675 42350 -12555
rect 42470 -12675 42515 -12555
rect 42635 -12675 42680 -12555
rect 42800 -12675 42845 -12555
rect 42965 -12675 43020 -12555
rect 43140 -12675 43185 -12555
rect 43305 -12675 43350 -12555
rect 43470 -12675 43515 -12555
rect 43635 -12675 43690 -12555
rect 43810 -12675 43855 -12555
rect 43975 -12675 44020 -12555
rect 44140 -12675 44185 -12555
rect 44305 -12675 44360 -12555
rect 44480 -12675 44525 -12555
rect 44645 -12675 44690 -12555
rect 44810 -12675 44855 -12555
rect 44975 -12675 45030 -12555
rect 45150 -12675 45195 -12555
rect 45315 -12675 45360 -12555
rect 45480 -12675 45525 -12555
rect 45645 -12675 45700 -12555
rect 45820 -12675 45865 -12555
rect 45985 -12675 46030 -12555
rect 46150 -12675 46195 -12555
rect 46315 -12675 46370 -12555
rect 46490 -12675 46535 -12555
rect 46655 -12675 46700 -12555
rect 46820 -12675 46865 -12555
rect 46985 -12675 47040 -12555
rect 47160 -12675 47205 -12555
rect 47325 -12675 47370 -12555
rect 47490 -12675 47535 -12555
rect 47655 -12675 47665 -12555
rect 42165 -12730 47665 -12675
rect 42165 -12850 42175 -12730
rect 42295 -12850 42350 -12730
rect 42470 -12850 42515 -12730
rect 42635 -12850 42680 -12730
rect 42800 -12850 42845 -12730
rect 42965 -12850 43020 -12730
rect 43140 -12850 43185 -12730
rect 43305 -12850 43350 -12730
rect 43470 -12850 43515 -12730
rect 43635 -12850 43690 -12730
rect 43810 -12850 43855 -12730
rect 43975 -12850 44020 -12730
rect 44140 -12850 44185 -12730
rect 44305 -12850 44360 -12730
rect 44480 -12850 44525 -12730
rect 44645 -12850 44690 -12730
rect 44810 -12850 44855 -12730
rect 44975 -12850 45030 -12730
rect 45150 -12850 45195 -12730
rect 45315 -12850 45360 -12730
rect 45480 -12850 45525 -12730
rect 45645 -12850 45700 -12730
rect 45820 -12850 45865 -12730
rect 45985 -12850 46030 -12730
rect 46150 -12850 46195 -12730
rect 46315 -12850 46370 -12730
rect 46490 -12850 46535 -12730
rect 46655 -12850 46700 -12730
rect 46820 -12850 46865 -12730
rect 46985 -12850 47040 -12730
rect 47160 -12850 47205 -12730
rect 47325 -12850 47370 -12730
rect 47490 -12850 47535 -12730
rect 47655 -12850 47665 -12730
rect 42165 -12895 47665 -12850
rect 42165 -13015 42175 -12895
rect 42295 -13015 42350 -12895
rect 42470 -13015 42515 -12895
rect 42635 -13015 42680 -12895
rect 42800 -13015 42845 -12895
rect 42965 -13015 43020 -12895
rect 43140 -13015 43185 -12895
rect 43305 -13015 43350 -12895
rect 43470 -13015 43515 -12895
rect 43635 -13015 43690 -12895
rect 43810 -13015 43855 -12895
rect 43975 -13015 44020 -12895
rect 44140 -13015 44185 -12895
rect 44305 -13015 44360 -12895
rect 44480 -13015 44525 -12895
rect 44645 -13015 44690 -12895
rect 44810 -13015 44855 -12895
rect 44975 -13015 45030 -12895
rect 45150 -13015 45195 -12895
rect 45315 -13015 45360 -12895
rect 45480 -13015 45525 -12895
rect 45645 -13015 45700 -12895
rect 45820 -13015 45865 -12895
rect 45985 -13015 46030 -12895
rect 46150 -13015 46195 -12895
rect 46315 -13015 46370 -12895
rect 46490 -13015 46535 -12895
rect 46655 -13015 46700 -12895
rect 46820 -13015 46865 -12895
rect 46985 -13015 47040 -12895
rect 47160 -13015 47205 -12895
rect 47325 -13015 47370 -12895
rect 47490 -13015 47535 -12895
rect 47655 -13015 47665 -12895
rect 42165 -13060 47665 -13015
rect 42165 -13180 42175 -13060
rect 42295 -13180 42350 -13060
rect 42470 -13180 42515 -13060
rect 42635 -13180 42680 -13060
rect 42800 -13180 42845 -13060
rect 42965 -13180 43020 -13060
rect 43140 -13180 43185 -13060
rect 43305 -13180 43350 -13060
rect 43470 -13180 43515 -13060
rect 43635 -13180 43690 -13060
rect 43810 -13180 43855 -13060
rect 43975 -13180 44020 -13060
rect 44140 -13180 44185 -13060
rect 44305 -13180 44360 -13060
rect 44480 -13180 44525 -13060
rect 44645 -13180 44690 -13060
rect 44810 -13180 44855 -13060
rect 44975 -13180 45030 -13060
rect 45150 -13180 45195 -13060
rect 45315 -13180 45360 -13060
rect 45480 -13180 45525 -13060
rect 45645 -13180 45700 -13060
rect 45820 -13180 45865 -13060
rect 45985 -13180 46030 -13060
rect 46150 -13180 46195 -13060
rect 46315 -13180 46370 -13060
rect 46490 -13180 46535 -13060
rect 46655 -13180 46700 -13060
rect 46820 -13180 46865 -13060
rect 46985 -13180 47040 -13060
rect 47160 -13180 47205 -13060
rect 47325 -13180 47370 -13060
rect 47490 -13180 47535 -13060
rect 47655 -13180 47665 -13060
rect 42165 -13225 47665 -13180
rect 42165 -13345 42175 -13225
rect 42295 -13345 42350 -13225
rect 42470 -13345 42515 -13225
rect 42635 -13345 42680 -13225
rect 42800 -13345 42845 -13225
rect 42965 -13345 43020 -13225
rect 43140 -13345 43185 -13225
rect 43305 -13345 43350 -13225
rect 43470 -13345 43515 -13225
rect 43635 -13345 43690 -13225
rect 43810 -13345 43855 -13225
rect 43975 -13345 44020 -13225
rect 44140 -13345 44185 -13225
rect 44305 -13345 44360 -13225
rect 44480 -13345 44525 -13225
rect 44645 -13345 44690 -13225
rect 44810 -13345 44855 -13225
rect 44975 -13345 45030 -13225
rect 45150 -13345 45195 -13225
rect 45315 -13345 45360 -13225
rect 45480 -13345 45525 -13225
rect 45645 -13345 45700 -13225
rect 45820 -13345 45865 -13225
rect 45985 -13345 46030 -13225
rect 46150 -13345 46195 -13225
rect 46315 -13345 46370 -13225
rect 46490 -13345 46535 -13225
rect 46655 -13345 46700 -13225
rect 46820 -13345 46865 -13225
rect 46985 -13345 47040 -13225
rect 47160 -13345 47205 -13225
rect 47325 -13345 47370 -13225
rect 47490 -13345 47535 -13225
rect 47655 -13345 47665 -13225
rect 42165 -13400 47665 -13345
rect 42165 -13520 42175 -13400
rect 42295 -13520 42350 -13400
rect 42470 -13520 42515 -13400
rect 42635 -13520 42680 -13400
rect 42800 -13520 42845 -13400
rect 42965 -13520 43020 -13400
rect 43140 -13520 43185 -13400
rect 43305 -13520 43350 -13400
rect 43470 -13520 43515 -13400
rect 43635 -13520 43690 -13400
rect 43810 -13520 43855 -13400
rect 43975 -13520 44020 -13400
rect 44140 -13520 44185 -13400
rect 44305 -13520 44360 -13400
rect 44480 -13520 44525 -13400
rect 44645 -13520 44690 -13400
rect 44810 -13520 44855 -13400
rect 44975 -13520 45030 -13400
rect 45150 -13520 45195 -13400
rect 45315 -13520 45360 -13400
rect 45480 -13520 45525 -13400
rect 45645 -13520 45700 -13400
rect 45820 -13520 45865 -13400
rect 45985 -13520 46030 -13400
rect 46150 -13520 46195 -13400
rect 46315 -13520 46370 -13400
rect 46490 -13520 46535 -13400
rect 46655 -13520 46700 -13400
rect 46820 -13520 46865 -13400
rect 46985 -13520 47040 -13400
rect 47160 -13520 47205 -13400
rect 47325 -13520 47370 -13400
rect 47490 -13520 47535 -13400
rect 47655 -13520 47665 -13400
rect 42165 -13565 47665 -13520
rect 42165 -13685 42175 -13565
rect 42295 -13685 42350 -13565
rect 42470 -13685 42515 -13565
rect 42635 -13685 42680 -13565
rect 42800 -13685 42845 -13565
rect 42965 -13685 43020 -13565
rect 43140 -13685 43185 -13565
rect 43305 -13685 43350 -13565
rect 43470 -13685 43515 -13565
rect 43635 -13685 43690 -13565
rect 43810 -13685 43855 -13565
rect 43975 -13685 44020 -13565
rect 44140 -13685 44185 -13565
rect 44305 -13685 44360 -13565
rect 44480 -13685 44525 -13565
rect 44645 -13685 44690 -13565
rect 44810 -13685 44855 -13565
rect 44975 -13685 45030 -13565
rect 45150 -13685 45195 -13565
rect 45315 -13685 45360 -13565
rect 45480 -13685 45525 -13565
rect 45645 -13685 45700 -13565
rect 45820 -13685 45865 -13565
rect 45985 -13685 46030 -13565
rect 46150 -13685 46195 -13565
rect 46315 -13685 46370 -13565
rect 46490 -13685 46535 -13565
rect 46655 -13685 46700 -13565
rect 46820 -13685 46865 -13565
rect 46985 -13685 47040 -13565
rect 47160 -13685 47205 -13565
rect 47325 -13685 47370 -13565
rect 47490 -13685 47535 -13565
rect 47655 -13685 47665 -13565
rect 42165 -13730 47665 -13685
rect 42165 -13850 42175 -13730
rect 42295 -13850 42350 -13730
rect 42470 -13850 42515 -13730
rect 42635 -13850 42680 -13730
rect 42800 -13850 42845 -13730
rect 42965 -13850 43020 -13730
rect 43140 -13850 43185 -13730
rect 43305 -13850 43350 -13730
rect 43470 -13850 43515 -13730
rect 43635 -13850 43690 -13730
rect 43810 -13850 43855 -13730
rect 43975 -13850 44020 -13730
rect 44140 -13850 44185 -13730
rect 44305 -13850 44360 -13730
rect 44480 -13850 44525 -13730
rect 44645 -13850 44690 -13730
rect 44810 -13850 44855 -13730
rect 44975 -13850 45030 -13730
rect 45150 -13850 45195 -13730
rect 45315 -13850 45360 -13730
rect 45480 -13850 45525 -13730
rect 45645 -13850 45700 -13730
rect 45820 -13850 45865 -13730
rect 45985 -13850 46030 -13730
rect 46150 -13850 46195 -13730
rect 46315 -13850 46370 -13730
rect 46490 -13850 46535 -13730
rect 46655 -13850 46700 -13730
rect 46820 -13850 46865 -13730
rect 46985 -13850 47040 -13730
rect 47160 -13850 47205 -13730
rect 47325 -13850 47370 -13730
rect 47490 -13850 47535 -13730
rect 47655 -13850 47665 -13730
rect 42165 -13895 47665 -13850
rect 42165 -14015 42175 -13895
rect 42295 -14015 42350 -13895
rect 42470 -14015 42515 -13895
rect 42635 -14015 42680 -13895
rect 42800 -14015 42845 -13895
rect 42965 -14015 43020 -13895
rect 43140 -14015 43185 -13895
rect 43305 -14015 43350 -13895
rect 43470 -14015 43515 -13895
rect 43635 -14015 43690 -13895
rect 43810 -14015 43855 -13895
rect 43975 -14015 44020 -13895
rect 44140 -14015 44185 -13895
rect 44305 -14015 44360 -13895
rect 44480 -14015 44525 -13895
rect 44645 -14015 44690 -13895
rect 44810 -14015 44855 -13895
rect 44975 -14015 45030 -13895
rect 45150 -14015 45195 -13895
rect 45315 -14015 45360 -13895
rect 45480 -14015 45525 -13895
rect 45645 -14015 45700 -13895
rect 45820 -14015 45865 -13895
rect 45985 -14015 46030 -13895
rect 46150 -14015 46195 -13895
rect 46315 -14015 46370 -13895
rect 46490 -14015 46535 -13895
rect 46655 -14015 46700 -13895
rect 46820 -14015 46865 -13895
rect 46985 -14015 47040 -13895
rect 47160 -14015 47205 -13895
rect 47325 -14015 47370 -13895
rect 47490 -14015 47535 -13895
rect 47655 -14015 47665 -13895
rect 42165 -14070 47665 -14015
rect 42165 -14190 42175 -14070
rect 42295 -14190 42350 -14070
rect 42470 -14190 42515 -14070
rect 42635 -14190 42680 -14070
rect 42800 -14190 42845 -14070
rect 42965 -14190 43020 -14070
rect 43140 -14190 43185 -14070
rect 43305 -14190 43350 -14070
rect 43470 -14190 43515 -14070
rect 43635 -14190 43690 -14070
rect 43810 -14190 43855 -14070
rect 43975 -14190 44020 -14070
rect 44140 -14190 44185 -14070
rect 44305 -14190 44360 -14070
rect 44480 -14190 44525 -14070
rect 44645 -14190 44690 -14070
rect 44810 -14190 44855 -14070
rect 44975 -14190 45030 -14070
rect 45150 -14190 45195 -14070
rect 45315 -14190 45360 -14070
rect 45480 -14190 45525 -14070
rect 45645 -14190 45700 -14070
rect 45820 -14190 45865 -14070
rect 45985 -14190 46030 -14070
rect 46150 -14190 46195 -14070
rect 46315 -14190 46370 -14070
rect 46490 -14190 46535 -14070
rect 46655 -14190 46700 -14070
rect 46820 -14190 46865 -14070
rect 46985 -14190 47040 -14070
rect 47160 -14190 47205 -14070
rect 47325 -14190 47370 -14070
rect 47490 -14190 47535 -14070
rect 47655 -14190 47665 -14070
rect 42165 -14235 47665 -14190
rect 42165 -14355 42175 -14235
rect 42295 -14355 42350 -14235
rect 42470 -14355 42515 -14235
rect 42635 -14355 42680 -14235
rect 42800 -14355 42845 -14235
rect 42965 -14355 43020 -14235
rect 43140 -14355 43185 -14235
rect 43305 -14355 43350 -14235
rect 43470 -14355 43515 -14235
rect 43635 -14355 43690 -14235
rect 43810 -14355 43855 -14235
rect 43975 -14355 44020 -14235
rect 44140 -14355 44185 -14235
rect 44305 -14355 44360 -14235
rect 44480 -14355 44525 -14235
rect 44645 -14355 44690 -14235
rect 44810 -14355 44855 -14235
rect 44975 -14355 45030 -14235
rect 45150 -14355 45195 -14235
rect 45315 -14355 45360 -14235
rect 45480 -14355 45525 -14235
rect 45645 -14355 45700 -14235
rect 45820 -14355 45865 -14235
rect 45985 -14355 46030 -14235
rect 46150 -14355 46195 -14235
rect 46315 -14355 46370 -14235
rect 46490 -14355 46535 -14235
rect 46655 -14355 46700 -14235
rect 46820 -14355 46865 -14235
rect 46985 -14355 47040 -14235
rect 47160 -14355 47205 -14235
rect 47325 -14355 47370 -14235
rect 47490 -14355 47535 -14235
rect 47655 -14355 47665 -14235
rect 42165 -14400 47665 -14355
rect 42165 -14520 42175 -14400
rect 42295 -14520 42350 -14400
rect 42470 -14520 42515 -14400
rect 42635 -14520 42680 -14400
rect 42800 -14520 42845 -14400
rect 42965 -14520 43020 -14400
rect 43140 -14520 43185 -14400
rect 43305 -14520 43350 -14400
rect 43470 -14520 43515 -14400
rect 43635 -14520 43690 -14400
rect 43810 -14520 43855 -14400
rect 43975 -14520 44020 -14400
rect 44140 -14520 44185 -14400
rect 44305 -14520 44360 -14400
rect 44480 -14520 44525 -14400
rect 44645 -14520 44690 -14400
rect 44810 -14520 44855 -14400
rect 44975 -14520 45030 -14400
rect 45150 -14520 45195 -14400
rect 45315 -14520 45360 -14400
rect 45480 -14520 45525 -14400
rect 45645 -14520 45700 -14400
rect 45820 -14520 45865 -14400
rect 45985 -14520 46030 -14400
rect 46150 -14520 46195 -14400
rect 46315 -14520 46370 -14400
rect 46490 -14520 46535 -14400
rect 46655 -14520 46700 -14400
rect 46820 -14520 46865 -14400
rect 46985 -14520 47040 -14400
rect 47160 -14520 47205 -14400
rect 47325 -14520 47370 -14400
rect 47490 -14520 47535 -14400
rect 47655 -14520 47665 -14400
rect 42165 -14565 47665 -14520
rect 42165 -14685 42175 -14565
rect 42295 -14685 42350 -14565
rect 42470 -14685 42515 -14565
rect 42635 -14685 42680 -14565
rect 42800 -14685 42845 -14565
rect 42965 -14685 43020 -14565
rect 43140 -14685 43185 -14565
rect 43305 -14685 43350 -14565
rect 43470 -14685 43515 -14565
rect 43635 -14685 43690 -14565
rect 43810 -14685 43855 -14565
rect 43975 -14685 44020 -14565
rect 44140 -14685 44185 -14565
rect 44305 -14685 44360 -14565
rect 44480 -14685 44525 -14565
rect 44645 -14685 44690 -14565
rect 44810 -14685 44855 -14565
rect 44975 -14685 45030 -14565
rect 45150 -14685 45195 -14565
rect 45315 -14685 45360 -14565
rect 45480 -14685 45525 -14565
rect 45645 -14685 45700 -14565
rect 45820 -14685 45865 -14565
rect 45985 -14685 46030 -14565
rect 46150 -14685 46195 -14565
rect 46315 -14685 46370 -14565
rect 46490 -14685 46535 -14565
rect 46655 -14685 46700 -14565
rect 46820 -14685 46865 -14565
rect 46985 -14685 47040 -14565
rect 47160 -14685 47205 -14565
rect 47325 -14685 47370 -14565
rect 47490 -14685 47535 -14565
rect 47655 -14685 47665 -14565
rect 42165 -14740 47665 -14685
rect 42165 -14860 42175 -14740
rect 42295 -14860 42350 -14740
rect 42470 -14860 42515 -14740
rect 42635 -14860 42680 -14740
rect 42800 -14860 42845 -14740
rect 42965 -14860 43020 -14740
rect 43140 -14860 43185 -14740
rect 43305 -14860 43350 -14740
rect 43470 -14860 43515 -14740
rect 43635 -14860 43690 -14740
rect 43810 -14860 43855 -14740
rect 43975 -14860 44020 -14740
rect 44140 -14860 44185 -14740
rect 44305 -14860 44360 -14740
rect 44480 -14860 44525 -14740
rect 44645 -14860 44690 -14740
rect 44810 -14860 44855 -14740
rect 44975 -14860 45030 -14740
rect 45150 -14860 45195 -14740
rect 45315 -14860 45360 -14740
rect 45480 -14860 45525 -14740
rect 45645 -14860 45700 -14740
rect 45820 -14860 45865 -14740
rect 45985 -14860 46030 -14740
rect 46150 -14860 46195 -14740
rect 46315 -14860 46370 -14740
rect 46490 -14860 46535 -14740
rect 46655 -14860 46700 -14740
rect 46820 -14860 46865 -14740
rect 46985 -14860 47040 -14740
rect 47160 -14860 47205 -14740
rect 47325 -14860 47370 -14740
rect 47490 -14860 47535 -14740
rect 47655 -14860 47665 -14740
rect 42165 -14905 47665 -14860
rect 42165 -15025 42175 -14905
rect 42295 -15025 42350 -14905
rect 42470 -15025 42515 -14905
rect 42635 -15025 42680 -14905
rect 42800 -15025 42845 -14905
rect 42965 -15025 43020 -14905
rect 43140 -15025 43185 -14905
rect 43305 -15025 43350 -14905
rect 43470 -15025 43515 -14905
rect 43635 -15025 43690 -14905
rect 43810 -15025 43855 -14905
rect 43975 -15025 44020 -14905
rect 44140 -15025 44185 -14905
rect 44305 -15025 44360 -14905
rect 44480 -15025 44525 -14905
rect 44645 -15025 44690 -14905
rect 44810 -15025 44855 -14905
rect 44975 -15025 45030 -14905
rect 45150 -15025 45195 -14905
rect 45315 -15025 45360 -14905
rect 45480 -15025 45525 -14905
rect 45645 -15025 45700 -14905
rect 45820 -15025 45865 -14905
rect 45985 -15025 46030 -14905
rect 46150 -15025 46195 -14905
rect 46315 -15025 46370 -14905
rect 46490 -15025 46535 -14905
rect 46655 -15025 46700 -14905
rect 46820 -15025 46865 -14905
rect 46985 -15025 47040 -14905
rect 47160 -15025 47205 -14905
rect 47325 -15025 47370 -14905
rect 47490 -15025 47535 -14905
rect 47655 -15025 47665 -14905
rect 42165 -15070 47665 -15025
rect 42165 -15190 42175 -15070
rect 42295 -15190 42350 -15070
rect 42470 -15190 42515 -15070
rect 42635 -15190 42680 -15070
rect 42800 -15190 42845 -15070
rect 42965 -15190 43020 -15070
rect 43140 -15190 43185 -15070
rect 43305 -15190 43350 -15070
rect 43470 -15190 43515 -15070
rect 43635 -15190 43690 -15070
rect 43810 -15190 43855 -15070
rect 43975 -15190 44020 -15070
rect 44140 -15190 44185 -15070
rect 44305 -15190 44360 -15070
rect 44480 -15190 44525 -15070
rect 44645 -15190 44690 -15070
rect 44810 -15190 44855 -15070
rect 44975 -15190 45030 -15070
rect 45150 -15190 45195 -15070
rect 45315 -15190 45360 -15070
rect 45480 -15190 45525 -15070
rect 45645 -15190 45700 -15070
rect 45820 -15190 45865 -15070
rect 45985 -15190 46030 -15070
rect 46150 -15190 46195 -15070
rect 46315 -15190 46370 -15070
rect 46490 -15190 46535 -15070
rect 46655 -15190 46700 -15070
rect 46820 -15190 46865 -15070
rect 46985 -15190 47040 -15070
rect 47160 -15190 47205 -15070
rect 47325 -15190 47370 -15070
rect 47490 -15190 47535 -15070
rect 47655 -15190 47665 -15070
rect 42165 -15235 47665 -15190
rect 42165 -15355 42175 -15235
rect 42295 -15355 42350 -15235
rect 42470 -15355 42515 -15235
rect 42635 -15355 42680 -15235
rect 42800 -15355 42845 -15235
rect 42965 -15355 43020 -15235
rect 43140 -15355 43185 -15235
rect 43305 -15355 43350 -15235
rect 43470 -15355 43515 -15235
rect 43635 -15355 43690 -15235
rect 43810 -15355 43855 -15235
rect 43975 -15355 44020 -15235
rect 44140 -15355 44185 -15235
rect 44305 -15355 44360 -15235
rect 44480 -15355 44525 -15235
rect 44645 -15355 44690 -15235
rect 44810 -15355 44855 -15235
rect 44975 -15355 45030 -15235
rect 45150 -15355 45195 -15235
rect 45315 -15355 45360 -15235
rect 45480 -15355 45525 -15235
rect 45645 -15355 45700 -15235
rect 45820 -15355 45865 -15235
rect 45985 -15355 46030 -15235
rect 46150 -15355 46195 -15235
rect 46315 -15355 46370 -15235
rect 46490 -15355 46535 -15235
rect 46655 -15355 46700 -15235
rect 46820 -15355 46865 -15235
rect 46985 -15355 47040 -15235
rect 47160 -15355 47205 -15235
rect 47325 -15355 47370 -15235
rect 47490 -15355 47535 -15235
rect 47655 -15355 47665 -15235
rect 42165 -15410 47665 -15355
rect 42165 -15530 42175 -15410
rect 42295 -15530 42350 -15410
rect 42470 -15530 42515 -15410
rect 42635 -15530 42680 -15410
rect 42800 -15530 42845 -15410
rect 42965 -15530 43020 -15410
rect 43140 -15530 43185 -15410
rect 43305 -15530 43350 -15410
rect 43470 -15530 43515 -15410
rect 43635 -15530 43690 -15410
rect 43810 -15530 43855 -15410
rect 43975 -15530 44020 -15410
rect 44140 -15530 44185 -15410
rect 44305 -15530 44360 -15410
rect 44480 -15530 44525 -15410
rect 44645 -15530 44690 -15410
rect 44810 -15530 44855 -15410
rect 44975 -15530 45030 -15410
rect 45150 -15530 45195 -15410
rect 45315 -15530 45360 -15410
rect 45480 -15530 45525 -15410
rect 45645 -15530 45700 -15410
rect 45820 -15530 45865 -15410
rect 45985 -15530 46030 -15410
rect 46150 -15530 46195 -15410
rect 46315 -15530 46370 -15410
rect 46490 -15530 46535 -15410
rect 46655 -15530 46700 -15410
rect 46820 -15530 46865 -15410
rect 46985 -15530 47040 -15410
rect 47160 -15530 47205 -15410
rect 47325 -15530 47370 -15410
rect 47490 -15530 47535 -15410
rect 47655 -15530 47665 -15410
rect 42165 -15540 47665 -15530
rect 47855 -10050 53355 -10040
rect 47855 -10170 47865 -10050
rect 47985 -10170 48040 -10050
rect 48160 -10170 48205 -10050
rect 48325 -10170 48370 -10050
rect 48490 -10170 48535 -10050
rect 48655 -10170 48710 -10050
rect 48830 -10170 48875 -10050
rect 48995 -10170 49040 -10050
rect 49160 -10170 49205 -10050
rect 49325 -10170 49380 -10050
rect 49500 -10170 49545 -10050
rect 49665 -10170 49710 -10050
rect 49830 -10170 49875 -10050
rect 49995 -10170 50050 -10050
rect 50170 -10170 50215 -10050
rect 50335 -10170 50380 -10050
rect 50500 -10170 50545 -10050
rect 50665 -10170 50720 -10050
rect 50840 -10170 50885 -10050
rect 51005 -10170 51050 -10050
rect 51170 -10170 51215 -10050
rect 51335 -10170 51390 -10050
rect 51510 -10170 51555 -10050
rect 51675 -10170 51720 -10050
rect 51840 -10170 51885 -10050
rect 52005 -10170 52060 -10050
rect 52180 -10170 52225 -10050
rect 52345 -10170 52390 -10050
rect 52510 -10170 52555 -10050
rect 52675 -10170 52730 -10050
rect 52850 -10170 52895 -10050
rect 53015 -10170 53060 -10050
rect 53180 -10170 53225 -10050
rect 53345 -10170 53355 -10050
rect 47855 -10215 53355 -10170
rect 47855 -10335 47865 -10215
rect 47985 -10335 48040 -10215
rect 48160 -10335 48205 -10215
rect 48325 -10335 48370 -10215
rect 48490 -10335 48535 -10215
rect 48655 -10335 48710 -10215
rect 48830 -10335 48875 -10215
rect 48995 -10335 49040 -10215
rect 49160 -10335 49205 -10215
rect 49325 -10335 49380 -10215
rect 49500 -10335 49545 -10215
rect 49665 -10335 49710 -10215
rect 49830 -10335 49875 -10215
rect 49995 -10335 50050 -10215
rect 50170 -10335 50215 -10215
rect 50335 -10335 50380 -10215
rect 50500 -10335 50545 -10215
rect 50665 -10335 50720 -10215
rect 50840 -10335 50885 -10215
rect 51005 -10335 51050 -10215
rect 51170 -10335 51215 -10215
rect 51335 -10335 51390 -10215
rect 51510 -10335 51555 -10215
rect 51675 -10335 51720 -10215
rect 51840 -10335 51885 -10215
rect 52005 -10335 52060 -10215
rect 52180 -10335 52225 -10215
rect 52345 -10335 52390 -10215
rect 52510 -10335 52555 -10215
rect 52675 -10335 52730 -10215
rect 52850 -10335 52895 -10215
rect 53015 -10335 53060 -10215
rect 53180 -10335 53225 -10215
rect 53345 -10335 53355 -10215
rect 47855 -10380 53355 -10335
rect 47855 -10500 47865 -10380
rect 47985 -10500 48040 -10380
rect 48160 -10500 48205 -10380
rect 48325 -10500 48370 -10380
rect 48490 -10500 48535 -10380
rect 48655 -10500 48710 -10380
rect 48830 -10500 48875 -10380
rect 48995 -10500 49040 -10380
rect 49160 -10500 49205 -10380
rect 49325 -10500 49380 -10380
rect 49500 -10500 49545 -10380
rect 49665 -10500 49710 -10380
rect 49830 -10500 49875 -10380
rect 49995 -10500 50050 -10380
rect 50170 -10500 50215 -10380
rect 50335 -10500 50380 -10380
rect 50500 -10500 50545 -10380
rect 50665 -10500 50720 -10380
rect 50840 -10500 50885 -10380
rect 51005 -10500 51050 -10380
rect 51170 -10500 51215 -10380
rect 51335 -10500 51390 -10380
rect 51510 -10500 51555 -10380
rect 51675 -10500 51720 -10380
rect 51840 -10500 51885 -10380
rect 52005 -10500 52060 -10380
rect 52180 -10500 52225 -10380
rect 52345 -10500 52390 -10380
rect 52510 -10500 52555 -10380
rect 52675 -10500 52730 -10380
rect 52850 -10500 52895 -10380
rect 53015 -10500 53060 -10380
rect 53180 -10500 53225 -10380
rect 53345 -10500 53355 -10380
rect 47855 -10545 53355 -10500
rect 47855 -10665 47865 -10545
rect 47985 -10665 48040 -10545
rect 48160 -10665 48205 -10545
rect 48325 -10665 48370 -10545
rect 48490 -10665 48535 -10545
rect 48655 -10665 48710 -10545
rect 48830 -10665 48875 -10545
rect 48995 -10665 49040 -10545
rect 49160 -10665 49205 -10545
rect 49325 -10665 49380 -10545
rect 49500 -10665 49545 -10545
rect 49665 -10665 49710 -10545
rect 49830 -10665 49875 -10545
rect 49995 -10665 50050 -10545
rect 50170 -10665 50215 -10545
rect 50335 -10665 50380 -10545
rect 50500 -10665 50545 -10545
rect 50665 -10665 50720 -10545
rect 50840 -10665 50885 -10545
rect 51005 -10665 51050 -10545
rect 51170 -10665 51215 -10545
rect 51335 -10665 51390 -10545
rect 51510 -10665 51555 -10545
rect 51675 -10665 51720 -10545
rect 51840 -10665 51885 -10545
rect 52005 -10665 52060 -10545
rect 52180 -10665 52225 -10545
rect 52345 -10665 52390 -10545
rect 52510 -10665 52555 -10545
rect 52675 -10665 52730 -10545
rect 52850 -10665 52895 -10545
rect 53015 -10665 53060 -10545
rect 53180 -10665 53225 -10545
rect 53345 -10665 53355 -10545
rect 47855 -10720 53355 -10665
rect 47855 -10840 47865 -10720
rect 47985 -10840 48040 -10720
rect 48160 -10840 48205 -10720
rect 48325 -10840 48370 -10720
rect 48490 -10840 48535 -10720
rect 48655 -10840 48710 -10720
rect 48830 -10840 48875 -10720
rect 48995 -10840 49040 -10720
rect 49160 -10840 49205 -10720
rect 49325 -10840 49380 -10720
rect 49500 -10840 49545 -10720
rect 49665 -10840 49710 -10720
rect 49830 -10840 49875 -10720
rect 49995 -10840 50050 -10720
rect 50170 -10840 50215 -10720
rect 50335 -10840 50380 -10720
rect 50500 -10840 50545 -10720
rect 50665 -10840 50720 -10720
rect 50840 -10840 50885 -10720
rect 51005 -10840 51050 -10720
rect 51170 -10840 51215 -10720
rect 51335 -10840 51390 -10720
rect 51510 -10840 51555 -10720
rect 51675 -10840 51720 -10720
rect 51840 -10840 51885 -10720
rect 52005 -10840 52060 -10720
rect 52180 -10840 52225 -10720
rect 52345 -10840 52390 -10720
rect 52510 -10840 52555 -10720
rect 52675 -10840 52730 -10720
rect 52850 -10840 52895 -10720
rect 53015 -10840 53060 -10720
rect 53180 -10840 53225 -10720
rect 53345 -10840 53355 -10720
rect 47855 -10885 53355 -10840
rect 47855 -11005 47865 -10885
rect 47985 -11005 48040 -10885
rect 48160 -11005 48205 -10885
rect 48325 -11005 48370 -10885
rect 48490 -11005 48535 -10885
rect 48655 -11005 48710 -10885
rect 48830 -11005 48875 -10885
rect 48995 -11005 49040 -10885
rect 49160 -11005 49205 -10885
rect 49325 -11005 49380 -10885
rect 49500 -11005 49545 -10885
rect 49665 -11005 49710 -10885
rect 49830 -11005 49875 -10885
rect 49995 -11005 50050 -10885
rect 50170 -11005 50215 -10885
rect 50335 -11005 50380 -10885
rect 50500 -11005 50545 -10885
rect 50665 -11005 50720 -10885
rect 50840 -11005 50885 -10885
rect 51005 -11005 51050 -10885
rect 51170 -11005 51215 -10885
rect 51335 -11005 51390 -10885
rect 51510 -11005 51555 -10885
rect 51675 -11005 51720 -10885
rect 51840 -11005 51885 -10885
rect 52005 -11005 52060 -10885
rect 52180 -11005 52225 -10885
rect 52345 -11005 52390 -10885
rect 52510 -11005 52555 -10885
rect 52675 -11005 52730 -10885
rect 52850 -11005 52895 -10885
rect 53015 -11005 53060 -10885
rect 53180 -11005 53225 -10885
rect 53345 -11005 53355 -10885
rect 47855 -11050 53355 -11005
rect 47855 -11170 47865 -11050
rect 47985 -11170 48040 -11050
rect 48160 -11170 48205 -11050
rect 48325 -11170 48370 -11050
rect 48490 -11170 48535 -11050
rect 48655 -11170 48710 -11050
rect 48830 -11170 48875 -11050
rect 48995 -11170 49040 -11050
rect 49160 -11170 49205 -11050
rect 49325 -11170 49380 -11050
rect 49500 -11170 49545 -11050
rect 49665 -11170 49710 -11050
rect 49830 -11170 49875 -11050
rect 49995 -11170 50050 -11050
rect 50170 -11170 50215 -11050
rect 50335 -11170 50380 -11050
rect 50500 -11170 50545 -11050
rect 50665 -11170 50720 -11050
rect 50840 -11170 50885 -11050
rect 51005 -11170 51050 -11050
rect 51170 -11170 51215 -11050
rect 51335 -11170 51390 -11050
rect 51510 -11170 51555 -11050
rect 51675 -11170 51720 -11050
rect 51840 -11170 51885 -11050
rect 52005 -11170 52060 -11050
rect 52180 -11170 52225 -11050
rect 52345 -11170 52390 -11050
rect 52510 -11170 52555 -11050
rect 52675 -11170 52730 -11050
rect 52850 -11170 52895 -11050
rect 53015 -11170 53060 -11050
rect 53180 -11170 53225 -11050
rect 53345 -11170 53355 -11050
rect 47855 -11215 53355 -11170
rect 47855 -11335 47865 -11215
rect 47985 -11335 48040 -11215
rect 48160 -11335 48205 -11215
rect 48325 -11335 48370 -11215
rect 48490 -11335 48535 -11215
rect 48655 -11335 48710 -11215
rect 48830 -11335 48875 -11215
rect 48995 -11335 49040 -11215
rect 49160 -11335 49205 -11215
rect 49325 -11335 49380 -11215
rect 49500 -11335 49545 -11215
rect 49665 -11335 49710 -11215
rect 49830 -11335 49875 -11215
rect 49995 -11335 50050 -11215
rect 50170 -11335 50215 -11215
rect 50335 -11335 50380 -11215
rect 50500 -11335 50545 -11215
rect 50665 -11335 50720 -11215
rect 50840 -11335 50885 -11215
rect 51005 -11335 51050 -11215
rect 51170 -11335 51215 -11215
rect 51335 -11335 51390 -11215
rect 51510 -11335 51555 -11215
rect 51675 -11335 51720 -11215
rect 51840 -11335 51885 -11215
rect 52005 -11335 52060 -11215
rect 52180 -11335 52225 -11215
rect 52345 -11335 52390 -11215
rect 52510 -11335 52555 -11215
rect 52675 -11335 52730 -11215
rect 52850 -11335 52895 -11215
rect 53015 -11335 53060 -11215
rect 53180 -11335 53225 -11215
rect 53345 -11335 53355 -11215
rect 47855 -11390 53355 -11335
rect 47855 -11510 47865 -11390
rect 47985 -11510 48040 -11390
rect 48160 -11510 48205 -11390
rect 48325 -11510 48370 -11390
rect 48490 -11510 48535 -11390
rect 48655 -11510 48710 -11390
rect 48830 -11510 48875 -11390
rect 48995 -11510 49040 -11390
rect 49160 -11510 49205 -11390
rect 49325 -11510 49380 -11390
rect 49500 -11510 49545 -11390
rect 49665 -11510 49710 -11390
rect 49830 -11510 49875 -11390
rect 49995 -11510 50050 -11390
rect 50170 -11510 50215 -11390
rect 50335 -11510 50380 -11390
rect 50500 -11510 50545 -11390
rect 50665 -11510 50720 -11390
rect 50840 -11510 50885 -11390
rect 51005 -11510 51050 -11390
rect 51170 -11510 51215 -11390
rect 51335 -11510 51390 -11390
rect 51510 -11510 51555 -11390
rect 51675 -11510 51720 -11390
rect 51840 -11510 51885 -11390
rect 52005 -11510 52060 -11390
rect 52180 -11510 52225 -11390
rect 52345 -11510 52390 -11390
rect 52510 -11510 52555 -11390
rect 52675 -11510 52730 -11390
rect 52850 -11510 52895 -11390
rect 53015 -11510 53060 -11390
rect 53180 -11510 53225 -11390
rect 53345 -11510 53355 -11390
rect 47855 -11555 53355 -11510
rect 47855 -11675 47865 -11555
rect 47985 -11675 48040 -11555
rect 48160 -11675 48205 -11555
rect 48325 -11675 48370 -11555
rect 48490 -11675 48535 -11555
rect 48655 -11675 48710 -11555
rect 48830 -11675 48875 -11555
rect 48995 -11675 49040 -11555
rect 49160 -11675 49205 -11555
rect 49325 -11675 49380 -11555
rect 49500 -11675 49545 -11555
rect 49665 -11675 49710 -11555
rect 49830 -11675 49875 -11555
rect 49995 -11675 50050 -11555
rect 50170 -11675 50215 -11555
rect 50335 -11675 50380 -11555
rect 50500 -11675 50545 -11555
rect 50665 -11675 50720 -11555
rect 50840 -11675 50885 -11555
rect 51005 -11675 51050 -11555
rect 51170 -11675 51215 -11555
rect 51335 -11675 51390 -11555
rect 51510 -11675 51555 -11555
rect 51675 -11675 51720 -11555
rect 51840 -11675 51885 -11555
rect 52005 -11675 52060 -11555
rect 52180 -11675 52225 -11555
rect 52345 -11675 52390 -11555
rect 52510 -11675 52555 -11555
rect 52675 -11675 52730 -11555
rect 52850 -11675 52895 -11555
rect 53015 -11675 53060 -11555
rect 53180 -11675 53225 -11555
rect 53345 -11675 53355 -11555
rect 47855 -11720 53355 -11675
rect 47855 -11840 47865 -11720
rect 47985 -11840 48040 -11720
rect 48160 -11840 48205 -11720
rect 48325 -11840 48370 -11720
rect 48490 -11840 48535 -11720
rect 48655 -11840 48710 -11720
rect 48830 -11840 48875 -11720
rect 48995 -11840 49040 -11720
rect 49160 -11840 49205 -11720
rect 49325 -11840 49380 -11720
rect 49500 -11840 49545 -11720
rect 49665 -11840 49710 -11720
rect 49830 -11840 49875 -11720
rect 49995 -11840 50050 -11720
rect 50170 -11840 50215 -11720
rect 50335 -11840 50380 -11720
rect 50500 -11840 50545 -11720
rect 50665 -11840 50720 -11720
rect 50840 -11840 50885 -11720
rect 51005 -11840 51050 -11720
rect 51170 -11840 51215 -11720
rect 51335 -11840 51390 -11720
rect 51510 -11840 51555 -11720
rect 51675 -11840 51720 -11720
rect 51840 -11840 51885 -11720
rect 52005 -11840 52060 -11720
rect 52180 -11840 52225 -11720
rect 52345 -11840 52390 -11720
rect 52510 -11840 52555 -11720
rect 52675 -11840 52730 -11720
rect 52850 -11840 52895 -11720
rect 53015 -11840 53060 -11720
rect 53180 -11840 53225 -11720
rect 53345 -11840 53355 -11720
rect 47855 -11885 53355 -11840
rect 47855 -12005 47865 -11885
rect 47985 -12005 48040 -11885
rect 48160 -12005 48205 -11885
rect 48325 -12005 48370 -11885
rect 48490 -12005 48535 -11885
rect 48655 -12005 48710 -11885
rect 48830 -12005 48875 -11885
rect 48995 -12005 49040 -11885
rect 49160 -12005 49205 -11885
rect 49325 -12005 49380 -11885
rect 49500 -12005 49545 -11885
rect 49665 -12005 49710 -11885
rect 49830 -12005 49875 -11885
rect 49995 -12005 50050 -11885
rect 50170 -12005 50215 -11885
rect 50335 -12005 50380 -11885
rect 50500 -12005 50545 -11885
rect 50665 -12005 50720 -11885
rect 50840 -12005 50885 -11885
rect 51005 -12005 51050 -11885
rect 51170 -12005 51215 -11885
rect 51335 -12005 51390 -11885
rect 51510 -12005 51555 -11885
rect 51675 -12005 51720 -11885
rect 51840 -12005 51885 -11885
rect 52005 -12005 52060 -11885
rect 52180 -12005 52225 -11885
rect 52345 -12005 52390 -11885
rect 52510 -12005 52555 -11885
rect 52675 -12005 52730 -11885
rect 52850 -12005 52895 -11885
rect 53015 -12005 53060 -11885
rect 53180 -12005 53225 -11885
rect 53345 -12005 53355 -11885
rect 47855 -12060 53355 -12005
rect 47855 -12180 47865 -12060
rect 47985 -12180 48040 -12060
rect 48160 -12180 48205 -12060
rect 48325 -12180 48370 -12060
rect 48490 -12180 48535 -12060
rect 48655 -12180 48710 -12060
rect 48830 -12180 48875 -12060
rect 48995 -12180 49040 -12060
rect 49160 -12180 49205 -12060
rect 49325 -12180 49380 -12060
rect 49500 -12180 49545 -12060
rect 49665 -12180 49710 -12060
rect 49830 -12180 49875 -12060
rect 49995 -12180 50050 -12060
rect 50170 -12180 50215 -12060
rect 50335 -12180 50380 -12060
rect 50500 -12180 50545 -12060
rect 50665 -12180 50720 -12060
rect 50840 -12180 50885 -12060
rect 51005 -12180 51050 -12060
rect 51170 -12180 51215 -12060
rect 51335 -12180 51390 -12060
rect 51510 -12180 51555 -12060
rect 51675 -12180 51720 -12060
rect 51840 -12180 51885 -12060
rect 52005 -12180 52060 -12060
rect 52180 -12180 52225 -12060
rect 52345 -12180 52390 -12060
rect 52510 -12180 52555 -12060
rect 52675 -12180 52730 -12060
rect 52850 -12180 52895 -12060
rect 53015 -12180 53060 -12060
rect 53180 -12180 53225 -12060
rect 53345 -12180 53355 -12060
rect 47855 -12225 53355 -12180
rect 47855 -12345 47865 -12225
rect 47985 -12345 48040 -12225
rect 48160 -12345 48205 -12225
rect 48325 -12345 48370 -12225
rect 48490 -12345 48535 -12225
rect 48655 -12345 48710 -12225
rect 48830 -12345 48875 -12225
rect 48995 -12345 49040 -12225
rect 49160 -12345 49205 -12225
rect 49325 -12345 49380 -12225
rect 49500 -12345 49545 -12225
rect 49665 -12345 49710 -12225
rect 49830 -12345 49875 -12225
rect 49995 -12345 50050 -12225
rect 50170 -12345 50215 -12225
rect 50335 -12345 50380 -12225
rect 50500 -12345 50545 -12225
rect 50665 -12345 50720 -12225
rect 50840 -12345 50885 -12225
rect 51005 -12345 51050 -12225
rect 51170 -12345 51215 -12225
rect 51335 -12345 51390 -12225
rect 51510 -12345 51555 -12225
rect 51675 -12345 51720 -12225
rect 51840 -12345 51885 -12225
rect 52005 -12345 52060 -12225
rect 52180 -12345 52225 -12225
rect 52345 -12345 52390 -12225
rect 52510 -12345 52555 -12225
rect 52675 -12345 52730 -12225
rect 52850 -12345 52895 -12225
rect 53015 -12345 53060 -12225
rect 53180 -12345 53225 -12225
rect 53345 -12345 53355 -12225
rect 47855 -12390 53355 -12345
rect 47855 -12510 47865 -12390
rect 47985 -12510 48040 -12390
rect 48160 -12510 48205 -12390
rect 48325 -12510 48370 -12390
rect 48490 -12510 48535 -12390
rect 48655 -12510 48710 -12390
rect 48830 -12510 48875 -12390
rect 48995 -12510 49040 -12390
rect 49160 -12510 49205 -12390
rect 49325 -12510 49380 -12390
rect 49500 -12510 49545 -12390
rect 49665 -12510 49710 -12390
rect 49830 -12510 49875 -12390
rect 49995 -12510 50050 -12390
rect 50170 -12510 50215 -12390
rect 50335 -12510 50380 -12390
rect 50500 -12510 50545 -12390
rect 50665 -12510 50720 -12390
rect 50840 -12510 50885 -12390
rect 51005 -12510 51050 -12390
rect 51170 -12510 51215 -12390
rect 51335 -12510 51390 -12390
rect 51510 -12510 51555 -12390
rect 51675 -12510 51720 -12390
rect 51840 -12510 51885 -12390
rect 52005 -12510 52060 -12390
rect 52180 -12510 52225 -12390
rect 52345 -12510 52390 -12390
rect 52510 -12510 52555 -12390
rect 52675 -12510 52730 -12390
rect 52850 -12510 52895 -12390
rect 53015 -12510 53060 -12390
rect 53180 -12510 53225 -12390
rect 53345 -12510 53355 -12390
rect 47855 -12555 53355 -12510
rect 47855 -12675 47865 -12555
rect 47985 -12675 48040 -12555
rect 48160 -12675 48205 -12555
rect 48325 -12675 48370 -12555
rect 48490 -12675 48535 -12555
rect 48655 -12675 48710 -12555
rect 48830 -12675 48875 -12555
rect 48995 -12675 49040 -12555
rect 49160 -12675 49205 -12555
rect 49325 -12675 49380 -12555
rect 49500 -12675 49545 -12555
rect 49665 -12675 49710 -12555
rect 49830 -12675 49875 -12555
rect 49995 -12675 50050 -12555
rect 50170 -12675 50215 -12555
rect 50335 -12675 50380 -12555
rect 50500 -12675 50545 -12555
rect 50665 -12675 50720 -12555
rect 50840 -12675 50885 -12555
rect 51005 -12675 51050 -12555
rect 51170 -12675 51215 -12555
rect 51335 -12675 51390 -12555
rect 51510 -12675 51555 -12555
rect 51675 -12675 51720 -12555
rect 51840 -12675 51885 -12555
rect 52005 -12675 52060 -12555
rect 52180 -12675 52225 -12555
rect 52345 -12675 52390 -12555
rect 52510 -12675 52555 -12555
rect 52675 -12675 52730 -12555
rect 52850 -12675 52895 -12555
rect 53015 -12675 53060 -12555
rect 53180 -12675 53225 -12555
rect 53345 -12675 53355 -12555
rect 47855 -12730 53355 -12675
rect 47855 -12850 47865 -12730
rect 47985 -12850 48040 -12730
rect 48160 -12850 48205 -12730
rect 48325 -12850 48370 -12730
rect 48490 -12850 48535 -12730
rect 48655 -12850 48710 -12730
rect 48830 -12850 48875 -12730
rect 48995 -12850 49040 -12730
rect 49160 -12850 49205 -12730
rect 49325 -12850 49380 -12730
rect 49500 -12850 49545 -12730
rect 49665 -12850 49710 -12730
rect 49830 -12850 49875 -12730
rect 49995 -12850 50050 -12730
rect 50170 -12850 50215 -12730
rect 50335 -12850 50380 -12730
rect 50500 -12850 50545 -12730
rect 50665 -12850 50720 -12730
rect 50840 -12850 50885 -12730
rect 51005 -12850 51050 -12730
rect 51170 -12850 51215 -12730
rect 51335 -12850 51390 -12730
rect 51510 -12850 51555 -12730
rect 51675 -12850 51720 -12730
rect 51840 -12850 51885 -12730
rect 52005 -12850 52060 -12730
rect 52180 -12850 52225 -12730
rect 52345 -12850 52390 -12730
rect 52510 -12850 52555 -12730
rect 52675 -12850 52730 -12730
rect 52850 -12850 52895 -12730
rect 53015 -12850 53060 -12730
rect 53180 -12850 53225 -12730
rect 53345 -12850 53355 -12730
rect 47855 -12895 53355 -12850
rect 47855 -13015 47865 -12895
rect 47985 -13015 48040 -12895
rect 48160 -13015 48205 -12895
rect 48325 -13015 48370 -12895
rect 48490 -13015 48535 -12895
rect 48655 -13015 48710 -12895
rect 48830 -13015 48875 -12895
rect 48995 -13015 49040 -12895
rect 49160 -13015 49205 -12895
rect 49325 -13015 49380 -12895
rect 49500 -13015 49545 -12895
rect 49665 -13015 49710 -12895
rect 49830 -13015 49875 -12895
rect 49995 -13015 50050 -12895
rect 50170 -13015 50215 -12895
rect 50335 -13015 50380 -12895
rect 50500 -13015 50545 -12895
rect 50665 -13015 50720 -12895
rect 50840 -13015 50885 -12895
rect 51005 -13015 51050 -12895
rect 51170 -13015 51215 -12895
rect 51335 -13015 51390 -12895
rect 51510 -13015 51555 -12895
rect 51675 -13015 51720 -12895
rect 51840 -13015 51885 -12895
rect 52005 -13015 52060 -12895
rect 52180 -13015 52225 -12895
rect 52345 -13015 52390 -12895
rect 52510 -13015 52555 -12895
rect 52675 -13015 52730 -12895
rect 52850 -13015 52895 -12895
rect 53015 -13015 53060 -12895
rect 53180 -13015 53225 -12895
rect 53345 -13015 53355 -12895
rect 47855 -13060 53355 -13015
rect 47855 -13180 47865 -13060
rect 47985 -13180 48040 -13060
rect 48160 -13180 48205 -13060
rect 48325 -13180 48370 -13060
rect 48490 -13180 48535 -13060
rect 48655 -13180 48710 -13060
rect 48830 -13180 48875 -13060
rect 48995 -13180 49040 -13060
rect 49160 -13180 49205 -13060
rect 49325 -13180 49380 -13060
rect 49500 -13180 49545 -13060
rect 49665 -13180 49710 -13060
rect 49830 -13180 49875 -13060
rect 49995 -13180 50050 -13060
rect 50170 -13180 50215 -13060
rect 50335 -13180 50380 -13060
rect 50500 -13180 50545 -13060
rect 50665 -13180 50720 -13060
rect 50840 -13180 50885 -13060
rect 51005 -13180 51050 -13060
rect 51170 -13180 51215 -13060
rect 51335 -13180 51390 -13060
rect 51510 -13180 51555 -13060
rect 51675 -13180 51720 -13060
rect 51840 -13180 51885 -13060
rect 52005 -13180 52060 -13060
rect 52180 -13180 52225 -13060
rect 52345 -13180 52390 -13060
rect 52510 -13180 52555 -13060
rect 52675 -13180 52730 -13060
rect 52850 -13180 52895 -13060
rect 53015 -13180 53060 -13060
rect 53180 -13180 53225 -13060
rect 53345 -13180 53355 -13060
rect 47855 -13225 53355 -13180
rect 47855 -13345 47865 -13225
rect 47985 -13345 48040 -13225
rect 48160 -13345 48205 -13225
rect 48325 -13345 48370 -13225
rect 48490 -13345 48535 -13225
rect 48655 -13345 48710 -13225
rect 48830 -13345 48875 -13225
rect 48995 -13345 49040 -13225
rect 49160 -13345 49205 -13225
rect 49325 -13345 49380 -13225
rect 49500 -13345 49545 -13225
rect 49665 -13345 49710 -13225
rect 49830 -13345 49875 -13225
rect 49995 -13345 50050 -13225
rect 50170 -13345 50215 -13225
rect 50335 -13345 50380 -13225
rect 50500 -13345 50545 -13225
rect 50665 -13345 50720 -13225
rect 50840 -13345 50885 -13225
rect 51005 -13345 51050 -13225
rect 51170 -13345 51215 -13225
rect 51335 -13345 51390 -13225
rect 51510 -13345 51555 -13225
rect 51675 -13345 51720 -13225
rect 51840 -13345 51885 -13225
rect 52005 -13345 52060 -13225
rect 52180 -13345 52225 -13225
rect 52345 -13345 52390 -13225
rect 52510 -13345 52555 -13225
rect 52675 -13345 52730 -13225
rect 52850 -13345 52895 -13225
rect 53015 -13345 53060 -13225
rect 53180 -13345 53225 -13225
rect 53345 -13345 53355 -13225
rect 47855 -13400 53355 -13345
rect 47855 -13520 47865 -13400
rect 47985 -13520 48040 -13400
rect 48160 -13520 48205 -13400
rect 48325 -13520 48370 -13400
rect 48490 -13520 48535 -13400
rect 48655 -13520 48710 -13400
rect 48830 -13520 48875 -13400
rect 48995 -13520 49040 -13400
rect 49160 -13520 49205 -13400
rect 49325 -13520 49380 -13400
rect 49500 -13520 49545 -13400
rect 49665 -13520 49710 -13400
rect 49830 -13520 49875 -13400
rect 49995 -13520 50050 -13400
rect 50170 -13520 50215 -13400
rect 50335 -13520 50380 -13400
rect 50500 -13520 50545 -13400
rect 50665 -13520 50720 -13400
rect 50840 -13520 50885 -13400
rect 51005 -13520 51050 -13400
rect 51170 -13520 51215 -13400
rect 51335 -13520 51390 -13400
rect 51510 -13520 51555 -13400
rect 51675 -13520 51720 -13400
rect 51840 -13520 51885 -13400
rect 52005 -13520 52060 -13400
rect 52180 -13520 52225 -13400
rect 52345 -13520 52390 -13400
rect 52510 -13520 52555 -13400
rect 52675 -13520 52730 -13400
rect 52850 -13520 52895 -13400
rect 53015 -13520 53060 -13400
rect 53180 -13520 53225 -13400
rect 53345 -13520 53355 -13400
rect 47855 -13565 53355 -13520
rect 47855 -13685 47865 -13565
rect 47985 -13685 48040 -13565
rect 48160 -13685 48205 -13565
rect 48325 -13685 48370 -13565
rect 48490 -13685 48535 -13565
rect 48655 -13685 48710 -13565
rect 48830 -13685 48875 -13565
rect 48995 -13685 49040 -13565
rect 49160 -13685 49205 -13565
rect 49325 -13685 49380 -13565
rect 49500 -13685 49545 -13565
rect 49665 -13685 49710 -13565
rect 49830 -13685 49875 -13565
rect 49995 -13685 50050 -13565
rect 50170 -13685 50215 -13565
rect 50335 -13685 50380 -13565
rect 50500 -13685 50545 -13565
rect 50665 -13685 50720 -13565
rect 50840 -13685 50885 -13565
rect 51005 -13685 51050 -13565
rect 51170 -13685 51215 -13565
rect 51335 -13685 51390 -13565
rect 51510 -13685 51555 -13565
rect 51675 -13685 51720 -13565
rect 51840 -13685 51885 -13565
rect 52005 -13685 52060 -13565
rect 52180 -13685 52225 -13565
rect 52345 -13685 52390 -13565
rect 52510 -13685 52555 -13565
rect 52675 -13685 52730 -13565
rect 52850 -13685 52895 -13565
rect 53015 -13685 53060 -13565
rect 53180 -13685 53225 -13565
rect 53345 -13685 53355 -13565
rect 47855 -13730 53355 -13685
rect 47855 -13850 47865 -13730
rect 47985 -13850 48040 -13730
rect 48160 -13850 48205 -13730
rect 48325 -13850 48370 -13730
rect 48490 -13850 48535 -13730
rect 48655 -13850 48710 -13730
rect 48830 -13850 48875 -13730
rect 48995 -13850 49040 -13730
rect 49160 -13850 49205 -13730
rect 49325 -13850 49380 -13730
rect 49500 -13850 49545 -13730
rect 49665 -13850 49710 -13730
rect 49830 -13850 49875 -13730
rect 49995 -13850 50050 -13730
rect 50170 -13850 50215 -13730
rect 50335 -13850 50380 -13730
rect 50500 -13850 50545 -13730
rect 50665 -13850 50720 -13730
rect 50840 -13850 50885 -13730
rect 51005 -13850 51050 -13730
rect 51170 -13850 51215 -13730
rect 51335 -13850 51390 -13730
rect 51510 -13850 51555 -13730
rect 51675 -13850 51720 -13730
rect 51840 -13850 51885 -13730
rect 52005 -13850 52060 -13730
rect 52180 -13850 52225 -13730
rect 52345 -13850 52390 -13730
rect 52510 -13850 52555 -13730
rect 52675 -13850 52730 -13730
rect 52850 -13850 52895 -13730
rect 53015 -13850 53060 -13730
rect 53180 -13850 53225 -13730
rect 53345 -13850 53355 -13730
rect 47855 -13895 53355 -13850
rect 47855 -14015 47865 -13895
rect 47985 -14015 48040 -13895
rect 48160 -14015 48205 -13895
rect 48325 -14015 48370 -13895
rect 48490 -14015 48535 -13895
rect 48655 -14015 48710 -13895
rect 48830 -14015 48875 -13895
rect 48995 -14015 49040 -13895
rect 49160 -14015 49205 -13895
rect 49325 -14015 49380 -13895
rect 49500 -14015 49545 -13895
rect 49665 -14015 49710 -13895
rect 49830 -14015 49875 -13895
rect 49995 -14015 50050 -13895
rect 50170 -14015 50215 -13895
rect 50335 -14015 50380 -13895
rect 50500 -14015 50545 -13895
rect 50665 -14015 50720 -13895
rect 50840 -14015 50885 -13895
rect 51005 -14015 51050 -13895
rect 51170 -14015 51215 -13895
rect 51335 -14015 51390 -13895
rect 51510 -14015 51555 -13895
rect 51675 -14015 51720 -13895
rect 51840 -14015 51885 -13895
rect 52005 -14015 52060 -13895
rect 52180 -14015 52225 -13895
rect 52345 -14015 52390 -13895
rect 52510 -14015 52555 -13895
rect 52675 -14015 52730 -13895
rect 52850 -14015 52895 -13895
rect 53015 -14015 53060 -13895
rect 53180 -14015 53225 -13895
rect 53345 -14015 53355 -13895
rect 47855 -14070 53355 -14015
rect 47855 -14190 47865 -14070
rect 47985 -14190 48040 -14070
rect 48160 -14190 48205 -14070
rect 48325 -14190 48370 -14070
rect 48490 -14190 48535 -14070
rect 48655 -14190 48710 -14070
rect 48830 -14190 48875 -14070
rect 48995 -14190 49040 -14070
rect 49160 -14190 49205 -14070
rect 49325 -14190 49380 -14070
rect 49500 -14190 49545 -14070
rect 49665 -14190 49710 -14070
rect 49830 -14190 49875 -14070
rect 49995 -14190 50050 -14070
rect 50170 -14190 50215 -14070
rect 50335 -14190 50380 -14070
rect 50500 -14190 50545 -14070
rect 50665 -14190 50720 -14070
rect 50840 -14190 50885 -14070
rect 51005 -14190 51050 -14070
rect 51170 -14190 51215 -14070
rect 51335 -14190 51390 -14070
rect 51510 -14190 51555 -14070
rect 51675 -14190 51720 -14070
rect 51840 -14190 51885 -14070
rect 52005 -14190 52060 -14070
rect 52180 -14190 52225 -14070
rect 52345 -14190 52390 -14070
rect 52510 -14190 52555 -14070
rect 52675 -14190 52730 -14070
rect 52850 -14190 52895 -14070
rect 53015 -14190 53060 -14070
rect 53180 -14190 53225 -14070
rect 53345 -14190 53355 -14070
rect 47855 -14235 53355 -14190
rect 47855 -14355 47865 -14235
rect 47985 -14355 48040 -14235
rect 48160 -14355 48205 -14235
rect 48325 -14355 48370 -14235
rect 48490 -14355 48535 -14235
rect 48655 -14355 48710 -14235
rect 48830 -14355 48875 -14235
rect 48995 -14355 49040 -14235
rect 49160 -14355 49205 -14235
rect 49325 -14355 49380 -14235
rect 49500 -14355 49545 -14235
rect 49665 -14355 49710 -14235
rect 49830 -14355 49875 -14235
rect 49995 -14355 50050 -14235
rect 50170 -14355 50215 -14235
rect 50335 -14355 50380 -14235
rect 50500 -14355 50545 -14235
rect 50665 -14355 50720 -14235
rect 50840 -14355 50885 -14235
rect 51005 -14355 51050 -14235
rect 51170 -14355 51215 -14235
rect 51335 -14355 51390 -14235
rect 51510 -14355 51555 -14235
rect 51675 -14355 51720 -14235
rect 51840 -14355 51885 -14235
rect 52005 -14355 52060 -14235
rect 52180 -14355 52225 -14235
rect 52345 -14355 52390 -14235
rect 52510 -14355 52555 -14235
rect 52675 -14355 52730 -14235
rect 52850 -14355 52895 -14235
rect 53015 -14355 53060 -14235
rect 53180 -14355 53225 -14235
rect 53345 -14355 53355 -14235
rect 47855 -14400 53355 -14355
rect 47855 -14520 47865 -14400
rect 47985 -14520 48040 -14400
rect 48160 -14520 48205 -14400
rect 48325 -14520 48370 -14400
rect 48490 -14520 48535 -14400
rect 48655 -14520 48710 -14400
rect 48830 -14520 48875 -14400
rect 48995 -14520 49040 -14400
rect 49160 -14520 49205 -14400
rect 49325 -14520 49380 -14400
rect 49500 -14520 49545 -14400
rect 49665 -14520 49710 -14400
rect 49830 -14520 49875 -14400
rect 49995 -14520 50050 -14400
rect 50170 -14520 50215 -14400
rect 50335 -14520 50380 -14400
rect 50500 -14520 50545 -14400
rect 50665 -14520 50720 -14400
rect 50840 -14520 50885 -14400
rect 51005 -14520 51050 -14400
rect 51170 -14520 51215 -14400
rect 51335 -14520 51390 -14400
rect 51510 -14520 51555 -14400
rect 51675 -14520 51720 -14400
rect 51840 -14520 51885 -14400
rect 52005 -14520 52060 -14400
rect 52180 -14520 52225 -14400
rect 52345 -14520 52390 -14400
rect 52510 -14520 52555 -14400
rect 52675 -14520 52730 -14400
rect 52850 -14520 52895 -14400
rect 53015 -14520 53060 -14400
rect 53180 -14520 53225 -14400
rect 53345 -14520 53355 -14400
rect 47855 -14565 53355 -14520
rect 47855 -14685 47865 -14565
rect 47985 -14685 48040 -14565
rect 48160 -14685 48205 -14565
rect 48325 -14685 48370 -14565
rect 48490 -14685 48535 -14565
rect 48655 -14685 48710 -14565
rect 48830 -14685 48875 -14565
rect 48995 -14685 49040 -14565
rect 49160 -14685 49205 -14565
rect 49325 -14685 49380 -14565
rect 49500 -14685 49545 -14565
rect 49665 -14685 49710 -14565
rect 49830 -14685 49875 -14565
rect 49995 -14685 50050 -14565
rect 50170 -14685 50215 -14565
rect 50335 -14685 50380 -14565
rect 50500 -14685 50545 -14565
rect 50665 -14685 50720 -14565
rect 50840 -14685 50885 -14565
rect 51005 -14685 51050 -14565
rect 51170 -14685 51215 -14565
rect 51335 -14685 51390 -14565
rect 51510 -14685 51555 -14565
rect 51675 -14685 51720 -14565
rect 51840 -14685 51885 -14565
rect 52005 -14685 52060 -14565
rect 52180 -14685 52225 -14565
rect 52345 -14685 52390 -14565
rect 52510 -14685 52555 -14565
rect 52675 -14685 52730 -14565
rect 52850 -14685 52895 -14565
rect 53015 -14685 53060 -14565
rect 53180 -14685 53225 -14565
rect 53345 -14685 53355 -14565
rect 47855 -14740 53355 -14685
rect 47855 -14860 47865 -14740
rect 47985 -14860 48040 -14740
rect 48160 -14860 48205 -14740
rect 48325 -14860 48370 -14740
rect 48490 -14860 48535 -14740
rect 48655 -14860 48710 -14740
rect 48830 -14860 48875 -14740
rect 48995 -14860 49040 -14740
rect 49160 -14860 49205 -14740
rect 49325 -14860 49380 -14740
rect 49500 -14860 49545 -14740
rect 49665 -14860 49710 -14740
rect 49830 -14860 49875 -14740
rect 49995 -14860 50050 -14740
rect 50170 -14860 50215 -14740
rect 50335 -14860 50380 -14740
rect 50500 -14860 50545 -14740
rect 50665 -14860 50720 -14740
rect 50840 -14860 50885 -14740
rect 51005 -14860 51050 -14740
rect 51170 -14860 51215 -14740
rect 51335 -14860 51390 -14740
rect 51510 -14860 51555 -14740
rect 51675 -14860 51720 -14740
rect 51840 -14860 51885 -14740
rect 52005 -14860 52060 -14740
rect 52180 -14860 52225 -14740
rect 52345 -14860 52390 -14740
rect 52510 -14860 52555 -14740
rect 52675 -14860 52730 -14740
rect 52850 -14860 52895 -14740
rect 53015 -14860 53060 -14740
rect 53180 -14860 53225 -14740
rect 53345 -14860 53355 -14740
rect 47855 -14905 53355 -14860
rect 47855 -15025 47865 -14905
rect 47985 -15025 48040 -14905
rect 48160 -15025 48205 -14905
rect 48325 -15025 48370 -14905
rect 48490 -15025 48535 -14905
rect 48655 -15025 48710 -14905
rect 48830 -15025 48875 -14905
rect 48995 -15025 49040 -14905
rect 49160 -15025 49205 -14905
rect 49325 -15025 49380 -14905
rect 49500 -15025 49545 -14905
rect 49665 -15025 49710 -14905
rect 49830 -15025 49875 -14905
rect 49995 -15025 50050 -14905
rect 50170 -15025 50215 -14905
rect 50335 -15025 50380 -14905
rect 50500 -15025 50545 -14905
rect 50665 -15025 50720 -14905
rect 50840 -15025 50885 -14905
rect 51005 -15025 51050 -14905
rect 51170 -15025 51215 -14905
rect 51335 -15025 51390 -14905
rect 51510 -15025 51555 -14905
rect 51675 -15025 51720 -14905
rect 51840 -15025 51885 -14905
rect 52005 -15025 52060 -14905
rect 52180 -15025 52225 -14905
rect 52345 -15025 52390 -14905
rect 52510 -15025 52555 -14905
rect 52675 -15025 52730 -14905
rect 52850 -15025 52895 -14905
rect 53015 -15025 53060 -14905
rect 53180 -15025 53225 -14905
rect 53345 -15025 53355 -14905
rect 47855 -15070 53355 -15025
rect 47855 -15190 47865 -15070
rect 47985 -15190 48040 -15070
rect 48160 -15190 48205 -15070
rect 48325 -15190 48370 -15070
rect 48490 -15190 48535 -15070
rect 48655 -15190 48710 -15070
rect 48830 -15190 48875 -15070
rect 48995 -15190 49040 -15070
rect 49160 -15190 49205 -15070
rect 49325 -15190 49380 -15070
rect 49500 -15190 49545 -15070
rect 49665 -15190 49710 -15070
rect 49830 -15190 49875 -15070
rect 49995 -15190 50050 -15070
rect 50170 -15190 50215 -15070
rect 50335 -15190 50380 -15070
rect 50500 -15190 50545 -15070
rect 50665 -15190 50720 -15070
rect 50840 -15190 50885 -15070
rect 51005 -15190 51050 -15070
rect 51170 -15190 51215 -15070
rect 51335 -15190 51390 -15070
rect 51510 -15190 51555 -15070
rect 51675 -15190 51720 -15070
rect 51840 -15190 51885 -15070
rect 52005 -15190 52060 -15070
rect 52180 -15190 52225 -15070
rect 52345 -15190 52390 -15070
rect 52510 -15190 52555 -15070
rect 52675 -15190 52730 -15070
rect 52850 -15190 52895 -15070
rect 53015 -15190 53060 -15070
rect 53180 -15190 53225 -15070
rect 53345 -15190 53355 -15070
rect 47855 -15235 53355 -15190
rect 47855 -15355 47865 -15235
rect 47985 -15355 48040 -15235
rect 48160 -15355 48205 -15235
rect 48325 -15355 48370 -15235
rect 48490 -15355 48535 -15235
rect 48655 -15355 48710 -15235
rect 48830 -15355 48875 -15235
rect 48995 -15355 49040 -15235
rect 49160 -15355 49205 -15235
rect 49325 -15355 49380 -15235
rect 49500 -15355 49545 -15235
rect 49665 -15355 49710 -15235
rect 49830 -15355 49875 -15235
rect 49995 -15355 50050 -15235
rect 50170 -15355 50215 -15235
rect 50335 -15355 50380 -15235
rect 50500 -15355 50545 -15235
rect 50665 -15355 50720 -15235
rect 50840 -15355 50885 -15235
rect 51005 -15355 51050 -15235
rect 51170 -15355 51215 -15235
rect 51335 -15355 51390 -15235
rect 51510 -15355 51555 -15235
rect 51675 -15355 51720 -15235
rect 51840 -15355 51885 -15235
rect 52005 -15355 52060 -15235
rect 52180 -15355 52225 -15235
rect 52345 -15355 52390 -15235
rect 52510 -15355 52555 -15235
rect 52675 -15355 52730 -15235
rect 52850 -15355 52895 -15235
rect 53015 -15355 53060 -15235
rect 53180 -15355 53225 -15235
rect 53345 -15355 53355 -15235
rect 47855 -15410 53355 -15355
rect 47855 -15530 47865 -15410
rect 47985 -15530 48040 -15410
rect 48160 -15530 48205 -15410
rect 48325 -15530 48370 -15410
rect 48490 -15530 48535 -15410
rect 48655 -15530 48710 -15410
rect 48830 -15530 48875 -15410
rect 48995 -15530 49040 -15410
rect 49160 -15530 49205 -15410
rect 49325 -15530 49380 -15410
rect 49500 -15530 49545 -15410
rect 49665 -15530 49710 -15410
rect 49830 -15530 49875 -15410
rect 49995 -15530 50050 -15410
rect 50170 -15530 50215 -15410
rect 50335 -15530 50380 -15410
rect 50500 -15530 50545 -15410
rect 50665 -15530 50720 -15410
rect 50840 -15530 50885 -15410
rect 51005 -15530 51050 -15410
rect 51170 -15530 51215 -15410
rect 51335 -15530 51390 -15410
rect 51510 -15530 51555 -15410
rect 51675 -15530 51720 -15410
rect 51840 -15530 51885 -15410
rect 52005 -15530 52060 -15410
rect 52180 -15530 52225 -15410
rect 52345 -15530 52390 -15410
rect 52510 -15530 52555 -15410
rect 52675 -15530 52730 -15410
rect 52850 -15530 52895 -15410
rect 53015 -15530 53060 -15410
rect 53180 -15530 53225 -15410
rect 53345 -15530 53355 -15410
rect 47855 -15540 53355 -15530
<< mimcapcontact >>
rect 30795 7080 30915 7200
rect 30960 7080 31080 7200
rect 31125 7080 31245 7200
rect 31290 7080 31410 7200
rect 31465 7080 31585 7200
rect 31630 7080 31750 7200
rect 31795 7080 31915 7200
rect 31960 7080 32080 7200
rect 32135 7080 32255 7200
rect 32300 7080 32420 7200
rect 32465 7080 32585 7200
rect 32630 7080 32750 7200
rect 32805 7080 32925 7200
rect 32970 7080 33090 7200
rect 33135 7080 33255 7200
rect 33300 7080 33420 7200
rect 33475 7080 33595 7200
rect 33640 7080 33760 7200
rect 33805 7080 33925 7200
rect 33970 7080 34090 7200
rect 34145 7080 34265 7200
rect 34310 7080 34430 7200
rect 34475 7080 34595 7200
rect 34640 7080 34760 7200
rect 34815 7080 34935 7200
rect 34980 7080 35100 7200
rect 35145 7080 35265 7200
rect 35310 7080 35430 7200
rect 35485 7080 35605 7200
rect 35650 7080 35770 7200
rect 35815 7080 35935 7200
rect 35980 7080 36100 7200
rect 36155 7080 36275 7200
rect 30795 6905 30915 7025
rect 30960 6905 31080 7025
rect 31125 6905 31245 7025
rect 31290 6905 31410 7025
rect 31465 6905 31585 7025
rect 31630 6905 31750 7025
rect 31795 6905 31915 7025
rect 31960 6905 32080 7025
rect 32135 6905 32255 7025
rect 32300 6905 32420 7025
rect 32465 6905 32585 7025
rect 32630 6905 32750 7025
rect 32805 6905 32925 7025
rect 32970 6905 33090 7025
rect 33135 6905 33255 7025
rect 33300 6905 33420 7025
rect 33475 6905 33595 7025
rect 33640 6905 33760 7025
rect 33805 6905 33925 7025
rect 33970 6905 34090 7025
rect 34145 6905 34265 7025
rect 34310 6905 34430 7025
rect 34475 6905 34595 7025
rect 34640 6905 34760 7025
rect 34815 6905 34935 7025
rect 34980 6905 35100 7025
rect 35145 6905 35265 7025
rect 35310 6905 35430 7025
rect 35485 6905 35605 7025
rect 35650 6905 35770 7025
rect 35815 6905 35935 7025
rect 35980 6905 36100 7025
rect 36155 6905 36275 7025
rect 30795 6740 30915 6860
rect 30960 6740 31080 6860
rect 31125 6740 31245 6860
rect 31290 6740 31410 6860
rect 31465 6740 31585 6860
rect 31630 6740 31750 6860
rect 31795 6740 31915 6860
rect 31960 6740 32080 6860
rect 32135 6740 32255 6860
rect 32300 6740 32420 6860
rect 32465 6740 32585 6860
rect 32630 6740 32750 6860
rect 32805 6740 32925 6860
rect 32970 6740 33090 6860
rect 33135 6740 33255 6860
rect 33300 6740 33420 6860
rect 33475 6740 33595 6860
rect 33640 6740 33760 6860
rect 33805 6740 33925 6860
rect 33970 6740 34090 6860
rect 34145 6740 34265 6860
rect 34310 6740 34430 6860
rect 34475 6740 34595 6860
rect 34640 6740 34760 6860
rect 34815 6740 34935 6860
rect 34980 6740 35100 6860
rect 35145 6740 35265 6860
rect 35310 6740 35430 6860
rect 35485 6740 35605 6860
rect 35650 6740 35770 6860
rect 35815 6740 35935 6860
rect 35980 6740 36100 6860
rect 36155 6740 36275 6860
rect 30795 6575 30915 6695
rect 30960 6575 31080 6695
rect 31125 6575 31245 6695
rect 31290 6575 31410 6695
rect 31465 6575 31585 6695
rect 31630 6575 31750 6695
rect 31795 6575 31915 6695
rect 31960 6575 32080 6695
rect 32135 6575 32255 6695
rect 32300 6575 32420 6695
rect 32465 6575 32585 6695
rect 32630 6575 32750 6695
rect 32805 6575 32925 6695
rect 32970 6575 33090 6695
rect 33135 6575 33255 6695
rect 33300 6575 33420 6695
rect 33475 6575 33595 6695
rect 33640 6575 33760 6695
rect 33805 6575 33925 6695
rect 33970 6575 34090 6695
rect 34145 6575 34265 6695
rect 34310 6575 34430 6695
rect 34475 6575 34595 6695
rect 34640 6575 34760 6695
rect 34815 6575 34935 6695
rect 34980 6575 35100 6695
rect 35145 6575 35265 6695
rect 35310 6575 35430 6695
rect 35485 6575 35605 6695
rect 35650 6575 35770 6695
rect 35815 6575 35935 6695
rect 35980 6575 36100 6695
rect 36155 6575 36275 6695
rect 30795 6410 30915 6530
rect 30960 6410 31080 6530
rect 31125 6410 31245 6530
rect 31290 6410 31410 6530
rect 31465 6410 31585 6530
rect 31630 6410 31750 6530
rect 31795 6410 31915 6530
rect 31960 6410 32080 6530
rect 32135 6410 32255 6530
rect 32300 6410 32420 6530
rect 32465 6410 32585 6530
rect 32630 6410 32750 6530
rect 32805 6410 32925 6530
rect 32970 6410 33090 6530
rect 33135 6410 33255 6530
rect 33300 6410 33420 6530
rect 33475 6410 33595 6530
rect 33640 6410 33760 6530
rect 33805 6410 33925 6530
rect 33970 6410 34090 6530
rect 34145 6410 34265 6530
rect 34310 6410 34430 6530
rect 34475 6410 34595 6530
rect 34640 6410 34760 6530
rect 34815 6410 34935 6530
rect 34980 6410 35100 6530
rect 35145 6410 35265 6530
rect 35310 6410 35430 6530
rect 35485 6410 35605 6530
rect 35650 6410 35770 6530
rect 35815 6410 35935 6530
rect 35980 6410 36100 6530
rect 36155 6410 36275 6530
rect 30795 6235 30915 6355
rect 30960 6235 31080 6355
rect 31125 6235 31245 6355
rect 31290 6235 31410 6355
rect 31465 6235 31585 6355
rect 31630 6235 31750 6355
rect 31795 6235 31915 6355
rect 31960 6235 32080 6355
rect 32135 6235 32255 6355
rect 32300 6235 32420 6355
rect 32465 6235 32585 6355
rect 32630 6235 32750 6355
rect 32805 6235 32925 6355
rect 32970 6235 33090 6355
rect 33135 6235 33255 6355
rect 33300 6235 33420 6355
rect 33475 6235 33595 6355
rect 33640 6235 33760 6355
rect 33805 6235 33925 6355
rect 33970 6235 34090 6355
rect 34145 6235 34265 6355
rect 34310 6235 34430 6355
rect 34475 6235 34595 6355
rect 34640 6235 34760 6355
rect 34815 6235 34935 6355
rect 34980 6235 35100 6355
rect 35145 6235 35265 6355
rect 35310 6235 35430 6355
rect 35485 6235 35605 6355
rect 35650 6235 35770 6355
rect 35815 6235 35935 6355
rect 35980 6235 36100 6355
rect 36155 6235 36275 6355
rect 30795 6070 30915 6190
rect 30960 6070 31080 6190
rect 31125 6070 31245 6190
rect 31290 6070 31410 6190
rect 31465 6070 31585 6190
rect 31630 6070 31750 6190
rect 31795 6070 31915 6190
rect 31960 6070 32080 6190
rect 32135 6070 32255 6190
rect 32300 6070 32420 6190
rect 32465 6070 32585 6190
rect 32630 6070 32750 6190
rect 32805 6070 32925 6190
rect 32970 6070 33090 6190
rect 33135 6070 33255 6190
rect 33300 6070 33420 6190
rect 33475 6070 33595 6190
rect 33640 6070 33760 6190
rect 33805 6070 33925 6190
rect 33970 6070 34090 6190
rect 34145 6070 34265 6190
rect 34310 6070 34430 6190
rect 34475 6070 34595 6190
rect 34640 6070 34760 6190
rect 34815 6070 34935 6190
rect 34980 6070 35100 6190
rect 35145 6070 35265 6190
rect 35310 6070 35430 6190
rect 35485 6070 35605 6190
rect 35650 6070 35770 6190
rect 35815 6070 35935 6190
rect 35980 6070 36100 6190
rect 36155 6070 36275 6190
rect 30795 5905 30915 6025
rect 30960 5905 31080 6025
rect 31125 5905 31245 6025
rect 31290 5905 31410 6025
rect 31465 5905 31585 6025
rect 31630 5905 31750 6025
rect 31795 5905 31915 6025
rect 31960 5905 32080 6025
rect 32135 5905 32255 6025
rect 32300 5905 32420 6025
rect 32465 5905 32585 6025
rect 32630 5905 32750 6025
rect 32805 5905 32925 6025
rect 32970 5905 33090 6025
rect 33135 5905 33255 6025
rect 33300 5905 33420 6025
rect 33475 5905 33595 6025
rect 33640 5905 33760 6025
rect 33805 5905 33925 6025
rect 33970 5905 34090 6025
rect 34145 5905 34265 6025
rect 34310 5905 34430 6025
rect 34475 5905 34595 6025
rect 34640 5905 34760 6025
rect 34815 5905 34935 6025
rect 34980 5905 35100 6025
rect 35145 5905 35265 6025
rect 35310 5905 35430 6025
rect 35485 5905 35605 6025
rect 35650 5905 35770 6025
rect 35815 5905 35935 6025
rect 35980 5905 36100 6025
rect 36155 5905 36275 6025
rect 30795 5740 30915 5860
rect 30960 5740 31080 5860
rect 31125 5740 31245 5860
rect 31290 5740 31410 5860
rect 31465 5740 31585 5860
rect 31630 5740 31750 5860
rect 31795 5740 31915 5860
rect 31960 5740 32080 5860
rect 32135 5740 32255 5860
rect 32300 5740 32420 5860
rect 32465 5740 32585 5860
rect 32630 5740 32750 5860
rect 32805 5740 32925 5860
rect 32970 5740 33090 5860
rect 33135 5740 33255 5860
rect 33300 5740 33420 5860
rect 33475 5740 33595 5860
rect 33640 5740 33760 5860
rect 33805 5740 33925 5860
rect 33970 5740 34090 5860
rect 34145 5740 34265 5860
rect 34310 5740 34430 5860
rect 34475 5740 34595 5860
rect 34640 5740 34760 5860
rect 34815 5740 34935 5860
rect 34980 5740 35100 5860
rect 35145 5740 35265 5860
rect 35310 5740 35430 5860
rect 35485 5740 35605 5860
rect 35650 5740 35770 5860
rect 35815 5740 35935 5860
rect 35980 5740 36100 5860
rect 36155 5740 36275 5860
rect 30795 5565 30915 5685
rect 30960 5565 31080 5685
rect 31125 5565 31245 5685
rect 31290 5565 31410 5685
rect 31465 5565 31585 5685
rect 31630 5565 31750 5685
rect 31795 5565 31915 5685
rect 31960 5565 32080 5685
rect 32135 5565 32255 5685
rect 32300 5565 32420 5685
rect 32465 5565 32585 5685
rect 32630 5565 32750 5685
rect 32805 5565 32925 5685
rect 32970 5565 33090 5685
rect 33135 5565 33255 5685
rect 33300 5565 33420 5685
rect 33475 5565 33595 5685
rect 33640 5565 33760 5685
rect 33805 5565 33925 5685
rect 33970 5565 34090 5685
rect 34145 5565 34265 5685
rect 34310 5565 34430 5685
rect 34475 5565 34595 5685
rect 34640 5565 34760 5685
rect 34815 5565 34935 5685
rect 34980 5565 35100 5685
rect 35145 5565 35265 5685
rect 35310 5565 35430 5685
rect 35485 5565 35605 5685
rect 35650 5565 35770 5685
rect 35815 5565 35935 5685
rect 35980 5565 36100 5685
rect 36155 5565 36275 5685
rect 30795 5400 30915 5520
rect 30960 5400 31080 5520
rect 31125 5400 31245 5520
rect 31290 5400 31410 5520
rect 31465 5400 31585 5520
rect 31630 5400 31750 5520
rect 31795 5400 31915 5520
rect 31960 5400 32080 5520
rect 32135 5400 32255 5520
rect 32300 5400 32420 5520
rect 32465 5400 32585 5520
rect 32630 5400 32750 5520
rect 32805 5400 32925 5520
rect 32970 5400 33090 5520
rect 33135 5400 33255 5520
rect 33300 5400 33420 5520
rect 33475 5400 33595 5520
rect 33640 5400 33760 5520
rect 33805 5400 33925 5520
rect 33970 5400 34090 5520
rect 34145 5400 34265 5520
rect 34310 5400 34430 5520
rect 34475 5400 34595 5520
rect 34640 5400 34760 5520
rect 34815 5400 34935 5520
rect 34980 5400 35100 5520
rect 35145 5400 35265 5520
rect 35310 5400 35430 5520
rect 35485 5400 35605 5520
rect 35650 5400 35770 5520
rect 35815 5400 35935 5520
rect 35980 5400 36100 5520
rect 36155 5400 36275 5520
rect 30795 5235 30915 5355
rect 30960 5235 31080 5355
rect 31125 5235 31245 5355
rect 31290 5235 31410 5355
rect 31465 5235 31585 5355
rect 31630 5235 31750 5355
rect 31795 5235 31915 5355
rect 31960 5235 32080 5355
rect 32135 5235 32255 5355
rect 32300 5235 32420 5355
rect 32465 5235 32585 5355
rect 32630 5235 32750 5355
rect 32805 5235 32925 5355
rect 32970 5235 33090 5355
rect 33135 5235 33255 5355
rect 33300 5235 33420 5355
rect 33475 5235 33595 5355
rect 33640 5235 33760 5355
rect 33805 5235 33925 5355
rect 33970 5235 34090 5355
rect 34145 5235 34265 5355
rect 34310 5235 34430 5355
rect 34475 5235 34595 5355
rect 34640 5235 34760 5355
rect 34815 5235 34935 5355
rect 34980 5235 35100 5355
rect 35145 5235 35265 5355
rect 35310 5235 35430 5355
rect 35485 5235 35605 5355
rect 35650 5235 35770 5355
rect 35815 5235 35935 5355
rect 35980 5235 36100 5355
rect 36155 5235 36275 5355
rect 30795 5070 30915 5190
rect 30960 5070 31080 5190
rect 31125 5070 31245 5190
rect 31290 5070 31410 5190
rect 31465 5070 31585 5190
rect 31630 5070 31750 5190
rect 31795 5070 31915 5190
rect 31960 5070 32080 5190
rect 32135 5070 32255 5190
rect 32300 5070 32420 5190
rect 32465 5070 32585 5190
rect 32630 5070 32750 5190
rect 32805 5070 32925 5190
rect 32970 5070 33090 5190
rect 33135 5070 33255 5190
rect 33300 5070 33420 5190
rect 33475 5070 33595 5190
rect 33640 5070 33760 5190
rect 33805 5070 33925 5190
rect 33970 5070 34090 5190
rect 34145 5070 34265 5190
rect 34310 5070 34430 5190
rect 34475 5070 34595 5190
rect 34640 5070 34760 5190
rect 34815 5070 34935 5190
rect 34980 5070 35100 5190
rect 35145 5070 35265 5190
rect 35310 5070 35430 5190
rect 35485 5070 35605 5190
rect 35650 5070 35770 5190
rect 35815 5070 35935 5190
rect 35980 5070 36100 5190
rect 36155 5070 36275 5190
rect 30795 4895 30915 5015
rect 30960 4895 31080 5015
rect 31125 4895 31245 5015
rect 31290 4895 31410 5015
rect 31465 4895 31585 5015
rect 31630 4895 31750 5015
rect 31795 4895 31915 5015
rect 31960 4895 32080 5015
rect 32135 4895 32255 5015
rect 32300 4895 32420 5015
rect 32465 4895 32585 5015
rect 32630 4895 32750 5015
rect 32805 4895 32925 5015
rect 32970 4895 33090 5015
rect 33135 4895 33255 5015
rect 33300 4895 33420 5015
rect 33475 4895 33595 5015
rect 33640 4895 33760 5015
rect 33805 4895 33925 5015
rect 33970 4895 34090 5015
rect 34145 4895 34265 5015
rect 34310 4895 34430 5015
rect 34475 4895 34595 5015
rect 34640 4895 34760 5015
rect 34815 4895 34935 5015
rect 34980 4895 35100 5015
rect 35145 4895 35265 5015
rect 35310 4895 35430 5015
rect 35485 4895 35605 5015
rect 35650 4895 35770 5015
rect 35815 4895 35935 5015
rect 35980 4895 36100 5015
rect 36155 4895 36275 5015
rect 30795 4730 30915 4850
rect 30960 4730 31080 4850
rect 31125 4730 31245 4850
rect 31290 4730 31410 4850
rect 31465 4730 31585 4850
rect 31630 4730 31750 4850
rect 31795 4730 31915 4850
rect 31960 4730 32080 4850
rect 32135 4730 32255 4850
rect 32300 4730 32420 4850
rect 32465 4730 32585 4850
rect 32630 4730 32750 4850
rect 32805 4730 32925 4850
rect 32970 4730 33090 4850
rect 33135 4730 33255 4850
rect 33300 4730 33420 4850
rect 33475 4730 33595 4850
rect 33640 4730 33760 4850
rect 33805 4730 33925 4850
rect 33970 4730 34090 4850
rect 34145 4730 34265 4850
rect 34310 4730 34430 4850
rect 34475 4730 34595 4850
rect 34640 4730 34760 4850
rect 34815 4730 34935 4850
rect 34980 4730 35100 4850
rect 35145 4730 35265 4850
rect 35310 4730 35430 4850
rect 35485 4730 35605 4850
rect 35650 4730 35770 4850
rect 35815 4730 35935 4850
rect 35980 4730 36100 4850
rect 36155 4730 36275 4850
rect 30795 4565 30915 4685
rect 30960 4565 31080 4685
rect 31125 4565 31245 4685
rect 31290 4565 31410 4685
rect 31465 4565 31585 4685
rect 31630 4565 31750 4685
rect 31795 4565 31915 4685
rect 31960 4565 32080 4685
rect 32135 4565 32255 4685
rect 32300 4565 32420 4685
rect 32465 4565 32585 4685
rect 32630 4565 32750 4685
rect 32805 4565 32925 4685
rect 32970 4565 33090 4685
rect 33135 4565 33255 4685
rect 33300 4565 33420 4685
rect 33475 4565 33595 4685
rect 33640 4565 33760 4685
rect 33805 4565 33925 4685
rect 33970 4565 34090 4685
rect 34145 4565 34265 4685
rect 34310 4565 34430 4685
rect 34475 4565 34595 4685
rect 34640 4565 34760 4685
rect 34815 4565 34935 4685
rect 34980 4565 35100 4685
rect 35145 4565 35265 4685
rect 35310 4565 35430 4685
rect 35485 4565 35605 4685
rect 35650 4565 35770 4685
rect 35815 4565 35935 4685
rect 35980 4565 36100 4685
rect 36155 4565 36275 4685
rect 30795 4400 30915 4520
rect 30960 4400 31080 4520
rect 31125 4400 31245 4520
rect 31290 4400 31410 4520
rect 31465 4400 31585 4520
rect 31630 4400 31750 4520
rect 31795 4400 31915 4520
rect 31960 4400 32080 4520
rect 32135 4400 32255 4520
rect 32300 4400 32420 4520
rect 32465 4400 32585 4520
rect 32630 4400 32750 4520
rect 32805 4400 32925 4520
rect 32970 4400 33090 4520
rect 33135 4400 33255 4520
rect 33300 4400 33420 4520
rect 33475 4400 33595 4520
rect 33640 4400 33760 4520
rect 33805 4400 33925 4520
rect 33970 4400 34090 4520
rect 34145 4400 34265 4520
rect 34310 4400 34430 4520
rect 34475 4400 34595 4520
rect 34640 4400 34760 4520
rect 34815 4400 34935 4520
rect 34980 4400 35100 4520
rect 35145 4400 35265 4520
rect 35310 4400 35430 4520
rect 35485 4400 35605 4520
rect 35650 4400 35770 4520
rect 35815 4400 35935 4520
rect 35980 4400 36100 4520
rect 36155 4400 36275 4520
rect 30795 4225 30915 4345
rect 30960 4225 31080 4345
rect 31125 4225 31245 4345
rect 31290 4225 31410 4345
rect 31465 4225 31585 4345
rect 31630 4225 31750 4345
rect 31795 4225 31915 4345
rect 31960 4225 32080 4345
rect 32135 4225 32255 4345
rect 32300 4225 32420 4345
rect 32465 4225 32585 4345
rect 32630 4225 32750 4345
rect 32805 4225 32925 4345
rect 32970 4225 33090 4345
rect 33135 4225 33255 4345
rect 33300 4225 33420 4345
rect 33475 4225 33595 4345
rect 33640 4225 33760 4345
rect 33805 4225 33925 4345
rect 33970 4225 34090 4345
rect 34145 4225 34265 4345
rect 34310 4225 34430 4345
rect 34475 4225 34595 4345
rect 34640 4225 34760 4345
rect 34815 4225 34935 4345
rect 34980 4225 35100 4345
rect 35145 4225 35265 4345
rect 35310 4225 35430 4345
rect 35485 4225 35605 4345
rect 35650 4225 35770 4345
rect 35815 4225 35935 4345
rect 35980 4225 36100 4345
rect 36155 4225 36275 4345
rect 30795 4060 30915 4180
rect 30960 4060 31080 4180
rect 31125 4060 31245 4180
rect 31290 4060 31410 4180
rect 31465 4060 31585 4180
rect 31630 4060 31750 4180
rect 31795 4060 31915 4180
rect 31960 4060 32080 4180
rect 32135 4060 32255 4180
rect 32300 4060 32420 4180
rect 32465 4060 32585 4180
rect 32630 4060 32750 4180
rect 32805 4060 32925 4180
rect 32970 4060 33090 4180
rect 33135 4060 33255 4180
rect 33300 4060 33420 4180
rect 33475 4060 33595 4180
rect 33640 4060 33760 4180
rect 33805 4060 33925 4180
rect 33970 4060 34090 4180
rect 34145 4060 34265 4180
rect 34310 4060 34430 4180
rect 34475 4060 34595 4180
rect 34640 4060 34760 4180
rect 34815 4060 34935 4180
rect 34980 4060 35100 4180
rect 35145 4060 35265 4180
rect 35310 4060 35430 4180
rect 35485 4060 35605 4180
rect 35650 4060 35770 4180
rect 35815 4060 35935 4180
rect 35980 4060 36100 4180
rect 36155 4060 36275 4180
rect 30795 3895 30915 4015
rect 30960 3895 31080 4015
rect 31125 3895 31245 4015
rect 31290 3895 31410 4015
rect 31465 3895 31585 4015
rect 31630 3895 31750 4015
rect 31795 3895 31915 4015
rect 31960 3895 32080 4015
rect 32135 3895 32255 4015
rect 32300 3895 32420 4015
rect 32465 3895 32585 4015
rect 32630 3895 32750 4015
rect 32805 3895 32925 4015
rect 32970 3895 33090 4015
rect 33135 3895 33255 4015
rect 33300 3895 33420 4015
rect 33475 3895 33595 4015
rect 33640 3895 33760 4015
rect 33805 3895 33925 4015
rect 33970 3895 34090 4015
rect 34145 3895 34265 4015
rect 34310 3895 34430 4015
rect 34475 3895 34595 4015
rect 34640 3895 34760 4015
rect 34815 3895 34935 4015
rect 34980 3895 35100 4015
rect 35145 3895 35265 4015
rect 35310 3895 35430 4015
rect 35485 3895 35605 4015
rect 35650 3895 35770 4015
rect 35815 3895 35935 4015
rect 35980 3895 36100 4015
rect 36155 3895 36275 4015
rect 30795 3730 30915 3850
rect 30960 3730 31080 3850
rect 31125 3730 31245 3850
rect 31290 3730 31410 3850
rect 31465 3730 31585 3850
rect 31630 3730 31750 3850
rect 31795 3730 31915 3850
rect 31960 3730 32080 3850
rect 32135 3730 32255 3850
rect 32300 3730 32420 3850
rect 32465 3730 32585 3850
rect 32630 3730 32750 3850
rect 32805 3730 32925 3850
rect 32970 3730 33090 3850
rect 33135 3730 33255 3850
rect 33300 3730 33420 3850
rect 33475 3730 33595 3850
rect 33640 3730 33760 3850
rect 33805 3730 33925 3850
rect 33970 3730 34090 3850
rect 34145 3730 34265 3850
rect 34310 3730 34430 3850
rect 34475 3730 34595 3850
rect 34640 3730 34760 3850
rect 34815 3730 34935 3850
rect 34980 3730 35100 3850
rect 35145 3730 35265 3850
rect 35310 3730 35430 3850
rect 35485 3730 35605 3850
rect 35650 3730 35770 3850
rect 35815 3730 35935 3850
rect 35980 3730 36100 3850
rect 36155 3730 36275 3850
rect 30795 3555 30915 3675
rect 30960 3555 31080 3675
rect 31125 3555 31245 3675
rect 31290 3555 31410 3675
rect 31465 3555 31585 3675
rect 31630 3555 31750 3675
rect 31795 3555 31915 3675
rect 31960 3555 32080 3675
rect 32135 3555 32255 3675
rect 32300 3555 32420 3675
rect 32465 3555 32585 3675
rect 32630 3555 32750 3675
rect 32805 3555 32925 3675
rect 32970 3555 33090 3675
rect 33135 3555 33255 3675
rect 33300 3555 33420 3675
rect 33475 3555 33595 3675
rect 33640 3555 33760 3675
rect 33805 3555 33925 3675
rect 33970 3555 34090 3675
rect 34145 3555 34265 3675
rect 34310 3555 34430 3675
rect 34475 3555 34595 3675
rect 34640 3555 34760 3675
rect 34815 3555 34935 3675
rect 34980 3555 35100 3675
rect 35145 3555 35265 3675
rect 35310 3555 35430 3675
rect 35485 3555 35605 3675
rect 35650 3555 35770 3675
rect 35815 3555 35935 3675
rect 35980 3555 36100 3675
rect 36155 3555 36275 3675
rect 30795 3390 30915 3510
rect 30960 3390 31080 3510
rect 31125 3390 31245 3510
rect 31290 3390 31410 3510
rect 31465 3390 31585 3510
rect 31630 3390 31750 3510
rect 31795 3390 31915 3510
rect 31960 3390 32080 3510
rect 32135 3390 32255 3510
rect 32300 3390 32420 3510
rect 32465 3390 32585 3510
rect 32630 3390 32750 3510
rect 32805 3390 32925 3510
rect 32970 3390 33090 3510
rect 33135 3390 33255 3510
rect 33300 3390 33420 3510
rect 33475 3390 33595 3510
rect 33640 3390 33760 3510
rect 33805 3390 33925 3510
rect 33970 3390 34090 3510
rect 34145 3390 34265 3510
rect 34310 3390 34430 3510
rect 34475 3390 34595 3510
rect 34640 3390 34760 3510
rect 34815 3390 34935 3510
rect 34980 3390 35100 3510
rect 35145 3390 35265 3510
rect 35310 3390 35430 3510
rect 35485 3390 35605 3510
rect 35650 3390 35770 3510
rect 35815 3390 35935 3510
rect 35980 3390 36100 3510
rect 36155 3390 36275 3510
rect 30795 3225 30915 3345
rect 30960 3225 31080 3345
rect 31125 3225 31245 3345
rect 31290 3225 31410 3345
rect 31465 3225 31585 3345
rect 31630 3225 31750 3345
rect 31795 3225 31915 3345
rect 31960 3225 32080 3345
rect 32135 3225 32255 3345
rect 32300 3225 32420 3345
rect 32465 3225 32585 3345
rect 32630 3225 32750 3345
rect 32805 3225 32925 3345
rect 32970 3225 33090 3345
rect 33135 3225 33255 3345
rect 33300 3225 33420 3345
rect 33475 3225 33595 3345
rect 33640 3225 33760 3345
rect 33805 3225 33925 3345
rect 33970 3225 34090 3345
rect 34145 3225 34265 3345
rect 34310 3225 34430 3345
rect 34475 3225 34595 3345
rect 34640 3225 34760 3345
rect 34815 3225 34935 3345
rect 34980 3225 35100 3345
rect 35145 3225 35265 3345
rect 35310 3225 35430 3345
rect 35485 3225 35605 3345
rect 35650 3225 35770 3345
rect 35815 3225 35935 3345
rect 35980 3225 36100 3345
rect 36155 3225 36275 3345
rect 30795 3060 30915 3180
rect 30960 3060 31080 3180
rect 31125 3060 31245 3180
rect 31290 3060 31410 3180
rect 31465 3060 31585 3180
rect 31630 3060 31750 3180
rect 31795 3060 31915 3180
rect 31960 3060 32080 3180
rect 32135 3060 32255 3180
rect 32300 3060 32420 3180
rect 32465 3060 32585 3180
rect 32630 3060 32750 3180
rect 32805 3060 32925 3180
rect 32970 3060 33090 3180
rect 33135 3060 33255 3180
rect 33300 3060 33420 3180
rect 33475 3060 33595 3180
rect 33640 3060 33760 3180
rect 33805 3060 33925 3180
rect 33970 3060 34090 3180
rect 34145 3060 34265 3180
rect 34310 3060 34430 3180
rect 34475 3060 34595 3180
rect 34640 3060 34760 3180
rect 34815 3060 34935 3180
rect 34980 3060 35100 3180
rect 35145 3060 35265 3180
rect 35310 3060 35430 3180
rect 35485 3060 35605 3180
rect 35650 3060 35770 3180
rect 35815 3060 35935 3180
rect 35980 3060 36100 3180
rect 36155 3060 36275 3180
rect 30795 2885 30915 3005
rect 30960 2885 31080 3005
rect 31125 2885 31245 3005
rect 31290 2885 31410 3005
rect 31465 2885 31585 3005
rect 31630 2885 31750 3005
rect 31795 2885 31915 3005
rect 31960 2885 32080 3005
rect 32135 2885 32255 3005
rect 32300 2885 32420 3005
rect 32465 2885 32585 3005
rect 32630 2885 32750 3005
rect 32805 2885 32925 3005
rect 32970 2885 33090 3005
rect 33135 2885 33255 3005
rect 33300 2885 33420 3005
rect 33475 2885 33595 3005
rect 33640 2885 33760 3005
rect 33805 2885 33925 3005
rect 33970 2885 34090 3005
rect 34145 2885 34265 3005
rect 34310 2885 34430 3005
rect 34475 2885 34595 3005
rect 34640 2885 34760 3005
rect 34815 2885 34935 3005
rect 34980 2885 35100 3005
rect 35145 2885 35265 3005
rect 35310 2885 35430 3005
rect 35485 2885 35605 3005
rect 35650 2885 35770 3005
rect 35815 2885 35935 3005
rect 35980 2885 36100 3005
rect 36155 2885 36275 3005
rect 30795 2720 30915 2840
rect 30960 2720 31080 2840
rect 31125 2720 31245 2840
rect 31290 2720 31410 2840
rect 31465 2720 31585 2840
rect 31630 2720 31750 2840
rect 31795 2720 31915 2840
rect 31960 2720 32080 2840
rect 32135 2720 32255 2840
rect 32300 2720 32420 2840
rect 32465 2720 32585 2840
rect 32630 2720 32750 2840
rect 32805 2720 32925 2840
rect 32970 2720 33090 2840
rect 33135 2720 33255 2840
rect 33300 2720 33420 2840
rect 33475 2720 33595 2840
rect 33640 2720 33760 2840
rect 33805 2720 33925 2840
rect 33970 2720 34090 2840
rect 34145 2720 34265 2840
rect 34310 2720 34430 2840
rect 34475 2720 34595 2840
rect 34640 2720 34760 2840
rect 34815 2720 34935 2840
rect 34980 2720 35100 2840
rect 35145 2720 35265 2840
rect 35310 2720 35430 2840
rect 35485 2720 35605 2840
rect 35650 2720 35770 2840
rect 35815 2720 35935 2840
rect 35980 2720 36100 2840
rect 36155 2720 36275 2840
rect 30795 2555 30915 2675
rect 30960 2555 31080 2675
rect 31125 2555 31245 2675
rect 31290 2555 31410 2675
rect 31465 2555 31585 2675
rect 31630 2555 31750 2675
rect 31795 2555 31915 2675
rect 31960 2555 32080 2675
rect 32135 2555 32255 2675
rect 32300 2555 32420 2675
rect 32465 2555 32585 2675
rect 32630 2555 32750 2675
rect 32805 2555 32925 2675
rect 32970 2555 33090 2675
rect 33135 2555 33255 2675
rect 33300 2555 33420 2675
rect 33475 2555 33595 2675
rect 33640 2555 33760 2675
rect 33805 2555 33925 2675
rect 33970 2555 34090 2675
rect 34145 2555 34265 2675
rect 34310 2555 34430 2675
rect 34475 2555 34595 2675
rect 34640 2555 34760 2675
rect 34815 2555 34935 2675
rect 34980 2555 35100 2675
rect 35145 2555 35265 2675
rect 35310 2555 35430 2675
rect 35485 2555 35605 2675
rect 35650 2555 35770 2675
rect 35815 2555 35935 2675
rect 35980 2555 36100 2675
rect 36155 2555 36275 2675
rect 30795 2390 30915 2510
rect 30960 2390 31080 2510
rect 31125 2390 31245 2510
rect 31290 2390 31410 2510
rect 31465 2390 31585 2510
rect 31630 2390 31750 2510
rect 31795 2390 31915 2510
rect 31960 2390 32080 2510
rect 32135 2390 32255 2510
rect 32300 2390 32420 2510
rect 32465 2390 32585 2510
rect 32630 2390 32750 2510
rect 32805 2390 32925 2510
rect 32970 2390 33090 2510
rect 33135 2390 33255 2510
rect 33300 2390 33420 2510
rect 33475 2390 33595 2510
rect 33640 2390 33760 2510
rect 33805 2390 33925 2510
rect 33970 2390 34090 2510
rect 34145 2390 34265 2510
rect 34310 2390 34430 2510
rect 34475 2390 34595 2510
rect 34640 2390 34760 2510
rect 34815 2390 34935 2510
rect 34980 2390 35100 2510
rect 35145 2390 35265 2510
rect 35310 2390 35430 2510
rect 35485 2390 35605 2510
rect 35650 2390 35770 2510
rect 35815 2390 35935 2510
rect 35980 2390 36100 2510
rect 36155 2390 36275 2510
rect 30795 2215 30915 2335
rect 30960 2215 31080 2335
rect 31125 2215 31245 2335
rect 31290 2215 31410 2335
rect 31465 2215 31585 2335
rect 31630 2215 31750 2335
rect 31795 2215 31915 2335
rect 31960 2215 32080 2335
rect 32135 2215 32255 2335
rect 32300 2215 32420 2335
rect 32465 2215 32585 2335
rect 32630 2215 32750 2335
rect 32805 2215 32925 2335
rect 32970 2215 33090 2335
rect 33135 2215 33255 2335
rect 33300 2215 33420 2335
rect 33475 2215 33595 2335
rect 33640 2215 33760 2335
rect 33805 2215 33925 2335
rect 33970 2215 34090 2335
rect 34145 2215 34265 2335
rect 34310 2215 34430 2335
rect 34475 2215 34595 2335
rect 34640 2215 34760 2335
rect 34815 2215 34935 2335
rect 34980 2215 35100 2335
rect 35145 2215 35265 2335
rect 35310 2215 35430 2335
rect 35485 2215 35605 2335
rect 35650 2215 35770 2335
rect 35815 2215 35935 2335
rect 35980 2215 36100 2335
rect 36155 2215 36275 2335
rect 30795 2050 30915 2170
rect 30960 2050 31080 2170
rect 31125 2050 31245 2170
rect 31290 2050 31410 2170
rect 31465 2050 31585 2170
rect 31630 2050 31750 2170
rect 31795 2050 31915 2170
rect 31960 2050 32080 2170
rect 32135 2050 32255 2170
rect 32300 2050 32420 2170
rect 32465 2050 32585 2170
rect 32630 2050 32750 2170
rect 32805 2050 32925 2170
rect 32970 2050 33090 2170
rect 33135 2050 33255 2170
rect 33300 2050 33420 2170
rect 33475 2050 33595 2170
rect 33640 2050 33760 2170
rect 33805 2050 33925 2170
rect 33970 2050 34090 2170
rect 34145 2050 34265 2170
rect 34310 2050 34430 2170
rect 34475 2050 34595 2170
rect 34640 2050 34760 2170
rect 34815 2050 34935 2170
rect 34980 2050 35100 2170
rect 35145 2050 35265 2170
rect 35310 2050 35430 2170
rect 35485 2050 35605 2170
rect 35650 2050 35770 2170
rect 35815 2050 35935 2170
rect 35980 2050 36100 2170
rect 36155 2050 36275 2170
rect 30795 1885 30915 2005
rect 30960 1885 31080 2005
rect 31125 1885 31245 2005
rect 31290 1885 31410 2005
rect 31465 1885 31585 2005
rect 31630 1885 31750 2005
rect 31795 1885 31915 2005
rect 31960 1885 32080 2005
rect 32135 1885 32255 2005
rect 32300 1885 32420 2005
rect 32465 1885 32585 2005
rect 32630 1885 32750 2005
rect 32805 1885 32925 2005
rect 32970 1885 33090 2005
rect 33135 1885 33255 2005
rect 33300 1885 33420 2005
rect 33475 1885 33595 2005
rect 33640 1885 33760 2005
rect 33805 1885 33925 2005
rect 33970 1885 34090 2005
rect 34145 1885 34265 2005
rect 34310 1885 34430 2005
rect 34475 1885 34595 2005
rect 34640 1885 34760 2005
rect 34815 1885 34935 2005
rect 34980 1885 35100 2005
rect 35145 1885 35265 2005
rect 35310 1885 35430 2005
rect 35485 1885 35605 2005
rect 35650 1885 35770 2005
rect 35815 1885 35935 2005
rect 35980 1885 36100 2005
rect 36155 1885 36275 2005
rect 30795 1720 30915 1840
rect 30960 1720 31080 1840
rect 31125 1720 31245 1840
rect 31290 1720 31410 1840
rect 31465 1720 31585 1840
rect 31630 1720 31750 1840
rect 31795 1720 31915 1840
rect 31960 1720 32080 1840
rect 32135 1720 32255 1840
rect 32300 1720 32420 1840
rect 32465 1720 32585 1840
rect 32630 1720 32750 1840
rect 32805 1720 32925 1840
rect 32970 1720 33090 1840
rect 33135 1720 33255 1840
rect 33300 1720 33420 1840
rect 33475 1720 33595 1840
rect 33640 1720 33760 1840
rect 33805 1720 33925 1840
rect 33970 1720 34090 1840
rect 34145 1720 34265 1840
rect 34310 1720 34430 1840
rect 34475 1720 34595 1840
rect 34640 1720 34760 1840
rect 34815 1720 34935 1840
rect 34980 1720 35100 1840
rect 35145 1720 35265 1840
rect 35310 1720 35430 1840
rect 35485 1720 35605 1840
rect 35650 1720 35770 1840
rect 35815 1720 35935 1840
rect 35980 1720 36100 1840
rect 36155 1720 36275 1840
rect 36485 7080 36605 7200
rect 36650 7080 36770 7200
rect 36815 7080 36935 7200
rect 36980 7080 37100 7200
rect 37155 7080 37275 7200
rect 37320 7080 37440 7200
rect 37485 7080 37605 7200
rect 37650 7080 37770 7200
rect 37825 7080 37945 7200
rect 37990 7080 38110 7200
rect 38155 7080 38275 7200
rect 38320 7080 38440 7200
rect 38495 7080 38615 7200
rect 38660 7080 38780 7200
rect 38825 7080 38945 7200
rect 38990 7080 39110 7200
rect 39165 7080 39285 7200
rect 39330 7080 39450 7200
rect 39495 7080 39615 7200
rect 39660 7080 39780 7200
rect 39835 7080 39955 7200
rect 40000 7080 40120 7200
rect 40165 7080 40285 7200
rect 40330 7080 40450 7200
rect 40505 7080 40625 7200
rect 40670 7080 40790 7200
rect 40835 7080 40955 7200
rect 41000 7080 41120 7200
rect 41175 7080 41295 7200
rect 41340 7080 41460 7200
rect 41505 7080 41625 7200
rect 41670 7080 41790 7200
rect 41845 7080 41965 7200
rect 36485 6905 36605 7025
rect 36650 6905 36770 7025
rect 36815 6905 36935 7025
rect 36980 6905 37100 7025
rect 37155 6905 37275 7025
rect 37320 6905 37440 7025
rect 37485 6905 37605 7025
rect 37650 6905 37770 7025
rect 37825 6905 37945 7025
rect 37990 6905 38110 7025
rect 38155 6905 38275 7025
rect 38320 6905 38440 7025
rect 38495 6905 38615 7025
rect 38660 6905 38780 7025
rect 38825 6905 38945 7025
rect 38990 6905 39110 7025
rect 39165 6905 39285 7025
rect 39330 6905 39450 7025
rect 39495 6905 39615 7025
rect 39660 6905 39780 7025
rect 39835 6905 39955 7025
rect 40000 6905 40120 7025
rect 40165 6905 40285 7025
rect 40330 6905 40450 7025
rect 40505 6905 40625 7025
rect 40670 6905 40790 7025
rect 40835 6905 40955 7025
rect 41000 6905 41120 7025
rect 41175 6905 41295 7025
rect 41340 6905 41460 7025
rect 41505 6905 41625 7025
rect 41670 6905 41790 7025
rect 41845 6905 41965 7025
rect 36485 6740 36605 6860
rect 36650 6740 36770 6860
rect 36815 6740 36935 6860
rect 36980 6740 37100 6860
rect 37155 6740 37275 6860
rect 37320 6740 37440 6860
rect 37485 6740 37605 6860
rect 37650 6740 37770 6860
rect 37825 6740 37945 6860
rect 37990 6740 38110 6860
rect 38155 6740 38275 6860
rect 38320 6740 38440 6860
rect 38495 6740 38615 6860
rect 38660 6740 38780 6860
rect 38825 6740 38945 6860
rect 38990 6740 39110 6860
rect 39165 6740 39285 6860
rect 39330 6740 39450 6860
rect 39495 6740 39615 6860
rect 39660 6740 39780 6860
rect 39835 6740 39955 6860
rect 40000 6740 40120 6860
rect 40165 6740 40285 6860
rect 40330 6740 40450 6860
rect 40505 6740 40625 6860
rect 40670 6740 40790 6860
rect 40835 6740 40955 6860
rect 41000 6740 41120 6860
rect 41175 6740 41295 6860
rect 41340 6740 41460 6860
rect 41505 6740 41625 6860
rect 41670 6740 41790 6860
rect 41845 6740 41965 6860
rect 36485 6575 36605 6695
rect 36650 6575 36770 6695
rect 36815 6575 36935 6695
rect 36980 6575 37100 6695
rect 37155 6575 37275 6695
rect 37320 6575 37440 6695
rect 37485 6575 37605 6695
rect 37650 6575 37770 6695
rect 37825 6575 37945 6695
rect 37990 6575 38110 6695
rect 38155 6575 38275 6695
rect 38320 6575 38440 6695
rect 38495 6575 38615 6695
rect 38660 6575 38780 6695
rect 38825 6575 38945 6695
rect 38990 6575 39110 6695
rect 39165 6575 39285 6695
rect 39330 6575 39450 6695
rect 39495 6575 39615 6695
rect 39660 6575 39780 6695
rect 39835 6575 39955 6695
rect 40000 6575 40120 6695
rect 40165 6575 40285 6695
rect 40330 6575 40450 6695
rect 40505 6575 40625 6695
rect 40670 6575 40790 6695
rect 40835 6575 40955 6695
rect 41000 6575 41120 6695
rect 41175 6575 41295 6695
rect 41340 6575 41460 6695
rect 41505 6575 41625 6695
rect 41670 6575 41790 6695
rect 41845 6575 41965 6695
rect 36485 6410 36605 6530
rect 36650 6410 36770 6530
rect 36815 6410 36935 6530
rect 36980 6410 37100 6530
rect 37155 6410 37275 6530
rect 37320 6410 37440 6530
rect 37485 6410 37605 6530
rect 37650 6410 37770 6530
rect 37825 6410 37945 6530
rect 37990 6410 38110 6530
rect 38155 6410 38275 6530
rect 38320 6410 38440 6530
rect 38495 6410 38615 6530
rect 38660 6410 38780 6530
rect 38825 6410 38945 6530
rect 38990 6410 39110 6530
rect 39165 6410 39285 6530
rect 39330 6410 39450 6530
rect 39495 6410 39615 6530
rect 39660 6410 39780 6530
rect 39835 6410 39955 6530
rect 40000 6410 40120 6530
rect 40165 6410 40285 6530
rect 40330 6410 40450 6530
rect 40505 6410 40625 6530
rect 40670 6410 40790 6530
rect 40835 6410 40955 6530
rect 41000 6410 41120 6530
rect 41175 6410 41295 6530
rect 41340 6410 41460 6530
rect 41505 6410 41625 6530
rect 41670 6410 41790 6530
rect 41845 6410 41965 6530
rect 36485 6235 36605 6355
rect 36650 6235 36770 6355
rect 36815 6235 36935 6355
rect 36980 6235 37100 6355
rect 37155 6235 37275 6355
rect 37320 6235 37440 6355
rect 37485 6235 37605 6355
rect 37650 6235 37770 6355
rect 37825 6235 37945 6355
rect 37990 6235 38110 6355
rect 38155 6235 38275 6355
rect 38320 6235 38440 6355
rect 38495 6235 38615 6355
rect 38660 6235 38780 6355
rect 38825 6235 38945 6355
rect 38990 6235 39110 6355
rect 39165 6235 39285 6355
rect 39330 6235 39450 6355
rect 39495 6235 39615 6355
rect 39660 6235 39780 6355
rect 39835 6235 39955 6355
rect 40000 6235 40120 6355
rect 40165 6235 40285 6355
rect 40330 6235 40450 6355
rect 40505 6235 40625 6355
rect 40670 6235 40790 6355
rect 40835 6235 40955 6355
rect 41000 6235 41120 6355
rect 41175 6235 41295 6355
rect 41340 6235 41460 6355
rect 41505 6235 41625 6355
rect 41670 6235 41790 6355
rect 41845 6235 41965 6355
rect 36485 6070 36605 6190
rect 36650 6070 36770 6190
rect 36815 6070 36935 6190
rect 36980 6070 37100 6190
rect 37155 6070 37275 6190
rect 37320 6070 37440 6190
rect 37485 6070 37605 6190
rect 37650 6070 37770 6190
rect 37825 6070 37945 6190
rect 37990 6070 38110 6190
rect 38155 6070 38275 6190
rect 38320 6070 38440 6190
rect 38495 6070 38615 6190
rect 38660 6070 38780 6190
rect 38825 6070 38945 6190
rect 38990 6070 39110 6190
rect 39165 6070 39285 6190
rect 39330 6070 39450 6190
rect 39495 6070 39615 6190
rect 39660 6070 39780 6190
rect 39835 6070 39955 6190
rect 40000 6070 40120 6190
rect 40165 6070 40285 6190
rect 40330 6070 40450 6190
rect 40505 6070 40625 6190
rect 40670 6070 40790 6190
rect 40835 6070 40955 6190
rect 41000 6070 41120 6190
rect 41175 6070 41295 6190
rect 41340 6070 41460 6190
rect 41505 6070 41625 6190
rect 41670 6070 41790 6190
rect 41845 6070 41965 6190
rect 36485 5905 36605 6025
rect 36650 5905 36770 6025
rect 36815 5905 36935 6025
rect 36980 5905 37100 6025
rect 37155 5905 37275 6025
rect 37320 5905 37440 6025
rect 37485 5905 37605 6025
rect 37650 5905 37770 6025
rect 37825 5905 37945 6025
rect 37990 5905 38110 6025
rect 38155 5905 38275 6025
rect 38320 5905 38440 6025
rect 38495 5905 38615 6025
rect 38660 5905 38780 6025
rect 38825 5905 38945 6025
rect 38990 5905 39110 6025
rect 39165 5905 39285 6025
rect 39330 5905 39450 6025
rect 39495 5905 39615 6025
rect 39660 5905 39780 6025
rect 39835 5905 39955 6025
rect 40000 5905 40120 6025
rect 40165 5905 40285 6025
rect 40330 5905 40450 6025
rect 40505 5905 40625 6025
rect 40670 5905 40790 6025
rect 40835 5905 40955 6025
rect 41000 5905 41120 6025
rect 41175 5905 41295 6025
rect 41340 5905 41460 6025
rect 41505 5905 41625 6025
rect 41670 5905 41790 6025
rect 41845 5905 41965 6025
rect 36485 5740 36605 5860
rect 36650 5740 36770 5860
rect 36815 5740 36935 5860
rect 36980 5740 37100 5860
rect 37155 5740 37275 5860
rect 37320 5740 37440 5860
rect 37485 5740 37605 5860
rect 37650 5740 37770 5860
rect 37825 5740 37945 5860
rect 37990 5740 38110 5860
rect 38155 5740 38275 5860
rect 38320 5740 38440 5860
rect 38495 5740 38615 5860
rect 38660 5740 38780 5860
rect 38825 5740 38945 5860
rect 38990 5740 39110 5860
rect 39165 5740 39285 5860
rect 39330 5740 39450 5860
rect 39495 5740 39615 5860
rect 39660 5740 39780 5860
rect 39835 5740 39955 5860
rect 40000 5740 40120 5860
rect 40165 5740 40285 5860
rect 40330 5740 40450 5860
rect 40505 5740 40625 5860
rect 40670 5740 40790 5860
rect 40835 5740 40955 5860
rect 41000 5740 41120 5860
rect 41175 5740 41295 5860
rect 41340 5740 41460 5860
rect 41505 5740 41625 5860
rect 41670 5740 41790 5860
rect 41845 5740 41965 5860
rect 36485 5565 36605 5685
rect 36650 5565 36770 5685
rect 36815 5565 36935 5685
rect 36980 5565 37100 5685
rect 37155 5565 37275 5685
rect 37320 5565 37440 5685
rect 37485 5565 37605 5685
rect 37650 5565 37770 5685
rect 37825 5565 37945 5685
rect 37990 5565 38110 5685
rect 38155 5565 38275 5685
rect 38320 5565 38440 5685
rect 38495 5565 38615 5685
rect 38660 5565 38780 5685
rect 38825 5565 38945 5685
rect 38990 5565 39110 5685
rect 39165 5565 39285 5685
rect 39330 5565 39450 5685
rect 39495 5565 39615 5685
rect 39660 5565 39780 5685
rect 39835 5565 39955 5685
rect 40000 5565 40120 5685
rect 40165 5565 40285 5685
rect 40330 5565 40450 5685
rect 40505 5565 40625 5685
rect 40670 5565 40790 5685
rect 40835 5565 40955 5685
rect 41000 5565 41120 5685
rect 41175 5565 41295 5685
rect 41340 5565 41460 5685
rect 41505 5565 41625 5685
rect 41670 5565 41790 5685
rect 41845 5565 41965 5685
rect 36485 5400 36605 5520
rect 36650 5400 36770 5520
rect 36815 5400 36935 5520
rect 36980 5400 37100 5520
rect 37155 5400 37275 5520
rect 37320 5400 37440 5520
rect 37485 5400 37605 5520
rect 37650 5400 37770 5520
rect 37825 5400 37945 5520
rect 37990 5400 38110 5520
rect 38155 5400 38275 5520
rect 38320 5400 38440 5520
rect 38495 5400 38615 5520
rect 38660 5400 38780 5520
rect 38825 5400 38945 5520
rect 38990 5400 39110 5520
rect 39165 5400 39285 5520
rect 39330 5400 39450 5520
rect 39495 5400 39615 5520
rect 39660 5400 39780 5520
rect 39835 5400 39955 5520
rect 40000 5400 40120 5520
rect 40165 5400 40285 5520
rect 40330 5400 40450 5520
rect 40505 5400 40625 5520
rect 40670 5400 40790 5520
rect 40835 5400 40955 5520
rect 41000 5400 41120 5520
rect 41175 5400 41295 5520
rect 41340 5400 41460 5520
rect 41505 5400 41625 5520
rect 41670 5400 41790 5520
rect 41845 5400 41965 5520
rect 36485 5235 36605 5355
rect 36650 5235 36770 5355
rect 36815 5235 36935 5355
rect 36980 5235 37100 5355
rect 37155 5235 37275 5355
rect 37320 5235 37440 5355
rect 37485 5235 37605 5355
rect 37650 5235 37770 5355
rect 37825 5235 37945 5355
rect 37990 5235 38110 5355
rect 38155 5235 38275 5355
rect 38320 5235 38440 5355
rect 38495 5235 38615 5355
rect 38660 5235 38780 5355
rect 38825 5235 38945 5355
rect 38990 5235 39110 5355
rect 39165 5235 39285 5355
rect 39330 5235 39450 5355
rect 39495 5235 39615 5355
rect 39660 5235 39780 5355
rect 39835 5235 39955 5355
rect 40000 5235 40120 5355
rect 40165 5235 40285 5355
rect 40330 5235 40450 5355
rect 40505 5235 40625 5355
rect 40670 5235 40790 5355
rect 40835 5235 40955 5355
rect 41000 5235 41120 5355
rect 41175 5235 41295 5355
rect 41340 5235 41460 5355
rect 41505 5235 41625 5355
rect 41670 5235 41790 5355
rect 41845 5235 41965 5355
rect 36485 5070 36605 5190
rect 36650 5070 36770 5190
rect 36815 5070 36935 5190
rect 36980 5070 37100 5190
rect 37155 5070 37275 5190
rect 37320 5070 37440 5190
rect 37485 5070 37605 5190
rect 37650 5070 37770 5190
rect 37825 5070 37945 5190
rect 37990 5070 38110 5190
rect 38155 5070 38275 5190
rect 38320 5070 38440 5190
rect 38495 5070 38615 5190
rect 38660 5070 38780 5190
rect 38825 5070 38945 5190
rect 38990 5070 39110 5190
rect 39165 5070 39285 5190
rect 39330 5070 39450 5190
rect 39495 5070 39615 5190
rect 39660 5070 39780 5190
rect 39835 5070 39955 5190
rect 40000 5070 40120 5190
rect 40165 5070 40285 5190
rect 40330 5070 40450 5190
rect 40505 5070 40625 5190
rect 40670 5070 40790 5190
rect 40835 5070 40955 5190
rect 41000 5070 41120 5190
rect 41175 5070 41295 5190
rect 41340 5070 41460 5190
rect 41505 5070 41625 5190
rect 41670 5070 41790 5190
rect 41845 5070 41965 5190
rect 36485 4895 36605 5015
rect 36650 4895 36770 5015
rect 36815 4895 36935 5015
rect 36980 4895 37100 5015
rect 37155 4895 37275 5015
rect 37320 4895 37440 5015
rect 37485 4895 37605 5015
rect 37650 4895 37770 5015
rect 37825 4895 37945 5015
rect 37990 4895 38110 5015
rect 38155 4895 38275 5015
rect 38320 4895 38440 5015
rect 38495 4895 38615 5015
rect 38660 4895 38780 5015
rect 38825 4895 38945 5015
rect 38990 4895 39110 5015
rect 39165 4895 39285 5015
rect 39330 4895 39450 5015
rect 39495 4895 39615 5015
rect 39660 4895 39780 5015
rect 39835 4895 39955 5015
rect 40000 4895 40120 5015
rect 40165 4895 40285 5015
rect 40330 4895 40450 5015
rect 40505 4895 40625 5015
rect 40670 4895 40790 5015
rect 40835 4895 40955 5015
rect 41000 4895 41120 5015
rect 41175 4895 41295 5015
rect 41340 4895 41460 5015
rect 41505 4895 41625 5015
rect 41670 4895 41790 5015
rect 41845 4895 41965 5015
rect 36485 4730 36605 4850
rect 36650 4730 36770 4850
rect 36815 4730 36935 4850
rect 36980 4730 37100 4850
rect 37155 4730 37275 4850
rect 37320 4730 37440 4850
rect 37485 4730 37605 4850
rect 37650 4730 37770 4850
rect 37825 4730 37945 4850
rect 37990 4730 38110 4850
rect 38155 4730 38275 4850
rect 38320 4730 38440 4850
rect 38495 4730 38615 4850
rect 38660 4730 38780 4850
rect 38825 4730 38945 4850
rect 38990 4730 39110 4850
rect 39165 4730 39285 4850
rect 39330 4730 39450 4850
rect 39495 4730 39615 4850
rect 39660 4730 39780 4850
rect 39835 4730 39955 4850
rect 40000 4730 40120 4850
rect 40165 4730 40285 4850
rect 40330 4730 40450 4850
rect 40505 4730 40625 4850
rect 40670 4730 40790 4850
rect 40835 4730 40955 4850
rect 41000 4730 41120 4850
rect 41175 4730 41295 4850
rect 41340 4730 41460 4850
rect 41505 4730 41625 4850
rect 41670 4730 41790 4850
rect 41845 4730 41965 4850
rect 36485 4565 36605 4685
rect 36650 4565 36770 4685
rect 36815 4565 36935 4685
rect 36980 4565 37100 4685
rect 37155 4565 37275 4685
rect 37320 4565 37440 4685
rect 37485 4565 37605 4685
rect 37650 4565 37770 4685
rect 37825 4565 37945 4685
rect 37990 4565 38110 4685
rect 38155 4565 38275 4685
rect 38320 4565 38440 4685
rect 38495 4565 38615 4685
rect 38660 4565 38780 4685
rect 38825 4565 38945 4685
rect 38990 4565 39110 4685
rect 39165 4565 39285 4685
rect 39330 4565 39450 4685
rect 39495 4565 39615 4685
rect 39660 4565 39780 4685
rect 39835 4565 39955 4685
rect 40000 4565 40120 4685
rect 40165 4565 40285 4685
rect 40330 4565 40450 4685
rect 40505 4565 40625 4685
rect 40670 4565 40790 4685
rect 40835 4565 40955 4685
rect 41000 4565 41120 4685
rect 41175 4565 41295 4685
rect 41340 4565 41460 4685
rect 41505 4565 41625 4685
rect 41670 4565 41790 4685
rect 41845 4565 41965 4685
rect 36485 4400 36605 4520
rect 36650 4400 36770 4520
rect 36815 4400 36935 4520
rect 36980 4400 37100 4520
rect 37155 4400 37275 4520
rect 37320 4400 37440 4520
rect 37485 4400 37605 4520
rect 37650 4400 37770 4520
rect 37825 4400 37945 4520
rect 37990 4400 38110 4520
rect 38155 4400 38275 4520
rect 38320 4400 38440 4520
rect 38495 4400 38615 4520
rect 38660 4400 38780 4520
rect 38825 4400 38945 4520
rect 38990 4400 39110 4520
rect 39165 4400 39285 4520
rect 39330 4400 39450 4520
rect 39495 4400 39615 4520
rect 39660 4400 39780 4520
rect 39835 4400 39955 4520
rect 40000 4400 40120 4520
rect 40165 4400 40285 4520
rect 40330 4400 40450 4520
rect 40505 4400 40625 4520
rect 40670 4400 40790 4520
rect 40835 4400 40955 4520
rect 41000 4400 41120 4520
rect 41175 4400 41295 4520
rect 41340 4400 41460 4520
rect 41505 4400 41625 4520
rect 41670 4400 41790 4520
rect 41845 4400 41965 4520
rect 36485 4225 36605 4345
rect 36650 4225 36770 4345
rect 36815 4225 36935 4345
rect 36980 4225 37100 4345
rect 37155 4225 37275 4345
rect 37320 4225 37440 4345
rect 37485 4225 37605 4345
rect 37650 4225 37770 4345
rect 37825 4225 37945 4345
rect 37990 4225 38110 4345
rect 38155 4225 38275 4345
rect 38320 4225 38440 4345
rect 38495 4225 38615 4345
rect 38660 4225 38780 4345
rect 38825 4225 38945 4345
rect 38990 4225 39110 4345
rect 39165 4225 39285 4345
rect 39330 4225 39450 4345
rect 39495 4225 39615 4345
rect 39660 4225 39780 4345
rect 39835 4225 39955 4345
rect 40000 4225 40120 4345
rect 40165 4225 40285 4345
rect 40330 4225 40450 4345
rect 40505 4225 40625 4345
rect 40670 4225 40790 4345
rect 40835 4225 40955 4345
rect 41000 4225 41120 4345
rect 41175 4225 41295 4345
rect 41340 4225 41460 4345
rect 41505 4225 41625 4345
rect 41670 4225 41790 4345
rect 41845 4225 41965 4345
rect 36485 4060 36605 4180
rect 36650 4060 36770 4180
rect 36815 4060 36935 4180
rect 36980 4060 37100 4180
rect 37155 4060 37275 4180
rect 37320 4060 37440 4180
rect 37485 4060 37605 4180
rect 37650 4060 37770 4180
rect 37825 4060 37945 4180
rect 37990 4060 38110 4180
rect 38155 4060 38275 4180
rect 38320 4060 38440 4180
rect 38495 4060 38615 4180
rect 38660 4060 38780 4180
rect 38825 4060 38945 4180
rect 38990 4060 39110 4180
rect 39165 4060 39285 4180
rect 39330 4060 39450 4180
rect 39495 4060 39615 4180
rect 39660 4060 39780 4180
rect 39835 4060 39955 4180
rect 40000 4060 40120 4180
rect 40165 4060 40285 4180
rect 40330 4060 40450 4180
rect 40505 4060 40625 4180
rect 40670 4060 40790 4180
rect 40835 4060 40955 4180
rect 41000 4060 41120 4180
rect 41175 4060 41295 4180
rect 41340 4060 41460 4180
rect 41505 4060 41625 4180
rect 41670 4060 41790 4180
rect 41845 4060 41965 4180
rect 36485 3895 36605 4015
rect 36650 3895 36770 4015
rect 36815 3895 36935 4015
rect 36980 3895 37100 4015
rect 37155 3895 37275 4015
rect 37320 3895 37440 4015
rect 37485 3895 37605 4015
rect 37650 3895 37770 4015
rect 37825 3895 37945 4015
rect 37990 3895 38110 4015
rect 38155 3895 38275 4015
rect 38320 3895 38440 4015
rect 38495 3895 38615 4015
rect 38660 3895 38780 4015
rect 38825 3895 38945 4015
rect 38990 3895 39110 4015
rect 39165 3895 39285 4015
rect 39330 3895 39450 4015
rect 39495 3895 39615 4015
rect 39660 3895 39780 4015
rect 39835 3895 39955 4015
rect 40000 3895 40120 4015
rect 40165 3895 40285 4015
rect 40330 3895 40450 4015
rect 40505 3895 40625 4015
rect 40670 3895 40790 4015
rect 40835 3895 40955 4015
rect 41000 3895 41120 4015
rect 41175 3895 41295 4015
rect 41340 3895 41460 4015
rect 41505 3895 41625 4015
rect 41670 3895 41790 4015
rect 41845 3895 41965 4015
rect 36485 3730 36605 3850
rect 36650 3730 36770 3850
rect 36815 3730 36935 3850
rect 36980 3730 37100 3850
rect 37155 3730 37275 3850
rect 37320 3730 37440 3850
rect 37485 3730 37605 3850
rect 37650 3730 37770 3850
rect 37825 3730 37945 3850
rect 37990 3730 38110 3850
rect 38155 3730 38275 3850
rect 38320 3730 38440 3850
rect 38495 3730 38615 3850
rect 38660 3730 38780 3850
rect 38825 3730 38945 3850
rect 38990 3730 39110 3850
rect 39165 3730 39285 3850
rect 39330 3730 39450 3850
rect 39495 3730 39615 3850
rect 39660 3730 39780 3850
rect 39835 3730 39955 3850
rect 40000 3730 40120 3850
rect 40165 3730 40285 3850
rect 40330 3730 40450 3850
rect 40505 3730 40625 3850
rect 40670 3730 40790 3850
rect 40835 3730 40955 3850
rect 41000 3730 41120 3850
rect 41175 3730 41295 3850
rect 41340 3730 41460 3850
rect 41505 3730 41625 3850
rect 41670 3730 41790 3850
rect 41845 3730 41965 3850
rect 36485 3555 36605 3675
rect 36650 3555 36770 3675
rect 36815 3555 36935 3675
rect 36980 3555 37100 3675
rect 37155 3555 37275 3675
rect 37320 3555 37440 3675
rect 37485 3555 37605 3675
rect 37650 3555 37770 3675
rect 37825 3555 37945 3675
rect 37990 3555 38110 3675
rect 38155 3555 38275 3675
rect 38320 3555 38440 3675
rect 38495 3555 38615 3675
rect 38660 3555 38780 3675
rect 38825 3555 38945 3675
rect 38990 3555 39110 3675
rect 39165 3555 39285 3675
rect 39330 3555 39450 3675
rect 39495 3555 39615 3675
rect 39660 3555 39780 3675
rect 39835 3555 39955 3675
rect 40000 3555 40120 3675
rect 40165 3555 40285 3675
rect 40330 3555 40450 3675
rect 40505 3555 40625 3675
rect 40670 3555 40790 3675
rect 40835 3555 40955 3675
rect 41000 3555 41120 3675
rect 41175 3555 41295 3675
rect 41340 3555 41460 3675
rect 41505 3555 41625 3675
rect 41670 3555 41790 3675
rect 41845 3555 41965 3675
rect 36485 3390 36605 3510
rect 36650 3390 36770 3510
rect 36815 3390 36935 3510
rect 36980 3390 37100 3510
rect 37155 3390 37275 3510
rect 37320 3390 37440 3510
rect 37485 3390 37605 3510
rect 37650 3390 37770 3510
rect 37825 3390 37945 3510
rect 37990 3390 38110 3510
rect 38155 3390 38275 3510
rect 38320 3390 38440 3510
rect 38495 3390 38615 3510
rect 38660 3390 38780 3510
rect 38825 3390 38945 3510
rect 38990 3390 39110 3510
rect 39165 3390 39285 3510
rect 39330 3390 39450 3510
rect 39495 3390 39615 3510
rect 39660 3390 39780 3510
rect 39835 3390 39955 3510
rect 40000 3390 40120 3510
rect 40165 3390 40285 3510
rect 40330 3390 40450 3510
rect 40505 3390 40625 3510
rect 40670 3390 40790 3510
rect 40835 3390 40955 3510
rect 41000 3390 41120 3510
rect 41175 3390 41295 3510
rect 41340 3390 41460 3510
rect 41505 3390 41625 3510
rect 41670 3390 41790 3510
rect 41845 3390 41965 3510
rect 36485 3225 36605 3345
rect 36650 3225 36770 3345
rect 36815 3225 36935 3345
rect 36980 3225 37100 3345
rect 37155 3225 37275 3345
rect 37320 3225 37440 3345
rect 37485 3225 37605 3345
rect 37650 3225 37770 3345
rect 37825 3225 37945 3345
rect 37990 3225 38110 3345
rect 38155 3225 38275 3345
rect 38320 3225 38440 3345
rect 38495 3225 38615 3345
rect 38660 3225 38780 3345
rect 38825 3225 38945 3345
rect 38990 3225 39110 3345
rect 39165 3225 39285 3345
rect 39330 3225 39450 3345
rect 39495 3225 39615 3345
rect 39660 3225 39780 3345
rect 39835 3225 39955 3345
rect 40000 3225 40120 3345
rect 40165 3225 40285 3345
rect 40330 3225 40450 3345
rect 40505 3225 40625 3345
rect 40670 3225 40790 3345
rect 40835 3225 40955 3345
rect 41000 3225 41120 3345
rect 41175 3225 41295 3345
rect 41340 3225 41460 3345
rect 41505 3225 41625 3345
rect 41670 3225 41790 3345
rect 41845 3225 41965 3345
rect 36485 3060 36605 3180
rect 36650 3060 36770 3180
rect 36815 3060 36935 3180
rect 36980 3060 37100 3180
rect 37155 3060 37275 3180
rect 37320 3060 37440 3180
rect 37485 3060 37605 3180
rect 37650 3060 37770 3180
rect 37825 3060 37945 3180
rect 37990 3060 38110 3180
rect 38155 3060 38275 3180
rect 38320 3060 38440 3180
rect 38495 3060 38615 3180
rect 38660 3060 38780 3180
rect 38825 3060 38945 3180
rect 38990 3060 39110 3180
rect 39165 3060 39285 3180
rect 39330 3060 39450 3180
rect 39495 3060 39615 3180
rect 39660 3060 39780 3180
rect 39835 3060 39955 3180
rect 40000 3060 40120 3180
rect 40165 3060 40285 3180
rect 40330 3060 40450 3180
rect 40505 3060 40625 3180
rect 40670 3060 40790 3180
rect 40835 3060 40955 3180
rect 41000 3060 41120 3180
rect 41175 3060 41295 3180
rect 41340 3060 41460 3180
rect 41505 3060 41625 3180
rect 41670 3060 41790 3180
rect 41845 3060 41965 3180
rect 36485 2885 36605 3005
rect 36650 2885 36770 3005
rect 36815 2885 36935 3005
rect 36980 2885 37100 3005
rect 37155 2885 37275 3005
rect 37320 2885 37440 3005
rect 37485 2885 37605 3005
rect 37650 2885 37770 3005
rect 37825 2885 37945 3005
rect 37990 2885 38110 3005
rect 38155 2885 38275 3005
rect 38320 2885 38440 3005
rect 38495 2885 38615 3005
rect 38660 2885 38780 3005
rect 38825 2885 38945 3005
rect 38990 2885 39110 3005
rect 39165 2885 39285 3005
rect 39330 2885 39450 3005
rect 39495 2885 39615 3005
rect 39660 2885 39780 3005
rect 39835 2885 39955 3005
rect 40000 2885 40120 3005
rect 40165 2885 40285 3005
rect 40330 2885 40450 3005
rect 40505 2885 40625 3005
rect 40670 2885 40790 3005
rect 40835 2885 40955 3005
rect 41000 2885 41120 3005
rect 41175 2885 41295 3005
rect 41340 2885 41460 3005
rect 41505 2885 41625 3005
rect 41670 2885 41790 3005
rect 41845 2885 41965 3005
rect 36485 2720 36605 2840
rect 36650 2720 36770 2840
rect 36815 2720 36935 2840
rect 36980 2720 37100 2840
rect 37155 2720 37275 2840
rect 37320 2720 37440 2840
rect 37485 2720 37605 2840
rect 37650 2720 37770 2840
rect 37825 2720 37945 2840
rect 37990 2720 38110 2840
rect 38155 2720 38275 2840
rect 38320 2720 38440 2840
rect 38495 2720 38615 2840
rect 38660 2720 38780 2840
rect 38825 2720 38945 2840
rect 38990 2720 39110 2840
rect 39165 2720 39285 2840
rect 39330 2720 39450 2840
rect 39495 2720 39615 2840
rect 39660 2720 39780 2840
rect 39835 2720 39955 2840
rect 40000 2720 40120 2840
rect 40165 2720 40285 2840
rect 40330 2720 40450 2840
rect 40505 2720 40625 2840
rect 40670 2720 40790 2840
rect 40835 2720 40955 2840
rect 41000 2720 41120 2840
rect 41175 2720 41295 2840
rect 41340 2720 41460 2840
rect 41505 2720 41625 2840
rect 41670 2720 41790 2840
rect 41845 2720 41965 2840
rect 36485 2555 36605 2675
rect 36650 2555 36770 2675
rect 36815 2555 36935 2675
rect 36980 2555 37100 2675
rect 37155 2555 37275 2675
rect 37320 2555 37440 2675
rect 37485 2555 37605 2675
rect 37650 2555 37770 2675
rect 37825 2555 37945 2675
rect 37990 2555 38110 2675
rect 38155 2555 38275 2675
rect 38320 2555 38440 2675
rect 38495 2555 38615 2675
rect 38660 2555 38780 2675
rect 38825 2555 38945 2675
rect 38990 2555 39110 2675
rect 39165 2555 39285 2675
rect 39330 2555 39450 2675
rect 39495 2555 39615 2675
rect 39660 2555 39780 2675
rect 39835 2555 39955 2675
rect 40000 2555 40120 2675
rect 40165 2555 40285 2675
rect 40330 2555 40450 2675
rect 40505 2555 40625 2675
rect 40670 2555 40790 2675
rect 40835 2555 40955 2675
rect 41000 2555 41120 2675
rect 41175 2555 41295 2675
rect 41340 2555 41460 2675
rect 41505 2555 41625 2675
rect 41670 2555 41790 2675
rect 41845 2555 41965 2675
rect 36485 2390 36605 2510
rect 36650 2390 36770 2510
rect 36815 2390 36935 2510
rect 36980 2390 37100 2510
rect 37155 2390 37275 2510
rect 37320 2390 37440 2510
rect 37485 2390 37605 2510
rect 37650 2390 37770 2510
rect 37825 2390 37945 2510
rect 37990 2390 38110 2510
rect 38155 2390 38275 2510
rect 38320 2390 38440 2510
rect 38495 2390 38615 2510
rect 38660 2390 38780 2510
rect 38825 2390 38945 2510
rect 38990 2390 39110 2510
rect 39165 2390 39285 2510
rect 39330 2390 39450 2510
rect 39495 2390 39615 2510
rect 39660 2390 39780 2510
rect 39835 2390 39955 2510
rect 40000 2390 40120 2510
rect 40165 2390 40285 2510
rect 40330 2390 40450 2510
rect 40505 2390 40625 2510
rect 40670 2390 40790 2510
rect 40835 2390 40955 2510
rect 41000 2390 41120 2510
rect 41175 2390 41295 2510
rect 41340 2390 41460 2510
rect 41505 2390 41625 2510
rect 41670 2390 41790 2510
rect 41845 2390 41965 2510
rect 36485 2215 36605 2335
rect 36650 2215 36770 2335
rect 36815 2215 36935 2335
rect 36980 2215 37100 2335
rect 37155 2215 37275 2335
rect 37320 2215 37440 2335
rect 37485 2215 37605 2335
rect 37650 2215 37770 2335
rect 37825 2215 37945 2335
rect 37990 2215 38110 2335
rect 38155 2215 38275 2335
rect 38320 2215 38440 2335
rect 38495 2215 38615 2335
rect 38660 2215 38780 2335
rect 38825 2215 38945 2335
rect 38990 2215 39110 2335
rect 39165 2215 39285 2335
rect 39330 2215 39450 2335
rect 39495 2215 39615 2335
rect 39660 2215 39780 2335
rect 39835 2215 39955 2335
rect 40000 2215 40120 2335
rect 40165 2215 40285 2335
rect 40330 2215 40450 2335
rect 40505 2215 40625 2335
rect 40670 2215 40790 2335
rect 40835 2215 40955 2335
rect 41000 2215 41120 2335
rect 41175 2215 41295 2335
rect 41340 2215 41460 2335
rect 41505 2215 41625 2335
rect 41670 2215 41790 2335
rect 41845 2215 41965 2335
rect 36485 2050 36605 2170
rect 36650 2050 36770 2170
rect 36815 2050 36935 2170
rect 36980 2050 37100 2170
rect 37155 2050 37275 2170
rect 37320 2050 37440 2170
rect 37485 2050 37605 2170
rect 37650 2050 37770 2170
rect 37825 2050 37945 2170
rect 37990 2050 38110 2170
rect 38155 2050 38275 2170
rect 38320 2050 38440 2170
rect 38495 2050 38615 2170
rect 38660 2050 38780 2170
rect 38825 2050 38945 2170
rect 38990 2050 39110 2170
rect 39165 2050 39285 2170
rect 39330 2050 39450 2170
rect 39495 2050 39615 2170
rect 39660 2050 39780 2170
rect 39835 2050 39955 2170
rect 40000 2050 40120 2170
rect 40165 2050 40285 2170
rect 40330 2050 40450 2170
rect 40505 2050 40625 2170
rect 40670 2050 40790 2170
rect 40835 2050 40955 2170
rect 41000 2050 41120 2170
rect 41175 2050 41295 2170
rect 41340 2050 41460 2170
rect 41505 2050 41625 2170
rect 41670 2050 41790 2170
rect 41845 2050 41965 2170
rect 36485 1885 36605 2005
rect 36650 1885 36770 2005
rect 36815 1885 36935 2005
rect 36980 1885 37100 2005
rect 37155 1885 37275 2005
rect 37320 1885 37440 2005
rect 37485 1885 37605 2005
rect 37650 1885 37770 2005
rect 37825 1885 37945 2005
rect 37990 1885 38110 2005
rect 38155 1885 38275 2005
rect 38320 1885 38440 2005
rect 38495 1885 38615 2005
rect 38660 1885 38780 2005
rect 38825 1885 38945 2005
rect 38990 1885 39110 2005
rect 39165 1885 39285 2005
rect 39330 1885 39450 2005
rect 39495 1885 39615 2005
rect 39660 1885 39780 2005
rect 39835 1885 39955 2005
rect 40000 1885 40120 2005
rect 40165 1885 40285 2005
rect 40330 1885 40450 2005
rect 40505 1885 40625 2005
rect 40670 1885 40790 2005
rect 40835 1885 40955 2005
rect 41000 1885 41120 2005
rect 41175 1885 41295 2005
rect 41340 1885 41460 2005
rect 41505 1885 41625 2005
rect 41670 1885 41790 2005
rect 41845 1885 41965 2005
rect 36485 1720 36605 1840
rect 36650 1720 36770 1840
rect 36815 1720 36935 1840
rect 36980 1720 37100 1840
rect 37155 1720 37275 1840
rect 37320 1720 37440 1840
rect 37485 1720 37605 1840
rect 37650 1720 37770 1840
rect 37825 1720 37945 1840
rect 37990 1720 38110 1840
rect 38155 1720 38275 1840
rect 38320 1720 38440 1840
rect 38495 1720 38615 1840
rect 38660 1720 38780 1840
rect 38825 1720 38945 1840
rect 38990 1720 39110 1840
rect 39165 1720 39285 1840
rect 39330 1720 39450 1840
rect 39495 1720 39615 1840
rect 39660 1720 39780 1840
rect 39835 1720 39955 1840
rect 40000 1720 40120 1840
rect 40165 1720 40285 1840
rect 40330 1720 40450 1840
rect 40505 1720 40625 1840
rect 40670 1720 40790 1840
rect 40835 1720 40955 1840
rect 41000 1720 41120 1840
rect 41175 1720 41295 1840
rect 41340 1720 41460 1840
rect 41505 1720 41625 1840
rect 41670 1720 41790 1840
rect 41845 1720 41965 1840
rect 42175 7080 42295 7200
rect 42340 7080 42460 7200
rect 42505 7080 42625 7200
rect 42670 7080 42790 7200
rect 42845 7080 42965 7200
rect 43010 7080 43130 7200
rect 43175 7080 43295 7200
rect 43340 7080 43460 7200
rect 43515 7080 43635 7200
rect 43680 7080 43800 7200
rect 43845 7080 43965 7200
rect 44010 7080 44130 7200
rect 44185 7080 44305 7200
rect 44350 7080 44470 7200
rect 44515 7080 44635 7200
rect 44680 7080 44800 7200
rect 44855 7080 44975 7200
rect 45020 7080 45140 7200
rect 45185 7080 45305 7200
rect 45350 7080 45470 7200
rect 45525 7080 45645 7200
rect 45690 7080 45810 7200
rect 45855 7080 45975 7200
rect 46020 7080 46140 7200
rect 46195 7080 46315 7200
rect 46360 7080 46480 7200
rect 46525 7080 46645 7200
rect 46690 7080 46810 7200
rect 46865 7080 46985 7200
rect 47030 7080 47150 7200
rect 47195 7080 47315 7200
rect 47360 7080 47480 7200
rect 47535 7080 47655 7200
rect 42175 6905 42295 7025
rect 42340 6905 42460 7025
rect 42505 6905 42625 7025
rect 42670 6905 42790 7025
rect 42845 6905 42965 7025
rect 43010 6905 43130 7025
rect 43175 6905 43295 7025
rect 43340 6905 43460 7025
rect 43515 6905 43635 7025
rect 43680 6905 43800 7025
rect 43845 6905 43965 7025
rect 44010 6905 44130 7025
rect 44185 6905 44305 7025
rect 44350 6905 44470 7025
rect 44515 6905 44635 7025
rect 44680 6905 44800 7025
rect 44855 6905 44975 7025
rect 45020 6905 45140 7025
rect 45185 6905 45305 7025
rect 45350 6905 45470 7025
rect 45525 6905 45645 7025
rect 45690 6905 45810 7025
rect 45855 6905 45975 7025
rect 46020 6905 46140 7025
rect 46195 6905 46315 7025
rect 46360 6905 46480 7025
rect 46525 6905 46645 7025
rect 46690 6905 46810 7025
rect 46865 6905 46985 7025
rect 47030 6905 47150 7025
rect 47195 6905 47315 7025
rect 47360 6905 47480 7025
rect 47535 6905 47655 7025
rect 42175 6740 42295 6860
rect 42340 6740 42460 6860
rect 42505 6740 42625 6860
rect 42670 6740 42790 6860
rect 42845 6740 42965 6860
rect 43010 6740 43130 6860
rect 43175 6740 43295 6860
rect 43340 6740 43460 6860
rect 43515 6740 43635 6860
rect 43680 6740 43800 6860
rect 43845 6740 43965 6860
rect 44010 6740 44130 6860
rect 44185 6740 44305 6860
rect 44350 6740 44470 6860
rect 44515 6740 44635 6860
rect 44680 6740 44800 6860
rect 44855 6740 44975 6860
rect 45020 6740 45140 6860
rect 45185 6740 45305 6860
rect 45350 6740 45470 6860
rect 45525 6740 45645 6860
rect 45690 6740 45810 6860
rect 45855 6740 45975 6860
rect 46020 6740 46140 6860
rect 46195 6740 46315 6860
rect 46360 6740 46480 6860
rect 46525 6740 46645 6860
rect 46690 6740 46810 6860
rect 46865 6740 46985 6860
rect 47030 6740 47150 6860
rect 47195 6740 47315 6860
rect 47360 6740 47480 6860
rect 47535 6740 47655 6860
rect 42175 6575 42295 6695
rect 42340 6575 42460 6695
rect 42505 6575 42625 6695
rect 42670 6575 42790 6695
rect 42845 6575 42965 6695
rect 43010 6575 43130 6695
rect 43175 6575 43295 6695
rect 43340 6575 43460 6695
rect 43515 6575 43635 6695
rect 43680 6575 43800 6695
rect 43845 6575 43965 6695
rect 44010 6575 44130 6695
rect 44185 6575 44305 6695
rect 44350 6575 44470 6695
rect 44515 6575 44635 6695
rect 44680 6575 44800 6695
rect 44855 6575 44975 6695
rect 45020 6575 45140 6695
rect 45185 6575 45305 6695
rect 45350 6575 45470 6695
rect 45525 6575 45645 6695
rect 45690 6575 45810 6695
rect 45855 6575 45975 6695
rect 46020 6575 46140 6695
rect 46195 6575 46315 6695
rect 46360 6575 46480 6695
rect 46525 6575 46645 6695
rect 46690 6575 46810 6695
rect 46865 6575 46985 6695
rect 47030 6575 47150 6695
rect 47195 6575 47315 6695
rect 47360 6575 47480 6695
rect 47535 6575 47655 6695
rect 42175 6410 42295 6530
rect 42340 6410 42460 6530
rect 42505 6410 42625 6530
rect 42670 6410 42790 6530
rect 42845 6410 42965 6530
rect 43010 6410 43130 6530
rect 43175 6410 43295 6530
rect 43340 6410 43460 6530
rect 43515 6410 43635 6530
rect 43680 6410 43800 6530
rect 43845 6410 43965 6530
rect 44010 6410 44130 6530
rect 44185 6410 44305 6530
rect 44350 6410 44470 6530
rect 44515 6410 44635 6530
rect 44680 6410 44800 6530
rect 44855 6410 44975 6530
rect 45020 6410 45140 6530
rect 45185 6410 45305 6530
rect 45350 6410 45470 6530
rect 45525 6410 45645 6530
rect 45690 6410 45810 6530
rect 45855 6410 45975 6530
rect 46020 6410 46140 6530
rect 46195 6410 46315 6530
rect 46360 6410 46480 6530
rect 46525 6410 46645 6530
rect 46690 6410 46810 6530
rect 46865 6410 46985 6530
rect 47030 6410 47150 6530
rect 47195 6410 47315 6530
rect 47360 6410 47480 6530
rect 47535 6410 47655 6530
rect 42175 6235 42295 6355
rect 42340 6235 42460 6355
rect 42505 6235 42625 6355
rect 42670 6235 42790 6355
rect 42845 6235 42965 6355
rect 43010 6235 43130 6355
rect 43175 6235 43295 6355
rect 43340 6235 43460 6355
rect 43515 6235 43635 6355
rect 43680 6235 43800 6355
rect 43845 6235 43965 6355
rect 44010 6235 44130 6355
rect 44185 6235 44305 6355
rect 44350 6235 44470 6355
rect 44515 6235 44635 6355
rect 44680 6235 44800 6355
rect 44855 6235 44975 6355
rect 45020 6235 45140 6355
rect 45185 6235 45305 6355
rect 45350 6235 45470 6355
rect 45525 6235 45645 6355
rect 45690 6235 45810 6355
rect 45855 6235 45975 6355
rect 46020 6235 46140 6355
rect 46195 6235 46315 6355
rect 46360 6235 46480 6355
rect 46525 6235 46645 6355
rect 46690 6235 46810 6355
rect 46865 6235 46985 6355
rect 47030 6235 47150 6355
rect 47195 6235 47315 6355
rect 47360 6235 47480 6355
rect 47535 6235 47655 6355
rect 42175 6070 42295 6190
rect 42340 6070 42460 6190
rect 42505 6070 42625 6190
rect 42670 6070 42790 6190
rect 42845 6070 42965 6190
rect 43010 6070 43130 6190
rect 43175 6070 43295 6190
rect 43340 6070 43460 6190
rect 43515 6070 43635 6190
rect 43680 6070 43800 6190
rect 43845 6070 43965 6190
rect 44010 6070 44130 6190
rect 44185 6070 44305 6190
rect 44350 6070 44470 6190
rect 44515 6070 44635 6190
rect 44680 6070 44800 6190
rect 44855 6070 44975 6190
rect 45020 6070 45140 6190
rect 45185 6070 45305 6190
rect 45350 6070 45470 6190
rect 45525 6070 45645 6190
rect 45690 6070 45810 6190
rect 45855 6070 45975 6190
rect 46020 6070 46140 6190
rect 46195 6070 46315 6190
rect 46360 6070 46480 6190
rect 46525 6070 46645 6190
rect 46690 6070 46810 6190
rect 46865 6070 46985 6190
rect 47030 6070 47150 6190
rect 47195 6070 47315 6190
rect 47360 6070 47480 6190
rect 47535 6070 47655 6190
rect 42175 5905 42295 6025
rect 42340 5905 42460 6025
rect 42505 5905 42625 6025
rect 42670 5905 42790 6025
rect 42845 5905 42965 6025
rect 43010 5905 43130 6025
rect 43175 5905 43295 6025
rect 43340 5905 43460 6025
rect 43515 5905 43635 6025
rect 43680 5905 43800 6025
rect 43845 5905 43965 6025
rect 44010 5905 44130 6025
rect 44185 5905 44305 6025
rect 44350 5905 44470 6025
rect 44515 5905 44635 6025
rect 44680 5905 44800 6025
rect 44855 5905 44975 6025
rect 45020 5905 45140 6025
rect 45185 5905 45305 6025
rect 45350 5905 45470 6025
rect 45525 5905 45645 6025
rect 45690 5905 45810 6025
rect 45855 5905 45975 6025
rect 46020 5905 46140 6025
rect 46195 5905 46315 6025
rect 46360 5905 46480 6025
rect 46525 5905 46645 6025
rect 46690 5905 46810 6025
rect 46865 5905 46985 6025
rect 47030 5905 47150 6025
rect 47195 5905 47315 6025
rect 47360 5905 47480 6025
rect 47535 5905 47655 6025
rect 42175 5740 42295 5860
rect 42340 5740 42460 5860
rect 42505 5740 42625 5860
rect 42670 5740 42790 5860
rect 42845 5740 42965 5860
rect 43010 5740 43130 5860
rect 43175 5740 43295 5860
rect 43340 5740 43460 5860
rect 43515 5740 43635 5860
rect 43680 5740 43800 5860
rect 43845 5740 43965 5860
rect 44010 5740 44130 5860
rect 44185 5740 44305 5860
rect 44350 5740 44470 5860
rect 44515 5740 44635 5860
rect 44680 5740 44800 5860
rect 44855 5740 44975 5860
rect 45020 5740 45140 5860
rect 45185 5740 45305 5860
rect 45350 5740 45470 5860
rect 45525 5740 45645 5860
rect 45690 5740 45810 5860
rect 45855 5740 45975 5860
rect 46020 5740 46140 5860
rect 46195 5740 46315 5860
rect 46360 5740 46480 5860
rect 46525 5740 46645 5860
rect 46690 5740 46810 5860
rect 46865 5740 46985 5860
rect 47030 5740 47150 5860
rect 47195 5740 47315 5860
rect 47360 5740 47480 5860
rect 47535 5740 47655 5860
rect 42175 5565 42295 5685
rect 42340 5565 42460 5685
rect 42505 5565 42625 5685
rect 42670 5565 42790 5685
rect 42845 5565 42965 5685
rect 43010 5565 43130 5685
rect 43175 5565 43295 5685
rect 43340 5565 43460 5685
rect 43515 5565 43635 5685
rect 43680 5565 43800 5685
rect 43845 5565 43965 5685
rect 44010 5565 44130 5685
rect 44185 5565 44305 5685
rect 44350 5565 44470 5685
rect 44515 5565 44635 5685
rect 44680 5565 44800 5685
rect 44855 5565 44975 5685
rect 45020 5565 45140 5685
rect 45185 5565 45305 5685
rect 45350 5565 45470 5685
rect 45525 5565 45645 5685
rect 45690 5565 45810 5685
rect 45855 5565 45975 5685
rect 46020 5565 46140 5685
rect 46195 5565 46315 5685
rect 46360 5565 46480 5685
rect 46525 5565 46645 5685
rect 46690 5565 46810 5685
rect 46865 5565 46985 5685
rect 47030 5565 47150 5685
rect 47195 5565 47315 5685
rect 47360 5565 47480 5685
rect 47535 5565 47655 5685
rect 42175 5400 42295 5520
rect 42340 5400 42460 5520
rect 42505 5400 42625 5520
rect 42670 5400 42790 5520
rect 42845 5400 42965 5520
rect 43010 5400 43130 5520
rect 43175 5400 43295 5520
rect 43340 5400 43460 5520
rect 43515 5400 43635 5520
rect 43680 5400 43800 5520
rect 43845 5400 43965 5520
rect 44010 5400 44130 5520
rect 44185 5400 44305 5520
rect 44350 5400 44470 5520
rect 44515 5400 44635 5520
rect 44680 5400 44800 5520
rect 44855 5400 44975 5520
rect 45020 5400 45140 5520
rect 45185 5400 45305 5520
rect 45350 5400 45470 5520
rect 45525 5400 45645 5520
rect 45690 5400 45810 5520
rect 45855 5400 45975 5520
rect 46020 5400 46140 5520
rect 46195 5400 46315 5520
rect 46360 5400 46480 5520
rect 46525 5400 46645 5520
rect 46690 5400 46810 5520
rect 46865 5400 46985 5520
rect 47030 5400 47150 5520
rect 47195 5400 47315 5520
rect 47360 5400 47480 5520
rect 47535 5400 47655 5520
rect 42175 5235 42295 5355
rect 42340 5235 42460 5355
rect 42505 5235 42625 5355
rect 42670 5235 42790 5355
rect 42845 5235 42965 5355
rect 43010 5235 43130 5355
rect 43175 5235 43295 5355
rect 43340 5235 43460 5355
rect 43515 5235 43635 5355
rect 43680 5235 43800 5355
rect 43845 5235 43965 5355
rect 44010 5235 44130 5355
rect 44185 5235 44305 5355
rect 44350 5235 44470 5355
rect 44515 5235 44635 5355
rect 44680 5235 44800 5355
rect 44855 5235 44975 5355
rect 45020 5235 45140 5355
rect 45185 5235 45305 5355
rect 45350 5235 45470 5355
rect 45525 5235 45645 5355
rect 45690 5235 45810 5355
rect 45855 5235 45975 5355
rect 46020 5235 46140 5355
rect 46195 5235 46315 5355
rect 46360 5235 46480 5355
rect 46525 5235 46645 5355
rect 46690 5235 46810 5355
rect 46865 5235 46985 5355
rect 47030 5235 47150 5355
rect 47195 5235 47315 5355
rect 47360 5235 47480 5355
rect 47535 5235 47655 5355
rect 42175 5070 42295 5190
rect 42340 5070 42460 5190
rect 42505 5070 42625 5190
rect 42670 5070 42790 5190
rect 42845 5070 42965 5190
rect 43010 5070 43130 5190
rect 43175 5070 43295 5190
rect 43340 5070 43460 5190
rect 43515 5070 43635 5190
rect 43680 5070 43800 5190
rect 43845 5070 43965 5190
rect 44010 5070 44130 5190
rect 44185 5070 44305 5190
rect 44350 5070 44470 5190
rect 44515 5070 44635 5190
rect 44680 5070 44800 5190
rect 44855 5070 44975 5190
rect 45020 5070 45140 5190
rect 45185 5070 45305 5190
rect 45350 5070 45470 5190
rect 45525 5070 45645 5190
rect 45690 5070 45810 5190
rect 45855 5070 45975 5190
rect 46020 5070 46140 5190
rect 46195 5070 46315 5190
rect 46360 5070 46480 5190
rect 46525 5070 46645 5190
rect 46690 5070 46810 5190
rect 46865 5070 46985 5190
rect 47030 5070 47150 5190
rect 47195 5070 47315 5190
rect 47360 5070 47480 5190
rect 47535 5070 47655 5190
rect 42175 4895 42295 5015
rect 42340 4895 42460 5015
rect 42505 4895 42625 5015
rect 42670 4895 42790 5015
rect 42845 4895 42965 5015
rect 43010 4895 43130 5015
rect 43175 4895 43295 5015
rect 43340 4895 43460 5015
rect 43515 4895 43635 5015
rect 43680 4895 43800 5015
rect 43845 4895 43965 5015
rect 44010 4895 44130 5015
rect 44185 4895 44305 5015
rect 44350 4895 44470 5015
rect 44515 4895 44635 5015
rect 44680 4895 44800 5015
rect 44855 4895 44975 5015
rect 45020 4895 45140 5015
rect 45185 4895 45305 5015
rect 45350 4895 45470 5015
rect 45525 4895 45645 5015
rect 45690 4895 45810 5015
rect 45855 4895 45975 5015
rect 46020 4895 46140 5015
rect 46195 4895 46315 5015
rect 46360 4895 46480 5015
rect 46525 4895 46645 5015
rect 46690 4895 46810 5015
rect 46865 4895 46985 5015
rect 47030 4895 47150 5015
rect 47195 4895 47315 5015
rect 47360 4895 47480 5015
rect 47535 4895 47655 5015
rect 42175 4730 42295 4850
rect 42340 4730 42460 4850
rect 42505 4730 42625 4850
rect 42670 4730 42790 4850
rect 42845 4730 42965 4850
rect 43010 4730 43130 4850
rect 43175 4730 43295 4850
rect 43340 4730 43460 4850
rect 43515 4730 43635 4850
rect 43680 4730 43800 4850
rect 43845 4730 43965 4850
rect 44010 4730 44130 4850
rect 44185 4730 44305 4850
rect 44350 4730 44470 4850
rect 44515 4730 44635 4850
rect 44680 4730 44800 4850
rect 44855 4730 44975 4850
rect 45020 4730 45140 4850
rect 45185 4730 45305 4850
rect 45350 4730 45470 4850
rect 45525 4730 45645 4850
rect 45690 4730 45810 4850
rect 45855 4730 45975 4850
rect 46020 4730 46140 4850
rect 46195 4730 46315 4850
rect 46360 4730 46480 4850
rect 46525 4730 46645 4850
rect 46690 4730 46810 4850
rect 46865 4730 46985 4850
rect 47030 4730 47150 4850
rect 47195 4730 47315 4850
rect 47360 4730 47480 4850
rect 47535 4730 47655 4850
rect 42175 4565 42295 4685
rect 42340 4565 42460 4685
rect 42505 4565 42625 4685
rect 42670 4565 42790 4685
rect 42845 4565 42965 4685
rect 43010 4565 43130 4685
rect 43175 4565 43295 4685
rect 43340 4565 43460 4685
rect 43515 4565 43635 4685
rect 43680 4565 43800 4685
rect 43845 4565 43965 4685
rect 44010 4565 44130 4685
rect 44185 4565 44305 4685
rect 44350 4565 44470 4685
rect 44515 4565 44635 4685
rect 44680 4565 44800 4685
rect 44855 4565 44975 4685
rect 45020 4565 45140 4685
rect 45185 4565 45305 4685
rect 45350 4565 45470 4685
rect 45525 4565 45645 4685
rect 45690 4565 45810 4685
rect 45855 4565 45975 4685
rect 46020 4565 46140 4685
rect 46195 4565 46315 4685
rect 46360 4565 46480 4685
rect 46525 4565 46645 4685
rect 46690 4565 46810 4685
rect 46865 4565 46985 4685
rect 47030 4565 47150 4685
rect 47195 4565 47315 4685
rect 47360 4565 47480 4685
rect 47535 4565 47655 4685
rect 42175 4400 42295 4520
rect 42340 4400 42460 4520
rect 42505 4400 42625 4520
rect 42670 4400 42790 4520
rect 42845 4400 42965 4520
rect 43010 4400 43130 4520
rect 43175 4400 43295 4520
rect 43340 4400 43460 4520
rect 43515 4400 43635 4520
rect 43680 4400 43800 4520
rect 43845 4400 43965 4520
rect 44010 4400 44130 4520
rect 44185 4400 44305 4520
rect 44350 4400 44470 4520
rect 44515 4400 44635 4520
rect 44680 4400 44800 4520
rect 44855 4400 44975 4520
rect 45020 4400 45140 4520
rect 45185 4400 45305 4520
rect 45350 4400 45470 4520
rect 45525 4400 45645 4520
rect 45690 4400 45810 4520
rect 45855 4400 45975 4520
rect 46020 4400 46140 4520
rect 46195 4400 46315 4520
rect 46360 4400 46480 4520
rect 46525 4400 46645 4520
rect 46690 4400 46810 4520
rect 46865 4400 46985 4520
rect 47030 4400 47150 4520
rect 47195 4400 47315 4520
rect 47360 4400 47480 4520
rect 47535 4400 47655 4520
rect 42175 4225 42295 4345
rect 42340 4225 42460 4345
rect 42505 4225 42625 4345
rect 42670 4225 42790 4345
rect 42845 4225 42965 4345
rect 43010 4225 43130 4345
rect 43175 4225 43295 4345
rect 43340 4225 43460 4345
rect 43515 4225 43635 4345
rect 43680 4225 43800 4345
rect 43845 4225 43965 4345
rect 44010 4225 44130 4345
rect 44185 4225 44305 4345
rect 44350 4225 44470 4345
rect 44515 4225 44635 4345
rect 44680 4225 44800 4345
rect 44855 4225 44975 4345
rect 45020 4225 45140 4345
rect 45185 4225 45305 4345
rect 45350 4225 45470 4345
rect 45525 4225 45645 4345
rect 45690 4225 45810 4345
rect 45855 4225 45975 4345
rect 46020 4225 46140 4345
rect 46195 4225 46315 4345
rect 46360 4225 46480 4345
rect 46525 4225 46645 4345
rect 46690 4225 46810 4345
rect 46865 4225 46985 4345
rect 47030 4225 47150 4345
rect 47195 4225 47315 4345
rect 47360 4225 47480 4345
rect 47535 4225 47655 4345
rect 42175 4060 42295 4180
rect 42340 4060 42460 4180
rect 42505 4060 42625 4180
rect 42670 4060 42790 4180
rect 42845 4060 42965 4180
rect 43010 4060 43130 4180
rect 43175 4060 43295 4180
rect 43340 4060 43460 4180
rect 43515 4060 43635 4180
rect 43680 4060 43800 4180
rect 43845 4060 43965 4180
rect 44010 4060 44130 4180
rect 44185 4060 44305 4180
rect 44350 4060 44470 4180
rect 44515 4060 44635 4180
rect 44680 4060 44800 4180
rect 44855 4060 44975 4180
rect 45020 4060 45140 4180
rect 45185 4060 45305 4180
rect 45350 4060 45470 4180
rect 45525 4060 45645 4180
rect 45690 4060 45810 4180
rect 45855 4060 45975 4180
rect 46020 4060 46140 4180
rect 46195 4060 46315 4180
rect 46360 4060 46480 4180
rect 46525 4060 46645 4180
rect 46690 4060 46810 4180
rect 46865 4060 46985 4180
rect 47030 4060 47150 4180
rect 47195 4060 47315 4180
rect 47360 4060 47480 4180
rect 47535 4060 47655 4180
rect 42175 3895 42295 4015
rect 42340 3895 42460 4015
rect 42505 3895 42625 4015
rect 42670 3895 42790 4015
rect 42845 3895 42965 4015
rect 43010 3895 43130 4015
rect 43175 3895 43295 4015
rect 43340 3895 43460 4015
rect 43515 3895 43635 4015
rect 43680 3895 43800 4015
rect 43845 3895 43965 4015
rect 44010 3895 44130 4015
rect 44185 3895 44305 4015
rect 44350 3895 44470 4015
rect 44515 3895 44635 4015
rect 44680 3895 44800 4015
rect 44855 3895 44975 4015
rect 45020 3895 45140 4015
rect 45185 3895 45305 4015
rect 45350 3895 45470 4015
rect 45525 3895 45645 4015
rect 45690 3895 45810 4015
rect 45855 3895 45975 4015
rect 46020 3895 46140 4015
rect 46195 3895 46315 4015
rect 46360 3895 46480 4015
rect 46525 3895 46645 4015
rect 46690 3895 46810 4015
rect 46865 3895 46985 4015
rect 47030 3895 47150 4015
rect 47195 3895 47315 4015
rect 47360 3895 47480 4015
rect 47535 3895 47655 4015
rect 42175 3730 42295 3850
rect 42340 3730 42460 3850
rect 42505 3730 42625 3850
rect 42670 3730 42790 3850
rect 42845 3730 42965 3850
rect 43010 3730 43130 3850
rect 43175 3730 43295 3850
rect 43340 3730 43460 3850
rect 43515 3730 43635 3850
rect 43680 3730 43800 3850
rect 43845 3730 43965 3850
rect 44010 3730 44130 3850
rect 44185 3730 44305 3850
rect 44350 3730 44470 3850
rect 44515 3730 44635 3850
rect 44680 3730 44800 3850
rect 44855 3730 44975 3850
rect 45020 3730 45140 3850
rect 45185 3730 45305 3850
rect 45350 3730 45470 3850
rect 45525 3730 45645 3850
rect 45690 3730 45810 3850
rect 45855 3730 45975 3850
rect 46020 3730 46140 3850
rect 46195 3730 46315 3850
rect 46360 3730 46480 3850
rect 46525 3730 46645 3850
rect 46690 3730 46810 3850
rect 46865 3730 46985 3850
rect 47030 3730 47150 3850
rect 47195 3730 47315 3850
rect 47360 3730 47480 3850
rect 47535 3730 47655 3850
rect 42175 3555 42295 3675
rect 42340 3555 42460 3675
rect 42505 3555 42625 3675
rect 42670 3555 42790 3675
rect 42845 3555 42965 3675
rect 43010 3555 43130 3675
rect 43175 3555 43295 3675
rect 43340 3555 43460 3675
rect 43515 3555 43635 3675
rect 43680 3555 43800 3675
rect 43845 3555 43965 3675
rect 44010 3555 44130 3675
rect 44185 3555 44305 3675
rect 44350 3555 44470 3675
rect 44515 3555 44635 3675
rect 44680 3555 44800 3675
rect 44855 3555 44975 3675
rect 45020 3555 45140 3675
rect 45185 3555 45305 3675
rect 45350 3555 45470 3675
rect 45525 3555 45645 3675
rect 45690 3555 45810 3675
rect 45855 3555 45975 3675
rect 46020 3555 46140 3675
rect 46195 3555 46315 3675
rect 46360 3555 46480 3675
rect 46525 3555 46645 3675
rect 46690 3555 46810 3675
rect 46865 3555 46985 3675
rect 47030 3555 47150 3675
rect 47195 3555 47315 3675
rect 47360 3555 47480 3675
rect 47535 3555 47655 3675
rect 42175 3390 42295 3510
rect 42340 3390 42460 3510
rect 42505 3390 42625 3510
rect 42670 3390 42790 3510
rect 42845 3390 42965 3510
rect 43010 3390 43130 3510
rect 43175 3390 43295 3510
rect 43340 3390 43460 3510
rect 43515 3390 43635 3510
rect 43680 3390 43800 3510
rect 43845 3390 43965 3510
rect 44010 3390 44130 3510
rect 44185 3390 44305 3510
rect 44350 3390 44470 3510
rect 44515 3390 44635 3510
rect 44680 3390 44800 3510
rect 44855 3390 44975 3510
rect 45020 3390 45140 3510
rect 45185 3390 45305 3510
rect 45350 3390 45470 3510
rect 45525 3390 45645 3510
rect 45690 3390 45810 3510
rect 45855 3390 45975 3510
rect 46020 3390 46140 3510
rect 46195 3390 46315 3510
rect 46360 3390 46480 3510
rect 46525 3390 46645 3510
rect 46690 3390 46810 3510
rect 46865 3390 46985 3510
rect 47030 3390 47150 3510
rect 47195 3390 47315 3510
rect 47360 3390 47480 3510
rect 47535 3390 47655 3510
rect 42175 3225 42295 3345
rect 42340 3225 42460 3345
rect 42505 3225 42625 3345
rect 42670 3225 42790 3345
rect 42845 3225 42965 3345
rect 43010 3225 43130 3345
rect 43175 3225 43295 3345
rect 43340 3225 43460 3345
rect 43515 3225 43635 3345
rect 43680 3225 43800 3345
rect 43845 3225 43965 3345
rect 44010 3225 44130 3345
rect 44185 3225 44305 3345
rect 44350 3225 44470 3345
rect 44515 3225 44635 3345
rect 44680 3225 44800 3345
rect 44855 3225 44975 3345
rect 45020 3225 45140 3345
rect 45185 3225 45305 3345
rect 45350 3225 45470 3345
rect 45525 3225 45645 3345
rect 45690 3225 45810 3345
rect 45855 3225 45975 3345
rect 46020 3225 46140 3345
rect 46195 3225 46315 3345
rect 46360 3225 46480 3345
rect 46525 3225 46645 3345
rect 46690 3225 46810 3345
rect 46865 3225 46985 3345
rect 47030 3225 47150 3345
rect 47195 3225 47315 3345
rect 47360 3225 47480 3345
rect 47535 3225 47655 3345
rect 42175 3060 42295 3180
rect 42340 3060 42460 3180
rect 42505 3060 42625 3180
rect 42670 3060 42790 3180
rect 42845 3060 42965 3180
rect 43010 3060 43130 3180
rect 43175 3060 43295 3180
rect 43340 3060 43460 3180
rect 43515 3060 43635 3180
rect 43680 3060 43800 3180
rect 43845 3060 43965 3180
rect 44010 3060 44130 3180
rect 44185 3060 44305 3180
rect 44350 3060 44470 3180
rect 44515 3060 44635 3180
rect 44680 3060 44800 3180
rect 44855 3060 44975 3180
rect 45020 3060 45140 3180
rect 45185 3060 45305 3180
rect 45350 3060 45470 3180
rect 45525 3060 45645 3180
rect 45690 3060 45810 3180
rect 45855 3060 45975 3180
rect 46020 3060 46140 3180
rect 46195 3060 46315 3180
rect 46360 3060 46480 3180
rect 46525 3060 46645 3180
rect 46690 3060 46810 3180
rect 46865 3060 46985 3180
rect 47030 3060 47150 3180
rect 47195 3060 47315 3180
rect 47360 3060 47480 3180
rect 47535 3060 47655 3180
rect 42175 2885 42295 3005
rect 42340 2885 42460 3005
rect 42505 2885 42625 3005
rect 42670 2885 42790 3005
rect 42845 2885 42965 3005
rect 43010 2885 43130 3005
rect 43175 2885 43295 3005
rect 43340 2885 43460 3005
rect 43515 2885 43635 3005
rect 43680 2885 43800 3005
rect 43845 2885 43965 3005
rect 44010 2885 44130 3005
rect 44185 2885 44305 3005
rect 44350 2885 44470 3005
rect 44515 2885 44635 3005
rect 44680 2885 44800 3005
rect 44855 2885 44975 3005
rect 45020 2885 45140 3005
rect 45185 2885 45305 3005
rect 45350 2885 45470 3005
rect 45525 2885 45645 3005
rect 45690 2885 45810 3005
rect 45855 2885 45975 3005
rect 46020 2885 46140 3005
rect 46195 2885 46315 3005
rect 46360 2885 46480 3005
rect 46525 2885 46645 3005
rect 46690 2885 46810 3005
rect 46865 2885 46985 3005
rect 47030 2885 47150 3005
rect 47195 2885 47315 3005
rect 47360 2885 47480 3005
rect 47535 2885 47655 3005
rect 42175 2720 42295 2840
rect 42340 2720 42460 2840
rect 42505 2720 42625 2840
rect 42670 2720 42790 2840
rect 42845 2720 42965 2840
rect 43010 2720 43130 2840
rect 43175 2720 43295 2840
rect 43340 2720 43460 2840
rect 43515 2720 43635 2840
rect 43680 2720 43800 2840
rect 43845 2720 43965 2840
rect 44010 2720 44130 2840
rect 44185 2720 44305 2840
rect 44350 2720 44470 2840
rect 44515 2720 44635 2840
rect 44680 2720 44800 2840
rect 44855 2720 44975 2840
rect 45020 2720 45140 2840
rect 45185 2720 45305 2840
rect 45350 2720 45470 2840
rect 45525 2720 45645 2840
rect 45690 2720 45810 2840
rect 45855 2720 45975 2840
rect 46020 2720 46140 2840
rect 46195 2720 46315 2840
rect 46360 2720 46480 2840
rect 46525 2720 46645 2840
rect 46690 2720 46810 2840
rect 46865 2720 46985 2840
rect 47030 2720 47150 2840
rect 47195 2720 47315 2840
rect 47360 2720 47480 2840
rect 47535 2720 47655 2840
rect 42175 2555 42295 2675
rect 42340 2555 42460 2675
rect 42505 2555 42625 2675
rect 42670 2555 42790 2675
rect 42845 2555 42965 2675
rect 43010 2555 43130 2675
rect 43175 2555 43295 2675
rect 43340 2555 43460 2675
rect 43515 2555 43635 2675
rect 43680 2555 43800 2675
rect 43845 2555 43965 2675
rect 44010 2555 44130 2675
rect 44185 2555 44305 2675
rect 44350 2555 44470 2675
rect 44515 2555 44635 2675
rect 44680 2555 44800 2675
rect 44855 2555 44975 2675
rect 45020 2555 45140 2675
rect 45185 2555 45305 2675
rect 45350 2555 45470 2675
rect 45525 2555 45645 2675
rect 45690 2555 45810 2675
rect 45855 2555 45975 2675
rect 46020 2555 46140 2675
rect 46195 2555 46315 2675
rect 46360 2555 46480 2675
rect 46525 2555 46645 2675
rect 46690 2555 46810 2675
rect 46865 2555 46985 2675
rect 47030 2555 47150 2675
rect 47195 2555 47315 2675
rect 47360 2555 47480 2675
rect 47535 2555 47655 2675
rect 42175 2390 42295 2510
rect 42340 2390 42460 2510
rect 42505 2390 42625 2510
rect 42670 2390 42790 2510
rect 42845 2390 42965 2510
rect 43010 2390 43130 2510
rect 43175 2390 43295 2510
rect 43340 2390 43460 2510
rect 43515 2390 43635 2510
rect 43680 2390 43800 2510
rect 43845 2390 43965 2510
rect 44010 2390 44130 2510
rect 44185 2390 44305 2510
rect 44350 2390 44470 2510
rect 44515 2390 44635 2510
rect 44680 2390 44800 2510
rect 44855 2390 44975 2510
rect 45020 2390 45140 2510
rect 45185 2390 45305 2510
rect 45350 2390 45470 2510
rect 45525 2390 45645 2510
rect 45690 2390 45810 2510
rect 45855 2390 45975 2510
rect 46020 2390 46140 2510
rect 46195 2390 46315 2510
rect 46360 2390 46480 2510
rect 46525 2390 46645 2510
rect 46690 2390 46810 2510
rect 46865 2390 46985 2510
rect 47030 2390 47150 2510
rect 47195 2390 47315 2510
rect 47360 2390 47480 2510
rect 47535 2390 47655 2510
rect 42175 2215 42295 2335
rect 42340 2215 42460 2335
rect 42505 2215 42625 2335
rect 42670 2215 42790 2335
rect 42845 2215 42965 2335
rect 43010 2215 43130 2335
rect 43175 2215 43295 2335
rect 43340 2215 43460 2335
rect 43515 2215 43635 2335
rect 43680 2215 43800 2335
rect 43845 2215 43965 2335
rect 44010 2215 44130 2335
rect 44185 2215 44305 2335
rect 44350 2215 44470 2335
rect 44515 2215 44635 2335
rect 44680 2215 44800 2335
rect 44855 2215 44975 2335
rect 45020 2215 45140 2335
rect 45185 2215 45305 2335
rect 45350 2215 45470 2335
rect 45525 2215 45645 2335
rect 45690 2215 45810 2335
rect 45855 2215 45975 2335
rect 46020 2215 46140 2335
rect 46195 2215 46315 2335
rect 46360 2215 46480 2335
rect 46525 2215 46645 2335
rect 46690 2215 46810 2335
rect 46865 2215 46985 2335
rect 47030 2215 47150 2335
rect 47195 2215 47315 2335
rect 47360 2215 47480 2335
rect 47535 2215 47655 2335
rect 42175 2050 42295 2170
rect 42340 2050 42460 2170
rect 42505 2050 42625 2170
rect 42670 2050 42790 2170
rect 42845 2050 42965 2170
rect 43010 2050 43130 2170
rect 43175 2050 43295 2170
rect 43340 2050 43460 2170
rect 43515 2050 43635 2170
rect 43680 2050 43800 2170
rect 43845 2050 43965 2170
rect 44010 2050 44130 2170
rect 44185 2050 44305 2170
rect 44350 2050 44470 2170
rect 44515 2050 44635 2170
rect 44680 2050 44800 2170
rect 44855 2050 44975 2170
rect 45020 2050 45140 2170
rect 45185 2050 45305 2170
rect 45350 2050 45470 2170
rect 45525 2050 45645 2170
rect 45690 2050 45810 2170
rect 45855 2050 45975 2170
rect 46020 2050 46140 2170
rect 46195 2050 46315 2170
rect 46360 2050 46480 2170
rect 46525 2050 46645 2170
rect 46690 2050 46810 2170
rect 46865 2050 46985 2170
rect 47030 2050 47150 2170
rect 47195 2050 47315 2170
rect 47360 2050 47480 2170
rect 47535 2050 47655 2170
rect 42175 1885 42295 2005
rect 42340 1885 42460 2005
rect 42505 1885 42625 2005
rect 42670 1885 42790 2005
rect 42845 1885 42965 2005
rect 43010 1885 43130 2005
rect 43175 1885 43295 2005
rect 43340 1885 43460 2005
rect 43515 1885 43635 2005
rect 43680 1885 43800 2005
rect 43845 1885 43965 2005
rect 44010 1885 44130 2005
rect 44185 1885 44305 2005
rect 44350 1885 44470 2005
rect 44515 1885 44635 2005
rect 44680 1885 44800 2005
rect 44855 1885 44975 2005
rect 45020 1885 45140 2005
rect 45185 1885 45305 2005
rect 45350 1885 45470 2005
rect 45525 1885 45645 2005
rect 45690 1885 45810 2005
rect 45855 1885 45975 2005
rect 46020 1885 46140 2005
rect 46195 1885 46315 2005
rect 46360 1885 46480 2005
rect 46525 1885 46645 2005
rect 46690 1885 46810 2005
rect 46865 1885 46985 2005
rect 47030 1885 47150 2005
rect 47195 1885 47315 2005
rect 47360 1885 47480 2005
rect 47535 1885 47655 2005
rect 42175 1720 42295 1840
rect 42340 1720 42460 1840
rect 42505 1720 42625 1840
rect 42670 1720 42790 1840
rect 42845 1720 42965 1840
rect 43010 1720 43130 1840
rect 43175 1720 43295 1840
rect 43340 1720 43460 1840
rect 43515 1720 43635 1840
rect 43680 1720 43800 1840
rect 43845 1720 43965 1840
rect 44010 1720 44130 1840
rect 44185 1720 44305 1840
rect 44350 1720 44470 1840
rect 44515 1720 44635 1840
rect 44680 1720 44800 1840
rect 44855 1720 44975 1840
rect 45020 1720 45140 1840
rect 45185 1720 45305 1840
rect 45350 1720 45470 1840
rect 45525 1720 45645 1840
rect 45690 1720 45810 1840
rect 45855 1720 45975 1840
rect 46020 1720 46140 1840
rect 46195 1720 46315 1840
rect 46360 1720 46480 1840
rect 46525 1720 46645 1840
rect 46690 1720 46810 1840
rect 46865 1720 46985 1840
rect 47030 1720 47150 1840
rect 47195 1720 47315 1840
rect 47360 1720 47480 1840
rect 47535 1720 47655 1840
rect 47865 7080 47985 7200
rect 48030 7080 48150 7200
rect 48195 7080 48315 7200
rect 48360 7080 48480 7200
rect 48535 7080 48655 7200
rect 48700 7080 48820 7200
rect 48865 7080 48985 7200
rect 49030 7080 49150 7200
rect 49205 7080 49325 7200
rect 49370 7080 49490 7200
rect 49535 7080 49655 7200
rect 49700 7080 49820 7200
rect 49875 7080 49995 7200
rect 50040 7080 50160 7200
rect 50205 7080 50325 7200
rect 50370 7080 50490 7200
rect 50545 7080 50665 7200
rect 50710 7080 50830 7200
rect 50875 7080 50995 7200
rect 51040 7080 51160 7200
rect 51215 7080 51335 7200
rect 51380 7080 51500 7200
rect 51545 7080 51665 7200
rect 51710 7080 51830 7200
rect 51885 7080 52005 7200
rect 52050 7080 52170 7200
rect 52215 7080 52335 7200
rect 52380 7080 52500 7200
rect 52555 7080 52675 7200
rect 52720 7080 52840 7200
rect 52885 7080 53005 7200
rect 53050 7080 53170 7200
rect 53225 7080 53345 7200
rect 47865 6905 47985 7025
rect 48030 6905 48150 7025
rect 48195 6905 48315 7025
rect 48360 6905 48480 7025
rect 48535 6905 48655 7025
rect 48700 6905 48820 7025
rect 48865 6905 48985 7025
rect 49030 6905 49150 7025
rect 49205 6905 49325 7025
rect 49370 6905 49490 7025
rect 49535 6905 49655 7025
rect 49700 6905 49820 7025
rect 49875 6905 49995 7025
rect 50040 6905 50160 7025
rect 50205 6905 50325 7025
rect 50370 6905 50490 7025
rect 50545 6905 50665 7025
rect 50710 6905 50830 7025
rect 50875 6905 50995 7025
rect 51040 6905 51160 7025
rect 51215 6905 51335 7025
rect 51380 6905 51500 7025
rect 51545 6905 51665 7025
rect 51710 6905 51830 7025
rect 51885 6905 52005 7025
rect 52050 6905 52170 7025
rect 52215 6905 52335 7025
rect 52380 6905 52500 7025
rect 52555 6905 52675 7025
rect 52720 6905 52840 7025
rect 52885 6905 53005 7025
rect 53050 6905 53170 7025
rect 53225 6905 53345 7025
rect 47865 6740 47985 6860
rect 48030 6740 48150 6860
rect 48195 6740 48315 6860
rect 48360 6740 48480 6860
rect 48535 6740 48655 6860
rect 48700 6740 48820 6860
rect 48865 6740 48985 6860
rect 49030 6740 49150 6860
rect 49205 6740 49325 6860
rect 49370 6740 49490 6860
rect 49535 6740 49655 6860
rect 49700 6740 49820 6860
rect 49875 6740 49995 6860
rect 50040 6740 50160 6860
rect 50205 6740 50325 6860
rect 50370 6740 50490 6860
rect 50545 6740 50665 6860
rect 50710 6740 50830 6860
rect 50875 6740 50995 6860
rect 51040 6740 51160 6860
rect 51215 6740 51335 6860
rect 51380 6740 51500 6860
rect 51545 6740 51665 6860
rect 51710 6740 51830 6860
rect 51885 6740 52005 6860
rect 52050 6740 52170 6860
rect 52215 6740 52335 6860
rect 52380 6740 52500 6860
rect 52555 6740 52675 6860
rect 52720 6740 52840 6860
rect 52885 6740 53005 6860
rect 53050 6740 53170 6860
rect 53225 6740 53345 6860
rect 47865 6575 47985 6695
rect 48030 6575 48150 6695
rect 48195 6575 48315 6695
rect 48360 6575 48480 6695
rect 48535 6575 48655 6695
rect 48700 6575 48820 6695
rect 48865 6575 48985 6695
rect 49030 6575 49150 6695
rect 49205 6575 49325 6695
rect 49370 6575 49490 6695
rect 49535 6575 49655 6695
rect 49700 6575 49820 6695
rect 49875 6575 49995 6695
rect 50040 6575 50160 6695
rect 50205 6575 50325 6695
rect 50370 6575 50490 6695
rect 50545 6575 50665 6695
rect 50710 6575 50830 6695
rect 50875 6575 50995 6695
rect 51040 6575 51160 6695
rect 51215 6575 51335 6695
rect 51380 6575 51500 6695
rect 51545 6575 51665 6695
rect 51710 6575 51830 6695
rect 51885 6575 52005 6695
rect 52050 6575 52170 6695
rect 52215 6575 52335 6695
rect 52380 6575 52500 6695
rect 52555 6575 52675 6695
rect 52720 6575 52840 6695
rect 52885 6575 53005 6695
rect 53050 6575 53170 6695
rect 53225 6575 53345 6695
rect 47865 6410 47985 6530
rect 48030 6410 48150 6530
rect 48195 6410 48315 6530
rect 48360 6410 48480 6530
rect 48535 6410 48655 6530
rect 48700 6410 48820 6530
rect 48865 6410 48985 6530
rect 49030 6410 49150 6530
rect 49205 6410 49325 6530
rect 49370 6410 49490 6530
rect 49535 6410 49655 6530
rect 49700 6410 49820 6530
rect 49875 6410 49995 6530
rect 50040 6410 50160 6530
rect 50205 6410 50325 6530
rect 50370 6410 50490 6530
rect 50545 6410 50665 6530
rect 50710 6410 50830 6530
rect 50875 6410 50995 6530
rect 51040 6410 51160 6530
rect 51215 6410 51335 6530
rect 51380 6410 51500 6530
rect 51545 6410 51665 6530
rect 51710 6410 51830 6530
rect 51885 6410 52005 6530
rect 52050 6410 52170 6530
rect 52215 6410 52335 6530
rect 52380 6410 52500 6530
rect 52555 6410 52675 6530
rect 52720 6410 52840 6530
rect 52885 6410 53005 6530
rect 53050 6410 53170 6530
rect 53225 6410 53345 6530
rect 47865 6235 47985 6355
rect 48030 6235 48150 6355
rect 48195 6235 48315 6355
rect 48360 6235 48480 6355
rect 48535 6235 48655 6355
rect 48700 6235 48820 6355
rect 48865 6235 48985 6355
rect 49030 6235 49150 6355
rect 49205 6235 49325 6355
rect 49370 6235 49490 6355
rect 49535 6235 49655 6355
rect 49700 6235 49820 6355
rect 49875 6235 49995 6355
rect 50040 6235 50160 6355
rect 50205 6235 50325 6355
rect 50370 6235 50490 6355
rect 50545 6235 50665 6355
rect 50710 6235 50830 6355
rect 50875 6235 50995 6355
rect 51040 6235 51160 6355
rect 51215 6235 51335 6355
rect 51380 6235 51500 6355
rect 51545 6235 51665 6355
rect 51710 6235 51830 6355
rect 51885 6235 52005 6355
rect 52050 6235 52170 6355
rect 52215 6235 52335 6355
rect 52380 6235 52500 6355
rect 52555 6235 52675 6355
rect 52720 6235 52840 6355
rect 52885 6235 53005 6355
rect 53050 6235 53170 6355
rect 53225 6235 53345 6355
rect 47865 6070 47985 6190
rect 48030 6070 48150 6190
rect 48195 6070 48315 6190
rect 48360 6070 48480 6190
rect 48535 6070 48655 6190
rect 48700 6070 48820 6190
rect 48865 6070 48985 6190
rect 49030 6070 49150 6190
rect 49205 6070 49325 6190
rect 49370 6070 49490 6190
rect 49535 6070 49655 6190
rect 49700 6070 49820 6190
rect 49875 6070 49995 6190
rect 50040 6070 50160 6190
rect 50205 6070 50325 6190
rect 50370 6070 50490 6190
rect 50545 6070 50665 6190
rect 50710 6070 50830 6190
rect 50875 6070 50995 6190
rect 51040 6070 51160 6190
rect 51215 6070 51335 6190
rect 51380 6070 51500 6190
rect 51545 6070 51665 6190
rect 51710 6070 51830 6190
rect 51885 6070 52005 6190
rect 52050 6070 52170 6190
rect 52215 6070 52335 6190
rect 52380 6070 52500 6190
rect 52555 6070 52675 6190
rect 52720 6070 52840 6190
rect 52885 6070 53005 6190
rect 53050 6070 53170 6190
rect 53225 6070 53345 6190
rect 47865 5905 47985 6025
rect 48030 5905 48150 6025
rect 48195 5905 48315 6025
rect 48360 5905 48480 6025
rect 48535 5905 48655 6025
rect 48700 5905 48820 6025
rect 48865 5905 48985 6025
rect 49030 5905 49150 6025
rect 49205 5905 49325 6025
rect 49370 5905 49490 6025
rect 49535 5905 49655 6025
rect 49700 5905 49820 6025
rect 49875 5905 49995 6025
rect 50040 5905 50160 6025
rect 50205 5905 50325 6025
rect 50370 5905 50490 6025
rect 50545 5905 50665 6025
rect 50710 5905 50830 6025
rect 50875 5905 50995 6025
rect 51040 5905 51160 6025
rect 51215 5905 51335 6025
rect 51380 5905 51500 6025
rect 51545 5905 51665 6025
rect 51710 5905 51830 6025
rect 51885 5905 52005 6025
rect 52050 5905 52170 6025
rect 52215 5905 52335 6025
rect 52380 5905 52500 6025
rect 52555 5905 52675 6025
rect 52720 5905 52840 6025
rect 52885 5905 53005 6025
rect 53050 5905 53170 6025
rect 53225 5905 53345 6025
rect 47865 5740 47985 5860
rect 48030 5740 48150 5860
rect 48195 5740 48315 5860
rect 48360 5740 48480 5860
rect 48535 5740 48655 5860
rect 48700 5740 48820 5860
rect 48865 5740 48985 5860
rect 49030 5740 49150 5860
rect 49205 5740 49325 5860
rect 49370 5740 49490 5860
rect 49535 5740 49655 5860
rect 49700 5740 49820 5860
rect 49875 5740 49995 5860
rect 50040 5740 50160 5860
rect 50205 5740 50325 5860
rect 50370 5740 50490 5860
rect 50545 5740 50665 5860
rect 50710 5740 50830 5860
rect 50875 5740 50995 5860
rect 51040 5740 51160 5860
rect 51215 5740 51335 5860
rect 51380 5740 51500 5860
rect 51545 5740 51665 5860
rect 51710 5740 51830 5860
rect 51885 5740 52005 5860
rect 52050 5740 52170 5860
rect 52215 5740 52335 5860
rect 52380 5740 52500 5860
rect 52555 5740 52675 5860
rect 52720 5740 52840 5860
rect 52885 5740 53005 5860
rect 53050 5740 53170 5860
rect 53225 5740 53345 5860
rect 47865 5565 47985 5685
rect 48030 5565 48150 5685
rect 48195 5565 48315 5685
rect 48360 5565 48480 5685
rect 48535 5565 48655 5685
rect 48700 5565 48820 5685
rect 48865 5565 48985 5685
rect 49030 5565 49150 5685
rect 49205 5565 49325 5685
rect 49370 5565 49490 5685
rect 49535 5565 49655 5685
rect 49700 5565 49820 5685
rect 49875 5565 49995 5685
rect 50040 5565 50160 5685
rect 50205 5565 50325 5685
rect 50370 5565 50490 5685
rect 50545 5565 50665 5685
rect 50710 5565 50830 5685
rect 50875 5565 50995 5685
rect 51040 5565 51160 5685
rect 51215 5565 51335 5685
rect 51380 5565 51500 5685
rect 51545 5565 51665 5685
rect 51710 5565 51830 5685
rect 51885 5565 52005 5685
rect 52050 5565 52170 5685
rect 52215 5565 52335 5685
rect 52380 5565 52500 5685
rect 52555 5565 52675 5685
rect 52720 5565 52840 5685
rect 52885 5565 53005 5685
rect 53050 5565 53170 5685
rect 53225 5565 53345 5685
rect 47865 5400 47985 5520
rect 48030 5400 48150 5520
rect 48195 5400 48315 5520
rect 48360 5400 48480 5520
rect 48535 5400 48655 5520
rect 48700 5400 48820 5520
rect 48865 5400 48985 5520
rect 49030 5400 49150 5520
rect 49205 5400 49325 5520
rect 49370 5400 49490 5520
rect 49535 5400 49655 5520
rect 49700 5400 49820 5520
rect 49875 5400 49995 5520
rect 50040 5400 50160 5520
rect 50205 5400 50325 5520
rect 50370 5400 50490 5520
rect 50545 5400 50665 5520
rect 50710 5400 50830 5520
rect 50875 5400 50995 5520
rect 51040 5400 51160 5520
rect 51215 5400 51335 5520
rect 51380 5400 51500 5520
rect 51545 5400 51665 5520
rect 51710 5400 51830 5520
rect 51885 5400 52005 5520
rect 52050 5400 52170 5520
rect 52215 5400 52335 5520
rect 52380 5400 52500 5520
rect 52555 5400 52675 5520
rect 52720 5400 52840 5520
rect 52885 5400 53005 5520
rect 53050 5400 53170 5520
rect 53225 5400 53345 5520
rect 47865 5235 47985 5355
rect 48030 5235 48150 5355
rect 48195 5235 48315 5355
rect 48360 5235 48480 5355
rect 48535 5235 48655 5355
rect 48700 5235 48820 5355
rect 48865 5235 48985 5355
rect 49030 5235 49150 5355
rect 49205 5235 49325 5355
rect 49370 5235 49490 5355
rect 49535 5235 49655 5355
rect 49700 5235 49820 5355
rect 49875 5235 49995 5355
rect 50040 5235 50160 5355
rect 50205 5235 50325 5355
rect 50370 5235 50490 5355
rect 50545 5235 50665 5355
rect 50710 5235 50830 5355
rect 50875 5235 50995 5355
rect 51040 5235 51160 5355
rect 51215 5235 51335 5355
rect 51380 5235 51500 5355
rect 51545 5235 51665 5355
rect 51710 5235 51830 5355
rect 51885 5235 52005 5355
rect 52050 5235 52170 5355
rect 52215 5235 52335 5355
rect 52380 5235 52500 5355
rect 52555 5235 52675 5355
rect 52720 5235 52840 5355
rect 52885 5235 53005 5355
rect 53050 5235 53170 5355
rect 53225 5235 53345 5355
rect 47865 5070 47985 5190
rect 48030 5070 48150 5190
rect 48195 5070 48315 5190
rect 48360 5070 48480 5190
rect 48535 5070 48655 5190
rect 48700 5070 48820 5190
rect 48865 5070 48985 5190
rect 49030 5070 49150 5190
rect 49205 5070 49325 5190
rect 49370 5070 49490 5190
rect 49535 5070 49655 5190
rect 49700 5070 49820 5190
rect 49875 5070 49995 5190
rect 50040 5070 50160 5190
rect 50205 5070 50325 5190
rect 50370 5070 50490 5190
rect 50545 5070 50665 5190
rect 50710 5070 50830 5190
rect 50875 5070 50995 5190
rect 51040 5070 51160 5190
rect 51215 5070 51335 5190
rect 51380 5070 51500 5190
rect 51545 5070 51665 5190
rect 51710 5070 51830 5190
rect 51885 5070 52005 5190
rect 52050 5070 52170 5190
rect 52215 5070 52335 5190
rect 52380 5070 52500 5190
rect 52555 5070 52675 5190
rect 52720 5070 52840 5190
rect 52885 5070 53005 5190
rect 53050 5070 53170 5190
rect 53225 5070 53345 5190
rect 47865 4895 47985 5015
rect 48030 4895 48150 5015
rect 48195 4895 48315 5015
rect 48360 4895 48480 5015
rect 48535 4895 48655 5015
rect 48700 4895 48820 5015
rect 48865 4895 48985 5015
rect 49030 4895 49150 5015
rect 49205 4895 49325 5015
rect 49370 4895 49490 5015
rect 49535 4895 49655 5015
rect 49700 4895 49820 5015
rect 49875 4895 49995 5015
rect 50040 4895 50160 5015
rect 50205 4895 50325 5015
rect 50370 4895 50490 5015
rect 50545 4895 50665 5015
rect 50710 4895 50830 5015
rect 50875 4895 50995 5015
rect 51040 4895 51160 5015
rect 51215 4895 51335 5015
rect 51380 4895 51500 5015
rect 51545 4895 51665 5015
rect 51710 4895 51830 5015
rect 51885 4895 52005 5015
rect 52050 4895 52170 5015
rect 52215 4895 52335 5015
rect 52380 4895 52500 5015
rect 52555 4895 52675 5015
rect 52720 4895 52840 5015
rect 52885 4895 53005 5015
rect 53050 4895 53170 5015
rect 53225 4895 53345 5015
rect 47865 4730 47985 4850
rect 48030 4730 48150 4850
rect 48195 4730 48315 4850
rect 48360 4730 48480 4850
rect 48535 4730 48655 4850
rect 48700 4730 48820 4850
rect 48865 4730 48985 4850
rect 49030 4730 49150 4850
rect 49205 4730 49325 4850
rect 49370 4730 49490 4850
rect 49535 4730 49655 4850
rect 49700 4730 49820 4850
rect 49875 4730 49995 4850
rect 50040 4730 50160 4850
rect 50205 4730 50325 4850
rect 50370 4730 50490 4850
rect 50545 4730 50665 4850
rect 50710 4730 50830 4850
rect 50875 4730 50995 4850
rect 51040 4730 51160 4850
rect 51215 4730 51335 4850
rect 51380 4730 51500 4850
rect 51545 4730 51665 4850
rect 51710 4730 51830 4850
rect 51885 4730 52005 4850
rect 52050 4730 52170 4850
rect 52215 4730 52335 4850
rect 52380 4730 52500 4850
rect 52555 4730 52675 4850
rect 52720 4730 52840 4850
rect 52885 4730 53005 4850
rect 53050 4730 53170 4850
rect 53225 4730 53345 4850
rect 47865 4565 47985 4685
rect 48030 4565 48150 4685
rect 48195 4565 48315 4685
rect 48360 4565 48480 4685
rect 48535 4565 48655 4685
rect 48700 4565 48820 4685
rect 48865 4565 48985 4685
rect 49030 4565 49150 4685
rect 49205 4565 49325 4685
rect 49370 4565 49490 4685
rect 49535 4565 49655 4685
rect 49700 4565 49820 4685
rect 49875 4565 49995 4685
rect 50040 4565 50160 4685
rect 50205 4565 50325 4685
rect 50370 4565 50490 4685
rect 50545 4565 50665 4685
rect 50710 4565 50830 4685
rect 50875 4565 50995 4685
rect 51040 4565 51160 4685
rect 51215 4565 51335 4685
rect 51380 4565 51500 4685
rect 51545 4565 51665 4685
rect 51710 4565 51830 4685
rect 51885 4565 52005 4685
rect 52050 4565 52170 4685
rect 52215 4565 52335 4685
rect 52380 4565 52500 4685
rect 52555 4565 52675 4685
rect 52720 4565 52840 4685
rect 52885 4565 53005 4685
rect 53050 4565 53170 4685
rect 53225 4565 53345 4685
rect 47865 4400 47985 4520
rect 48030 4400 48150 4520
rect 48195 4400 48315 4520
rect 48360 4400 48480 4520
rect 48535 4400 48655 4520
rect 48700 4400 48820 4520
rect 48865 4400 48985 4520
rect 49030 4400 49150 4520
rect 49205 4400 49325 4520
rect 49370 4400 49490 4520
rect 49535 4400 49655 4520
rect 49700 4400 49820 4520
rect 49875 4400 49995 4520
rect 50040 4400 50160 4520
rect 50205 4400 50325 4520
rect 50370 4400 50490 4520
rect 50545 4400 50665 4520
rect 50710 4400 50830 4520
rect 50875 4400 50995 4520
rect 51040 4400 51160 4520
rect 51215 4400 51335 4520
rect 51380 4400 51500 4520
rect 51545 4400 51665 4520
rect 51710 4400 51830 4520
rect 51885 4400 52005 4520
rect 52050 4400 52170 4520
rect 52215 4400 52335 4520
rect 52380 4400 52500 4520
rect 52555 4400 52675 4520
rect 52720 4400 52840 4520
rect 52885 4400 53005 4520
rect 53050 4400 53170 4520
rect 53225 4400 53345 4520
rect 47865 4225 47985 4345
rect 48030 4225 48150 4345
rect 48195 4225 48315 4345
rect 48360 4225 48480 4345
rect 48535 4225 48655 4345
rect 48700 4225 48820 4345
rect 48865 4225 48985 4345
rect 49030 4225 49150 4345
rect 49205 4225 49325 4345
rect 49370 4225 49490 4345
rect 49535 4225 49655 4345
rect 49700 4225 49820 4345
rect 49875 4225 49995 4345
rect 50040 4225 50160 4345
rect 50205 4225 50325 4345
rect 50370 4225 50490 4345
rect 50545 4225 50665 4345
rect 50710 4225 50830 4345
rect 50875 4225 50995 4345
rect 51040 4225 51160 4345
rect 51215 4225 51335 4345
rect 51380 4225 51500 4345
rect 51545 4225 51665 4345
rect 51710 4225 51830 4345
rect 51885 4225 52005 4345
rect 52050 4225 52170 4345
rect 52215 4225 52335 4345
rect 52380 4225 52500 4345
rect 52555 4225 52675 4345
rect 52720 4225 52840 4345
rect 52885 4225 53005 4345
rect 53050 4225 53170 4345
rect 53225 4225 53345 4345
rect 47865 4060 47985 4180
rect 48030 4060 48150 4180
rect 48195 4060 48315 4180
rect 48360 4060 48480 4180
rect 48535 4060 48655 4180
rect 48700 4060 48820 4180
rect 48865 4060 48985 4180
rect 49030 4060 49150 4180
rect 49205 4060 49325 4180
rect 49370 4060 49490 4180
rect 49535 4060 49655 4180
rect 49700 4060 49820 4180
rect 49875 4060 49995 4180
rect 50040 4060 50160 4180
rect 50205 4060 50325 4180
rect 50370 4060 50490 4180
rect 50545 4060 50665 4180
rect 50710 4060 50830 4180
rect 50875 4060 50995 4180
rect 51040 4060 51160 4180
rect 51215 4060 51335 4180
rect 51380 4060 51500 4180
rect 51545 4060 51665 4180
rect 51710 4060 51830 4180
rect 51885 4060 52005 4180
rect 52050 4060 52170 4180
rect 52215 4060 52335 4180
rect 52380 4060 52500 4180
rect 52555 4060 52675 4180
rect 52720 4060 52840 4180
rect 52885 4060 53005 4180
rect 53050 4060 53170 4180
rect 53225 4060 53345 4180
rect 47865 3895 47985 4015
rect 48030 3895 48150 4015
rect 48195 3895 48315 4015
rect 48360 3895 48480 4015
rect 48535 3895 48655 4015
rect 48700 3895 48820 4015
rect 48865 3895 48985 4015
rect 49030 3895 49150 4015
rect 49205 3895 49325 4015
rect 49370 3895 49490 4015
rect 49535 3895 49655 4015
rect 49700 3895 49820 4015
rect 49875 3895 49995 4015
rect 50040 3895 50160 4015
rect 50205 3895 50325 4015
rect 50370 3895 50490 4015
rect 50545 3895 50665 4015
rect 50710 3895 50830 4015
rect 50875 3895 50995 4015
rect 51040 3895 51160 4015
rect 51215 3895 51335 4015
rect 51380 3895 51500 4015
rect 51545 3895 51665 4015
rect 51710 3895 51830 4015
rect 51885 3895 52005 4015
rect 52050 3895 52170 4015
rect 52215 3895 52335 4015
rect 52380 3895 52500 4015
rect 52555 3895 52675 4015
rect 52720 3895 52840 4015
rect 52885 3895 53005 4015
rect 53050 3895 53170 4015
rect 53225 3895 53345 4015
rect 47865 3730 47985 3850
rect 48030 3730 48150 3850
rect 48195 3730 48315 3850
rect 48360 3730 48480 3850
rect 48535 3730 48655 3850
rect 48700 3730 48820 3850
rect 48865 3730 48985 3850
rect 49030 3730 49150 3850
rect 49205 3730 49325 3850
rect 49370 3730 49490 3850
rect 49535 3730 49655 3850
rect 49700 3730 49820 3850
rect 49875 3730 49995 3850
rect 50040 3730 50160 3850
rect 50205 3730 50325 3850
rect 50370 3730 50490 3850
rect 50545 3730 50665 3850
rect 50710 3730 50830 3850
rect 50875 3730 50995 3850
rect 51040 3730 51160 3850
rect 51215 3730 51335 3850
rect 51380 3730 51500 3850
rect 51545 3730 51665 3850
rect 51710 3730 51830 3850
rect 51885 3730 52005 3850
rect 52050 3730 52170 3850
rect 52215 3730 52335 3850
rect 52380 3730 52500 3850
rect 52555 3730 52675 3850
rect 52720 3730 52840 3850
rect 52885 3730 53005 3850
rect 53050 3730 53170 3850
rect 53225 3730 53345 3850
rect 47865 3555 47985 3675
rect 48030 3555 48150 3675
rect 48195 3555 48315 3675
rect 48360 3555 48480 3675
rect 48535 3555 48655 3675
rect 48700 3555 48820 3675
rect 48865 3555 48985 3675
rect 49030 3555 49150 3675
rect 49205 3555 49325 3675
rect 49370 3555 49490 3675
rect 49535 3555 49655 3675
rect 49700 3555 49820 3675
rect 49875 3555 49995 3675
rect 50040 3555 50160 3675
rect 50205 3555 50325 3675
rect 50370 3555 50490 3675
rect 50545 3555 50665 3675
rect 50710 3555 50830 3675
rect 50875 3555 50995 3675
rect 51040 3555 51160 3675
rect 51215 3555 51335 3675
rect 51380 3555 51500 3675
rect 51545 3555 51665 3675
rect 51710 3555 51830 3675
rect 51885 3555 52005 3675
rect 52050 3555 52170 3675
rect 52215 3555 52335 3675
rect 52380 3555 52500 3675
rect 52555 3555 52675 3675
rect 52720 3555 52840 3675
rect 52885 3555 53005 3675
rect 53050 3555 53170 3675
rect 53225 3555 53345 3675
rect 47865 3390 47985 3510
rect 48030 3390 48150 3510
rect 48195 3390 48315 3510
rect 48360 3390 48480 3510
rect 48535 3390 48655 3510
rect 48700 3390 48820 3510
rect 48865 3390 48985 3510
rect 49030 3390 49150 3510
rect 49205 3390 49325 3510
rect 49370 3390 49490 3510
rect 49535 3390 49655 3510
rect 49700 3390 49820 3510
rect 49875 3390 49995 3510
rect 50040 3390 50160 3510
rect 50205 3390 50325 3510
rect 50370 3390 50490 3510
rect 50545 3390 50665 3510
rect 50710 3390 50830 3510
rect 50875 3390 50995 3510
rect 51040 3390 51160 3510
rect 51215 3390 51335 3510
rect 51380 3390 51500 3510
rect 51545 3390 51665 3510
rect 51710 3390 51830 3510
rect 51885 3390 52005 3510
rect 52050 3390 52170 3510
rect 52215 3390 52335 3510
rect 52380 3390 52500 3510
rect 52555 3390 52675 3510
rect 52720 3390 52840 3510
rect 52885 3390 53005 3510
rect 53050 3390 53170 3510
rect 53225 3390 53345 3510
rect 47865 3225 47985 3345
rect 48030 3225 48150 3345
rect 48195 3225 48315 3345
rect 48360 3225 48480 3345
rect 48535 3225 48655 3345
rect 48700 3225 48820 3345
rect 48865 3225 48985 3345
rect 49030 3225 49150 3345
rect 49205 3225 49325 3345
rect 49370 3225 49490 3345
rect 49535 3225 49655 3345
rect 49700 3225 49820 3345
rect 49875 3225 49995 3345
rect 50040 3225 50160 3345
rect 50205 3225 50325 3345
rect 50370 3225 50490 3345
rect 50545 3225 50665 3345
rect 50710 3225 50830 3345
rect 50875 3225 50995 3345
rect 51040 3225 51160 3345
rect 51215 3225 51335 3345
rect 51380 3225 51500 3345
rect 51545 3225 51665 3345
rect 51710 3225 51830 3345
rect 51885 3225 52005 3345
rect 52050 3225 52170 3345
rect 52215 3225 52335 3345
rect 52380 3225 52500 3345
rect 52555 3225 52675 3345
rect 52720 3225 52840 3345
rect 52885 3225 53005 3345
rect 53050 3225 53170 3345
rect 53225 3225 53345 3345
rect 47865 3060 47985 3180
rect 48030 3060 48150 3180
rect 48195 3060 48315 3180
rect 48360 3060 48480 3180
rect 48535 3060 48655 3180
rect 48700 3060 48820 3180
rect 48865 3060 48985 3180
rect 49030 3060 49150 3180
rect 49205 3060 49325 3180
rect 49370 3060 49490 3180
rect 49535 3060 49655 3180
rect 49700 3060 49820 3180
rect 49875 3060 49995 3180
rect 50040 3060 50160 3180
rect 50205 3060 50325 3180
rect 50370 3060 50490 3180
rect 50545 3060 50665 3180
rect 50710 3060 50830 3180
rect 50875 3060 50995 3180
rect 51040 3060 51160 3180
rect 51215 3060 51335 3180
rect 51380 3060 51500 3180
rect 51545 3060 51665 3180
rect 51710 3060 51830 3180
rect 51885 3060 52005 3180
rect 52050 3060 52170 3180
rect 52215 3060 52335 3180
rect 52380 3060 52500 3180
rect 52555 3060 52675 3180
rect 52720 3060 52840 3180
rect 52885 3060 53005 3180
rect 53050 3060 53170 3180
rect 53225 3060 53345 3180
rect 47865 2885 47985 3005
rect 48030 2885 48150 3005
rect 48195 2885 48315 3005
rect 48360 2885 48480 3005
rect 48535 2885 48655 3005
rect 48700 2885 48820 3005
rect 48865 2885 48985 3005
rect 49030 2885 49150 3005
rect 49205 2885 49325 3005
rect 49370 2885 49490 3005
rect 49535 2885 49655 3005
rect 49700 2885 49820 3005
rect 49875 2885 49995 3005
rect 50040 2885 50160 3005
rect 50205 2885 50325 3005
rect 50370 2885 50490 3005
rect 50545 2885 50665 3005
rect 50710 2885 50830 3005
rect 50875 2885 50995 3005
rect 51040 2885 51160 3005
rect 51215 2885 51335 3005
rect 51380 2885 51500 3005
rect 51545 2885 51665 3005
rect 51710 2885 51830 3005
rect 51885 2885 52005 3005
rect 52050 2885 52170 3005
rect 52215 2885 52335 3005
rect 52380 2885 52500 3005
rect 52555 2885 52675 3005
rect 52720 2885 52840 3005
rect 52885 2885 53005 3005
rect 53050 2885 53170 3005
rect 53225 2885 53345 3005
rect 47865 2720 47985 2840
rect 48030 2720 48150 2840
rect 48195 2720 48315 2840
rect 48360 2720 48480 2840
rect 48535 2720 48655 2840
rect 48700 2720 48820 2840
rect 48865 2720 48985 2840
rect 49030 2720 49150 2840
rect 49205 2720 49325 2840
rect 49370 2720 49490 2840
rect 49535 2720 49655 2840
rect 49700 2720 49820 2840
rect 49875 2720 49995 2840
rect 50040 2720 50160 2840
rect 50205 2720 50325 2840
rect 50370 2720 50490 2840
rect 50545 2720 50665 2840
rect 50710 2720 50830 2840
rect 50875 2720 50995 2840
rect 51040 2720 51160 2840
rect 51215 2720 51335 2840
rect 51380 2720 51500 2840
rect 51545 2720 51665 2840
rect 51710 2720 51830 2840
rect 51885 2720 52005 2840
rect 52050 2720 52170 2840
rect 52215 2720 52335 2840
rect 52380 2720 52500 2840
rect 52555 2720 52675 2840
rect 52720 2720 52840 2840
rect 52885 2720 53005 2840
rect 53050 2720 53170 2840
rect 53225 2720 53345 2840
rect 47865 2555 47985 2675
rect 48030 2555 48150 2675
rect 48195 2555 48315 2675
rect 48360 2555 48480 2675
rect 48535 2555 48655 2675
rect 48700 2555 48820 2675
rect 48865 2555 48985 2675
rect 49030 2555 49150 2675
rect 49205 2555 49325 2675
rect 49370 2555 49490 2675
rect 49535 2555 49655 2675
rect 49700 2555 49820 2675
rect 49875 2555 49995 2675
rect 50040 2555 50160 2675
rect 50205 2555 50325 2675
rect 50370 2555 50490 2675
rect 50545 2555 50665 2675
rect 50710 2555 50830 2675
rect 50875 2555 50995 2675
rect 51040 2555 51160 2675
rect 51215 2555 51335 2675
rect 51380 2555 51500 2675
rect 51545 2555 51665 2675
rect 51710 2555 51830 2675
rect 51885 2555 52005 2675
rect 52050 2555 52170 2675
rect 52215 2555 52335 2675
rect 52380 2555 52500 2675
rect 52555 2555 52675 2675
rect 52720 2555 52840 2675
rect 52885 2555 53005 2675
rect 53050 2555 53170 2675
rect 53225 2555 53345 2675
rect 47865 2390 47985 2510
rect 48030 2390 48150 2510
rect 48195 2390 48315 2510
rect 48360 2390 48480 2510
rect 48535 2390 48655 2510
rect 48700 2390 48820 2510
rect 48865 2390 48985 2510
rect 49030 2390 49150 2510
rect 49205 2390 49325 2510
rect 49370 2390 49490 2510
rect 49535 2390 49655 2510
rect 49700 2390 49820 2510
rect 49875 2390 49995 2510
rect 50040 2390 50160 2510
rect 50205 2390 50325 2510
rect 50370 2390 50490 2510
rect 50545 2390 50665 2510
rect 50710 2390 50830 2510
rect 50875 2390 50995 2510
rect 51040 2390 51160 2510
rect 51215 2390 51335 2510
rect 51380 2390 51500 2510
rect 51545 2390 51665 2510
rect 51710 2390 51830 2510
rect 51885 2390 52005 2510
rect 52050 2390 52170 2510
rect 52215 2390 52335 2510
rect 52380 2390 52500 2510
rect 52555 2390 52675 2510
rect 52720 2390 52840 2510
rect 52885 2390 53005 2510
rect 53050 2390 53170 2510
rect 53225 2390 53345 2510
rect 47865 2215 47985 2335
rect 48030 2215 48150 2335
rect 48195 2215 48315 2335
rect 48360 2215 48480 2335
rect 48535 2215 48655 2335
rect 48700 2215 48820 2335
rect 48865 2215 48985 2335
rect 49030 2215 49150 2335
rect 49205 2215 49325 2335
rect 49370 2215 49490 2335
rect 49535 2215 49655 2335
rect 49700 2215 49820 2335
rect 49875 2215 49995 2335
rect 50040 2215 50160 2335
rect 50205 2215 50325 2335
rect 50370 2215 50490 2335
rect 50545 2215 50665 2335
rect 50710 2215 50830 2335
rect 50875 2215 50995 2335
rect 51040 2215 51160 2335
rect 51215 2215 51335 2335
rect 51380 2215 51500 2335
rect 51545 2215 51665 2335
rect 51710 2215 51830 2335
rect 51885 2215 52005 2335
rect 52050 2215 52170 2335
rect 52215 2215 52335 2335
rect 52380 2215 52500 2335
rect 52555 2215 52675 2335
rect 52720 2215 52840 2335
rect 52885 2215 53005 2335
rect 53050 2215 53170 2335
rect 53225 2215 53345 2335
rect 47865 2050 47985 2170
rect 48030 2050 48150 2170
rect 48195 2050 48315 2170
rect 48360 2050 48480 2170
rect 48535 2050 48655 2170
rect 48700 2050 48820 2170
rect 48865 2050 48985 2170
rect 49030 2050 49150 2170
rect 49205 2050 49325 2170
rect 49370 2050 49490 2170
rect 49535 2050 49655 2170
rect 49700 2050 49820 2170
rect 49875 2050 49995 2170
rect 50040 2050 50160 2170
rect 50205 2050 50325 2170
rect 50370 2050 50490 2170
rect 50545 2050 50665 2170
rect 50710 2050 50830 2170
rect 50875 2050 50995 2170
rect 51040 2050 51160 2170
rect 51215 2050 51335 2170
rect 51380 2050 51500 2170
rect 51545 2050 51665 2170
rect 51710 2050 51830 2170
rect 51885 2050 52005 2170
rect 52050 2050 52170 2170
rect 52215 2050 52335 2170
rect 52380 2050 52500 2170
rect 52555 2050 52675 2170
rect 52720 2050 52840 2170
rect 52885 2050 53005 2170
rect 53050 2050 53170 2170
rect 53225 2050 53345 2170
rect 47865 1885 47985 2005
rect 48030 1885 48150 2005
rect 48195 1885 48315 2005
rect 48360 1885 48480 2005
rect 48535 1885 48655 2005
rect 48700 1885 48820 2005
rect 48865 1885 48985 2005
rect 49030 1885 49150 2005
rect 49205 1885 49325 2005
rect 49370 1885 49490 2005
rect 49535 1885 49655 2005
rect 49700 1885 49820 2005
rect 49875 1885 49995 2005
rect 50040 1885 50160 2005
rect 50205 1885 50325 2005
rect 50370 1885 50490 2005
rect 50545 1885 50665 2005
rect 50710 1885 50830 2005
rect 50875 1885 50995 2005
rect 51040 1885 51160 2005
rect 51215 1885 51335 2005
rect 51380 1885 51500 2005
rect 51545 1885 51665 2005
rect 51710 1885 51830 2005
rect 51885 1885 52005 2005
rect 52050 1885 52170 2005
rect 52215 1885 52335 2005
rect 52380 1885 52500 2005
rect 52555 1885 52675 2005
rect 52720 1885 52840 2005
rect 52885 1885 53005 2005
rect 53050 1885 53170 2005
rect 53225 1885 53345 2005
rect 47865 1720 47985 1840
rect 48030 1720 48150 1840
rect 48195 1720 48315 1840
rect 48360 1720 48480 1840
rect 48535 1720 48655 1840
rect 48700 1720 48820 1840
rect 48865 1720 48985 1840
rect 49030 1720 49150 1840
rect 49205 1720 49325 1840
rect 49370 1720 49490 1840
rect 49535 1720 49655 1840
rect 49700 1720 49820 1840
rect 49875 1720 49995 1840
rect 50040 1720 50160 1840
rect 50205 1720 50325 1840
rect 50370 1720 50490 1840
rect 50545 1720 50665 1840
rect 50710 1720 50830 1840
rect 50875 1720 50995 1840
rect 51040 1720 51160 1840
rect 51215 1720 51335 1840
rect 51380 1720 51500 1840
rect 51545 1720 51665 1840
rect 51710 1720 51830 1840
rect 51885 1720 52005 1840
rect 52050 1720 52170 1840
rect 52215 1720 52335 1840
rect 52380 1720 52500 1840
rect 52555 1720 52675 1840
rect 52720 1720 52840 1840
rect 52885 1720 53005 1840
rect 53050 1720 53170 1840
rect 53225 1720 53345 1840
rect 30795 1300 30915 1420
rect 30970 1300 31090 1420
rect 31135 1300 31255 1420
rect 31300 1300 31420 1420
rect 31465 1300 31585 1420
rect 31640 1300 31760 1420
rect 31805 1300 31925 1420
rect 31970 1300 32090 1420
rect 32135 1300 32255 1420
rect 32310 1300 32430 1420
rect 32475 1300 32595 1420
rect 32640 1300 32760 1420
rect 32805 1300 32925 1420
rect 32980 1300 33100 1420
rect 33145 1300 33265 1420
rect 33310 1300 33430 1420
rect 33475 1300 33595 1420
rect 33650 1300 33770 1420
rect 33815 1300 33935 1420
rect 33980 1300 34100 1420
rect 34145 1300 34265 1420
rect 34320 1300 34440 1420
rect 34485 1300 34605 1420
rect 34650 1300 34770 1420
rect 34815 1300 34935 1420
rect 34990 1300 35110 1420
rect 35155 1300 35275 1420
rect 35320 1300 35440 1420
rect 35485 1300 35605 1420
rect 35660 1300 35780 1420
rect 35825 1300 35945 1420
rect 35990 1300 36110 1420
rect 36155 1300 36275 1420
rect 30795 1135 30915 1255
rect 30970 1135 31090 1255
rect 31135 1135 31255 1255
rect 31300 1135 31420 1255
rect 31465 1135 31585 1255
rect 31640 1135 31760 1255
rect 31805 1135 31925 1255
rect 31970 1135 32090 1255
rect 32135 1135 32255 1255
rect 32310 1135 32430 1255
rect 32475 1135 32595 1255
rect 32640 1135 32760 1255
rect 32805 1135 32925 1255
rect 32980 1135 33100 1255
rect 33145 1135 33265 1255
rect 33310 1135 33430 1255
rect 33475 1135 33595 1255
rect 33650 1135 33770 1255
rect 33815 1135 33935 1255
rect 33980 1135 34100 1255
rect 34145 1135 34265 1255
rect 34320 1135 34440 1255
rect 34485 1135 34605 1255
rect 34650 1135 34770 1255
rect 34815 1135 34935 1255
rect 34990 1135 35110 1255
rect 35155 1135 35275 1255
rect 35320 1135 35440 1255
rect 35485 1135 35605 1255
rect 35660 1135 35780 1255
rect 35825 1135 35945 1255
rect 35990 1135 36110 1255
rect 36155 1135 36275 1255
rect 30795 970 30915 1090
rect 30970 970 31090 1090
rect 31135 970 31255 1090
rect 31300 970 31420 1090
rect 31465 970 31585 1090
rect 31640 970 31760 1090
rect 31805 970 31925 1090
rect 31970 970 32090 1090
rect 32135 970 32255 1090
rect 32310 970 32430 1090
rect 32475 970 32595 1090
rect 32640 970 32760 1090
rect 32805 970 32925 1090
rect 32980 970 33100 1090
rect 33145 970 33265 1090
rect 33310 970 33430 1090
rect 33475 970 33595 1090
rect 33650 970 33770 1090
rect 33815 970 33935 1090
rect 33980 970 34100 1090
rect 34145 970 34265 1090
rect 34320 970 34440 1090
rect 34485 970 34605 1090
rect 34650 970 34770 1090
rect 34815 970 34935 1090
rect 34990 970 35110 1090
rect 35155 970 35275 1090
rect 35320 970 35440 1090
rect 35485 970 35605 1090
rect 35660 970 35780 1090
rect 35825 970 35945 1090
rect 35990 970 36110 1090
rect 36155 970 36275 1090
rect 30795 805 30915 925
rect 30970 805 31090 925
rect 31135 805 31255 925
rect 31300 805 31420 925
rect 31465 805 31585 925
rect 31640 805 31760 925
rect 31805 805 31925 925
rect 31970 805 32090 925
rect 32135 805 32255 925
rect 32310 805 32430 925
rect 32475 805 32595 925
rect 32640 805 32760 925
rect 32805 805 32925 925
rect 32980 805 33100 925
rect 33145 805 33265 925
rect 33310 805 33430 925
rect 33475 805 33595 925
rect 33650 805 33770 925
rect 33815 805 33935 925
rect 33980 805 34100 925
rect 34145 805 34265 925
rect 34320 805 34440 925
rect 34485 805 34605 925
rect 34650 805 34770 925
rect 34815 805 34935 925
rect 34990 805 35110 925
rect 35155 805 35275 925
rect 35320 805 35440 925
rect 35485 805 35605 925
rect 35660 805 35780 925
rect 35825 805 35945 925
rect 35990 805 36110 925
rect 36155 805 36275 925
rect 30795 630 30915 750
rect 30970 630 31090 750
rect 31135 630 31255 750
rect 31300 630 31420 750
rect 31465 630 31585 750
rect 31640 630 31760 750
rect 31805 630 31925 750
rect 31970 630 32090 750
rect 32135 630 32255 750
rect 32310 630 32430 750
rect 32475 630 32595 750
rect 32640 630 32760 750
rect 32805 630 32925 750
rect 32980 630 33100 750
rect 33145 630 33265 750
rect 33310 630 33430 750
rect 33475 630 33595 750
rect 33650 630 33770 750
rect 33815 630 33935 750
rect 33980 630 34100 750
rect 34145 630 34265 750
rect 34320 630 34440 750
rect 34485 630 34605 750
rect 34650 630 34770 750
rect 34815 630 34935 750
rect 34990 630 35110 750
rect 35155 630 35275 750
rect 35320 630 35440 750
rect 35485 630 35605 750
rect 35660 630 35780 750
rect 35825 630 35945 750
rect 35990 630 36110 750
rect 36155 630 36275 750
rect 30795 465 30915 585
rect 30970 465 31090 585
rect 31135 465 31255 585
rect 31300 465 31420 585
rect 31465 465 31585 585
rect 31640 465 31760 585
rect 31805 465 31925 585
rect 31970 465 32090 585
rect 32135 465 32255 585
rect 32310 465 32430 585
rect 32475 465 32595 585
rect 32640 465 32760 585
rect 32805 465 32925 585
rect 32980 465 33100 585
rect 33145 465 33265 585
rect 33310 465 33430 585
rect 33475 465 33595 585
rect 33650 465 33770 585
rect 33815 465 33935 585
rect 33980 465 34100 585
rect 34145 465 34265 585
rect 34320 465 34440 585
rect 34485 465 34605 585
rect 34650 465 34770 585
rect 34815 465 34935 585
rect 34990 465 35110 585
rect 35155 465 35275 585
rect 35320 465 35440 585
rect 35485 465 35605 585
rect 35660 465 35780 585
rect 35825 465 35945 585
rect 35990 465 36110 585
rect 36155 465 36275 585
rect 30795 300 30915 420
rect 30970 300 31090 420
rect 31135 300 31255 420
rect 31300 300 31420 420
rect 31465 300 31585 420
rect 31640 300 31760 420
rect 31805 300 31925 420
rect 31970 300 32090 420
rect 32135 300 32255 420
rect 32310 300 32430 420
rect 32475 300 32595 420
rect 32640 300 32760 420
rect 32805 300 32925 420
rect 32980 300 33100 420
rect 33145 300 33265 420
rect 33310 300 33430 420
rect 33475 300 33595 420
rect 33650 300 33770 420
rect 33815 300 33935 420
rect 33980 300 34100 420
rect 34145 300 34265 420
rect 34320 300 34440 420
rect 34485 300 34605 420
rect 34650 300 34770 420
rect 34815 300 34935 420
rect 34990 300 35110 420
rect 35155 300 35275 420
rect 35320 300 35440 420
rect 35485 300 35605 420
rect 35660 300 35780 420
rect 35825 300 35945 420
rect 35990 300 36110 420
rect 36155 300 36275 420
rect 30795 135 30915 255
rect 30970 135 31090 255
rect 31135 135 31255 255
rect 31300 135 31420 255
rect 31465 135 31585 255
rect 31640 135 31760 255
rect 31805 135 31925 255
rect 31970 135 32090 255
rect 32135 135 32255 255
rect 32310 135 32430 255
rect 32475 135 32595 255
rect 32640 135 32760 255
rect 32805 135 32925 255
rect 32980 135 33100 255
rect 33145 135 33265 255
rect 33310 135 33430 255
rect 33475 135 33595 255
rect 33650 135 33770 255
rect 33815 135 33935 255
rect 33980 135 34100 255
rect 34145 135 34265 255
rect 34320 135 34440 255
rect 34485 135 34605 255
rect 34650 135 34770 255
rect 34815 135 34935 255
rect 34990 135 35110 255
rect 35155 135 35275 255
rect 35320 135 35440 255
rect 35485 135 35605 255
rect 35660 135 35780 255
rect 35825 135 35945 255
rect 35990 135 36110 255
rect 36155 135 36275 255
rect 30795 -40 30915 80
rect 30970 -40 31090 80
rect 31135 -40 31255 80
rect 31300 -40 31420 80
rect 31465 -40 31585 80
rect 31640 -40 31760 80
rect 31805 -40 31925 80
rect 31970 -40 32090 80
rect 32135 -40 32255 80
rect 32310 -40 32430 80
rect 32475 -40 32595 80
rect 32640 -40 32760 80
rect 32805 -40 32925 80
rect 32980 -40 33100 80
rect 33145 -40 33265 80
rect 33310 -40 33430 80
rect 33475 -40 33595 80
rect 33650 -40 33770 80
rect 33815 -40 33935 80
rect 33980 -40 34100 80
rect 34145 -40 34265 80
rect 34320 -40 34440 80
rect 34485 -40 34605 80
rect 34650 -40 34770 80
rect 34815 -40 34935 80
rect 34990 -40 35110 80
rect 35155 -40 35275 80
rect 35320 -40 35440 80
rect 35485 -40 35605 80
rect 35660 -40 35780 80
rect 35825 -40 35945 80
rect 35990 -40 36110 80
rect 36155 -40 36275 80
rect 30795 -205 30915 -85
rect 30970 -205 31090 -85
rect 31135 -205 31255 -85
rect 31300 -205 31420 -85
rect 31465 -205 31585 -85
rect 31640 -205 31760 -85
rect 31805 -205 31925 -85
rect 31970 -205 32090 -85
rect 32135 -205 32255 -85
rect 32310 -205 32430 -85
rect 32475 -205 32595 -85
rect 32640 -205 32760 -85
rect 32805 -205 32925 -85
rect 32980 -205 33100 -85
rect 33145 -205 33265 -85
rect 33310 -205 33430 -85
rect 33475 -205 33595 -85
rect 33650 -205 33770 -85
rect 33815 -205 33935 -85
rect 33980 -205 34100 -85
rect 34145 -205 34265 -85
rect 34320 -205 34440 -85
rect 34485 -205 34605 -85
rect 34650 -205 34770 -85
rect 34815 -205 34935 -85
rect 34990 -205 35110 -85
rect 35155 -205 35275 -85
rect 35320 -205 35440 -85
rect 35485 -205 35605 -85
rect 35660 -205 35780 -85
rect 35825 -205 35945 -85
rect 35990 -205 36110 -85
rect 36155 -205 36275 -85
rect 30795 -370 30915 -250
rect 30970 -370 31090 -250
rect 31135 -370 31255 -250
rect 31300 -370 31420 -250
rect 31465 -370 31585 -250
rect 31640 -370 31760 -250
rect 31805 -370 31925 -250
rect 31970 -370 32090 -250
rect 32135 -370 32255 -250
rect 32310 -370 32430 -250
rect 32475 -370 32595 -250
rect 32640 -370 32760 -250
rect 32805 -370 32925 -250
rect 32980 -370 33100 -250
rect 33145 -370 33265 -250
rect 33310 -370 33430 -250
rect 33475 -370 33595 -250
rect 33650 -370 33770 -250
rect 33815 -370 33935 -250
rect 33980 -370 34100 -250
rect 34145 -370 34265 -250
rect 34320 -370 34440 -250
rect 34485 -370 34605 -250
rect 34650 -370 34770 -250
rect 34815 -370 34935 -250
rect 34990 -370 35110 -250
rect 35155 -370 35275 -250
rect 35320 -370 35440 -250
rect 35485 -370 35605 -250
rect 35660 -370 35780 -250
rect 35825 -370 35945 -250
rect 35990 -370 36110 -250
rect 36155 -370 36275 -250
rect 30795 -535 30915 -415
rect 30970 -535 31090 -415
rect 31135 -535 31255 -415
rect 31300 -535 31420 -415
rect 31465 -535 31585 -415
rect 31640 -535 31760 -415
rect 31805 -535 31925 -415
rect 31970 -535 32090 -415
rect 32135 -535 32255 -415
rect 32310 -535 32430 -415
rect 32475 -535 32595 -415
rect 32640 -535 32760 -415
rect 32805 -535 32925 -415
rect 32980 -535 33100 -415
rect 33145 -535 33265 -415
rect 33310 -535 33430 -415
rect 33475 -535 33595 -415
rect 33650 -535 33770 -415
rect 33815 -535 33935 -415
rect 33980 -535 34100 -415
rect 34145 -535 34265 -415
rect 34320 -535 34440 -415
rect 34485 -535 34605 -415
rect 34650 -535 34770 -415
rect 34815 -535 34935 -415
rect 34990 -535 35110 -415
rect 35155 -535 35275 -415
rect 35320 -535 35440 -415
rect 35485 -535 35605 -415
rect 35660 -535 35780 -415
rect 35825 -535 35945 -415
rect 35990 -535 36110 -415
rect 36155 -535 36275 -415
rect 30795 -710 30915 -590
rect 30970 -710 31090 -590
rect 31135 -710 31255 -590
rect 31300 -710 31420 -590
rect 31465 -710 31585 -590
rect 31640 -710 31760 -590
rect 31805 -710 31925 -590
rect 31970 -710 32090 -590
rect 32135 -710 32255 -590
rect 32310 -710 32430 -590
rect 32475 -710 32595 -590
rect 32640 -710 32760 -590
rect 32805 -710 32925 -590
rect 32980 -710 33100 -590
rect 33145 -710 33265 -590
rect 33310 -710 33430 -590
rect 33475 -710 33595 -590
rect 33650 -710 33770 -590
rect 33815 -710 33935 -590
rect 33980 -710 34100 -590
rect 34145 -710 34265 -590
rect 34320 -710 34440 -590
rect 34485 -710 34605 -590
rect 34650 -710 34770 -590
rect 34815 -710 34935 -590
rect 34990 -710 35110 -590
rect 35155 -710 35275 -590
rect 35320 -710 35440 -590
rect 35485 -710 35605 -590
rect 35660 -710 35780 -590
rect 35825 -710 35945 -590
rect 35990 -710 36110 -590
rect 36155 -710 36275 -590
rect 30795 -875 30915 -755
rect 30970 -875 31090 -755
rect 31135 -875 31255 -755
rect 31300 -875 31420 -755
rect 31465 -875 31585 -755
rect 31640 -875 31760 -755
rect 31805 -875 31925 -755
rect 31970 -875 32090 -755
rect 32135 -875 32255 -755
rect 32310 -875 32430 -755
rect 32475 -875 32595 -755
rect 32640 -875 32760 -755
rect 32805 -875 32925 -755
rect 32980 -875 33100 -755
rect 33145 -875 33265 -755
rect 33310 -875 33430 -755
rect 33475 -875 33595 -755
rect 33650 -875 33770 -755
rect 33815 -875 33935 -755
rect 33980 -875 34100 -755
rect 34145 -875 34265 -755
rect 34320 -875 34440 -755
rect 34485 -875 34605 -755
rect 34650 -875 34770 -755
rect 34815 -875 34935 -755
rect 34990 -875 35110 -755
rect 35155 -875 35275 -755
rect 35320 -875 35440 -755
rect 35485 -875 35605 -755
rect 35660 -875 35780 -755
rect 35825 -875 35945 -755
rect 35990 -875 36110 -755
rect 36155 -875 36275 -755
rect 30795 -1040 30915 -920
rect 30970 -1040 31090 -920
rect 31135 -1040 31255 -920
rect 31300 -1040 31420 -920
rect 31465 -1040 31585 -920
rect 31640 -1040 31760 -920
rect 31805 -1040 31925 -920
rect 31970 -1040 32090 -920
rect 32135 -1040 32255 -920
rect 32310 -1040 32430 -920
rect 32475 -1040 32595 -920
rect 32640 -1040 32760 -920
rect 32805 -1040 32925 -920
rect 32980 -1040 33100 -920
rect 33145 -1040 33265 -920
rect 33310 -1040 33430 -920
rect 33475 -1040 33595 -920
rect 33650 -1040 33770 -920
rect 33815 -1040 33935 -920
rect 33980 -1040 34100 -920
rect 34145 -1040 34265 -920
rect 34320 -1040 34440 -920
rect 34485 -1040 34605 -920
rect 34650 -1040 34770 -920
rect 34815 -1040 34935 -920
rect 34990 -1040 35110 -920
rect 35155 -1040 35275 -920
rect 35320 -1040 35440 -920
rect 35485 -1040 35605 -920
rect 35660 -1040 35780 -920
rect 35825 -1040 35945 -920
rect 35990 -1040 36110 -920
rect 36155 -1040 36275 -920
rect 30795 -1205 30915 -1085
rect 30970 -1205 31090 -1085
rect 31135 -1205 31255 -1085
rect 31300 -1205 31420 -1085
rect 31465 -1205 31585 -1085
rect 31640 -1205 31760 -1085
rect 31805 -1205 31925 -1085
rect 31970 -1205 32090 -1085
rect 32135 -1205 32255 -1085
rect 32310 -1205 32430 -1085
rect 32475 -1205 32595 -1085
rect 32640 -1205 32760 -1085
rect 32805 -1205 32925 -1085
rect 32980 -1205 33100 -1085
rect 33145 -1205 33265 -1085
rect 33310 -1205 33430 -1085
rect 33475 -1205 33595 -1085
rect 33650 -1205 33770 -1085
rect 33815 -1205 33935 -1085
rect 33980 -1205 34100 -1085
rect 34145 -1205 34265 -1085
rect 34320 -1205 34440 -1085
rect 34485 -1205 34605 -1085
rect 34650 -1205 34770 -1085
rect 34815 -1205 34935 -1085
rect 34990 -1205 35110 -1085
rect 35155 -1205 35275 -1085
rect 35320 -1205 35440 -1085
rect 35485 -1205 35605 -1085
rect 35660 -1205 35780 -1085
rect 35825 -1205 35945 -1085
rect 35990 -1205 36110 -1085
rect 36155 -1205 36275 -1085
rect 30795 -1380 30915 -1260
rect 30970 -1380 31090 -1260
rect 31135 -1380 31255 -1260
rect 31300 -1380 31420 -1260
rect 31465 -1380 31585 -1260
rect 31640 -1380 31760 -1260
rect 31805 -1380 31925 -1260
rect 31970 -1380 32090 -1260
rect 32135 -1380 32255 -1260
rect 32310 -1380 32430 -1260
rect 32475 -1380 32595 -1260
rect 32640 -1380 32760 -1260
rect 32805 -1380 32925 -1260
rect 32980 -1380 33100 -1260
rect 33145 -1380 33265 -1260
rect 33310 -1380 33430 -1260
rect 33475 -1380 33595 -1260
rect 33650 -1380 33770 -1260
rect 33815 -1380 33935 -1260
rect 33980 -1380 34100 -1260
rect 34145 -1380 34265 -1260
rect 34320 -1380 34440 -1260
rect 34485 -1380 34605 -1260
rect 34650 -1380 34770 -1260
rect 34815 -1380 34935 -1260
rect 34990 -1380 35110 -1260
rect 35155 -1380 35275 -1260
rect 35320 -1380 35440 -1260
rect 35485 -1380 35605 -1260
rect 35660 -1380 35780 -1260
rect 35825 -1380 35945 -1260
rect 35990 -1380 36110 -1260
rect 36155 -1380 36275 -1260
rect 30795 -1545 30915 -1425
rect 30970 -1545 31090 -1425
rect 31135 -1545 31255 -1425
rect 31300 -1545 31420 -1425
rect 31465 -1545 31585 -1425
rect 31640 -1545 31760 -1425
rect 31805 -1545 31925 -1425
rect 31970 -1545 32090 -1425
rect 32135 -1545 32255 -1425
rect 32310 -1545 32430 -1425
rect 32475 -1545 32595 -1425
rect 32640 -1545 32760 -1425
rect 32805 -1545 32925 -1425
rect 32980 -1545 33100 -1425
rect 33145 -1545 33265 -1425
rect 33310 -1545 33430 -1425
rect 33475 -1545 33595 -1425
rect 33650 -1545 33770 -1425
rect 33815 -1545 33935 -1425
rect 33980 -1545 34100 -1425
rect 34145 -1545 34265 -1425
rect 34320 -1545 34440 -1425
rect 34485 -1545 34605 -1425
rect 34650 -1545 34770 -1425
rect 34815 -1545 34935 -1425
rect 34990 -1545 35110 -1425
rect 35155 -1545 35275 -1425
rect 35320 -1545 35440 -1425
rect 35485 -1545 35605 -1425
rect 35660 -1545 35780 -1425
rect 35825 -1545 35945 -1425
rect 35990 -1545 36110 -1425
rect 36155 -1545 36275 -1425
rect 30795 -1710 30915 -1590
rect 30970 -1710 31090 -1590
rect 31135 -1710 31255 -1590
rect 31300 -1710 31420 -1590
rect 31465 -1710 31585 -1590
rect 31640 -1710 31760 -1590
rect 31805 -1710 31925 -1590
rect 31970 -1710 32090 -1590
rect 32135 -1710 32255 -1590
rect 32310 -1710 32430 -1590
rect 32475 -1710 32595 -1590
rect 32640 -1710 32760 -1590
rect 32805 -1710 32925 -1590
rect 32980 -1710 33100 -1590
rect 33145 -1710 33265 -1590
rect 33310 -1710 33430 -1590
rect 33475 -1710 33595 -1590
rect 33650 -1710 33770 -1590
rect 33815 -1710 33935 -1590
rect 33980 -1710 34100 -1590
rect 34145 -1710 34265 -1590
rect 34320 -1710 34440 -1590
rect 34485 -1710 34605 -1590
rect 34650 -1710 34770 -1590
rect 34815 -1710 34935 -1590
rect 34990 -1710 35110 -1590
rect 35155 -1710 35275 -1590
rect 35320 -1710 35440 -1590
rect 35485 -1710 35605 -1590
rect 35660 -1710 35780 -1590
rect 35825 -1710 35945 -1590
rect 35990 -1710 36110 -1590
rect 36155 -1710 36275 -1590
rect 30795 -1875 30915 -1755
rect 30970 -1875 31090 -1755
rect 31135 -1875 31255 -1755
rect 31300 -1875 31420 -1755
rect 31465 -1875 31585 -1755
rect 31640 -1875 31760 -1755
rect 31805 -1875 31925 -1755
rect 31970 -1875 32090 -1755
rect 32135 -1875 32255 -1755
rect 32310 -1875 32430 -1755
rect 32475 -1875 32595 -1755
rect 32640 -1875 32760 -1755
rect 32805 -1875 32925 -1755
rect 32980 -1875 33100 -1755
rect 33145 -1875 33265 -1755
rect 33310 -1875 33430 -1755
rect 33475 -1875 33595 -1755
rect 33650 -1875 33770 -1755
rect 33815 -1875 33935 -1755
rect 33980 -1875 34100 -1755
rect 34145 -1875 34265 -1755
rect 34320 -1875 34440 -1755
rect 34485 -1875 34605 -1755
rect 34650 -1875 34770 -1755
rect 34815 -1875 34935 -1755
rect 34990 -1875 35110 -1755
rect 35155 -1875 35275 -1755
rect 35320 -1875 35440 -1755
rect 35485 -1875 35605 -1755
rect 35660 -1875 35780 -1755
rect 35825 -1875 35945 -1755
rect 35990 -1875 36110 -1755
rect 36155 -1875 36275 -1755
rect 30795 -2050 30915 -1930
rect 30970 -2050 31090 -1930
rect 31135 -2050 31255 -1930
rect 31300 -2050 31420 -1930
rect 31465 -2050 31585 -1930
rect 31640 -2050 31760 -1930
rect 31805 -2050 31925 -1930
rect 31970 -2050 32090 -1930
rect 32135 -2050 32255 -1930
rect 32310 -2050 32430 -1930
rect 32475 -2050 32595 -1930
rect 32640 -2050 32760 -1930
rect 32805 -2050 32925 -1930
rect 32980 -2050 33100 -1930
rect 33145 -2050 33265 -1930
rect 33310 -2050 33430 -1930
rect 33475 -2050 33595 -1930
rect 33650 -2050 33770 -1930
rect 33815 -2050 33935 -1930
rect 33980 -2050 34100 -1930
rect 34145 -2050 34265 -1930
rect 34320 -2050 34440 -1930
rect 34485 -2050 34605 -1930
rect 34650 -2050 34770 -1930
rect 34815 -2050 34935 -1930
rect 34990 -2050 35110 -1930
rect 35155 -2050 35275 -1930
rect 35320 -2050 35440 -1930
rect 35485 -2050 35605 -1930
rect 35660 -2050 35780 -1930
rect 35825 -2050 35945 -1930
rect 35990 -2050 36110 -1930
rect 36155 -2050 36275 -1930
rect 30795 -2215 30915 -2095
rect 30970 -2215 31090 -2095
rect 31135 -2215 31255 -2095
rect 31300 -2215 31420 -2095
rect 31465 -2215 31585 -2095
rect 31640 -2215 31760 -2095
rect 31805 -2215 31925 -2095
rect 31970 -2215 32090 -2095
rect 32135 -2215 32255 -2095
rect 32310 -2215 32430 -2095
rect 32475 -2215 32595 -2095
rect 32640 -2215 32760 -2095
rect 32805 -2215 32925 -2095
rect 32980 -2215 33100 -2095
rect 33145 -2215 33265 -2095
rect 33310 -2215 33430 -2095
rect 33475 -2215 33595 -2095
rect 33650 -2215 33770 -2095
rect 33815 -2215 33935 -2095
rect 33980 -2215 34100 -2095
rect 34145 -2215 34265 -2095
rect 34320 -2215 34440 -2095
rect 34485 -2215 34605 -2095
rect 34650 -2215 34770 -2095
rect 34815 -2215 34935 -2095
rect 34990 -2215 35110 -2095
rect 35155 -2215 35275 -2095
rect 35320 -2215 35440 -2095
rect 35485 -2215 35605 -2095
rect 35660 -2215 35780 -2095
rect 35825 -2215 35945 -2095
rect 35990 -2215 36110 -2095
rect 36155 -2215 36275 -2095
rect 30795 -2380 30915 -2260
rect 30970 -2380 31090 -2260
rect 31135 -2380 31255 -2260
rect 31300 -2380 31420 -2260
rect 31465 -2380 31585 -2260
rect 31640 -2380 31760 -2260
rect 31805 -2380 31925 -2260
rect 31970 -2380 32090 -2260
rect 32135 -2380 32255 -2260
rect 32310 -2380 32430 -2260
rect 32475 -2380 32595 -2260
rect 32640 -2380 32760 -2260
rect 32805 -2380 32925 -2260
rect 32980 -2380 33100 -2260
rect 33145 -2380 33265 -2260
rect 33310 -2380 33430 -2260
rect 33475 -2380 33595 -2260
rect 33650 -2380 33770 -2260
rect 33815 -2380 33935 -2260
rect 33980 -2380 34100 -2260
rect 34145 -2380 34265 -2260
rect 34320 -2380 34440 -2260
rect 34485 -2380 34605 -2260
rect 34650 -2380 34770 -2260
rect 34815 -2380 34935 -2260
rect 34990 -2380 35110 -2260
rect 35155 -2380 35275 -2260
rect 35320 -2380 35440 -2260
rect 35485 -2380 35605 -2260
rect 35660 -2380 35780 -2260
rect 35825 -2380 35945 -2260
rect 35990 -2380 36110 -2260
rect 36155 -2380 36275 -2260
rect 30795 -2545 30915 -2425
rect 30970 -2545 31090 -2425
rect 31135 -2545 31255 -2425
rect 31300 -2545 31420 -2425
rect 31465 -2545 31585 -2425
rect 31640 -2545 31760 -2425
rect 31805 -2545 31925 -2425
rect 31970 -2545 32090 -2425
rect 32135 -2545 32255 -2425
rect 32310 -2545 32430 -2425
rect 32475 -2545 32595 -2425
rect 32640 -2545 32760 -2425
rect 32805 -2545 32925 -2425
rect 32980 -2545 33100 -2425
rect 33145 -2545 33265 -2425
rect 33310 -2545 33430 -2425
rect 33475 -2545 33595 -2425
rect 33650 -2545 33770 -2425
rect 33815 -2545 33935 -2425
rect 33980 -2545 34100 -2425
rect 34145 -2545 34265 -2425
rect 34320 -2545 34440 -2425
rect 34485 -2545 34605 -2425
rect 34650 -2545 34770 -2425
rect 34815 -2545 34935 -2425
rect 34990 -2545 35110 -2425
rect 35155 -2545 35275 -2425
rect 35320 -2545 35440 -2425
rect 35485 -2545 35605 -2425
rect 35660 -2545 35780 -2425
rect 35825 -2545 35945 -2425
rect 35990 -2545 36110 -2425
rect 36155 -2545 36275 -2425
rect 30795 -2720 30915 -2600
rect 30970 -2720 31090 -2600
rect 31135 -2720 31255 -2600
rect 31300 -2720 31420 -2600
rect 31465 -2720 31585 -2600
rect 31640 -2720 31760 -2600
rect 31805 -2720 31925 -2600
rect 31970 -2720 32090 -2600
rect 32135 -2720 32255 -2600
rect 32310 -2720 32430 -2600
rect 32475 -2720 32595 -2600
rect 32640 -2720 32760 -2600
rect 32805 -2720 32925 -2600
rect 32980 -2720 33100 -2600
rect 33145 -2720 33265 -2600
rect 33310 -2720 33430 -2600
rect 33475 -2720 33595 -2600
rect 33650 -2720 33770 -2600
rect 33815 -2720 33935 -2600
rect 33980 -2720 34100 -2600
rect 34145 -2720 34265 -2600
rect 34320 -2720 34440 -2600
rect 34485 -2720 34605 -2600
rect 34650 -2720 34770 -2600
rect 34815 -2720 34935 -2600
rect 34990 -2720 35110 -2600
rect 35155 -2720 35275 -2600
rect 35320 -2720 35440 -2600
rect 35485 -2720 35605 -2600
rect 35660 -2720 35780 -2600
rect 35825 -2720 35945 -2600
rect 35990 -2720 36110 -2600
rect 36155 -2720 36275 -2600
rect 30795 -2885 30915 -2765
rect 30970 -2885 31090 -2765
rect 31135 -2885 31255 -2765
rect 31300 -2885 31420 -2765
rect 31465 -2885 31585 -2765
rect 31640 -2885 31760 -2765
rect 31805 -2885 31925 -2765
rect 31970 -2885 32090 -2765
rect 32135 -2885 32255 -2765
rect 32310 -2885 32430 -2765
rect 32475 -2885 32595 -2765
rect 32640 -2885 32760 -2765
rect 32805 -2885 32925 -2765
rect 32980 -2885 33100 -2765
rect 33145 -2885 33265 -2765
rect 33310 -2885 33430 -2765
rect 33475 -2885 33595 -2765
rect 33650 -2885 33770 -2765
rect 33815 -2885 33935 -2765
rect 33980 -2885 34100 -2765
rect 34145 -2885 34265 -2765
rect 34320 -2885 34440 -2765
rect 34485 -2885 34605 -2765
rect 34650 -2885 34770 -2765
rect 34815 -2885 34935 -2765
rect 34990 -2885 35110 -2765
rect 35155 -2885 35275 -2765
rect 35320 -2885 35440 -2765
rect 35485 -2885 35605 -2765
rect 35660 -2885 35780 -2765
rect 35825 -2885 35945 -2765
rect 35990 -2885 36110 -2765
rect 36155 -2885 36275 -2765
rect 30795 -3050 30915 -2930
rect 30970 -3050 31090 -2930
rect 31135 -3050 31255 -2930
rect 31300 -3050 31420 -2930
rect 31465 -3050 31585 -2930
rect 31640 -3050 31760 -2930
rect 31805 -3050 31925 -2930
rect 31970 -3050 32090 -2930
rect 32135 -3050 32255 -2930
rect 32310 -3050 32430 -2930
rect 32475 -3050 32595 -2930
rect 32640 -3050 32760 -2930
rect 32805 -3050 32925 -2930
rect 32980 -3050 33100 -2930
rect 33145 -3050 33265 -2930
rect 33310 -3050 33430 -2930
rect 33475 -3050 33595 -2930
rect 33650 -3050 33770 -2930
rect 33815 -3050 33935 -2930
rect 33980 -3050 34100 -2930
rect 34145 -3050 34265 -2930
rect 34320 -3050 34440 -2930
rect 34485 -3050 34605 -2930
rect 34650 -3050 34770 -2930
rect 34815 -3050 34935 -2930
rect 34990 -3050 35110 -2930
rect 35155 -3050 35275 -2930
rect 35320 -3050 35440 -2930
rect 35485 -3050 35605 -2930
rect 35660 -3050 35780 -2930
rect 35825 -3050 35945 -2930
rect 35990 -3050 36110 -2930
rect 36155 -3050 36275 -2930
rect 30795 -3215 30915 -3095
rect 30970 -3215 31090 -3095
rect 31135 -3215 31255 -3095
rect 31300 -3215 31420 -3095
rect 31465 -3215 31585 -3095
rect 31640 -3215 31760 -3095
rect 31805 -3215 31925 -3095
rect 31970 -3215 32090 -3095
rect 32135 -3215 32255 -3095
rect 32310 -3215 32430 -3095
rect 32475 -3215 32595 -3095
rect 32640 -3215 32760 -3095
rect 32805 -3215 32925 -3095
rect 32980 -3215 33100 -3095
rect 33145 -3215 33265 -3095
rect 33310 -3215 33430 -3095
rect 33475 -3215 33595 -3095
rect 33650 -3215 33770 -3095
rect 33815 -3215 33935 -3095
rect 33980 -3215 34100 -3095
rect 34145 -3215 34265 -3095
rect 34320 -3215 34440 -3095
rect 34485 -3215 34605 -3095
rect 34650 -3215 34770 -3095
rect 34815 -3215 34935 -3095
rect 34990 -3215 35110 -3095
rect 35155 -3215 35275 -3095
rect 35320 -3215 35440 -3095
rect 35485 -3215 35605 -3095
rect 35660 -3215 35780 -3095
rect 35825 -3215 35945 -3095
rect 35990 -3215 36110 -3095
rect 36155 -3215 36275 -3095
rect 30795 -3390 30915 -3270
rect 30970 -3390 31090 -3270
rect 31135 -3390 31255 -3270
rect 31300 -3390 31420 -3270
rect 31465 -3390 31585 -3270
rect 31640 -3390 31760 -3270
rect 31805 -3390 31925 -3270
rect 31970 -3390 32090 -3270
rect 32135 -3390 32255 -3270
rect 32310 -3390 32430 -3270
rect 32475 -3390 32595 -3270
rect 32640 -3390 32760 -3270
rect 32805 -3390 32925 -3270
rect 32980 -3390 33100 -3270
rect 33145 -3390 33265 -3270
rect 33310 -3390 33430 -3270
rect 33475 -3390 33595 -3270
rect 33650 -3390 33770 -3270
rect 33815 -3390 33935 -3270
rect 33980 -3390 34100 -3270
rect 34145 -3390 34265 -3270
rect 34320 -3390 34440 -3270
rect 34485 -3390 34605 -3270
rect 34650 -3390 34770 -3270
rect 34815 -3390 34935 -3270
rect 34990 -3390 35110 -3270
rect 35155 -3390 35275 -3270
rect 35320 -3390 35440 -3270
rect 35485 -3390 35605 -3270
rect 35660 -3390 35780 -3270
rect 35825 -3390 35945 -3270
rect 35990 -3390 36110 -3270
rect 36155 -3390 36275 -3270
rect 30795 -3555 30915 -3435
rect 30970 -3555 31090 -3435
rect 31135 -3555 31255 -3435
rect 31300 -3555 31420 -3435
rect 31465 -3555 31585 -3435
rect 31640 -3555 31760 -3435
rect 31805 -3555 31925 -3435
rect 31970 -3555 32090 -3435
rect 32135 -3555 32255 -3435
rect 32310 -3555 32430 -3435
rect 32475 -3555 32595 -3435
rect 32640 -3555 32760 -3435
rect 32805 -3555 32925 -3435
rect 32980 -3555 33100 -3435
rect 33145 -3555 33265 -3435
rect 33310 -3555 33430 -3435
rect 33475 -3555 33595 -3435
rect 33650 -3555 33770 -3435
rect 33815 -3555 33935 -3435
rect 33980 -3555 34100 -3435
rect 34145 -3555 34265 -3435
rect 34320 -3555 34440 -3435
rect 34485 -3555 34605 -3435
rect 34650 -3555 34770 -3435
rect 34815 -3555 34935 -3435
rect 34990 -3555 35110 -3435
rect 35155 -3555 35275 -3435
rect 35320 -3555 35440 -3435
rect 35485 -3555 35605 -3435
rect 35660 -3555 35780 -3435
rect 35825 -3555 35945 -3435
rect 35990 -3555 36110 -3435
rect 36155 -3555 36275 -3435
rect 30795 -3720 30915 -3600
rect 30970 -3720 31090 -3600
rect 31135 -3720 31255 -3600
rect 31300 -3720 31420 -3600
rect 31465 -3720 31585 -3600
rect 31640 -3720 31760 -3600
rect 31805 -3720 31925 -3600
rect 31970 -3720 32090 -3600
rect 32135 -3720 32255 -3600
rect 32310 -3720 32430 -3600
rect 32475 -3720 32595 -3600
rect 32640 -3720 32760 -3600
rect 32805 -3720 32925 -3600
rect 32980 -3720 33100 -3600
rect 33145 -3720 33265 -3600
rect 33310 -3720 33430 -3600
rect 33475 -3720 33595 -3600
rect 33650 -3720 33770 -3600
rect 33815 -3720 33935 -3600
rect 33980 -3720 34100 -3600
rect 34145 -3720 34265 -3600
rect 34320 -3720 34440 -3600
rect 34485 -3720 34605 -3600
rect 34650 -3720 34770 -3600
rect 34815 -3720 34935 -3600
rect 34990 -3720 35110 -3600
rect 35155 -3720 35275 -3600
rect 35320 -3720 35440 -3600
rect 35485 -3720 35605 -3600
rect 35660 -3720 35780 -3600
rect 35825 -3720 35945 -3600
rect 35990 -3720 36110 -3600
rect 36155 -3720 36275 -3600
rect 30795 -3885 30915 -3765
rect 30970 -3885 31090 -3765
rect 31135 -3885 31255 -3765
rect 31300 -3885 31420 -3765
rect 31465 -3885 31585 -3765
rect 31640 -3885 31760 -3765
rect 31805 -3885 31925 -3765
rect 31970 -3885 32090 -3765
rect 32135 -3885 32255 -3765
rect 32310 -3885 32430 -3765
rect 32475 -3885 32595 -3765
rect 32640 -3885 32760 -3765
rect 32805 -3885 32925 -3765
rect 32980 -3885 33100 -3765
rect 33145 -3885 33265 -3765
rect 33310 -3885 33430 -3765
rect 33475 -3885 33595 -3765
rect 33650 -3885 33770 -3765
rect 33815 -3885 33935 -3765
rect 33980 -3885 34100 -3765
rect 34145 -3885 34265 -3765
rect 34320 -3885 34440 -3765
rect 34485 -3885 34605 -3765
rect 34650 -3885 34770 -3765
rect 34815 -3885 34935 -3765
rect 34990 -3885 35110 -3765
rect 35155 -3885 35275 -3765
rect 35320 -3885 35440 -3765
rect 35485 -3885 35605 -3765
rect 35660 -3885 35780 -3765
rect 35825 -3885 35945 -3765
rect 35990 -3885 36110 -3765
rect 36155 -3885 36275 -3765
rect 30795 -4060 30915 -3940
rect 30970 -4060 31090 -3940
rect 31135 -4060 31255 -3940
rect 31300 -4060 31420 -3940
rect 31465 -4060 31585 -3940
rect 31640 -4060 31760 -3940
rect 31805 -4060 31925 -3940
rect 31970 -4060 32090 -3940
rect 32135 -4060 32255 -3940
rect 32310 -4060 32430 -3940
rect 32475 -4060 32595 -3940
rect 32640 -4060 32760 -3940
rect 32805 -4060 32925 -3940
rect 32980 -4060 33100 -3940
rect 33145 -4060 33265 -3940
rect 33310 -4060 33430 -3940
rect 33475 -4060 33595 -3940
rect 33650 -4060 33770 -3940
rect 33815 -4060 33935 -3940
rect 33980 -4060 34100 -3940
rect 34145 -4060 34265 -3940
rect 34320 -4060 34440 -3940
rect 34485 -4060 34605 -3940
rect 34650 -4060 34770 -3940
rect 34815 -4060 34935 -3940
rect 34990 -4060 35110 -3940
rect 35155 -4060 35275 -3940
rect 35320 -4060 35440 -3940
rect 35485 -4060 35605 -3940
rect 35660 -4060 35780 -3940
rect 35825 -4060 35945 -3940
rect 35990 -4060 36110 -3940
rect 36155 -4060 36275 -3940
rect 36485 1300 36605 1420
rect 36660 1300 36780 1420
rect 36825 1300 36945 1420
rect 36990 1300 37110 1420
rect 37155 1300 37275 1420
rect 37330 1300 37450 1420
rect 37495 1300 37615 1420
rect 37660 1300 37780 1420
rect 37825 1300 37945 1420
rect 38000 1300 38120 1420
rect 38165 1300 38285 1420
rect 38330 1300 38450 1420
rect 38495 1300 38615 1420
rect 38670 1300 38790 1420
rect 38835 1300 38955 1420
rect 39000 1300 39120 1420
rect 39165 1300 39285 1420
rect 39340 1300 39460 1420
rect 39505 1300 39625 1420
rect 39670 1300 39790 1420
rect 39835 1300 39955 1420
rect 40010 1300 40130 1420
rect 40175 1300 40295 1420
rect 40340 1300 40460 1420
rect 40505 1300 40625 1420
rect 40680 1300 40800 1420
rect 40845 1300 40965 1420
rect 41010 1300 41130 1420
rect 41175 1300 41295 1420
rect 41350 1300 41470 1420
rect 41515 1300 41635 1420
rect 41680 1300 41800 1420
rect 41845 1300 41965 1420
rect 36485 1135 36605 1255
rect 36660 1135 36780 1255
rect 36825 1135 36945 1255
rect 36990 1135 37110 1255
rect 37155 1135 37275 1255
rect 37330 1135 37450 1255
rect 37495 1135 37615 1255
rect 37660 1135 37780 1255
rect 37825 1135 37945 1255
rect 38000 1135 38120 1255
rect 38165 1135 38285 1255
rect 38330 1135 38450 1255
rect 38495 1135 38615 1255
rect 38670 1135 38790 1255
rect 38835 1135 38955 1255
rect 39000 1135 39120 1255
rect 39165 1135 39285 1255
rect 39340 1135 39460 1255
rect 39505 1135 39625 1255
rect 39670 1135 39790 1255
rect 39835 1135 39955 1255
rect 40010 1135 40130 1255
rect 40175 1135 40295 1255
rect 40340 1135 40460 1255
rect 40505 1135 40625 1255
rect 40680 1135 40800 1255
rect 40845 1135 40965 1255
rect 41010 1135 41130 1255
rect 41175 1135 41295 1255
rect 41350 1135 41470 1255
rect 41515 1135 41635 1255
rect 41680 1135 41800 1255
rect 41845 1135 41965 1255
rect 36485 970 36605 1090
rect 36660 970 36780 1090
rect 36825 970 36945 1090
rect 36990 970 37110 1090
rect 37155 970 37275 1090
rect 37330 970 37450 1090
rect 37495 970 37615 1090
rect 37660 970 37780 1090
rect 37825 970 37945 1090
rect 38000 970 38120 1090
rect 38165 970 38285 1090
rect 38330 970 38450 1090
rect 38495 970 38615 1090
rect 38670 970 38790 1090
rect 38835 970 38955 1090
rect 39000 970 39120 1090
rect 39165 970 39285 1090
rect 39340 970 39460 1090
rect 39505 970 39625 1090
rect 39670 970 39790 1090
rect 39835 970 39955 1090
rect 40010 970 40130 1090
rect 40175 970 40295 1090
rect 40340 970 40460 1090
rect 40505 970 40625 1090
rect 40680 970 40800 1090
rect 40845 970 40965 1090
rect 41010 970 41130 1090
rect 41175 970 41295 1090
rect 41350 970 41470 1090
rect 41515 970 41635 1090
rect 41680 970 41800 1090
rect 41845 970 41965 1090
rect 36485 805 36605 925
rect 36660 805 36780 925
rect 36825 805 36945 925
rect 36990 805 37110 925
rect 37155 805 37275 925
rect 37330 805 37450 925
rect 37495 805 37615 925
rect 37660 805 37780 925
rect 37825 805 37945 925
rect 38000 805 38120 925
rect 38165 805 38285 925
rect 38330 805 38450 925
rect 38495 805 38615 925
rect 38670 805 38790 925
rect 38835 805 38955 925
rect 39000 805 39120 925
rect 39165 805 39285 925
rect 39340 805 39460 925
rect 39505 805 39625 925
rect 39670 805 39790 925
rect 39835 805 39955 925
rect 40010 805 40130 925
rect 40175 805 40295 925
rect 40340 805 40460 925
rect 40505 805 40625 925
rect 40680 805 40800 925
rect 40845 805 40965 925
rect 41010 805 41130 925
rect 41175 805 41295 925
rect 41350 805 41470 925
rect 41515 805 41635 925
rect 41680 805 41800 925
rect 41845 805 41965 925
rect 36485 630 36605 750
rect 36660 630 36780 750
rect 36825 630 36945 750
rect 36990 630 37110 750
rect 37155 630 37275 750
rect 37330 630 37450 750
rect 37495 630 37615 750
rect 37660 630 37780 750
rect 37825 630 37945 750
rect 38000 630 38120 750
rect 38165 630 38285 750
rect 38330 630 38450 750
rect 38495 630 38615 750
rect 38670 630 38790 750
rect 38835 630 38955 750
rect 39000 630 39120 750
rect 39165 630 39285 750
rect 39340 630 39460 750
rect 39505 630 39625 750
rect 39670 630 39790 750
rect 39835 630 39955 750
rect 40010 630 40130 750
rect 40175 630 40295 750
rect 40340 630 40460 750
rect 40505 630 40625 750
rect 40680 630 40800 750
rect 40845 630 40965 750
rect 41010 630 41130 750
rect 41175 630 41295 750
rect 41350 630 41470 750
rect 41515 630 41635 750
rect 41680 630 41800 750
rect 41845 630 41965 750
rect 36485 465 36605 585
rect 36660 465 36780 585
rect 36825 465 36945 585
rect 36990 465 37110 585
rect 37155 465 37275 585
rect 37330 465 37450 585
rect 37495 465 37615 585
rect 37660 465 37780 585
rect 37825 465 37945 585
rect 38000 465 38120 585
rect 38165 465 38285 585
rect 38330 465 38450 585
rect 38495 465 38615 585
rect 38670 465 38790 585
rect 38835 465 38955 585
rect 39000 465 39120 585
rect 39165 465 39285 585
rect 39340 465 39460 585
rect 39505 465 39625 585
rect 39670 465 39790 585
rect 39835 465 39955 585
rect 40010 465 40130 585
rect 40175 465 40295 585
rect 40340 465 40460 585
rect 40505 465 40625 585
rect 40680 465 40800 585
rect 40845 465 40965 585
rect 41010 465 41130 585
rect 41175 465 41295 585
rect 41350 465 41470 585
rect 41515 465 41635 585
rect 41680 465 41800 585
rect 41845 465 41965 585
rect 36485 300 36605 420
rect 36660 300 36780 420
rect 36825 300 36945 420
rect 36990 300 37110 420
rect 37155 300 37275 420
rect 37330 300 37450 420
rect 37495 300 37615 420
rect 37660 300 37780 420
rect 37825 300 37945 420
rect 38000 300 38120 420
rect 38165 300 38285 420
rect 38330 300 38450 420
rect 38495 300 38615 420
rect 38670 300 38790 420
rect 38835 300 38955 420
rect 39000 300 39120 420
rect 39165 300 39285 420
rect 39340 300 39460 420
rect 39505 300 39625 420
rect 39670 300 39790 420
rect 39835 300 39955 420
rect 40010 300 40130 420
rect 40175 300 40295 420
rect 40340 300 40460 420
rect 40505 300 40625 420
rect 40680 300 40800 420
rect 40845 300 40965 420
rect 41010 300 41130 420
rect 41175 300 41295 420
rect 41350 300 41470 420
rect 41515 300 41635 420
rect 41680 300 41800 420
rect 41845 300 41965 420
rect 36485 135 36605 255
rect 36660 135 36780 255
rect 36825 135 36945 255
rect 36990 135 37110 255
rect 37155 135 37275 255
rect 37330 135 37450 255
rect 37495 135 37615 255
rect 37660 135 37780 255
rect 37825 135 37945 255
rect 38000 135 38120 255
rect 38165 135 38285 255
rect 38330 135 38450 255
rect 38495 135 38615 255
rect 38670 135 38790 255
rect 38835 135 38955 255
rect 39000 135 39120 255
rect 39165 135 39285 255
rect 39340 135 39460 255
rect 39505 135 39625 255
rect 39670 135 39790 255
rect 39835 135 39955 255
rect 40010 135 40130 255
rect 40175 135 40295 255
rect 40340 135 40460 255
rect 40505 135 40625 255
rect 40680 135 40800 255
rect 40845 135 40965 255
rect 41010 135 41130 255
rect 41175 135 41295 255
rect 41350 135 41470 255
rect 41515 135 41635 255
rect 41680 135 41800 255
rect 41845 135 41965 255
rect 36485 -40 36605 80
rect 36660 -40 36780 80
rect 36825 -40 36945 80
rect 36990 -40 37110 80
rect 37155 -40 37275 80
rect 37330 -40 37450 80
rect 37495 -40 37615 80
rect 37660 -40 37780 80
rect 37825 -40 37945 80
rect 38000 -40 38120 80
rect 38165 -40 38285 80
rect 38330 -40 38450 80
rect 38495 -40 38615 80
rect 38670 -40 38790 80
rect 38835 -40 38955 80
rect 39000 -40 39120 80
rect 39165 -40 39285 80
rect 39340 -40 39460 80
rect 39505 -40 39625 80
rect 39670 -40 39790 80
rect 39835 -40 39955 80
rect 40010 -40 40130 80
rect 40175 -40 40295 80
rect 40340 -40 40460 80
rect 40505 -40 40625 80
rect 40680 -40 40800 80
rect 40845 -40 40965 80
rect 41010 -40 41130 80
rect 41175 -40 41295 80
rect 41350 -40 41470 80
rect 41515 -40 41635 80
rect 41680 -40 41800 80
rect 41845 -40 41965 80
rect 36485 -205 36605 -85
rect 36660 -205 36780 -85
rect 36825 -205 36945 -85
rect 36990 -205 37110 -85
rect 37155 -205 37275 -85
rect 37330 -205 37450 -85
rect 37495 -205 37615 -85
rect 37660 -205 37780 -85
rect 37825 -205 37945 -85
rect 38000 -205 38120 -85
rect 38165 -205 38285 -85
rect 38330 -205 38450 -85
rect 38495 -205 38615 -85
rect 38670 -205 38790 -85
rect 38835 -205 38955 -85
rect 39000 -205 39120 -85
rect 39165 -205 39285 -85
rect 39340 -205 39460 -85
rect 39505 -205 39625 -85
rect 39670 -205 39790 -85
rect 39835 -205 39955 -85
rect 40010 -205 40130 -85
rect 40175 -205 40295 -85
rect 40340 -205 40460 -85
rect 40505 -205 40625 -85
rect 40680 -205 40800 -85
rect 40845 -205 40965 -85
rect 41010 -205 41130 -85
rect 41175 -205 41295 -85
rect 41350 -205 41470 -85
rect 41515 -205 41635 -85
rect 41680 -205 41800 -85
rect 41845 -205 41965 -85
rect 36485 -370 36605 -250
rect 36660 -370 36780 -250
rect 36825 -370 36945 -250
rect 36990 -370 37110 -250
rect 37155 -370 37275 -250
rect 37330 -370 37450 -250
rect 37495 -370 37615 -250
rect 37660 -370 37780 -250
rect 37825 -370 37945 -250
rect 38000 -370 38120 -250
rect 38165 -370 38285 -250
rect 38330 -370 38450 -250
rect 38495 -370 38615 -250
rect 38670 -370 38790 -250
rect 38835 -370 38955 -250
rect 39000 -370 39120 -250
rect 39165 -370 39285 -250
rect 39340 -370 39460 -250
rect 39505 -370 39625 -250
rect 39670 -370 39790 -250
rect 39835 -370 39955 -250
rect 40010 -370 40130 -250
rect 40175 -370 40295 -250
rect 40340 -370 40460 -250
rect 40505 -370 40625 -250
rect 40680 -370 40800 -250
rect 40845 -370 40965 -250
rect 41010 -370 41130 -250
rect 41175 -370 41295 -250
rect 41350 -370 41470 -250
rect 41515 -370 41635 -250
rect 41680 -370 41800 -250
rect 41845 -370 41965 -250
rect 36485 -535 36605 -415
rect 36660 -535 36780 -415
rect 36825 -535 36945 -415
rect 36990 -535 37110 -415
rect 37155 -535 37275 -415
rect 37330 -535 37450 -415
rect 37495 -535 37615 -415
rect 37660 -535 37780 -415
rect 37825 -535 37945 -415
rect 38000 -535 38120 -415
rect 38165 -535 38285 -415
rect 38330 -535 38450 -415
rect 38495 -535 38615 -415
rect 38670 -535 38790 -415
rect 38835 -535 38955 -415
rect 39000 -535 39120 -415
rect 39165 -535 39285 -415
rect 39340 -535 39460 -415
rect 39505 -535 39625 -415
rect 39670 -535 39790 -415
rect 39835 -535 39955 -415
rect 40010 -535 40130 -415
rect 40175 -535 40295 -415
rect 40340 -535 40460 -415
rect 40505 -535 40625 -415
rect 40680 -535 40800 -415
rect 40845 -535 40965 -415
rect 41010 -535 41130 -415
rect 41175 -535 41295 -415
rect 41350 -535 41470 -415
rect 41515 -535 41635 -415
rect 41680 -535 41800 -415
rect 41845 -535 41965 -415
rect 36485 -710 36605 -590
rect 36660 -710 36780 -590
rect 36825 -710 36945 -590
rect 36990 -710 37110 -590
rect 37155 -710 37275 -590
rect 37330 -710 37450 -590
rect 37495 -710 37615 -590
rect 37660 -710 37780 -590
rect 37825 -710 37945 -590
rect 38000 -710 38120 -590
rect 38165 -710 38285 -590
rect 38330 -710 38450 -590
rect 38495 -710 38615 -590
rect 38670 -710 38790 -590
rect 38835 -710 38955 -590
rect 39000 -710 39120 -590
rect 39165 -710 39285 -590
rect 39340 -710 39460 -590
rect 39505 -710 39625 -590
rect 39670 -710 39790 -590
rect 39835 -710 39955 -590
rect 40010 -710 40130 -590
rect 40175 -710 40295 -590
rect 40340 -710 40460 -590
rect 40505 -710 40625 -590
rect 40680 -710 40800 -590
rect 40845 -710 40965 -590
rect 41010 -710 41130 -590
rect 41175 -710 41295 -590
rect 41350 -710 41470 -590
rect 41515 -710 41635 -590
rect 41680 -710 41800 -590
rect 41845 -710 41965 -590
rect 36485 -875 36605 -755
rect 36660 -875 36780 -755
rect 36825 -875 36945 -755
rect 36990 -875 37110 -755
rect 37155 -875 37275 -755
rect 37330 -875 37450 -755
rect 37495 -875 37615 -755
rect 37660 -875 37780 -755
rect 37825 -875 37945 -755
rect 38000 -875 38120 -755
rect 38165 -875 38285 -755
rect 38330 -875 38450 -755
rect 38495 -875 38615 -755
rect 38670 -875 38790 -755
rect 38835 -875 38955 -755
rect 39000 -875 39120 -755
rect 39165 -875 39285 -755
rect 39340 -875 39460 -755
rect 39505 -875 39625 -755
rect 39670 -875 39790 -755
rect 39835 -875 39955 -755
rect 40010 -875 40130 -755
rect 40175 -875 40295 -755
rect 40340 -875 40460 -755
rect 40505 -875 40625 -755
rect 40680 -875 40800 -755
rect 40845 -875 40965 -755
rect 41010 -875 41130 -755
rect 41175 -875 41295 -755
rect 41350 -875 41470 -755
rect 41515 -875 41635 -755
rect 41680 -875 41800 -755
rect 41845 -875 41965 -755
rect 36485 -1040 36605 -920
rect 36660 -1040 36780 -920
rect 36825 -1040 36945 -920
rect 36990 -1040 37110 -920
rect 37155 -1040 37275 -920
rect 37330 -1040 37450 -920
rect 37495 -1040 37615 -920
rect 37660 -1040 37780 -920
rect 37825 -1040 37945 -920
rect 38000 -1040 38120 -920
rect 38165 -1040 38285 -920
rect 38330 -1040 38450 -920
rect 38495 -1040 38615 -920
rect 38670 -1040 38790 -920
rect 38835 -1040 38955 -920
rect 39000 -1040 39120 -920
rect 39165 -1040 39285 -920
rect 39340 -1040 39460 -920
rect 39505 -1040 39625 -920
rect 39670 -1040 39790 -920
rect 39835 -1040 39955 -920
rect 40010 -1040 40130 -920
rect 40175 -1040 40295 -920
rect 40340 -1040 40460 -920
rect 40505 -1040 40625 -920
rect 40680 -1040 40800 -920
rect 40845 -1040 40965 -920
rect 41010 -1040 41130 -920
rect 41175 -1040 41295 -920
rect 41350 -1040 41470 -920
rect 41515 -1040 41635 -920
rect 41680 -1040 41800 -920
rect 41845 -1040 41965 -920
rect 36485 -1205 36605 -1085
rect 36660 -1205 36780 -1085
rect 36825 -1205 36945 -1085
rect 36990 -1205 37110 -1085
rect 37155 -1205 37275 -1085
rect 37330 -1205 37450 -1085
rect 37495 -1205 37615 -1085
rect 37660 -1205 37780 -1085
rect 37825 -1205 37945 -1085
rect 38000 -1205 38120 -1085
rect 38165 -1205 38285 -1085
rect 38330 -1205 38450 -1085
rect 38495 -1205 38615 -1085
rect 38670 -1205 38790 -1085
rect 38835 -1205 38955 -1085
rect 39000 -1205 39120 -1085
rect 39165 -1205 39285 -1085
rect 39340 -1205 39460 -1085
rect 39505 -1205 39625 -1085
rect 39670 -1205 39790 -1085
rect 39835 -1205 39955 -1085
rect 40010 -1205 40130 -1085
rect 40175 -1205 40295 -1085
rect 40340 -1205 40460 -1085
rect 40505 -1205 40625 -1085
rect 40680 -1205 40800 -1085
rect 40845 -1205 40965 -1085
rect 41010 -1205 41130 -1085
rect 41175 -1205 41295 -1085
rect 41350 -1205 41470 -1085
rect 41515 -1205 41635 -1085
rect 41680 -1205 41800 -1085
rect 41845 -1205 41965 -1085
rect 36485 -1380 36605 -1260
rect 36660 -1380 36780 -1260
rect 36825 -1380 36945 -1260
rect 36990 -1380 37110 -1260
rect 37155 -1380 37275 -1260
rect 37330 -1380 37450 -1260
rect 37495 -1380 37615 -1260
rect 37660 -1380 37780 -1260
rect 37825 -1380 37945 -1260
rect 38000 -1380 38120 -1260
rect 38165 -1380 38285 -1260
rect 38330 -1380 38450 -1260
rect 38495 -1380 38615 -1260
rect 38670 -1380 38790 -1260
rect 38835 -1380 38955 -1260
rect 39000 -1380 39120 -1260
rect 39165 -1380 39285 -1260
rect 39340 -1380 39460 -1260
rect 39505 -1380 39625 -1260
rect 39670 -1380 39790 -1260
rect 39835 -1380 39955 -1260
rect 40010 -1380 40130 -1260
rect 40175 -1380 40295 -1260
rect 40340 -1380 40460 -1260
rect 40505 -1380 40625 -1260
rect 40680 -1380 40800 -1260
rect 40845 -1380 40965 -1260
rect 41010 -1380 41130 -1260
rect 41175 -1380 41295 -1260
rect 41350 -1380 41470 -1260
rect 41515 -1380 41635 -1260
rect 41680 -1380 41800 -1260
rect 41845 -1380 41965 -1260
rect 36485 -1545 36605 -1425
rect 36660 -1545 36780 -1425
rect 36825 -1545 36945 -1425
rect 36990 -1545 37110 -1425
rect 37155 -1545 37275 -1425
rect 37330 -1545 37450 -1425
rect 37495 -1545 37615 -1425
rect 37660 -1545 37780 -1425
rect 37825 -1545 37945 -1425
rect 38000 -1545 38120 -1425
rect 38165 -1545 38285 -1425
rect 38330 -1545 38450 -1425
rect 38495 -1545 38615 -1425
rect 38670 -1545 38790 -1425
rect 38835 -1545 38955 -1425
rect 39000 -1545 39120 -1425
rect 39165 -1545 39285 -1425
rect 39340 -1545 39460 -1425
rect 39505 -1545 39625 -1425
rect 39670 -1545 39790 -1425
rect 39835 -1545 39955 -1425
rect 40010 -1545 40130 -1425
rect 40175 -1545 40295 -1425
rect 40340 -1545 40460 -1425
rect 40505 -1545 40625 -1425
rect 40680 -1545 40800 -1425
rect 40845 -1545 40965 -1425
rect 41010 -1545 41130 -1425
rect 41175 -1545 41295 -1425
rect 41350 -1545 41470 -1425
rect 41515 -1545 41635 -1425
rect 41680 -1545 41800 -1425
rect 41845 -1545 41965 -1425
rect 36485 -1710 36605 -1590
rect 36660 -1710 36780 -1590
rect 36825 -1710 36945 -1590
rect 36990 -1710 37110 -1590
rect 37155 -1710 37275 -1590
rect 37330 -1710 37450 -1590
rect 37495 -1710 37615 -1590
rect 37660 -1710 37780 -1590
rect 37825 -1710 37945 -1590
rect 38000 -1710 38120 -1590
rect 38165 -1710 38285 -1590
rect 38330 -1710 38450 -1590
rect 38495 -1710 38615 -1590
rect 38670 -1710 38790 -1590
rect 38835 -1710 38955 -1590
rect 39000 -1710 39120 -1590
rect 39165 -1710 39285 -1590
rect 39340 -1710 39460 -1590
rect 39505 -1710 39625 -1590
rect 39670 -1710 39790 -1590
rect 39835 -1710 39955 -1590
rect 40010 -1710 40130 -1590
rect 40175 -1710 40295 -1590
rect 40340 -1710 40460 -1590
rect 40505 -1710 40625 -1590
rect 40680 -1710 40800 -1590
rect 40845 -1710 40965 -1590
rect 41010 -1710 41130 -1590
rect 41175 -1710 41295 -1590
rect 41350 -1710 41470 -1590
rect 41515 -1710 41635 -1590
rect 41680 -1710 41800 -1590
rect 41845 -1710 41965 -1590
rect 36485 -1875 36605 -1755
rect 36660 -1875 36780 -1755
rect 36825 -1875 36945 -1755
rect 36990 -1875 37110 -1755
rect 37155 -1875 37275 -1755
rect 37330 -1875 37450 -1755
rect 37495 -1875 37615 -1755
rect 37660 -1875 37780 -1755
rect 37825 -1875 37945 -1755
rect 38000 -1875 38120 -1755
rect 38165 -1875 38285 -1755
rect 38330 -1875 38450 -1755
rect 38495 -1875 38615 -1755
rect 38670 -1875 38790 -1755
rect 38835 -1875 38955 -1755
rect 39000 -1875 39120 -1755
rect 39165 -1875 39285 -1755
rect 39340 -1875 39460 -1755
rect 39505 -1875 39625 -1755
rect 39670 -1875 39790 -1755
rect 39835 -1875 39955 -1755
rect 40010 -1875 40130 -1755
rect 40175 -1875 40295 -1755
rect 40340 -1875 40460 -1755
rect 40505 -1875 40625 -1755
rect 40680 -1875 40800 -1755
rect 40845 -1875 40965 -1755
rect 41010 -1875 41130 -1755
rect 41175 -1875 41295 -1755
rect 41350 -1875 41470 -1755
rect 41515 -1875 41635 -1755
rect 41680 -1875 41800 -1755
rect 41845 -1875 41965 -1755
rect 36485 -2050 36605 -1930
rect 36660 -2050 36780 -1930
rect 36825 -2050 36945 -1930
rect 36990 -2050 37110 -1930
rect 37155 -2050 37275 -1930
rect 37330 -2050 37450 -1930
rect 37495 -2050 37615 -1930
rect 37660 -2050 37780 -1930
rect 37825 -2050 37945 -1930
rect 38000 -2050 38120 -1930
rect 38165 -2050 38285 -1930
rect 38330 -2050 38450 -1930
rect 38495 -2050 38615 -1930
rect 38670 -2050 38790 -1930
rect 38835 -2050 38955 -1930
rect 39000 -2050 39120 -1930
rect 39165 -2050 39285 -1930
rect 39340 -2050 39460 -1930
rect 39505 -2050 39625 -1930
rect 39670 -2050 39790 -1930
rect 39835 -2050 39955 -1930
rect 40010 -2050 40130 -1930
rect 40175 -2050 40295 -1930
rect 40340 -2050 40460 -1930
rect 40505 -2050 40625 -1930
rect 40680 -2050 40800 -1930
rect 40845 -2050 40965 -1930
rect 41010 -2050 41130 -1930
rect 41175 -2050 41295 -1930
rect 41350 -2050 41470 -1930
rect 41515 -2050 41635 -1930
rect 41680 -2050 41800 -1930
rect 41845 -2050 41965 -1930
rect 36485 -2215 36605 -2095
rect 36660 -2215 36780 -2095
rect 36825 -2215 36945 -2095
rect 36990 -2215 37110 -2095
rect 37155 -2215 37275 -2095
rect 37330 -2215 37450 -2095
rect 37495 -2215 37615 -2095
rect 37660 -2215 37780 -2095
rect 37825 -2215 37945 -2095
rect 38000 -2215 38120 -2095
rect 38165 -2215 38285 -2095
rect 38330 -2215 38450 -2095
rect 38495 -2215 38615 -2095
rect 38670 -2215 38790 -2095
rect 38835 -2215 38955 -2095
rect 39000 -2215 39120 -2095
rect 39165 -2215 39285 -2095
rect 39340 -2215 39460 -2095
rect 39505 -2215 39625 -2095
rect 39670 -2215 39790 -2095
rect 39835 -2215 39955 -2095
rect 40010 -2215 40130 -2095
rect 40175 -2215 40295 -2095
rect 40340 -2215 40460 -2095
rect 40505 -2215 40625 -2095
rect 40680 -2215 40800 -2095
rect 40845 -2215 40965 -2095
rect 41010 -2215 41130 -2095
rect 41175 -2215 41295 -2095
rect 41350 -2215 41470 -2095
rect 41515 -2215 41635 -2095
rect 41680 -2215 41800 -2095
rect 41845 -2215 41965 -2095
rect 36485 -2380 36605 -2260
rect 36660 -2380 36780 -2260
rect 36825 -2380 36945 -2260
rect 36990 -2380 37110 -2260
rect 37155 -2380 37275 -2260
rect 37330 -2380 37450 -2260
rect 37495 -2380 37615 -2260
rect 37660 -2380 37780 -2260
rect 37825 -2380 37945 -2260
rect 38000 -2380 38120 -2260
rect 38165 -2380 38285 -2260
rect 38330 -2380 38450 -2260
rect 38495 -2380 38615 -2260
rect 38670 -2380 38790 -2260
rect 38835 -2380 38955 -2260
rect 39000 -2380 39120 -2260
rect 39165 -2380 39285 -2260
rect 39340 -2380 39460 -2260
rect 39505 -2380 39625 -2260
rect 39670 -2380 39790 -2260
rect 39835 -2380 39955 -2260
rect 40010 -2380 40130 -2260
rect 40175 -2380 40295 -2260
rect 40340 -2380 40460 -2260
rect 40505 -2380 40625 -2260
rect 40680 -2380 40800 -2260
rect 40845 -2380 40965 -2260
rect 41010 -2380 41130 -2260
rect 41175 -2380 41295 -2260
rect 41350 -2380 41470 -2260
rect 41515 -2380 41635 -2260
rect 41680 -2380 41800 -2260
rect 41845 -2380 41965 -2260
rect 36485 -2545 36605 -2425
rect 36660 -2545 36780 -2425
rect 36825 -2545 36945 -2425
rect 36990 -2545 37110 -2425
rect 37155 -2545 37275 -2425
rect 37330 -2545 37450 -2425
rect 37495 -2545 37615 -2425
rect 37660 -2545 37780 -2425
rect 37825 -2545 37945 -2425
rect 38000 -2545 38120 -2425
rect 38165 -2545 38285 -2425
rect 38330 -2545 38450 -2425
rect 38495 -2545 38615 -2425
rect 38670 -2545 38790 -2425
rect 38835 -2545 38955 -2425
rect 39000 -2545 39120 -2425
rect 39165 -2545 39285 -2425
rect 39340 -2545 39460 -2425
rect 39505 -2545 39625 -2425
rect 39670 -2545 39790 -2425
rect 39835 -2545 39955 -2425
rect 40010 -2545 40130 -2425
rect 40175 -2545 40295 -2425
rect 40340 -2545 40460 -2425
rect 40505 -2545 40625 -2425
rect 40680 -2545 40800 -2425
rect 40845 -2545 40965 -2425
rect 41010 -2545 41130 -2425
rect 41175 -2545 41295 -2425
rect 41350 -2545 41470 -2425
rect 41515 -2545 41635 -2425
rect 41680 -2545 41800 -2425
rect 41845 -2545 41965 -2425
rect 36485 -2720 36605 -2600
rect 36660 -2720 36780 -2600
rect 36825 -2720 36945 -2600
rect 36990 -2720 37110 -2600
rect 37155 -2720 37275 -2600
rect 37330 -2720 37450 -2600
rect 37495 -2720 37615 -2600
rect 37660 -2720 37780 -2600
rect 37825 -2720 37945 -2600
rect 38000 -2720 38120 -2600
rect 38165 -2720 38285 -2600
rect 38330 -2720 38450 -2600
rect 38495 -2720 38615 -2600
rect 38670 -2720 38790 -2600
rect 38835 -2720 38955 -2600
rect 39000 -2720 39120 -2600
rect 39165 -2720 39285 -2600
rect 39340 -2720 39460 -2600
rect 39505 -2720 39625 -2600
rect 39670 -2720 39790 -2600
rect 39835 -2720 39955 -2600
rect 40010 -2720 40130 -2600
rect 40175 -2720 40295 -2600
rect 40340 -2720 40460 -2600
rect 40505 -2720 40625 -2600
rect 40680 -2720 40800 -2600
rect 40845 -2720 40965 -2600
rect 41010 -2720 41130 -2600
rect 41175 -2720 41295 -2600
rect 41350 -2720 41470 -2600
rect 41515 -2720 41635 -2600
rect 41680 -2720 41800 -2600
rect 41845 -2720 41965 -2600
rect 36485 -2885 36605 -2765
rect 36660 -2885 36780 -2765
rect 36825 -2885 36945 -2765
rect 36990 -2885 37110 -2765
rect 37155 -2885 37275 -2765
rect 37330 -2885 37450 -2765
rect 37495 -2885 37615 -2765
rect 37660 -2885 37780 -2765
rect 37825 -2885 37945 -2765
rect 38000 -2885 38120 -2765
rect 38165 -2885 38285 -2765
rect 38330 -2885 38450 -2765
rect 38495 -2885 38615 -2765
rect 38670 -2885 38790 -2765
rect 38835 -2885 38955 -2765
rect 39000 -2885 39120 -2765
rect 39165 -2885 39285 -2765
rect 39340 -2885 39460 -2765
rect 39505 -2885 39625 -2765
rect 39670 -2885 39790 -2765
rect 39835 -2885 39955 -2765
rect 40010 -2885 40130 -2765
rect 40175 -2885 40295 -2765
rect 40340 -2885 40460 -2765
rect 40505 -2885 40625 -2765
rect 40680 -2885 40800 -2765
rect 40845 -2885 40965 -2765
rect 41010 -2885 41130 -2765
rect 41175 -2885 41295 -2765
rect 41350 -2885 41470 -2765
rect 41515 -2885 41635 -2765
rect 41680 -2885 41800 -2765
rect 41845 -2885 41965 -2765
rect 36485 -3050 36605 -2930
rect 36660 -3050 36780 -2930
rect 36825 -3050 36945 -2930
rect 36990 -3050 37110 -2930
rect 37155 -3050 37275 -2930
rect 37330 -3050 37450 -2930
rect 37495 -3050 37615 -2930
rect 37660 -3050 37780 -2930
rect 37825 -3050 37945 -2930
rect 38000 -3050 38120 -2930
rect 38165 -3050 38285 -2930
rect 38330 -3050 38450 -2930
rect 38495 -3050 38615 -2930
rect 38670 -3050 38790 -2930
rect 38835 -3050 38955 -2930
rect 39000 -3050 39120 -2930
rect 39165 -3050 39285 -2930
rect 39340 -3050 39460 -2930
rect 39505 -3050 39625 -2930
rect 39670 -3050 39790 -2930
rect 39835 -3050 39955 -2930
rect 40010 -3050 40130 -2930
rect 40175 -3050 40295 -2930
rect 40340 -3050 40460 -2930
rect 40505 -3050 40625 -2930
rect 40680 -3050 40800 -2930
rect 40845 -3050 40965 -2930
rect 41010 -3050 41130 -2930
rect 41175 -3050 41295 -2930
rect 41350 -3050 41470 -2930
rect 41515 -3050 41635 -2930
rect 41680 -3050 41800 -2930
rect 41845 -3050 41965 -2930
rect 36485 -3215 36605 -3095
rect 36660 -3215 36780 -3095
rect 36825 -3215 36945 -3095
rect 36990 -3215 37110 -3095
rect 37155 -3215 37275 -3095
rect 37330 -3215 37450 -3095
rect 37495 -3215 37615 -3095
rect 37660 -3215 37780 -3095
rect 37825 -3215 37945 -3095
rect 38000 -3215 38120 -3095
rect 38165 -3215 38285 -3095
rect 38330 -3215 38450 -3095
rect 38495 -3215 38615 -3095
rect 38670 -3215 38790 -3095
rect 38835 -3215 38955 -3095
rect 39000 -3215 39120 -3095
rect 39165 -3215 39285 -3095
rect 39340 -3215 39460 -3095
rect 39505 -3215 39625 -3095
rect 39670 -3215 39790 -3095
rect 39835 -3215 39955 -3095
rect 40010 -3215 40130 -3095
rect 40175 -3215 40295 -3095
rect 40340 -3215 40460 -3095
rect 40505 -3215 40625 -3095
rect 40680 -3215 40800 -3095
rect 40845 -3215 40965 -3095
rect 41010 -3215 41130 -3095
rect 41175 -3215 41295 -3095
rect 41350 -3215 41470 -3095
rect 41515 -3215 41635 -3095
rect 41680 -3215 41800 -3095
rect 41845 -3215 41965 -3095
rect 36485 -3390 36605 -3270
rect 36660 -3390 36780 -3270
rect 36825 -3390 36945 -3270
rect 36990 -3390 37110 -3270
rect 37155 -3390 37275 -3270
rect 37330 -3390 37450 -3270
rect 37495 -3390 37615 -3270
rect 37660 -3390 37780 -3270
rect 37825 -3390 37945 -3270
rect 38000 -3390 38120 -3270
rect 38165 -3390 38285 -3270
rect 38330 -3390 38450 -3270
rect 38495 -3390 38615 -3270
rect 38670 -3390 38790 -3270
rect 38835 -3390 38955 -3270
rect 39000 -3390 39120 -3270
rect 39165 -3390 39285 -3270
rect 39340 -3390 39460 -3270
rect 39505 -3390 39625 -3270
rect 39670 -3390 39790 -3270
rect 39835 -3390 39955 -3270
rect 40010 -3390 40130 -3270
rect 40175 -3390 40295 -3270
rect 40340 -3390 40460 -3270
rect 40505 -3390 40625 -3270
rect 40680 -3390 40800 -3270
rect 40845 -3390 40965 -3270
rect 41010 -3390 41130 -3270
rect 41175 -3390 41295 -3270
rect 41350 -3390 41470 -3270
rect 41515 -3390 41635 -3270
rect 41680 -3390 41800 -3270
rect 41845 -3390 41965 -3270
rect 36485 -3555 36605 -3435
rect 36660 -3555 36780 -3435
rect 36825 -3555 36945 -3435
rect 36990 -3555 37110 -3435
rect 37155 -3555 37275 -3435
rect 37330 -3555 37450 -3435
rect 37495 -3555 37615 -3435
rect 37660 -3555 37780 -3435
rect 37825 -3555 37945 -3435
rect 38000 -3555 38120 -3435
rect 38165 -3555 38285 -3435
rect 38330 -3555 38450 -3435
rect 38495 -3555 38615 -3435
rect 38670 -3555 38790 -3435
rect 38835 -3555 38955 -3435
rect 39000 -3555 39120 -3435
rect 39165 -3555 39285 -3435
rect 39340 -3555 39460 -3435
rect 39505 -3555 39625 -3435
rect 39670 -3555 39790 -3435
rect 39835 -3555 39955 -3435
rect 40010 -3555 40130 -3435
rect 40175 -3555 40295 -3435
rect 40340 -3555 40460 -3435
rect 40505 -3555 40625 -3435
rect 40680 -3555 40800 -3435
rect 40845 -3555 40965 -3435
rect 41010 -3555 41130 -3435
rect 41175 -3555 41295 -3435
rect 41350 -3555 41470 -3435
rect 41515 -3555 41635 -3435
rect 41680 -3555 41800 -3435
rect 41845 -3555 41965 -3435
rect 36485 -3720 36605 -3600
rect 36660 -3720 36780 -3600
rect 36825 -3720 36945 -3600
rect 36990 -3720 37110 -3600
rect 37155 -3720 37275 -3600
rect 37330 -3720 37450 -3600
rect 37495 -3720 37615 -3600
rect 37660 -3720 37780 -3600
rect 37825 -3720 37945 -3600
rect 38000 -3720 38120 -3600
rect 38165 -3720 38285 -3600
rect 38330 -3720 38450 -3600
rect 38495 -3720 38615 -3600
rect 38670 -3720 38790 -3600
rect 38835 -3720 38955 -3600
rect 39000 -3720 39120 -3600
rect 39165 -3720 39285 -3600
rect 39340 -3720 39460 -3600
rect 39505 -3720 39625 -3600
rect 39670 -3720 39790 -3600
rect 39835 -3720 39955 -3600
rect 40010 -3720 40130 -3600
rect 40175 -3720 40295 -3600
rect 40340 -3720 40460 -3600
rect 40505 -3720 40625 -3600
rect 40680 -3720 40800 -3600
rect 40845 -3720 40965 -3600
rect 41010 -3720 41130 -3600
rect 41175 -3720 41295 -3600
rect 41350 -3720 41470 -3600
rect 41515 -3720 41635 -3600
rect 41680 -3720 41800 -3600
rect 41845 -3720 41965 -3600
rect 36485 -3885 36605 -3765
rect 36660 -3885 36780 -3765
rect 36825 -3885 36945 -3765
rect 36990 -3885 37110 -3765
rect 37155 -3885 37275 -3765
rect 37330 -3885 37450 -3765
rect 37495 -3885 37615 -3765
rect 37660 -3885 37780 -3765
rect 37825 -3885 37945 -3765
rect 38000 -3885 38120 -3765
rect 38165 -3885 38285 -3765
rect 38330 -3885 38450 -3765
rect 38495 -3885 38615 -3765
rect 38670 -3885 38790 -3765
rect 38835 -3885 38955 -3765
rect 39000 -3885 39120 -3765
rect 39165 -3885 39285 -3765
rect 39340 -3885 39460 -3765
rect 39505 -3885 39625 -3765
rect 39670 -3885 39790 -3765
rect 39835 -3885 39955 -3765
rect 40010 -3885 40130 -3765
rect 40175 -3885 40295 -3765
rect 40340 -3885 40460 -3765
rect 40505 -3885 40625 -3765
rect 40680 -3885 40800 -3765
rect 40845 -3885 40965 -3765
rect 41010 -3885 41130 -3765
rect 41175 -3885 41295 -3765
rect 41350 -3885 41470 -3765
rect 41515 -3885 41635 -3765
rect 41680 -3885 41800 -3765
rect 41845 -3885 41965 -3765
rect 36485 -4060 36605 -3940
rect 36660 -4060 36780 -3940
rect 36825 -4060 36945 -3940
rect 36990 -4060 37110 -3940
rect 37155 -4060 37275 -3940
rect 37330 -4060 37450 -3940
rect 37495 -4060 37615 -3940
rect 37660 -4060 37780 -3940
rect 37825 -4060 37945 -3940
rect 38000 -4060 38120 -3940
rect 38165 -4060 38285 -3940
rect 38330 -4060 38450 -3940
rect 38495 -4060 38615 -3940
rect 38670 -4060 38790 -3940
rect 38835 -4060 38955 -3940
rect 39000 -4060 39120 -3940
rect 39165 -4060 39285 -3940
rect 39340 -4060 39460 -3940
rect 39505 -4060 39625 -3940
rect 39670 -4060 39790 -3940
rect 39835 -4060 39955 -3940
rect 40010 -4060 40130 -3940
rect 40175 -4060 40295 -3940
rect 40340 -4060 40460 -3940
rect 40505 -4060 40625 -3940
rect 40680 -4060 40800 -3940
rect 40845 -4060 40965 -3940
rect 41010 -4060 41130 -3940
rect 41175 -4060 41295 -3940
rect 41350 -4060 41470 -3940
rect 41515 -4060 41635 -3940
rect 41680 -4060 41800 -3940
rect 41845 -4060 41965 -3940
rect 42175 1300 42295 1420
rect 42350 1300 42470 1420
rect 42515 1300 42635 1420
rect 42680 1300 42800 1420
rect 42845 1300 42965 1420
rect 43020 1300 43140 1420
rect 43185 1300 43305 1420
rect 43350 1300 43470 1420
rect 43515 1300 43635 1420
rect 43690 1300 43810 1420
rect 43855 1300 43975 1420
rect 44020 1300 44140 1420
rect 44185 1300 44305 1420
rect 44360 1300 44480 1420
rect 44525 1300 44645 1420
rect 44690 1300 44810 1420
rect 44855 1300 44975 1420
rect 45030 1300 45150 1420
rect 45195 1300 45315 1420
rect 45360 1300 45480 1420
rect 45525 1300 45645 1420
rect 45700 1300 45820 1420
rect 45865 1300 45985 1420
rect 46030 1300 46150 1420
rect 46195 1300 46315 1420
rect 46370 1300 46490 1420
rect 46535 1300 46655 1420
rect 46700 1300 46820 1420
rect 46865 1300 46985 1420
rect 47040 1300 47160 1420
rect 47205 1300 47325 1420
rect 47370 1300 47490 1420
rect 47535 1300 47655 1420
rect 42175 1135 42295 1255
rect 42350 1135 42470 1255
rect 42515 1135 42635 1255
rect 42680 1135 42800 1255
rect 42845 1135 42965 1255
rect 43020 1135 43140 1255
rect 43185 1135 43305 1255
rect 43350 1135 43470 1255
rect 43515 1135 43635 1255
rect 43690 1135 43810 1255
rect 43855 1135 43975 1255
rect 44020 1135 44140 1255
rect 44185 1135 44305 1255
rect 44360 1135 44480 1255
rect 44525 1135 44645 1255
rect 44690 1135 44810 1255
rect 44855 1135 44975 1255
rect 45030 1135 45150 1255
rect 45195 1135 45315 1255
rect 45360 1135 45480 1255
rect 45525 1135 45645 1255
rect 45700 1135 45820 1255
rect 45865 1135 45985 1255
rect 46030 1135 46150 1255
rect 46195 1135 46315 1255
rect 46370 1135 46490 1255
rect 46535 1135 46655 1255
rect 46700 1135 46820 1255
rect 46865 1135 46985 1255
rect 47040 1135 47160 1255
rect 47205 1135 47325 1255
rect 47370 1135 47490 1255
rect 47535 1135 47655 1255
rect 42175 970 42295 1090
rect 42350 970 42470 1090
rect 42515 970 42635 1090
rect 42680 970 42800 1090
rect 42845 970 42965 1090
rect 43020 970 43140 1090
rect 43185 970 43305 1090
rect 43350 970 43470 1090
rect 43515 970 43635 1090
rect 43690 970 43810 1090
rect 43855 970 43975 1090
rect 44020 970 44140 1090
rect 44185 970 44305 1090
rect 44360 970 44480 1090
rect 44525 970 44645 1090
rect 44690 970 44810 1090
rect 44855 970 44975 1090
rect 45030 970 45150 1090
rect 45195 970 45315 1090
rect 45360 970 45480 1090
rect 45525 970 45645 1090
rect 45700 970 45820 1090
rect 45865 970 45985 1090
rect 46030 970 46150 1090
rect 46195 970 46315 1090
rect 46370 970 46490 1090
rect 46535 970 46655 1090
rect 46700 970 46820 1090
rect 46865 970 46985 1090
rect 47040 970 47160 1090
rect 47205 970 47325 1090
rect 47370 970 47490 1090
rect 47535 970 47655 1090
rect 42175 805 42295 925
rect 42350 805 42470 925
rect 42515 805 42635 925
rect 42680 805 42800 925
rect 42845 805 42965 925
rect 43020 805 43140 925
rect 43185 805 43305 925
rect 43350 805 43470 925
rect 43515 805 43635 925
rect 43690 805 43810 925
rect 43855 805 43975 925
rect 44020 805 44140 925
rect 44185 805 44305 925
rect 44360 805 44480 925
rect 44525 805 44645 925
rect 44690 805 44810 925
rect 44855 805 44975 925
rect 45030 805 45150 925
rect 45195 805 45315 925
rect 45360 805 45480 925
rect 45525 805 45645 925
rect 45700 805 45820 925
rect 45865 805 45985 925
rect 46030 805 46150 925
rect 46195 805 46315 925
rect 46370 805 46490 925
rect 46535 805 46655 925
rect 46700 805 46820 925
rect 46865 805 46985 925
rect 47040 805 47160 925
rect 47205 805 47325 925
rect 47370 805 47490 925
rect 47535 805 47655 925
rect 42175 630 42295 750
rect 42350 630 42470 750
rect 42515 630 42635 750
rect 42680 630 42800 750
rect 42845 630 42965 750
rect 43020 630 43140 750
rect 43185 630 43305 750
rect 43350 630 43470 750
rect 43515 630 43635 750
rect 43690 630 43810 750
rect 43855 630 43975 750
rect 44020 630 44140 750
rect 44185 630 44305 750
rect 44360 630 44480 750
rect 44525 630 44645 750
rect 44690 630 44810 750
rect 44855 630 44975 750
rect 45030 630 45150 750
rect 45195 630 45315 750
rect 45360 630 45480 750
rect 45525 630 45645 750
rect 45700 630 45820 750
rect 45865 630 45985 750
rect 46030 630 46150 750
rect 46195 630 46315 750
rect 46370 630 46490 750
rect 46535 630 46655 750
rect 46700 630 46820 750
rect 46865 630 46985 750
rect 47040 630 47160 750
rect 47205 630 47325 750
rect 47370 630 47490 750
rect 47535 630 47655 750
rect 42175 465 42295 585
rect 42350 465 42470 585
rect 42515 465 42635 585
rect 42680 465 42800 585
rect 42845 465 42965 585
rect 43020 465 43140 585
rect 43185 465 43305 585
rect 43350 465 43470 585
rect 43515 465 43635 585
rect 43690 465 43810 585
rect 43855 465 43975 585
rect 44020 465 44140 585
rect 44185 465 44305 585
rect 44360 465 44480 585
rect 44525 465 44645 585
rect 44690 465 44810 585
rect 44855 465 44975 585
rect 45030 465 45150 585
rect 45195 465 45315 585
rect 45360 465 45480 585
rect 45525 465 45645 585
rect 45700 465 45820 585
rect 45865 465 45985 585
rect 46030 465 46150 585
rect 46195 465 46315 585
rect 46370 465 46490 585
rect 46535 465 46655 585
rect 46700 465 46820 585
rect 46865 465 46985 585
rect 47040 465 47160 585
rect 47205 465 47325 585
rect 47370 465 47490 585
rect 47535 465 47655 585
rect 42175 300 42295 420
rect 42350 300 42470 420
rect 42515 300 42635 420
rect 42680 300 42800 420
rect 42845 300 42965 420
rect 43020 300 43140 420
rect 43185 300 43305 420
rect 43350 300 43470 420
rect 43515 300 43635 420
rect 43690 300 43810 420
rect 43855 300 43975 420
rect 44020 300 44140 420
rect 44185 300 44305 420
rect 44360 300 44480 420
rect 44525 300 44645 420
rect 44690 300 44810 420
rect 44855 300 44975 420
rect 45030 300 45150 420
rect 45195 300 45315 420
rect 45360 300 45480 420
rect 45525 300 45645 420
rect 45700 300 45820 420
rect 45865 300 45985 420
rect 46030 300 46150 420
rect 46195 300 46315 420
rect 46370 300 46490 420
rect 46535 300 46655 420
rect 46700 300 46820 420
rect 46865 300 46985 420
rect 47040 300 47160 420
rect 47205 300 47325 420
rect 47370 300 47490 420
rect 47535 300 47655 420
rect 42175 135 42295 255
rect 42350 135 42470 255
rect 42515 135 42635 255
rect 42680 135 42800 255
rect 42845 135 42965 255
rect 43020 135 43140 255
rect 43185 135 43305 255
rect 43350 135 43470 255
rect 43515 135 43635 255
rect 43690 135 43810 255
rect 43855 135 43975 255
rect 44020 135 44140 255
rect 44185 135 44305 255
rect 44360 135 44480 255
rect 44525 135 44645 255
rect 44690 135 44810 255
rect 44855 135 44975 255
rect 45030 135 45150 255
rect 45195 135 45315 255
rect 45360 135 45480 255
rect 45525 135 45645 255
rect 45700 135 45820 255
rect 45865 135 45985 255
rect 46030 135 46150 255
rect 46195 135 46315 255
rect 46370 135 46490 255
rect 46535 135 46655 255
rect 46700 135 46820 255
rect 46865 135 46985 255
rect 47040 135 47160 255
rect 47205 135 47325 255
rect 47370 135 47490 255
rect 47535 135 47655 255
rect 42175 -40 42295 80
rect 42350 -40 42470 80
rect 42515 -40 42635 80
rect 42680 -40 42800 80
rect 42845 -40 42965 80
rect 43020 -40 43140 80
rect 43185 -40 43305 80
rect 43350 -40 43470 80
rect 43515 -40 43635 80
rect 43690 -40 43810 80
rect 43855 -40 43975 80
rect 44020 -40 44140 80
rect 44185 -40 44305 80
rect 44360 -40 44480 80
rect 44525 -40 44645 80
rect 44690 -40 44810 80
rect 44855 -40 44975 80
rect 45030 -40 45150 80
rect 45195 -40 45315 80
rect 45360 -40 45480 80
rect 45525 -40 45645 80
rect 45700 -40 45820 80
rect 45865 -40 45985 80
rect 46030 -40 46150 80
rect 46195 -40 46315 80
rect 46370 -40 46490 80
rect 46535 -40 46655 80
rect 46700 -40 46820 80
rect 46865 -40 46985 80
rect 47040 -40 47160 80
rect 47205 -40 47325 80
rect 47370 -40 47490 80
rect 47535 -40 47655 80
rect 42175 -205 42295 -85
rect 42350 -205 42470 -85
rect 42515 -205 42635 -85
rect 42680 -205 42800 -85
rect 42845 -205 42965 -85
rect 43020 -205 43140 -85
rect 43185 -205 43305 -85
rect 43350 -205 43470 -85
rect 43515 -205 43635 -85
rect 43690 -205 43810 -85
rect 43855 -205 43975 -85
rect 44020 -205 44140 -85
rect 44185 -205 44305 -85
rect 44360 -205 44480 -85
rect 44525 -205 44645 -85
rect 44690 -205 44810 -85
rect 44855 -205 44975 -85
rect 45030 -205 45150 -85
rect 45195 -205 45315 -85
rect 45360 -205 45480 -85
rect 45525 -205 45645 -85
rect 45700 -205 45820 -85
rect 45865 -205 45985 -85
rect 46030 -205 46150 -85
rect 46195 -205 46315 -85
rect 46370 -205 46490 -85
rect 46535 -205 46655 -85
rect 46700 -205 46820 -85
rect 46865 -205 46985 -85
rect 47040 -205 47160 -85
rect 47205 -205 47325 -85
rect 47370 -205 47490 -85
rect 47535 -205 47655 -85
rect 42175 -370 42295 -250
rect 42350 -370 42470 -250
rect 42515 -370 42635 -250
rect 42680 -370 42800 -250
rect 42845 -370 42965 -250
rect 43020 -370 43140 -250
rect 43185 -370 43305 -250
rect 43350 -370 43470 -250
rect 43515 -370 43635 -250
rect 43690 -370 43810 -250
rect 43855 -370 43975 -250
rect 44020 -370 44140 -250
rect 44185 -370 44305 -250
rect 44360 -370 44480 -250
rect 44525 -370 44645 -250
rect 44690 -370 44810 -250
rect 44855 -370 44975 -250
rect 45030 -370 45150 -250
rect 45195 -370 45315 -250
rect 45360 -370 45480 -250
rect 45525 -370 45645 -250
rect 45700 -370 45820 -250
rect 45865 -370 45985 -250
rect 46030 -370 46150 -250
rect 46195 -370 46315 -250
rect 46370 -370 46490 -250
rect 46535 -370 46655 -250
rect 46700 -370 46820 -250
rect 46865 -370 46985 -250
rect 47040 -370 47160 -250
rect 47205 -370 47325 -250
rect 47370 -370 47490 -250
rect 47535 -370 47655 -250
rect 42175 -535 42295 -415
rect 42350 -535 42470 -415
rect 42515 -535 42635 -415
rect 42680 -535 42800 -415
rect 42845 -535 42965 -415
rect 43020 -535 43140 -415
rect 43185 -535 43305 -415
rect 43350 -535 43470 -415
rect 43515 -535 43635 -415
rect 43690 -535 43810 -415
rect 43855 -535 43975 -415
rect 44020 -535 44140 -415
rect 44185 -535 44305 -415
rect 44360 -535 44480 -415
rect 44525 -535 44645 -415
rect 44690 -535 44810 -415
rect 44855 -535 44975 -415
rect 45030 -535 45150 -415
rect 45195 -535 45315 -415
rect 45360 -535 45480 -415
rect 45525 -535 45645 -415
rect 45700 -535 45820 -415
rect 45865 -535 45985 -415
rect 46030 -535 46150 -415
rect 46195 -535 46315 -415
rect 46370 -535 46490 -415
rect 46535 -535 46655 -415
rect 46700 -535 46820 -415
rect 46865 -535 46985 -415
rect 47040 -535 47160 -415
rect 47205 -535 47325 -415
rect 47370 -535 47490 -415
rect 47535 -535 47655 -415
rect 42175 -710 42295 -590
rect 42350 -710 42470 -590
rect 42515 -710 42635 -590
rect 42680 -710 42800 -590
rect 42845 -710 42965 -590
rect 43020 -710 43140 -590
rect 43185 -710 43305 -590
rect 43350 -710 43470 -590
rect 43515 -710 43635 -590
rect 43690 -710 43810 -590
rect 43855 -710 43975 -590
rect 44020 -710 44140 -590
rect 44185 -710 44305 -590
rect 44360 -710 44480 -590
rect 44525 -710 44645 -590
rect 44690 -710 44810 -590
rect 44855 -710 44975 -590
rect 45030 -710 45150 -590
rect 45195 -710 45315 -590
rect 45360 -710 45480 -590
rect 45525 -710 45645 -590
rect 45700 -710 45820 -590
rect 45865 -710 45985 -590
rect 46030 -710 46150 -590
rect 46195 -710 46315 -590
rect 46370 -710 46490 -590
rect 46535 -710 46655 -590
rect 46700 -710 46820 -590
rect 46865 -710 46985 -590
rect 47040 -710 47160 -590
rect 47205 -710 47325 -590
rect 47370 -710 47490 -590
rect 47535 -710 47655 -590
rect 42175 -875 42295 -755
rect 42350 -875 42470 -755
rect 42515 -875 42635 -755
rect 42680 -875 42800 -755
rect 42845 -875 42965 -755
rect 43020 -875 43140 -755
rect 43185 -875 43305 -755
rect 43350 -875 43470 -755
rect 43515 -875 43635 -755
rect 43690 -875 43810 -755
rect 43855 -875 43975 -755
rect 44020 -875 44140 -755
rect 44185 -875 44305 -755
rect 44360 -875 44480 -755
rect 44525 -875 44645 -755
rect 44690 -875 44810 -755
rect 44855 -875 44975 -755
rect 45030 -875 45150 -755
rect 45195 -875 45315 -755
rect 45360 -875 45480 -755
rect 45525 -875 45645 -755
rect 45700 -875 45820 -755
rect 45865 -875 45985 -755
rect 46030 -875 46150 -755
rect 46195 -875 46315 -755
rect 46370 -875 46490 -755
rect 46535 -875 46655 -755
rect 46700 -875 46820 -755
rect 46865 -875 46985 -755
rect 47040 -875 47160 -755
rect 47205 -875 47325 -755
rect 47370 -875 47490 -755
rect 47535 -875 47655 -755
rect 42175 -1040 42295 -920
rect 42350 -1040 42470 -920
rect 42515 -1040 42635 -920
rect 42680 -1040 42800 -920
rect 42845 -1040 42965 -920
rect 43020 -1040 43140 -920
rect 43185 -1040 43305 -920
rect 43350 -1040 43470 -920
rect 43515 -1040 43635 -920
rect 43690 -1040 43810 -920
rect 43855 -1040 43975 -920
rect 44020 -1040 44140 -920
rect 44185 -1040 44305 -920
rect 44360 -1040 44480 -920
rect 44525 -1040 44645 -920
rect 44690 -1040 44810 -920
rect 44855 -1040 44975 -920
rect 45030 -1040 45150 -920
rect 45195 -1040 45315 -920
rect 45360 -1040 45480 -920
rect 45525 -1040 45645 -920
rect 45700 -1040 45820 -920
rect 45865 -1040 45985 -920
rect 46030 -1040 46150 -920
rect 46195 -1040 46315 -920
rect 46370 -1040 46490 -920
rect 46535 -1040 46655 -920
rect 46700 -1040 46820 -920
rect 46865 -1040 46985 -920
rect 47040 -1040 47160 -920
rect 47205 -1040 47325 -920
rect 47370 -1040 47490 -920
rect 47535 -1040 47655 -920
rect 42175 -1205 42295 -1085
rect 42350 -1205 42470 -1085
rect 42515 -1205 42635 -1085
rect 42680 -1205 42800 -1085
rect 42845 -1205 42965 -1085
rect 43020 -1205 43140 -1085
rect 43185 -1205 43305 -1085
rect 43350 -1205 43470 -1085
rect 43515 -1205 43635 -1085
rect 43690 -1205 43810 -1085
rect 43855 -1205 43975 -1085
rect 44020 -1205 44140 -1085
rect 44185 -1205 44305 -1085
rect 44360 -1205 44480 -1085
rect 44525 -1205 44645 -1085
rect 44690 -1205 44810 -1085
rect 44855 -1205 44975 -1085
rect 45030 -1205 45150 -1085
rect 45195 -1205 45315 -1085
rect 45360 -1205 45480 -1085
rect 45525 -1205 45645 -1085
rect 45700 -1205 45820 -1085
rect 45865 -1205 45985 -1085
rect 46030 -1205 46150 -1085
rect 46195 -1205 46315 -1085
rect 46370 -1205 46490 -1085
rect 46535 -1205 46655 -1085
rect 46700 -1205 46820 -1085
rect 46865 -1205 46985 -1085
rect 47040 -1205 47160 -1085
rect 47205 -1205 47325 -1085
rect 47370 -1205 47490 -1085
rect 47535 -1205 47655 -1085
rect 42175 -1380 42295 -1260
rect 42350 -1380 42470 -1260
rect 42515 -1380 42635 -1260
rect 42680 -1380 42800 -1260
rect 42845 -1380 42965 -1260
rect 43020 -1380 43140 -1260
rect 43185 -1380 43305 -1260
rect 43350 -1380 43470 -1260
rect 43515 -1380 43635 -1260
rect 43690 -1380 43810 -1260
rect 43855 -1380 43975 -1260
rect 44020 -1380 44140 -1260
rect 44185 -1380 44305 -1260
rect 44360 -1380 44480 -1260
rect 44525 -1380 44645 -1260
rect 44690 -1380 44810 -1260
rect 44855 -1380 44975 -1260
rect 45030 -1380 45150 -1260
rect 45195 -1380 45315 -1260
rect 45360 -1380 45480 -1260
rect 45525 -1380 45645 -1260
rect 45700 -1380 45820 -1260
rect 45865 -1380 45985 -1260
rect 46030 -1380 46150 -1260
rect 46195 -1380 46315 -1260
rect 46370 -1380 46490 -1260
rect 46535 -1380 46655 -1260
rect 46700 -1380 46820 -1260
rect 46865 -1380 46985 -1260
rect 47040 -1380 47160 -1260
rect 47205 -1380 47325 -1260
rect 47370 -1380 47490 -1260
rect 47535 -1380 47655 -1260
rect 42175 -1545 42295 -1425
rect 42350 -1545 42470 -1425
rect 42515 -1545 42635 -1425
rect 42680 -1545 42800 -1425
rect 42845 -1545 42965 -1425
rect 43020 -1545 43140 -1425
rect 43185 -1545 43305 -1425
rect 43350 -1545 43470 -1425
rect 43515 -1545 43635 -1425
rect 43690 -1545 43810 -1425
rect 43855 -1545 43975 -1425
rect 44020 -1545 44140 -1425
rect 44185 -1545 44305 -1425
rect 44360 -1545 44480 -1425
rect 44525 -1545 44645 -1425
rect 44690 -1545 44810 -1425
rect 44855 -1545 44975 -1425
rect 45030 -1545 45150 -1425
rect 45195 -1545 45315 -1425
rect 45360 -1545 45480 -1425
rect 45525 -1545 45645 -1425
rect 45700 -1545 45820 -1425
rect 45865 -1545 45985 -1425
rect 46030 -1545 46150 -1425
rect 46195 -1545 46315 -1425
rect 46370 -1545 46490 -1425
rect 46535 -1545 46655 -1425
rect 46700 -1545 46820 -1425
rect 46865 -1545 46985 -1425
rect 47040 -1545 47160 -1425
rect 47205 -1545 47325 -1425
rect 47370 -1545 47490 -1425
rect 47535 -1545 47655 -1425
rect 42175 -1710 42295 -1590
rect 42350 -1710 42470 -1590
rect 42515 -1710 42635 -1590
rect 42680 -1710 42800 -1590
rect 42845 -1710 42965 -1590
rect 43020 -1710 43140 -1590
rect 43185 -1710 43305 -1590
rect 43350 -1710 43470 -1590
rect 43515 -1710 43635 -1590
rect 43690 -1710 43810 -1590
rect 43855 -1710 43975 -1590
rect 44020 -1710 44140 -1590
rect 44185 -1710 44305 -1590
rect 44360 -1710 44480 -1590
rect 44525 -1710 44645 -1590
rect 44690 -1710 44810 -1590
rect 44855 -1710 44975 -1590
rect 45030 -1710 45150 -1590
rect 45195 -1710 45315 -1590
rect 45360 -1710 45480 -1590
rect 45525 -1710 45645 -1590
rect 45700 -1710 45820 -1590
rect 45865 -1710 45985 -1590
rect 46030 -1710 46150 -1590
rect 46195 -1710 46315 -1590
rect 46370 -1710 46490 -1590
rect 46535 -1710 46655 -1590
rect 46700 -1710 46820 -1590
rect 46865 -1710 46985 -1590
rect 47040 -1710 47160 -1590
rect 47205 -1710 47325 -1590
rect 47370 -1710 47490 -1590
rect 47535 -1710 47655 -1590
rect 42175 -1875 42295 -1755
rect 42350 -1875 42470 -1755
rect 42515 -1875 42635 -1755
rect 42680 -1875 42800 -1755
rect 42845 -1875 42965 -1755
rect 43020 -1875 43140 -1755
rect 43185 -1875 43305 -1755
rect 43350 -1875 43470 -1755
rect 43515 -1875 43635 -1755
rect 43690 -1875 43810 -1755
rect 43855 -1875 43975 -1755
rect 44020 -1875 44140 -1755
rect 44185 -1875 44305 -1755
rect 44360 -1875 44480 -1755
rect 44525 -1875 44645 -1755
rect 44690 -1875 44810 -1755
rect 44855 -1875 44975 -1755
rect 45030 -1875 45150 -1755
rect 45195 -1875 45315 -1755
rect 45360 -1875 45480 -1755
rect 45525 -1875 45645 -1755
rect 45700 -1875 45820 -1755
rect 45865 -1875 45985 -1755
rect 46030 -1875 46150 -1755
rect 46195 -1875 46315 -1755
rect 46370 -1875 46490 -1755
rect 46535 -1875 46655 -1755
rect 46700 -1875 46820 -1755
rect 46865 -1875 46985 -1755
rect 47040 -1875 47160 -1755
rect 47205 -1875 47325 -1755
rect 47370 -1875 47490 -1755
rect 47535 -1875 47655 -1755
rect 42175 -2050 42295 -1930
rect 42350 -2050 42470 -1930
rect 42515 -2050 42635 -1930
rect 42680 -2050 42800 -1930
rect 42845 -2050 42965 -1930
rect 43020 -2050 43140 -1930
rect 43185 -2050 43305 -1930
rect 43350 -2050 43470 -1930
rect 43515 -2050 43635 -1930
rect 43690 -2050 43810 -1930
rect 43855 -2050 43975 -1930
rect 44020 -2050 44140 -1930
rect 44185 -2050 44305 -1930
rect 44360 -2050 44480 -1930
rect 44525 -2050 44645 -1930
rect 44690 -2050 44810 -1930
rect 44855 -2050 44975 -1930
rect 45030 -2050 45150 -1930
rect 45195 -2050 45315 -1930
rect 45360 -2050 45480 -1930
rect 45525 -2050 45645 -1930
rect 45700 -2050 45820 -1930
rect 45865 -2050 45985 -1930
rect 46030 -2050 46150 -1930
rect 46195 -2050 46315 -1930
rect 46370 -2050 46490 -1930
rect 46535 -2050 46655 -1930
rect 46700 -2050 46820 -1930
rect 46865 -2050 46985 -1930
rect 47040 -2050 47160 -1930
rect 47205 -2050 47325 -1930
rect 47370 -2050 47490 -1930
rect 47535 -2050 47655 -1930
rect 42175 -2215 42295 -2095
rect 42350 -2215 42470 -2095
rect 42515 -2215 42635 -2095
rect 42680 -2215 42800 -2095
rect 42845 -2215 42965 -2095
rect 43020 -2215 43140 -2095
rect 43185 -2215 43305 -2095
rect 43350 -2215 43470 -2095
rect 43515 -2215 43635 -2095
rect 43690 -2215 43810 -2095
rect 43855 -2215 43975 -2095
rect 44020 -2215 44140 -2095
rect 44185 -2215 44305 -2095
rect 44360 -2215 44480 -2095
rect 44525 -2215 44645 -2095
rect 44690 -2215 44810 -2095
rect 44855 -2215 44975 -2095
rect 45030 -2215 45150 -2095
rect 45195 -2215 45315 -2095
rect 45360 -2215 45480 -2095
rect 45525 -2215 45645 -2095
rect 45700 -2215 45820 -2095
rect 45865 -2215 45985 -2095
rect 46030 -2215 46150 -2095
rect 46195 -2215 46315 -2095
rect 46370 -2215 46490 -2095
rect 46535 -2215 46655 -2095
rect 46700 -2215 46820 -2095
rect 46865 -2215 46985 -2095
rect 47040 -2215 47160 -2095
rect 47205 -2215 47325 -2095
rect 47370 -2215 47490 -2095
rect 47535 -2215 47655 -2095
rect 42175 -2380 42295 -2260
rect 42350 -2380 42470 -2260
rect 42515 -2380 42635 -2260
rect 42680 -2380 42800 -2260
rect 42845 -2380 42965 -2260
rect 43020 -2380 43140 -2260
rect 43185 -2380 43305 -2260
rect 43350 -2380 43470 -2260
rect 43515 -2380 43635 -2260
rect 43690 -2380 43810 -2260
rect 43855 -2380 43975 -2260
rect 44020 -2380 44140 -2260
rect 44185 -2380 44305 -2260
rect 44360 -2380 44480 -2260
rect 44525 -2380 44645 -2260
rect 44690 -2380 44810 -2260
rect 44855 -2380 44975 -2260
rect 45030 -2380 45150 -2260
rect 45195 -2380 45315 -2260
rect 45360 -2380 45480 -2260
rect 45525 -2380 45645 -2260
rect 45700 -2380 45820 -2260
rect 45865 -2380 45985 -2260
rect 46030 -2380 46150 -2260
rect 46195 -2380 46315 -2260
rect 46370 -2380 46490 -2260
rect 46535 -2380 46655 -2260
rect 46700 -2380 46820 -2260
rect 46865 -2380 46985 -2260
rect 47040 -2380 47160 -2260
rect 47205 -2380 47325 -2260
rect 47370 -2380 47490 -2260
rect 47535 -2380 47655 -2260
rect 42175 -2545 42295 -2425
rect 42350 -2545 42470 -2425
rect 42515 -2545 42635 -2425
rect 42680 -2545 42800 -2425
rect 42845 -2545 42965 -2425
rect 43020 -2545 43140 -2425
rect 43185 -2545 43305 -2425
rect 43350 -2545 43470 -2425
rect 43515 -2545 43635 -2425
rect 43690 -2545 43810 -2425
rect 43855 -2545 43975 -2425
rect 44020 -2545 44140 -2425
rect 44185 -2545 44305 -2425
rect 44360 -2545 44480 -2425
rect 44525 -2545 44645 -2425
rect 44690 -2545 44810 -2425
rect 44855 -2545 44975 -2425
rect 45030 -2545 45150 -2425
rect 45195 -2545 45315 -2425
rect 45360 -2545 45480 -2425
rect 45525 -2545 45645 -2425
rect 45700 -2545 45820 -2425
rect 45865 -2545 45985 -2425
rect 46030 -2545 46150 -2425
rect 46195 -2545 46315 -2425
rect 46370 -2545 46490 -2425
rect 46535 -2545 46655 -2425
rect 46700 -2545 46820 -2425
rect 46865 -2545 46985 -2425
rect 47040 -2545 47160 -2425
rect 47205 -2545 47325 -2425
rect 47370 -2545 47490 -2425
rect 47535 -2545 47655 -2425
rect 42175 -2720 42295 -2600
rect 42350 -2720 42470 -2600
rect 42515 -2720 42635 -2600
rect 42680 -2720 42800 -2600
rect 42845 -2720 42965 -2600
rect 43020 -2720 43140 -2600
rect 43185 -2720 43305 -2600
rect 43350 -2720 43470 -2600
rect 43515 -2720 43635 -2600
rect 43690 -2720 43810 -2600
rect 43855 -2720 43975 -2600
rect 44020 -2720 44140 -2600
rect 44185 -2720 44305 -2600
rect 44360 -2720 44480 -2600
rect 44525 -2720 44645 -2600
rect 44690 -2720 44810 -2600
rect 44855 -2720 44975 -2600
rect 45030 -2720 45150 -2600
rect 45195 -2720 45315 -2600
rect 45360 -2720 45480 -2600
rect 45525 -2720 45645 -2600
rect 45700 -2720 45820 -2600
rect 45865 -2720 45985 -2600
rect 46030 -2720 46150 -2600
rect 46195 -2720 46315 -2600
rect 46370 -2720 46490 -2600
rect 46535 -2720 46655 -2600
rect 46700 -2720 46820 -2600
rect 46865 -2720 46985 -2600
rect 47040 -2720 47160 -2600
rect 47205 -2720 47325 -2600
rect 47370 -2720 47490 -2600
rect 47535 -2720 47655 -2600
rect 42175 -2885 42295 -2765
rect 42350 -2885 42470 -2765
rect 42515 -2885 42635 -2765
rect 42680 -2885 42800 -2765
rect 42845 -2885 42965 -2765
rect 43020 -2885 43140 -2765
rect 43185 -2885 43305 -2765
rect 43350 -2885 43470 -2765
rect 43515 -2885 43635 -2765
rect 43690 -2885 43810 -2765
rect 43855 -2885 43975 -2765
rect 44020 -2885 44140 -2765
rect 44185 -2885 44305 -2765
rect 44360 -2885 44480 -2765
rect 44525 -2885 44645 -2765
rect 44690 -2885 44810 -2765
rect 44855 -2885 44975 -2765
rect 45030 -2885 45150 -2765
rect 45195 -2885 45315 -2765
rect 45360 -2885 45480 -2765
rect 45525 -2885 45645 -2765
rect 45700 -2885 45820 -2765
rect 45865 -2885 45985 -2765
rect 46030 -2885 46150 -2765
rect 46195 -2885 46315 -2765
rect 46370 -2885 46490 -2765
rect 46535 -2885 46655 -2765
rect 46700 -2885 46820 -2765
rect 46865 -2885 46985 -2765
rect 47040 -2885 47160 -2765
rect 47205 -2885 47325 -2765
rect 47370 -2885 47490 -2765
rect 47535 -2885 47655 -2765
rect 42175 -3050 42295 -2930
rect 42350 -3050 42470 -2930
rect 42515 -3050 42635 -2930
rect 42680 -3050 42800 -2930
rect 42845 -3050 42965 -2930
rect 43020 -3050 43140 -2930
rect 43185 -3050 43305 -2930
rect 43350 -3050 43470 -2930
rect 43515 -3050 43635 -2930
rect 43690 -3050 43810 -2930
rect 43855 -3050 43975 -2930
rect 44020 -3050 44140 -2930
rect 44185 -3050 44305 -2930
rect 44360 -3050 44480 -2930
rect 44525 -3050 44645 -2930
rect 44690 -3050 44810 -2930
rect 44855 -3050 44975 -2930
rect 45030 -3050 45150 -2930
rect 45195 -3050 45315 -2930
rect 45360 -3050 45480 -2930
rect 45525 -3050 45645 -2930
rect 45700 -3050 45820 -2930
rect 45865 -3050 45985 -2930
rect 46030 -3050 46150 -2930
rect 46195 -3050 46315 -2930
rect 46370 -3050 46490 -2930
rect 46535 -3050 46655 -2930
rect 46700 -3050 46820 -2930
rect 46865 -3050 46985 -2930
rect 47040 -3050 47160 -2930
rect 47205 -3050 47325 -2930
rect 47370 -3050 47490 -2930
rect 47535 -3050 47655 -2930
rect 42175 -3215 42295 -3095
rect 42350 -3215 42470 -3095
rect 42515 -3215 42635 -3095
rect 42680 -3215 42800 -3095
rect 42845 -3215 42965 -3095
rect 43020 -3215 43140 -3095
rect 43185 -3215 43305 -3095
rect 43350 -3215 43470 -3095
rect 43515 -3215 43635 -3095
rect 43690 -3215 43810 -3095
rect 43855 -3215 43975 -3095
rect 44020 -3215 44140 -3095
rect 44185 -3215 44305 -3095
rect 44360 -3215 44480 -3095
rect 44525 -3215 44645 -3095
rect 44690 -3215 44810 -3095
rect 44855 -3215 44975 -3095
rect 45030 -3215 45150 -3095
rect 45195 -3215 45315 -3095
rect 45360 -3215 45480 -3095
rect 45525 -3215 45645 -3095
rect 45700 -3215 45820 -3095
rect 45865 -3215 45985 -3095
rect 46030 -3215 46150 -3095
rect 46195 -3215 46315 -3095
rect 46370 -3215 46490 -3095
rect 46535 -3215 46655 -3095
rect 46700 -3215 46820 -3095
rect 46865 -3215 46985 -3095
rect 47040 -3215 47160 -3095
rect 47205 -3215 47325 -3095
rect 47370 -3215 47490 -3095
rect 47535 -3215 47655 -3095
rect 42175 -3390 42295 -3270
rect 42350 -3390 42470 -3270
rect 42515 -3390 42635 -3270
rect 42680 -3390 42800 -3270
rect 42845 -3390 42965 -3270
rect 43020 -3390 43140 -3270
rect 43185 -3390 43305 -3270
rect 43350 -3390 43470 -3270
rect 43515 -3390 43635 -3270
rect 43690 -3390 43810 -3270
rect 43855 -3390 43975 -3270
rect 44020 -3390 44140 -3270
rect 44185 -3390 44305 -3270
rect 44360 -3390 44480 -3270
rect 44525 -3390 44645 -3270
rect 44690 -3390 44810 -3270
rect 44855 -3390 44975 -3270
rect 45030 -3390 45150 -3270
rect 45195 -3390 45315 -3270
rect 45360 -3390 45480 -3270
rect 45525 -3390 45645 -3270
rect 45700 -3390 45820 -3270
rect 45865 -3390 45985 -3270
rect 46030 -3390 46150 -3270
rect 46195 -3390 46315 -3270
rect 46370 -3390 46490 -3270
rect 46535 -3390 46655 -3270
rect 46700 -3390 46820 -3270
rect 46865 -3390 46985 -3270
rect 47040 -3390 47160 -3270
rect 47205 -3390 47325 -3270
rect 47370 -3390 47490 -3270
rect 47535 -3390 47655 -3270
rect 42175 -3555 42295 -3435
rect 42350 -3555 42470 -3435
rect 42515 -3555 42635 -3435
rect 42680 -3555 42800 -3435
rect 42845 -3555 42965 -3435
rect 43020 -3555 43140 -3435
rect 43185 -3555 43305 -3435
rect 43350 -3555 43470 -3435
rect 43515 -3555 43635 -3435
rect 43690 -3555 43810 -3435
rect 43855 -3555 43975 -3435
rect 44020 -3555 44140 -3435
rect 44185 -3555 44305 -3435
rect 44360 -3555 44480 -3435
rect 44525 -3555 44645 -3435
rect 44690 -3555 44810 -3435
rect 44855 -3555 44975 -3435
rect 45030 -3555 45150 -3435
rect 45195 -3555 45315 -3435
rect 45360 -3555 45480 -3435
rect 45525 -3555 45645 -3435
rect 45700 -3555 45820 -3435
rect 45865 -3555 45985 -3435
rect 46030 -3555 46150 -3435
rect 46195 -3555 46315 -3435
rect 46370 -3555 46490 -3435
rect 46535 -3555 46655 -3435
rect 46700 -3555 46820 -3435
rect 46865 -3555 46985 -3435
rect 47040 -3555 47160 -3435
rect 47205 -3555 47325 -3435
rect 47370 -3555 47490 -3435
rect 47535 -3555 47655 -3435
rect 42175 -3720 42295 -3600
rect 42350 -3720 42470 -3600
rect 42515 -3720 42635 -3600
rect 42680 -3720 42800 -3600
rect 42845 -3720 42965 -3600
rect 43020 -3720 43140 -3600
rect 43185 -3720 43305 -3600
rect 43350 -3720 43470 -3600
rect 43515 -3720 43635 -3600
rect 43690 -3720 43810 -3600
rect 43855 -3720 43975 -3600
rect 44020 -3720 44140 -3600
rect 44185 -3720 44305 -3600
rect 44360 -3720 44480 -3600
rect 44525 -3720 44645 -3600
rect 44690 -3720 44810 -3600
rect 44855 -3720 44975 -3600
rect 45030 -3720 45150 -3600
rect 45195 -3720 45315 -3600
rect 45360 -3720 45480 -3600
rect 45525 -3720 45645 -3600
rect 45700 -3720 45820 -3600
rect 45865 -3720 45985 -3600
rect 46030 -3720 46150 -3600
rect 46195 -3720 46315 -3600
rect 46370 -3720 46490 -3600
rect 46535 -3720 46655 -3600
rect 46700 -3720 46820 -3600
rect 46865 -3720 46985 -3600
rect 47040 -3720 47160 -3600
rect 47205 -3720 47325 -3600
rect 47370 -3720 47490 -3600
rect 47535 -3720 47655 -3600
rect 42175 -3885 42295 -3765
rect 42350 -3885 42470 -3765
rect 42515 -3885 42635 -3765
rect 42680 -3885 42800 -3765
rect 42845 -3885 42965 -3765
rect 43020 -3885 43140 -3765
rect 43185 -3885 43305 -3765
rect 43350 -3885 43470 -3765
rect 43515 -3885 43635 -3765
rect 43690 -3885 43810 -3765
rect 43855 -3885 43975 -3765
rect 44020 -3885 44140 -3765
rect 44185 -3885 44305 -3765
rect 44360 -3885 44480 -3765
rect 44525 -3885 44645 -3765
rect 44690 -3885 44810 -3765
rect 44855 -3885 44975 -3765
rect 45030 -3885 45150 -3765
rect 45195 -3885 45315 -3765
rect 45360 -3885 45480 -3765
rect 45525 -3885 45645 -3765
rect 45700 -3885 45820 -3765
rect 45865 -3885 45985 -3765
rect 46030 -3885 46150 -3765
rect 46195 -3885 46315 -3765
rect 46370 -3885 46490 -3765
rect 46535 -3885 46655 -3765
rect 46700 -3885 46820 -3765
rect 46865 -3885 46985 -3765
rect 47040 -3885 47160 -3765
rect 47205 -3885 47325 -3765
rect 47370 -3885 47490 -3765
rect 47535 -3885 47655 -3765
rect 42175 -4060 42295 -3940
rect 42350 -4060 42470 -3940
rect 42515 -4060 42635 -3940
rect 42680 -4060 42800 -3940
rect 42845 -4060 42965 -3940
rect 43020 -4060 43140 -3940
rect 43185 -4060 43305 -3940
rect 43350 -4060 43470 -3940
rect 43515 -4060 43635 -3940
rect 43690 -4060 43810 -3940
rect 43855 -4060 43975 -3940
rect 44020 -4060 44140 -3940
rect 44185 -4060 44305 -3940
rect 44360 -4060 44480 -3940
rect 44525 -4060 44645 -3940
rect 44690 -4060 44810 -3940
rect 44855 -4060 44975 -3940
rect 45030 -4060 45150 -3940
rect 45195 -4060 45315 -3940
rect 45360 -4060 45480 -3940
rect 45525 -4060 45645 -3940
rect 45700 -4060 45820 -3940
rect 45865 -4060 45985 -3940
rect 46030 -4060 46150 -3940
rect 46195 -4060 46315 -3940
rect 46370 -4060 46490 -3940
rect 46535 -4060 46655 -3940
rect 46700 -4060 46820 -3940
rect 46865 -4060 46985 -3940
rect 47040 -4060 47160 -3940
rect 47205 -4060 47325 -3940
rect 47370 -4060 47490 -3940
rect 47535 -4060 47655 -3940
rect 47865 1300 47985 1420
rect 48040 1300 48160 1420
rect 48205 1300 48325 1420
rect 48370 1300 48490 1420
rect 48535 1300 48655 1420
rect 48710 1300 48830 1420
rect 48875 1300 48995 1420
rect 49040 1300 49160 1420
rect 49205 1300 49325 1420
rect 49380 1300 49500 1420
rect 49545 1300 49665 1420
rect 49710 1300 49830 1420
rect 49875 1300 49995 1420
rect 50050 1300 50170 1420
rect 50215 1300 50335 1420
rect 50380 1300 50500 1420
rect 50545 1300 50665 1420
rect 50720 1300 50840 1420
rect 50885 1300 51005 1420
rect 51050 1300 51170 1420
rect 51215 1300 51335 1420
rect 51390 1300 51510 1420
rect 51555 1300 51675 1420
rect 51720 1300 51840 1420
rect 51885 1300 52005 1420
rect 52060 1300 52180 1420
rect 52225 1300 52345 1420
rect 52390 1300 52510 1420
rect 52555 1300 52675 1420
rect 52730 1300 52850 1420
rect 52895 1300 53015 1420
rect 53060 1300 53180 1420
rect 53225 1300 53345 1420
rect 47865 1135 47985 1255
rect 48040 1135 48160 1255
rect 48205 1135 48325 1255
rect 48370 1135 48490 1255
rect 48535 1135 48655 1255
rect 48710 1135 48830 1255
rect 48875 1135 48995 1255
rect 49040 1135 49160 1255
rect 49205 1135 49325 1255
rect 49380 1135 49500 1255
rect 49545 1135 49665 1255
rect 49710 1135 49830 1255
rect 49875 1135 49995 1255
rect 50050 1135 50170 1255
rect 50215 1135 50335 1255
rect 50380 1135 50500 1255
rect 50545 1135 50665 1255
rect 50720 1135 50840 1255
rect 50885 1135 51005 1255
rect 51050 1135 51170 1255
rect 51215 1135 51335 1255
rect 51390 1135 51510 1255
rect 51555 1135 51675 1255
rect 51720 1135 51840 1255
rect 51885 1135 52005 1255
rect 52060 1135 52180 1255
rect 52225 1135 52345 1255
rect 52390 1135 52510 1255
rect 52555 1135 52675 1255
rect 52730 1135 52850 1255
rect 52895 1135 53015 1255
rect 53060 1135 53180 1255
rect 53225 1135 53345 1255
rect 47865 970 47985 1090
rect 48040 970 48160 1090
rect 48205 970 48325 1090
rect 48370 970 48490 1090
rect 48535 970 48655 1090
rect 48710 970 48830 1090
rect 48875 970 48995 1090
rect 49040 970 49160 1090
rect 49205 970 49325 1090
rect 49380 970 49500 1090
rect 49545 970 49665 1090
rect 49710 970 49830 1090
rect 49875 970 49995 1090
rect 50050 970 50170 1090
rect 50215 970 50335 1090
rect 50380 970 50500 1090
rect 50545 970 50665 1090
rect 50720 970 50840 1090
rect 50885 970 51005 1090
rect 51050 970 51170 1090
rect 51215 970 51335 1090
rect 51390 970 51510 1090
rect 51555 970 51675 1090
rect 51720 970 51840 1090
rect 51885 970 52005 1090
rect 52060 970 52180 1090
rect 52225 970 52345 1090
rect 52390 970 52510 1090
rect 52555 970 52675 1090
rect 52730 970 52850 1090
rect 52895 970 53015 1090
rect 53060 970 53180 1090
rect 53225 970 53345 1090
rect 47865 805 47985 925
rect 48040 805 48160 925
rect 48205 805 48325 925
rect 48370 805 48490 925
rect 48535 805 48655 925
rect 48710 805 48830 925
rect 48875 805 48995 925
rect 49040 805 49160 925
rect 49205 805 49325 925
rect 49380 805 49500 925
rect 49545 805 49665 925
rect 49710 805 49830 925
rect 49875 805 49995 925
rect 50050 805 50170 925
rect 50215 805 50335 925
rect 50380 805 50500 925
rect 50545 805 50665 925
rect 50720 805 50840 925
rect 50885 805 51005 925
rect 51050 805 51170 925
rect 51215 805 51335 925
rect 51390 805 51510 925
rect 51555 805 51675 925
rect 51720 805 51840 925
rect 51885 805 52005 925
rect 52060 805 52180 925
rect 52225 805 52345 925
rect 52390 805 52510 925
rect 52555 805 52675 925
rect 52730 805 52850 925
rect 52895 805 53015 925
rect 53060 805 53180 925
rect 53225 805 53345 925
rect 47865 630 47985 750
rect 48040 630 48160 750
rect 48205 630 48325 750
rect 48370 630 48490 750
rect 48535 630 48655 750
rect 48710 630 48830 750
rect 48875 630 48995 750
rect 49040 630 49160 750
rect 49205 630 49325 750
rect 49380 630 49500 750
rect 49545 630 49665 750
rect 49710 630 49830 750
rect 49875 630 49995 750
rect 50050 630 50170 750
rect 50215 630 50335 750
rect 50380 630 50500 750
rect 50545 630 50665 750
rect 50720 630 50840 750
rect 50885 630 51005 750
rect 51050 630 51170 750
rect 51215 630 51335 750
rect 51390 630 51510 750
rect 51555 630 51675 750
rect 51720 630 51840 750
rect 51885 630 52005 750
rect 52060 630 52180 750
rect 52225 630 52345 750
rect 52390 630 52510 750
rect 52555 630 52675 750
rect 52730 630 52850 750
rect 52895 630 53015 750
rect 53060 630 53180 750
rect 53225 630 53345 750
rect 47865 465 47985 585
rect 48040 465 48160 585
rect 48205 465 48325 585
rect 48370 465 48490 585
rect 48535 465 48655 585
rect 48710 465 48830 585
rect 48875 465 48995 585
rect 49040 465 49160 585
rect 49205 465 49325 585
rect 49380 465 49500 585
rect 49545 465 49665 585
rect 49710 465 49830 585
rect 49875 465 49995 585
rect 50050 465 50170 585
rect 50215 465 50335 585
rect 50380 465 50500 585
rect 50545 465 50665 585
rect 50720 465 50840 585
rect 50885 465 51005 585
rect 51050 465 51170 585
rect 51215 465 51335 585
rect 51390 465 51510 585
rect 51555 465 51675 585
rect 51720 465 51840 585
rect 51885 465 52005 585
rect 52060 465 52180 585
rect 52225 465 52345 585
rect 52390 465 52510 585
rect 52555 465 52675 585
rect 52730 465 52850 585
rect 52895 465 53015 585
rect 53060 465 53180 585
rect 53225 465 53345 585
rect 47865 300 47985 420
rect 48040 300 48160 420
rect 48205 300 48325 420
rect 48370 300 48490 420
rect 48535 300 48655 420
rect 48710 300 48830 420
rect 48875 300 48995 420
rect 49040 300 49160 420
rect 49205 300 49325 420
rect 49380 300 49500 420
rect 49545 300 49665 420
rect 49710 300 49830 420
rect 49875 300 49995 420
rect 50050 300 50170 420
rect 50215 300 50335 420
rect 50380 300 50500 420
rect 50545 300 50665 420
rect 50720 300 50840 420
rect 50885 300 51005 420
rect 51050 300 51170 420
rect 51215 300 51335 420
rect 51390 300 51510 420
rect 51555 300 51675 420
rect 51720 300 51840 420
rect 51885 300 52005 420
rect 52060 300 52180 420
rect 52225 300 52345 420
rect 52390 300 52510 420
rect 52555 300 52675 420
rect 52730 300 52850 420
rect 52895 300 53015 420
rect 53060 300 53180 420
rect 53225 300 53345 420
rect 47865 135 47985 255
rect 48040 135 48160 255
rect 48205 135 48325 255
rect 48370 135 48490 255
rect 48535 135 48655 255
rect 48710 135 48830 255
rect 48875 135 48995 255
rect 49040 135 49160 255
rect 49205 135 49325 255
rect 49380 135 49500 255
rect 49545 135 49665 255
rect 49710 135 49830 255
rect 49875 135 49995 255
rect 50050 135 50170 255
rect 50215 135 50335 255
rect 50380 135 50500 255
rect 50545 135 50665 255
rect 50720 135 50840 255
rect 50885 135 51005 255
rect 51050 135 51170 255
rect 51215 135 51335 255
rect 51390 135 51510 255
rect 51555 135 51675 255
rect 51720 135 51840 255
rect 51885 135 52005 255
rect 52060 135 52180 255
rect 52225 135 52345 255
rect 52390 135 52510 255
rect 52555 135 52675 255
rect 52730 135 52850 255
rect 52895 135 53015 255
rect 53060 135 53180 255
rect 53225 135 53345 255
rect 47865 -40 47985 80
rect 48040 -40 48160 80
rect 48205 -40 48325 80
rect 48370 -40 48490 80
rect 48535 -40 48655 80
rect 48710 -40 48830 80
rect 48875 -40 48995 80
rect 49040 -40 49160 80
rect 49205 -40 49325 80
rect 49380 -40 49500 80
rect 49545 -40 49665 80
rect 49710 -40 49830 80
rect 49875 -40 49995 80
rect 50050 -40 50170 80
rect 50215 -40 50335 80
rect 50380 -40 50500 80
rect 50545 -40 50665 80
rect 50720 -40 50840 80
rect 50885 -40 51005 80
rect 51050 -40 51170 80
rect 51215 -40 51335 80
rect 51390 -40 51510 80
rect 51555 -40 51675 80
rect 51720 -40 51840 80
rect 51885 -40 52005 80
rect 52060 -40 52180 80
rect 52225 -40 52345 80
rect 52390 -40 52510 80
rect 52555 -40 52675 80
rect 52730 -40 52850 80
rect 52895 -40 53015 80
rect 53060 -40 53180 80
rect 53225 -40 53345 80
rect 47865 -205 47985 -85
rect 48040 -205 48160 -85
rect 48205 -205 48325 -85
rect 48370 -205 48490 -85
rect 48535 -205 48655 -85
rect 48710 -205 48830 -85
rect 48875 -205 48995 -85
rect 49040 -205 49160 -85
rect 49205 -205 49325 -85
rect 49380 -205 49500 -85
rect 49545 -205 49665 -85
rect 49710 -205 49830 -85
rect 49875 -205 49995 -85
rect 50050 -205 50170 -85
rect 50215 -205 50335 -85
rect 50380 -205 50500 -85
rect 50545 -205 50665 -85
rect 50720 -205 50840 -85
rect 50885 -205 51005 -85
rect 51050 -205 51170 -85
rect 51215 -205 51335 -85
rect 51390 -205 51510 -85
rect 51555 -205 51675 -85
rect 51720 -205 51840 -85
rect 51885 -205 52005 -85
rect 52060 -205 52180 -85
rect 52225 -205 52345 -85
rect 52390 -205 52510 -85
rect 52555 -205 52675 -85
rect 52730 -205 52850 -85
rect 52895 -205 53015 -85
rect 53060 -205 53180 -85
rect 53225 -205 53345 -85
rect 47865 -370 47985 -250
rect 48040 -370 48160 -250
rect 48205 -370 48325 -250
rect 48370 -370 48490 -250
rect 48535 -370 48655 -250
rect 48710 -370 48830 -250
rect 48875 -370 48995 -250
rect 49040 -370 49160 -250
rect 49205 -370 49325 -250
rect 49380 -370 49500 -250
rect 49545 -370 49665 -250
rect 49710 -370 49830 -250
rect 49875 -370 49995 -250
rect 50050 -370 50170 -250
rect 50215 -370 50335 -250
rect 50380 -370 50500 -250
rect 50545 -370 50665 -250
rect 50720 -370 50840 -250
rect 50885 -370 51005 -250
rect 51050 -370 51170 -250
rect 51215 -370 51335 -250
rect 51390 -370 51510 -250
rect 51555 -370 51675 -250
rect 51720 -370 51840 -250
rect 51885 -370 52005 -250
rect 52060 -370 52180 -250
rect 52225 -370 52345 -250
rect 52390 -370 52510 -250
rect 52555 -370 52675 -250
rect 52730 -370 52850 -250
rect 52895 -370 53015 -250
rect 53060 -370 53180 -250
rect 53225 -370 53345 -250
rect 47865 -535 47985 -415
rect 48040 -535 48160 -415
rect 48205 -535 48325 -415
rect 48370 -535 48490 -415
rect 48535 -535 48655 -415
rect 48710 -535 48830 -415
rect 48875 -535 48995 -415
rect 49040 -535 49160 -415
rect 49205 -535 49325 -415
rect 49380 -535 49500 -415
rect 49545 -535 49665 -415
rect 49710 -535 49830 -415
rect 49875 -535 49995 -415
rect 50050 -535 50170 -415
rect 50215 -535 50335 -415
rect 50380 -535 50500 -415
rect 50545 -535 50665 -415
rect 50720 -535 50840 -415
rect 50885 -535 51005 -415
rect 51050 -535 51170 -415
rect 51215 -535 51335 -415
rect 51390 -535 51510 -415
rect 51555 -535 51675 -415
rect 51720 -535 51840 -415
rect 51885 -535 52005 -415
rect 52060 -535 52180 -415
rect 52225 -535 52345 -415
rect 52390 -535 52510 -415
rect 52555 -535 52675 -415
rect 52730 -535 52850 -415
rect 52895 -535 53015 -415
rect 53060 -535 53180 -415
rect 53225 -535 53345 -415
rect 47865 -710 47985 -590
rect 48040 -710 48160 -590
rect 48205 -710 48325 -590
rect 48370 -710 48490 -590
rect 48535 -710 48655 -590
rect 48710 -710 48830 -590
rect 48875 -710 48995 -590
rect 49040 -710 49160 -590
rect 49205 -710 49325 -590
rect 49380 -710 49500 -590
rect 49545 -710 49665 -590
rect 49710 -710 49830 -590
rect 49875 -710 49995 -590
rect 50050 -710 50170 -590
rect 50215 -710 50335 -590
rect 50380 -710 50500 -590
rect 50545 -710 50665 -590
rect 50720 -710 50840 -590
rect 50885 -710 51005 -590
rect 51050 -710 51170 -590
rect 51215 -710 51335 -590
rect 51390 -710 51510 -590
rect 51555 -710 51675 -590
rect 51720 -710 51840 -590
rect 51885 -710 52005 -590
rect 52060 -710 52180 -590
rect 52225 -710 52345 -590
rect 52390 -710 52510 -590
rect 52555 -710 52675 -590
rect 52730 -710 52850 -590
rect 52895 -710 53015 -590
rect 53060 -710 53180 -590
rect 53225 -710 53345 -590
rect 47865 -875 47985 -755
rect 48040 -875 48160 -755
rect 48205 -875 48325 -755
rect 48370 -875 48490 -755
rect 48535 -875 48655 -755
rect 48710 -875 48830 -755
rect 48875 -875 48995 -755
rect 49040 -875 49160 -755
rect 49205 -875 49325 -755
rect 49380 -875 49500 -755
rect 49545 -875 49665 -755
rect 49710 -875 49830 -755
rect 49875 -875 49995 -755
rect 50050 -875 50170 -755
rect 50215 -875 50335 -755
rect 50380 -875 50500 -755
rect 50545 -875 50665 -755
rect 50720 -875 50840 -755
rect 50885 -875 51005 -755
rect 51050 -875 51170 -755
rect 51215 -875 51335 -755
rect 51390 -875 51510 -755
rect 51555 -875 51675 -755
rect 51720 -875 51840 -755
rect 51885 -875 52005 -755
rect 52060 -875 52180 -755
rect 52225 -875 52345 -755
rect 52390 -875 52510 -755
rect 52555 -875 52675 -755
rect 52730 -875 52850 -755
rect 52895 -875 53015 -755
rect 53060 -875 53180 -755
rect 53225 -875 53345 -755
rect 47865 -1040 47985 -920
rect 48040 -1040 48160 -920
rect 48205 -1040 48325 -920
rect 48370 -1040 48490 -920
rect 48535 -1040 48655 -920
rect 48710 -1040 48830 -920
rect 48875 -1040 48995 -920
rect 49040 -1040 49160 -920
rect 49205 -1040 49325 -920
rect 49380 -1040 49500 -920
rect 49545 -1040 49665 -920
rect 49710 -1040 49830 -920
rect 49875 -1040 49995 -920
rect 50050 -1040 50170 -920
rect 50215 -1040 50335 -920
rect 50380 -1040 50500 -920
rect 50545 -1040 50665 -920
rect 50720 -1040 50840 -920
rect 50885 -1040 51005 -920
rect 51050 -1040 51170 -920
rect 51215 -1040 51335 -920
rect 51390 -1040 51510 -920
rect 51555 -1040 51675 -920
rect 51720 -1040 51840 -920
rect 51885 -1040 52005 -920
rect 52060 -1040 52180 -920
rect 52225 -1040 52345 -920
rect 52390 -1040 52510 -920
rect 52555 -1040 52675 -920
rect 52730 -1040 52850 -920
rect 52895 -1040 53015 -920
rect 53060 -1040 53180 -920
rect 53225 -1040 53345 -920
rect 47865 -1205 47985 -1085
rect 48040 -1205 48160 -1085
rect 48205 -1205 48325 -1085
rect 48370 -1205 48490 -1085
rect 48535 -1205 48655 -1085
rect 48710 -1205 48830 -1085
rect 48875 -1205 48995 -1085
rect 49040 -1205 49160 -1085
rect 49205 -1205 49325 -1085
rect 49380 -1205 49500 -1085
rect 49545 -1205 49665 -1085
rect 49710 -1205 49830 -1085
rect 49875 -1205 49995 -1085
rect 50050 -1205 50170 -1085
rect 50215 -1205 50335 -1085
rect 50380 -1205 50500 -1085
rect 50545 -1205 50665 -1085
rect 50720 -1205 50840 -1085
rect 50885 -1205 51005 -1085
rect 51050 -1205 51170 -1085
rect 51215 -1205 51335 -1085
rect 51390 -1205 51510 -1085
rect 51555 -1205 51675 -1085
rect 51720 -1205 51840 -1085
rect 51885 -1205 52005 -1085
rect 52060 -1205 52180 -1085
rect 52225 -1205 52345 -1085
rect 52390 -1205 52510 -1085
rect 52555 -1205 52675 -1085
rect 52730 -1205 52850 -1085
rect 52895 -1205 53015 -1085
rect 53060 -1205 53180 -1085
rect 53225 -1205 53345 -1085
rect 47865 -1380 47985 -1260
rect 48040 -1380 48160 -1260
rect 48205 -1380 48325 -1260
rect 48370 -1380 48490 -1260
rect 48535 -1380 48655 -1260
rect 48710 -1380 48830 -1260
rect 48875 -1380 48995 -1260
rect 49040 -1380 49160 -1260
rect 49205 -1380 49325 -1260
rect 49380 -1380 49500 -1260
rect 49545 -1380 49665 -1260
rect 49710 -1380 49830 -1260
rect 49875 -1380 49995 -1260
rect 50050 -1380 50170 -1260
rect 50215 -1380 50335 -1260
rect 50380 -1380 50500 -1260
rect 50545 -1380 50665 -1260
rect 50720 -1380 50840 -1260
rect 50885 -1380 51005 -1260
rect 51050 -1380 51170 -1260
rect 51215 -1380 51335 -1260
rect 51390 -1380 51510 -1260
rect 51555 -1380 51675 -1260
rect 51720 -1380 51840 -1260
rect 51885 -1380 52005 -1260
rect 52060 -1380 52180 -1260
rect 52225 -1380 52345 -1260
rect 52390 -1380 52510 -1260
rect 52555 -1380 52675 -1260
rect 52730 -1380 52850 -1260
rect 52895 -1380 53015 -1260
rect 53060 -1380 53180 -1260
rect 53225 -1380 53345 -1260
rect 47865 -1545 47985 -1425
rect 48040 -1545 48160 -1425
rect 48205 -1545 48325 -1425
rect 48370 -1545 48490 -1425
rect 48535 -1545 48655 -1425
rect 48710 -1545 48830 -1425
rect 48875 -1545 48995 -1425
rect 49040 -1545 49160 -1425
rect 49205 -1545 49325 -1425
rect 49380 -1545 49500 -1425
rect 49545 -1545 49665 -1425
rect 49710 -1545 49830 -1425
rect 49875 -1545 49995 -1425
rect 50050 -1545 50170 -1425
rect 50215 -1545 50335 -1425
rect 50380 -1545 50500 -1425
rect 50545 -1545 50665 -1425
rect 50720 -1545 50840 -1425
rect 50885 -1545 51005 -1425
rect 51050 -1545 51170 -1425
rect 51215 -1545 51335 -1425
rect 51390 -1545 51510 -1425
rect 51555 -1545 51675 -1425
rect 51720 -1545 51840 -1425
rect 51885 -1545 52005 -1425
rect 52060 -1545 52180 -1425
rect 52225 -1545 52345 -1425
rect 52390 -1545 52510 -1425
rect 52555 -1545 52675 -1425
rect 52730 -1545 52850 -1425
rect 52895 -1545 53015 -1425
rect 53060 -1545 53180 -1425
rect 53225 -1545 53345 -1425
rect 47865 -1710 47985 -1590
rect 48040 -1710 48160 -1590
rect 48205 -1710 48325 -1590
rect 48370 -1710 48490 -1590
rect 48535 -1710 48655 -1590
rect 48710 -1710 48830 -1590
rect 48875 -1710 48995 -1590
rect 49040 -1710 49160 -1590
rect 49205 -1710 49325 -1590
rect 49380 -1710 49500 -1590
rect 49545 -1710 49665 -1590
rect 49710 -1710 49830 -1590
rect 49875 -1710 49995 -1590
rect 50050 -1710 50170 -1590
rect 50215 -1710 50335 -1590
rect 50380 -1710 50500 -1590
rect 50545 -1710 50665 -1590
rect 50720 -1710 50840 -1590
rect 50885 -1710 51005 -1590
rect 51050 -1710 51170 -1590
rect 51215 -1710 51335 -1590
rect 51390 -1710 51510 -1590
rect 51555 -1710 51675 -1590
rect 51720 -1710 51840 -1590
rect 51885 -1710 52005 -1590
rect 52060 -1710 52180 -1590
rect 52225 -1710 52345 -1590
rect 52390 -1710 52510 -1590
rect 52555 -1710 52675 -1590
rect 52730 -1710 52850 -1590
rect 52895 -1710 53015 -1590
rect 53060 -1710 53180 -1590
rect 53225 -1710 53345 -1590
rect 47865 -1875 47985 -1755
rect 48040 -1875 48160 -1755
rect 48205 -1875 48325 -1755
rect 48370 -1875 48490 -1755
rect 48535 -1875 48655 -1755
rect 48710 -1875 48830 -1755
rect 48875 -1875 48995 -1755
rect 49040 -1875 49160 -1755
rect 49205 -1875 49325 -1755
rect 49380 -1875 49500 -1755
rect 49545 -1875 49665 -1755
rect 49710 -1875 49830 -1755
rect 49875 -1875 49995 -1755
rect 50050 -1875 50170 -1755
rect 50215 -1875 50335 -1755
rect 50380 -1875 50500 -1755
rect 50545 -1875 50665 -1755
rect 50720 -1875 50840 -1755
rect 50885 -1875 51005 -1755
rect 51050 -1875 51170 -1755
rect 51215 -1875 51335 -1755
rect 51390 -1875 51510 -1755
rect 51555 -1875 51675 -1755
rect 51720 -1875 51840 -1755
rect 51885 -1875 52005 -1755
rect 52060 -1875 52180 -1755
rect 52225 -1875 52345 -1755
rect 52390 -1875 52510 -1755
rect 52555 -1875 52675 -1755
rect 52730 -1875 52850 -1755
rect 52895 -1875 53015 -1755
rect 53060 -1875 53180 -1755
rect 53225 -1875 53345 -1755
rect 47865 -2050 47985 -1930
rect 48040 -2050 48160 -1930
rect 48205 -2050 48325 -1930
rect 48370 -2050 48490 -1930
rect 48535 -2050 48655 -1930
rect 48710 -2050 48830 -1930
rect 48875 -2050 48995 -1930
rect 49040 -2050 49160 -1930
rect 49205 -2050 49325 -1930
rect 49380 -2050 49500 -1930
rect 49545 -2050 49665 -1930
rect 49710 -2050 49830 -1930
rect 49875 -2050 49995 -1930
rect 50050 -2050 50170 -1930
rect 50215 -2050 50335 -1930
rect 50380 -2050 50500 -1930
rect 50545 -2050 50665 -1930
rect 50720 -2050 50840 -1930
rect 50885 -2050 51005 -1930
rect 51050 -2050 51170 -1930
rect 51215 -2050 51335 -1930
rect 51390 -2050 51510 -1930
rect 51555 -2050 51675 -1930
rect 51720 -2050 51840 -1930
rect 51885 -2050 52005 -1930
rect 52060 -2050 52180 -1930
rect 52225 -2050 52345 -1930
rect 52390 -2050 52510 -1930
rect 52555 -2050 52675 -1930
rect 52730 -2050 52850 -1930
rect 52895 -2050 53015 -1930
rect 53060 -2050 53180 -1930
rect 53225 -2050 53345 -1930
rect 47865 -2215 47985 -2095
rect 48040 -2215 48160 -2095
rect 48205 -2215 48325 -2095
rect 48370 -2215 48490 -2095
rect 48535 -2215 48655 -2095
rect 48710 -2215 48830 -2095
rect 48875 -2215 48995 -2095
rect 49040 -2215 49160 -2095
rect 49205 -2215 49325 -2095
rect 49380 -2215 49500 -2095
rect 49545 -2215 49665 -2095
rect 49710 -2215 49830 -2095
rect 49875 -2215 49995 -2095
rect 50050 -2215 50170 -2095
rect 50215 -2215 50335 -2095
rect 50380 -2215 50500 -2095
rect 50545 -2215 50665 -2095
rect 50720 -2215 50840 -2095
rect 50885 -2215 51005 -2095
rect 51050 -2215 51170 -2095
rect 51215 -2215 51335 -2095
rect 51390 -2215 51510 -2095
rect 51555 -2215 51675 -2095
rect 51720 -2215 51840 -2095
rect 51885 -2215 52005 -2095
rect 52060 -2215 52180 -2095
rect 52225 -2215 52345 -2095
rect 52390 -2215 52510 -2095
rect 52555 -2215 52675 -2095
rect 52730 -2215 52850 -2095
rect 52895 -2215 53015 -2095
rect 53060 -2215 53180 -2095
rect 53225 -2215 53345 -2095
rect 47865 -2380 47985 -2260
rect 48040 -2380 48160 -2260
rect 48205 -2380 48325 -2260
rect 48370 -2380 48490 -2260
rect 48535 -2380 48655 -2260
rect 48710 -2380 48830 -2260
rect 48875 -2380 48995 -2260
rect 49040 -2380 49160 -2260
rect 49205 -2380 49325 -2260
rect 49380 -2380 49500 -2260
rect 49545 -2380 49665 -2260
rect 49710 -2380 49830 -2260
rect 49875 -2380 49995 -2260
rect 50050 -2380 50170 -2260
rect 50215 -2380 50335 -2260
rect 50380 -2380 50500 -2260
rect 50545 -2380 50665 -2260
rect 50720 -2380 50840 -2260
rect 50885 -2380 51005 -2260
rect 51050 -2380 51170 -2260
rect 51215 -2380 51335 -2260
rect 51390 -2380 51510 -2260
rect 51555 -2380 51675 -2260
rect 51720 -2380 51840 -2260
rect 51885 -2380 52005 -2260
rect 52060 -2380 52180 -2260
rect 52225 -2380 52345 -2260
rect 52390 -2380 52510 -2260
rect 52555 -2380 52675 -2260
rect 52730 -2380 52850 -2260
rect 52895 -2380 53015 -2260
rect 53060 -2380 53180 -2260
rect 53225 -2380 53345 -2260
rect 47865 -2545 47985 -2425
rect 48040 -2545 48160 -2425
rect 48205 -2545 48325 -2425
rect 48370 -2545 48490 -2425
rect 48535 -2545 48655 -2425
rect 48710 -2545 48830 -2425
rect 48875 -2545 48995 -2425
rect 49040 -2545 49160 -2425
rect 49205 -2545 49325 -2425
rect 49380 -2545 49500 -2425
rect 49545 -2545 49665 -2425
rect 49710 -2545 49830 -2425
rect 49875 -2545 49995 -2425
rect 50050 -2545 50170 -2425
rect 50215 -2545 50335 -2425
rect 50380 -2545 50500 -2425
rect 50545 -2545 50665 -2425
rect 50720 -2545 50840 -2425
rect 50885 -2545 51005 -2425
rect 51050 -2545 51170 -2425
rect 51215 -2545 51335 -2425
rect 51390 -2545 51510 -2425
rect 51555 -2545 51675 -2425
rect 51720 -2545 51840 -2425
rect 51885 -2545 52005 -2425
rect 52060 -2545 52180 -2425
rect 52225 -2545 52345 -2425
rect 52390 -2545 52510 -2425
rect 52555 -2545 52675 -2425
rect 52730 -2545 52850 -2425
rect 52895 -2545 53015 -2425
rect 53060 -2545 53180 -2425
rect 53225 -2545 53345 -2425
rect 47865 -2720 47985 -2600
rect 48040 -2720 48160 -2600
rect 48205 -2720 48325 -2600
rect 48370 -2720 48490 -2600
rect 48535 -2720 48655 -2600
rect 48710 -2720 48830 -2600
rect 48875 -2720 48995 -2600
rect 49040 -2720 49160 -2600
rect 49205 -2720 49325 -2600
rect 49380 -2720 49500 -2600
rect 49545 -2720 49665 -2600
rect 49710 -2720 49830 -2600
rect 49875 -2720 49995 -2600
rect 50050 -2720 50170 -2600
rect 50215 -2720 50335 -2600
rect 50380 -2720 50500 -2600
rect 50545 -2720 50665 -2600
rect 50720 -2720 50840 -2600
rect 50885 -2720 51005 -2600
rect 51050 -2720 51170 -2600
rect 51215 -2720 51335 -2600
rect 51390 -2720 51510 -2600
rect 51555 -2720 51675 -2600
rect 51720 -2720 51840 -2600
rect 51885 -2720 52005 -2600
rect 52060 -2720 52180 -2600
rect 52225 -2720 52345 -2600
rect 52390 -2720 52510 -2600
rect 52555 -2720 52675 -2600
rect 52730 -2720 52850 -2600
rect 52895 -2720 53015 -2600
rect 53060 -2720 53180 -2600
rect 53225 -2720 53345 -2600
rect 47865 -2885 47985 -2765
rect 48040 -2885 48160 -2765
rect 48205 -2885 48325 -2765
rect 48370 -2885 48490 -2765
rect 48535 -2885 48655 -2765
rect 48710 -2885 48830 -2765
rect 48875 -2885 48995 -2765
rect 49040 -2885 49160 -2765
rect 49205 -2885 49325 -2765
rect 49380 -2885 49500 -2765
rect 49545 -2885 49665 -2765
rect 49710 -2885 49830 -2765
rect 49875 -2885 49995 -2765
rect 50050 -2885 50170 -2765
rect 50215 -2885 50335 -2765
rect 50380 -2885 50500 -2765
rect 50545 -2885 50665 -2765
rect 50720 -2885 50840 -2765
rect 50885 -2885 51005 -2765
rect 51050 -2885 51170 -2765
rect 51215 -2885 51335 -2765
rect 51390 -2885 51510 -2765
rect 51555 -2885 51675 -2765
rect 51720 -2885 51840 -2765
rect 51885 -2885 52005 -2765
rect 52060 -2885 52180 -2765
rect 52225 -2885 52345 -2765
rect 52390 -2885 52510 -2765
rect 52555 -2885 52675 -2765
rect 52730 -2885 52850 -2765
rect 52895 -2885 53015 -2765
rect 53060 -2885 53180 -2765
rect 53225 -2885 53345 -2765
rect 47865 -3050 47985 -2930
rect 48040 -3050 48160 -2930
rect 48205 -3050 48325 -2930
rect 48370 -3050 48490 -2930
rect 48535 -3050 48655 -2930
rect 48710 -3050 48830 -2930
rect 48875 -3050 48995 -2930
rect 49040 -3050 49160 -2930
rect 49205 -3050 49325 -2930
rect 49380 -3050 49500 -2930
rect 49545 -3050 49665 -2930
rect 49710 -3050 49830 -2930
rect 49875 -3050 49995 -2930
rect 50050 -3050 50170 -2930
rect 50215 -3050 50335 -2930
rect 50380 -3050 50500 -2930
rect 50545 -3050 50665 -2930
rect 50720 -3050 50840 -2930
rect 50885 -3050 51005 -2930
rect 51050 -3050 51170 -2930
rect 51215 -3050 51335 -2930
rect 51390 -3050 51510 -2930
rect 51555 -3050 51675 -2930
rect 51720 -3050 51840 -2930
rect 51885 -3050 52005 -2930
rect 52060 -3050 52180 -2930
rect 52225 -3050 52345 -2930
rect 52390 -3050 52510 -2930
rect 52555 -3050 52675 -2930
rect 52730 -3050 52850 -2930
rect 52895 -3050 53015 -2930
rect 53060 -3050 53180 -2930
rect 53225 -3050 53345 -2930
rect 47865 -3215 47985 -3095
rect 48040 -3215 48160 -3095
rect 48205 -3215 48325 -3095
rect 48370 -3215 48490 -3095
rect 48535 -3215 48655 -3095
rect 48710 -3215 48830 -3095
rect 48875 -3215 48995 -3095
rect 49040 -3215 49160 -3095
rect 49205 -3215 49325 -3095
rect 49380 -3215 49500 -3095
rect 49545 -3215 49665 -3095
rect 49710 -3215 49830 -3095
rect 49875 -3215 49995 -3095
rect 50050 -3215 50170 -3095
rect 50215 -3215 50335 -3095
rect 50380 -3215 50500 -3095
rect 50545 -3215 50665 -3095
rect 50720 -3215 50840 -3095
rect 50885 -3215 51005 -3095
rect 51050 -3215 51170 -3095
rect 51215 -3215 51335 -3095
rect 51390 -3215 51510 -3095
rect 51555 -3215 51675 -3095
rect 51720 -3215 51840 -3095
rect 51885 -3215 52005 -3095
rect 52060 -3215 52180 -3095
rect 52225 -3215 52345 -3095
rect 52390 -3215 52510 -3095
rect 52555 -3215 52675 -3095
rect 52730 -3215 52850 -3095
rect 52895 -3215 53015 -3095
rect 53060 -3215 53180 -3095
rect 53225 -3215 53345 -3095
rect 47865 -3390 47985 -3270
rect 48040 -3390 48160 -3270
rect 48205 -3390 48325 -3270
rect 48370 -3390 48490 -3270
rect 48535 -3390 48655 -3270
rect 48710 -3390 48830 -3270
rect 48875 -3390 48995 -3270
rect 49040 -3390 49160 -3270
rect 49205 -3390 49325 -3270
rect 49380 -3390 49500 -3270
rect 49545 -3390 49665 -3270
rect 49710 -3390 49830 -3270
rect 49875 -3390 49995 -3270
rect 50050 -3390 50170 -3270
rect 50215 -3390 50335 -3270
rect 50380 -3390 50500 -3270
rect 50545 -3390 50665 -3270
rect 50720 -3390 50840 -3270
rect 50885 -3390 51005 -3270
rect 51050 -3390 51170 -3270
rect 51215 -3390 51335 -3270
rect 51390 -3390 51510 -3270
rect 51555 -3390 51675 -3270
rect 51720 -3390 51840 -3270
rect 51885 -3390 52005 -3270
rect 52060 -3390 52180 -3270
rect 52225 -3390 52345 -3270
rect 52390 -3390 52510 -3270
rect 52555 -3390 52675 -3270
rect 52730 -3390 52850 -3270
rect 52895 -3390 53015 -3270
rect 53060 -3390 53180 -3270
rect 53225 -3390 53345 -3270
rect 47865 -3555 47985 -3435
rect 48040 -3555 48160 -3435
rect 48205 -3555 48325 -3435
rect 48370 -3555 48490 -3435
rect 48535 -3555 48655 -3435
rect 48710 -3555 48830 -3435
rect 48875 -3555 48995 -3435
rect 49040 -3555 49160 -3435
rect 49205 -3555 49325 -3435
rect 49380 -3555 49500 -3435
rect 49545 -3555 49665 -3435
rect 49710 -3555 49830 -3435
rect 49875 -3555 49995 -3435
rect 50050 -3555 50170 -3435
rect 50215 -3555 50335 -3435
rect 50380 -3555 50500 -3435
rect 50545 -3555 50665 -3435
rect 50720 -3555 50840 -3435
rect 50885 -3555 51005 -3435
rect 51050 -3555 51170 -3435
rect 51215 -3555 51335 -3435
rect 51390 -3555 51510 -3435
rect 51555 -3555 51675 -3435
rect 51720 -3555 51840 -3435
rect 51885 -3555 52005 -3435
rect 52060 -3555 52180 -3435
rect 52225 -3555 52345 -3435
rect 52390 -3555 52510 -3435
rect 52555 -3555 52675 -3435
rect 52730 -3555 52850 -3435
rect 52895 -3555 53015 -3435
rect 53060 -3555 53180 -3435
rect 53225 -3555 53345 -3435
rect 47865 -3720 47985 -3600
rect 48040 -3720 48160 -3600
rect 48205 -3720 48325 -3600
rect 48370 -3720 48490 -3600
rect 48535 -3720 48655 -3600
rect 48710 -3720 48830 -3600
rect 48875 -3720 48995 -3600
rect 49040 -3720 49160 -3600
rect 49205 -3720 49325 -3600
rect 49380 -3720 49500 -3600
rect 49545 -3720 49665 -3600
rect 49710 -3720 49830 -3600
rect 49875 -3720 49995 -3600
rect 50050 -3720 50170 -3600
rect 50215 -3720 50335 -3600
rect 50380 -3720 50500 -3600
rect 50545 -3720 50665 -3600
rect 50720 -3720 50840 -3600
rect 50885 -3720 51005 -3600
rect 51050 -3720 51170 -3600
rect 51215 -3720 51335 -3600
rect 51390 -3720 51510 -3600
rect 51555 -3720 51675 -3600
rect 51720 -3720 51840 -3600
rect 51885 -3720 52005 -3600
rect 52060 -3720 52180 -3600
rect 52225 -3720 52345 -3600
rect 52390 -3720 52510 -3600
rect 52555 -3720 52675 -3600
rect 52730 -3720 52850 -3600
rect 52895 -3720 53015 -3600
rect 53060 -3720 53180 -3600
rect 53225 -3720 53345 -3600
rect 47865 -3885 47985 -3765
rect 48040 -3885 48160 -3765
rect 48205 -3885 48325 -3765
rect 48370 -3885 48490 -3765
rect 48535 -3885 48655 -3765
rect 48710 -3885 48830 -3765
rect 48875 -3885 48995 -3765
rect 49040 -3885 49160 -3765
rect 49205 -3885 49325 -3765
rect 49380 -3885 49500 -3765
rect 49545 -3885 49665 -3765
rect 49710 -3885 49830 -3765
rect 49875 -3885 49995 -3765
rect 50050 -3885 50170 -3765
rect 50215 -3885 50335 -3765
rect 50380 -3885 50500 -3765
rect 50545 -3885 50665 -3765
rect 50720 -3885 50840 -3765
rect 50885 -3885 51005 -3765
rect 51050 -3885 51170 -3765
rect 51215 -3885 51335 -3765
rect 51390 -3885 51510 -3765
rect 51555 -3885 51675 -3765
rect 51720 -3885 51840 -3765
rect 51885 -3885 52005 -3765
rect 52060 -3885 52180 -3765
rect 52225 -3885 52345 -3765
rect 52390 -3885 52510 -3765
rect 52555 -3885 52675 -3765
rect 52730 -3885 52850 -3765
rect 52895 -3885 53015 -3765
rect 53060 -3885 53180 -3765
rect 53225 -3885 53345 -3765
rect 47865 -4060 47985 -3940
rect 48040 -4060 48160 -3940
rect 48205 -4060 48325 -3940
rect 48370 -4060 48490 -3940
rect 48535 -4060 48655 -3940
rect 48710 -4060 48830 -3940
rect 48875 -4060 48995 -3940
rect 49040 -4060 49160 -3940
rect 49205 -4060 49325 -3940
rect 49380 -4060 49500 -3940
rect 49545 -4060 49665 -3940
rect 49710 -4060 49830 -3940
rect 49875 -4060 49995 -3940
rect 50050 -4060 50170 -3940
rect 50215 -4060 50335 -3940
rect 50380 -4060 50500 -3940
rect 50545 -4060 50665 -3940
rect 50720 -4060 50840 -3940
rect 50885 -4060 51005 -3940
rect 51050 -4060 51170 -3940
rect 51215 -4060 51335 -3940
rect 51390 -4060 51510 -3940
rect 51555 -4060 51675 -3940
rect 51720 -4060 51840 -3940
rect 51885 -4060 52005 -3940
rect 52060 -4060 52180 -3940
rect 52225 -4060 52345 -3940
rect 52390 -4060 52510 -3940
rect 52555 -4060 52675 -3940
rect 52730 -4060 52850 -3940
rect 52895 -4060 53015 -3940
rect 53060 -4060 53180 -3940
rect 53225 -4060 53345 -3940
rect 30795 -4390 30915 -4270
rect 30960 -4390 31080 -4270
rect 31125 -4390 31245 -4270
rect 31290 -4390 31410 -4270
rect 31465 -4390 31585 -4270
rect 31630 -4390 31750 -4270
rect 31795 -4390 31915 -4270
rect 31960 -4390 32080 -4270
rect 32135 -4390 32255 -4270
rect 32300 -4390 32420 -4270
rect 32465 -4390 32585 -4270
rect 32630 -4390 32750 -4270
rect 32805 -4390 32925 -4270
rect 32970 -4390 33090 -4270
rect 33135 -4390 33255 -4270
rect 33300 -4390 33420 -4270
rect 33475 -4390 33595 -4270
rect 33640 -4390 33760 -4270
rect 33805 -4390 33925 -4270
rect 33970 -4390 34090 -4270
rect 34145 -4390 34265 -4270
rect 34310 -4390 34430 -4270
rect 34475 -4390 34595 -4270
rect 34640 -4390 34760 -4270
rect 34815 -4390 34935 -4270
rect 34980 -4390 35100 -4270
rect 35145 -4390 35265 -4270
rect 35310 -4390 35430 -4270
rect 35485 -4390 35605 -4270
rect 35650 -4390 35770 -4270
rect 35815 -4390 35935 -4270
rect 35980 -4390 36100 -4270
rect 36155 -4390 36275 -4270
rect 30795 -4565 30915 -4445
rect 30960 -4565 31080 -4445
rect 31125 -4565 31245 -4445
rect 31290 -4565 31410 -4445
rect 31465 -4565 31585 -4445
rect 31630 -4565 31750 -4445
rect 31795 -4565 31915 -4445
rect 31960 -4565 32080 -4445
rect 32135 -4565 32255 -4445
rect 32300 -4565 32420 -4445
rect 32465 -4565 32585 -4445
rect 32630 -4565 32750 -4445
rect 32805 -4565 32925 -4445
rect 32970 -4565 33090 -4445
rect 33135 -4565 33255 -4445
rect 33300 -4565 33420 -4445
rect 33475 -4565 33595 -4445
rect 33640 -4565 33760 -4445
rect 33805 -4565 33925 -4445
rect 33970 -4565 34090 -4445
rect 34145 -4565 34265 -4445
rect 34310 -4565 34430 -4445
rect 34475 -4565 34595 -4445
rect 34640 -4565 34760 -4445
rect 34815 -4565 34935 -4445
rect 34980 -4565 35100 -4445
rect 35145 -4565 35265 -4445
rect 35310 -4565 35430 -4445
rect 35485 -4565 35605 -4445
rect 35650 -4565 35770 -4445
rect 35815 -4565 35935 -4445
rect 35980 -4565 36100 -4445
rect 36155 -4565 36275 -4445
rect 30795 -4730 30915 -4610
rect 30960 -4730 31080 -4610
rect 31125 -4730 31245 -4610
rect 31290 -4730 31410 -4610
rect 31465 -4730 31585 -4610
rect 31630 -4730 31750 -4610
rect 31795 -4730 31915 -4610
rect 31960 -4730 32080 -4610
rect 32135 -4730 32255 -4610
rect 32300 -4730 32420 -4610
rect 32465 -4730 32585 -4610
rect 32630 -4730 32750 -4610
rect 32805 -4730 32925 -4610
rect 32970 -4730 33090 -4610
rect 33135 -4730 33255 -4610
rect 33300 -4730 33420 -4610
rect 33475 -4730 33595 -4610
rect 33640 -4730 33760 -4610
rect 33805 -4730 33925 -4610
rect 33970 -4730 34090 -4610
rect 34145 -4730 34265 -4610
rect 34310 -4730 34430 -4610
rect 34475 -4730 34595 -4610
rect 34640 -4730 34760 -4610
rect 34815 -4730 34935 -4610
rect 34980 -4730 35100 -4610
rect 35145 -4730 35265 -4610
rect 35310 -4730 35430 -4610
rect 35485 -4730 35605 -4610
rect 35650 -4730 35770 -4610
rect 35815 -4730 35935 -4610
rect 35980 -4730 36100 -4610
rect 36155 -4730 36275 -4610
rect 30795 -4895 30915 -4775
rect 30960 -4895 31080 -4775
rect 31125 -4895 31245 -4775
rect 31290 -4895 31410 -4775
rect 31465 -4895 31585 -4775
rect 31630 -4895 31750 -4775
rect 31795 -4895 31915 -4775
rect 31960 -4895 32080 -4775
rect 32135 -4895 32255 -4775
rect 32300 -4895 32420 -4775
rect 32465 -4895 32585 -4775
rect 32630 -4895 32750 -4775
rect 32805 -4895 32925 -4775
rect 32970 -4895 33090 -4775
rect 33135 -4895 33255 -4775
rect 33300 -4895 33420 -4775
rect 33475 -4895 33595 -4775
rect 33640 -4895 33760 -4775
rect 33805 -4895 33925 -4775
rect 33970 -4895 34090 -4775
rect 34145 -4895 34265 -4775
rect 34310 -4895 34430 -4775
rect 34475 -4895 34595 -4775
rect 34640 -4895 34760 -4775
rect 34815 -4895 34935 -4775
rect 34980 -4895 35100 -4775
rect 35145 -4895 35265 -4775
rect 35310 -4895 35430 -4775
rect 35485 -4895 35605 -4775
rect 35650 -4895 35770 -4775
rect 35815 -4895 35935 -4775
rect 35980 -4895 36100 -4775
rect 36155 -4895 36275 -4775
rect 30795 -5060 30915 -4940
rect 30960 -5060 31080 -4940
rect 31125 -5060 31245 -4940
rect 31290 -5060 31410 -4940
rect 31465 -5060 31585 -4940
rect 31630 -5060 31750 -4940
rect 31795 -5060 31915 -4940
rect 31960 -5060 32080 -4940
rect 32135 -5060 32255 -4940
rect 32300 -5060 32420 -4940
rect 32465 -5060 32585 -4940
rect 32630 -5060 32750 -4940
rect 32805 -5060 32925 -4940
rect 32970 -5060 33090 -4940
rect 33135 -5060 33255 -4940
rect 33300 -5060 33420 -4940
rect 33475 -5060 33595 -4940
rect 33640 -5060 33760 -4940
rect 33805 -5060 33925 -4940
rect 33970 -5060 34090 -4940
rect 34145 -5060 34265 -4940
rect 34310 -5060 34430 -4940
rect 34475 -5060 34595 -4940
rect 34640 -5060 34760 -4940
rect 34815 -5060 34935 -4940
rect 34980 -5060 35100 -4940
rect 35145 -5060 35265 -4940
rect 35310 -5060 35430 -4940
rect 35485 -5060 35605 -4940
rect 35650 -5060 35770 -4940
rect 35815 -5060 35935 -4940
rect 35980 -5060 36100 -4940
rect 36155 -5060 36275 -4940
rect 30795 -5235 30915 -5115
rect 30960 -5235 31080 -5115
rect 31125 -5235 31245 -5115
rect 31290 -5235 31410 -5115
rect 31465 -5235 31585 -5115
rect 31630 -5235 31750 -5115
rect 31795 -5235 31915 -5115
rect 31960 -5235 32080 -5115
rect 32135 -5235 32255 -5115
rect 32300 -5235 32420 -5115
rect 32465 -5235 32585 -5115
rect 32630 -5235 32750 -5115
rect 32805 -5235 32925 -5115
rect 32970 -5235 33090 -5115
rect 33135 -5235 33255 -5115
rect 33300 -5235 33420 -5115
rect 33475 -5235 33595 -5115
rect 33640 -5235 33760 -5115
rect 33805 -5235 33925 -5115
rect 33970 -5235 34090 -5115
rect 34145 -5235 34265 -5115
rect 34310 -5235 34430 -5115
rect 34475 -5235 34595 -5115
rect 34640 -5235 34760 -5115
rect 34815 -5235 34935 -5115
rect 34980 -5235 35100 -5115
rect 35145 -5235 35265 -5115
rect 35310 -5235 35430 -5115
rect 35485 -5235 35605 -5115
rect 35650 -5235 35770 -5115
rect 35815 -5235 35935 -5115
rect 35980 -5235 36100 -5115
rect 36155 -5235 36275 -5115
rect 30795 -5400 30915 -5280
rect 30960 -5400 31080 -5280
rect 31125 -5400 31245 -5280
rect 31290 -5400 31410 -5280
rect 31465 -5400 31585 -5280
rect 31630 -5400 31750 -5280
rect 31795 -5400 31915 -5280
rect 31960 -5400 32080 -5280
rect 32135 -5400 32255 -5280
rect 32300 -5400 32420 -5280
rect 32465 -5400 32585 -5280
rect 32630 -5400 32750 -5280
rect 32805 -5400 32925 -5280
rect 32970 -5400 33090 -5280
rect 33135 -5400 33255 -5280
rect 33300 -5400 33420 -5280
rect 33475 -5400 33595 -5280
rect 33640 -5400 33760 -5280
rect 33805 -5400 33925 -5280
rect 33970 -5400 34090 -5280
rect 34145 -5400 34265 -5280
rect 34310 -5400 34430 -5280
rect 34475 -5400 34595 -5280
rect 34640 -5400 34760 -5280
rect 34815 -5400 34935 -5280
rect 34980 -5400 35100 -5280
rect 35145 -5400 35265 -5280
rect 35310 -5400 35430 -5280
rect 35485 -5400 35605 -5280
rect 35650 -5400 35770 -5280
rect 35815 -5400 35935 -5280
rect 35980 -5400 36100 -5280
rect 36155 -5400 36275 -5280
rect 30795 -5565 30915 -5445
rect 30960 -5565 31080 -5445
rect 31125 -5565 31245 -5445
rect 31290 -5565 31410 -5445
rect 31465 -5565 31585 -5445
rect 31630 -5565 31750 -5445
rect 31795 -5565 31915 -5445
rect 31960 -5565 32080 -5445
rect 32135 -5565 32255 -5445
rect 32300 -5565 32420 -5445
rect 32465 -5565 32585 -5445
rect 32630 -5565 32750 -5445
rect 32805 -5565 32925 -5445
rect 32970 -5565 33090 -5445
rect 33135 -5565 33255 -5445
rect 33300 -5565 33420 -5445
rect 33475 -5565 33595 -5445
rect 33640 -5565 33760 -5445
rect 33805 -5565 33925 -5445
rect 33970 -5565 34090 -5445
rect 34145 -5565 34265 -5445
rect 34310 -5565 34430 -5445
rect 34475 -5565 34595 -5445
rect 34640 -5565 34760 -5445
rect 34815 -5565 34935 -5445
rect 34980 -5565 35100 -5445
rect 35145 -5565 35265 -5445
rect 35310 -5565 35430 -5445
rect 35485 -5565 35605 -5445
rect 35650 -5565 35770 -5445
rect 35815 -5565 35935 -5445
rect 35980 -5565 36100 -5445
rect 36155 -5565 36275 -5445
rect 30795 -5730 30915 -5610
rect 30960 -5730 31080 -5610
rect 31125 -5730 31245 -5610
rect 31290 -5730 31410 -5610
rect 31465 -5730 31585 -5610
rect 31630 -5730 31750 -5610
rect 31795 -5730 31915 -5610
rect 31960 -5730 32080 -5610
rect 32135 -5730 32255 -5610
rect 32300 -5730 32420 -5610
rect 32465 -5730 32585 -5610
rect 32630 -5730 32750 -5610
rect 32805 -5730 32925 -5610
rect 32970 -5730 33090 -5610
rect 33135 -5730 33255 -5610
rect 33300 -5730 33420 -5610
rect 33475 -5730 33595 -5610
rect 33640 -5730 33760 -5610
rect 33805 -5730 33925 -5610
rect 33970 -5730 34090 -5610
rect 34145 -5730 34265 -5610
rect 34310 -5730 34430 -5610
rect 34475 -5730 34595 -5610
rect 34640 -5730 34760 -5610
rect 34815 -5730 34935 -5610
rect 34980 -5730 35100 -5610
rect 35145 -5730 35265 -5610
rect 35310 -5730 35430 -5610
rect 35485 -5730 35605 -5610
rect 35650 -5730 35770 -5610
rect 35815 -5730 35935 -5610
rect 35980 -5730 36100 -5610
rect 36155 -5730 36275 -5610
rect 30795 -5905 30915 -5785
rect 30960 -5905 31080 -5785
rect 31125 -5905 31245 -5785
rect 31290 -5905 31410 -5785
rect 31465 -5905 31585 -5785
rect 31630 -5905 31750 -5785
rect 31795 -5905 31915 -5785
rect 31960 -5905 32080 -5785
rect 32135 -5905 32255 -5785
rect 32300 -5905 32420 -5785
rect 32465 -5905 32585 -5785
rect 32630 -5905 32750 -5785
rect 32805 -5905 32925 -5785
rect 32970 -5905 33090 -5785
rect 33135 -5905 33255 -5785
rect 33300 -5905 33420 -5785
rect 33475 -5905 33595 -5785
rect 33640 -5905 33760 -5785
rect 33805 -5905 33925 -5785
rect 33970 -5905 34090 -5785
rect 34145 -5905 34265 -5785
rect 34310 -5905 34430 -5785
rect 34475 -5905 34595 -5785
rect 34640 -5905 34760 -5785
rect 34815 -5905 34935 -5785
rect 34980 -5905 35100 -5785
rect 35145 -5905 35265 -5785
rect 35310 -5905 35430 -5785
rect 35485 -5905 35605 -5785
rect 35650 -5905 35770 -5785
rect 35815 -5905 35935 -5785
rect 35980 -5905 36100 -5785
rect 36155 -5905 36275 -5785
rect 30795 -6070 30915 -5950
rect 30960 -6070 31080 -5950
rect 31125 -6070 31245 -5950
rect 31290 -6070 31410 -5950
rect 31465 -6070 31585 -5950
rect 31630 -6070 31750 -5950
rect 31795 -6070 31915 -5950
rect 31960 -6070 32080 -5950
rect 32135 -6070 32255 -5950
rect 32300 -6070 32420 -5950
rect 32465 -6070 32585 -5950
rect 32630 -6070 32750 -5950
rect 32805 -6070 32925 -5950
rect 32970 -6070 33090 -5950
rect 33135 -6070 33255 -5950
rect 33300 -6070 33420 -5950
rect 33475 -6070 33595 -5950
rect 33640 -6070 33760 -5950
rect 33805 -6070 33925 -5950
rect 33970 -6070 34090 -5950
rect 34145 -6070 34265 -5950
rect 34310 -6070 34430 -5950
rect 34475 -6070 34595 -5950
rect 34640 -6070 34760 -5950
rect 34815 -6070 34935 -5950
rect 34980 -6070 35100 -5950
rect 35145 -6070 35265 -5950
rect 35310 -6070 35430 -5950
rect 35485 -6070 35605 -5950
rect 35650 -6070 35770 -5950
rect 35815 -6070 35935 -5950
rect 35980 -6070 36100 -5950
rect 36155 -6070 36275 -5950
rect 30795 -6235 30915 -6115
rect 30960 -6235 31080 -6115
rect 31125 -6235 31245 -6115
rect 31290 -6235 31410 -6115
rect 31465 -6235 31585 -6115
rect 31630 -6235 31750 -6115
rect 31795 -6235 31915 -6115
rect 31960 -6235 32080 -6115
rect 32135 -6235 32255 -6115
rect 32300 -6235 32420 -6115
rect 32465 -6235 32585 -6115
rect 32630 -6235 32750 -6115
rect 32805 -6235 32925 -6115
rect 32970 -6235 33090 -6115
rect 33135 -6235 33255 -6115
rect 33300 -6235 33420 -6115
rect 33475 -6235 33595 -6115
rect 33640 -6235 33760 -6115
rect 33805 -6235 33925 -6115
rect 33970 -6235 34090 -6115
rect 34145 -6235 34265 -6115
rect 34310 -6235 34430 -6115
rect 34475 -6235 34595 -6115
rect 34640 -6235 34760 -6115
rect 34815 -6235 34935 -6115
rect 34980 -6235 35100 -6115
rect 35145 -6235 35265 -6115
rect 35310 -6235 35430 -6115
rect 35485 -6235 35605 -6115
rect 35650 -6235 35770 -6115
rect 35815 -6235 35935 -6115
rect 35980 -6235 36100 -6115
rect 36155 -6235 36275 -6115
rect 30795 -6400 30915 -6280
rect 30960 -6400 31080 -6280
rect 31125 -6400 31245 -6280
rect 31290 -6400 31410 -6280
rect 31465 -6400 31585 -6280
rect 31630 -6400 31750 -6280
rect 31795 -6400 31915 -6280
rect 31960 -6400 32080 -6280
rect 32135 -6400 32255 -6280
rect 32300 -6400 32420 -6280
rect 32465 -6400 32585 -6280
rect 32630 -6400 32750 -6280
rect 32805 -6400 32925 -6280
rect 32970 -6400 33090 -6280
rect 33135 -6400 33255 -6280
rect 33300 -6400 33420 -6280
rect 33475 -6400 33595 -6280
rect 33640 -6400 33760 -6280
rect 33805 -6400 33925 -6280
rect 33970 -6400 34090 -6280
rect 34145 -6400 34265 -6280
rect 34310 -6400 34430 -6280
rect 34475 -6400 34595 -6280
rect 34640 -6400 34760 -6280
rect 34815 -6400 34935 -6280
rect 34980 -6400 35100 -6280
rect 35145 -6400 35265 -6280
rect 35310 -6400 35430 -6280
rect 35485 -6400 35605 -6280
rect 35650 -6400 35770 -6280
rect 35815 -6400 35935 -6280
rect 35980 -6400 36100 -6280
rect 36155 -6400 36275 -6280
rect 30795 -6575 30915 -6455
rect 30960 -6575 31080 -6455
rect 31125 -6575 31245 -6455
rect 31290 -6575 31410 -6455
rect 31465 -6575 31585 -6455
rect 31630 -6575 31750 -6455
rect 31795 -6575 31915 -6455
rect 31960 -6575 32080 -6455
rect 32135 -6575 32255 -6455
rect 32300 -6575 32420 -6455
rect 32465 -6575 32585 -6455
rect 32630 -6575 32750 -6455
rect 32805 -6575 32925 -6455
rect 32970 -6575 33090 -6455
rect 33135 -6575 33255 -6455
rect 33300 -6575 33420 -6455
rect 33475 -6575 33595 -6455
rect 33640 -6575 33760 -6455
rect 33805 -6575 33925 -6455
rect 33970 -6575 34090 -6455
rect 34145 -6575 34265 -6455
rect 34310 -6575 34430 -6455
rect 34475 -6575 34595 -6455
rect 34640 -6575 34760 -6455
rect 34815 -6575 34935 -6455
rect 34980 -6575 35100 -6455
rect 35145 -6575 35265 -6455
rect 35310 -6575 35430 -6455
rect 35485 -6575 35605 -6455
rect 35650 -6575 35770 -6455
rect 35815 -6575 35935 -6455
rect 35980 -6575 36100 -6455
rect 36155 -6575 36275 -6455
rect 30795 -6740 30915 -6620
rect 30960 -6740 31080 -6620
rect 31125 -6740 31245 -6620
rect 31290 -6740 31410 -6620
rect 31465 -6740 31585 -6620
rect 31630 -6740 31750 -6620
rect 31795 -6740 31915 -6620
rect 31960 -6740 32080 -6620
rect 32135 -6740 32255 -6620
rect 32300 -6740 32420 -6620
rect 32465 -6740 32585 -6620
rect 32630 -6740 32750 -6620
rect 32805 -6740 32925 -6620
rect 32970 -6740 33090 -6620
rect 33135 -6740 33255 -6620
rect 33300 -6740 33420 -6620
rect 33475 -6740 33595 -6620
rect 33640 -6740 33760 -6620
rect 33805 -6740 33925 -6620
rect 33970 -6740 34090 -6620
rect 34145 -6740 34265 -6620
rect 34310 -6740 34430 -6620
rect 34475 -6740 34595 -6620
rect 34640 -6740 34760 -6620
rect 34815 -6740 34935 -6620
rect 34980 -6740 35100 -6620
rect 35145 -6740 35265 -6620
rect 35310 -6740 35430 -6620
rect 35485 -6740 35605 -6620
rect 35650 -6740 35770 -6620
rect 35815 -6740 35935 -6620
rect 35980 -6740 36100 -6620
rect 36155 -6740 36275 -6620
rect 30795 -6905 30915 -6785
rect 30960 -6905 31080 -6785
rect 31125 -6905 31245 -6785
rect 31290 -6905 31410 -6785
rect 31465 -6905 31585 -6785
rect 31630 -6905 31750 -6785
rect 31795 -6905 31915 -6785
rect 31960 -6905 32080 -6785
rect 32135 -6905 32255 -6785
rect 32300 -6905 32420 -6785
rect 32465 -6905 32585 -6785
rect 32630 -6905 32750 -6785
rect 32805 -6905 32925 -6785
rect 32970 -6905 33090 -6785
rect 33135 -6905 33255 -6785
rect 33300 -6905 33420 -6785
rect 33475 -6905 33595 -6785
rect 33640 -6905 33760 -6785
rect 33805 -6905 33925 -6785
rect 33970 -6905 34090 -6785
rect 34145 -6905 34265 -6785
rect 34310 -6905 34430 -6785
rect 34475 -6905 34595 -6785
rect 34640 -6905 34760 -6785
rect 34815 -6905 34935 -6785
rect 34980 -6905 35100 -6785
rect 35145 -6905 35265 -6785
rect 35310 -6905 35430 -6785
rect 35485 -6905 35605 -6785
rect 35650 -6905 35770 -6785
rect 35815 -6905 35935 -6785
rect 35980 -6905 36100 -6785
rect 36155 -6905 36275 -6785
rect 30795 -7070 30915 -6950
rect 30960 -7070 31080 -6950
rect 31125 -7070 31245 -6950
rect 31290 -7070 31410 -6950
rect 31465 -7070 31585 -6950
rect 31630 -7070 31750 -6950
rect 31795 -7070 31915 -6950
rect 31960 -7070 32080 -6950
rect 32135 -7070 32255 -6950
rect 32300 -7070 32420 -6950
rect 32465 -7070 32585 -6950
rect 32630 -7070 32750 -6950
rect 32805 -7070 32925 -6950
rect 32970 -7070 33090 -6950
rect 33135 -7070 33255 -6950
rect 33300 -7070 33420 -6950
rect 33475 -7070 33595 -6950
rect 33640 -7070 33760 -6950
rect 33805 -7070 33925 -6950
rect 33970 -7070 34090 -6950
rect 34145 -7070 34265 -6950
rect 34310 -7070 34430 -6950
rect 34475 -7070 34595 -6950
rect 34640 -7070 34760 -6950
rect 34815 -7070 34935 -6950
rect 34980 -7070 35100 -6950
rect 35145 -7070 35265 -6950
rect 35310 -7070 35430 -6950
rect 35485 -7070 35605 -6950
rect 35650 -7070 35770 -6950
rect 35815 -7070 35935 -6950
rect 35980 -7070 36100 -6950
rect 36155 -7070 36275 -6950
rect 30795 -7245 30915 -7125
rect 30960 -7245 31080 -7125
rect 31125 -7245 31245 -7125
rect 31290 -7245 31410 -7125
rect 31465 -7245 31585 -7125
rect 31630 -7245 31750 -7125
rect 31795 -7245 31915 -7125
rect 31960 -7245 32080 -7125
rect 32135 -7245 32255 -7125
rect 32300 -7245 32420 -7125
rect 32465 -7245 32585 -7125
rect 32630 -7245 32750 -7125
rect 32805 -7245 32925 -7125
rect 32970 -7245 33090 -7125
rect 33135 -7245 33255 -7125
rect 33300 -7245 33420 -7125
rect 33475 -7245 33595 -7125
rect 33640 -7245 33760 -7125
rect 33805 -7245 33925 -7125
rect 33970 -7245 34090 -7125
rect 34145 -7245 34265 -7125
rect 34310 -7245 34430 -7125
rect 34475 -7245 34595 -7125
rect 34640 -7245 34760 -7125
rect 34815 -7245 34935 -7125
rect 34980 -7245 35100 -7125
rect 35145 -7245 35265 -7125
rect 35310 -7245 35430 -7125
rect 35485 -7245 35605 -7125
rect 35650 -7245 35770 -7125
rect 35815 -7245 35935 -7125
rect 35980 -7245 36100 -7125
rect 36155 -7245 36275 -7125
rect 30795 -7410 30915 -7290
rect 30960 -7410 31080 -7290
rect 31125 -7410 31245 -7290
rect 31290 -7410 31410 -7290
rect 31465 -7410 31585 -7290
rect 31630 -7410 31750 -7290
rect 31795 -7410 31915 -7290
rect 31960 -7410 32080 -7290
rect 32135 -7410 32255 -7290
rect 32300 -7410 32420 -7290
rect 32465 -7410 32585 -7290
rect 32630 -7410 32750 -7290
rect 32805 -7410 32925 -7290
rect 32970 -7410 33090 -7290
rect 33135 -7410 33255 -7290
rect 33300 -7410 33420 -7290
rect 33475 -7410 33595 -7290
rect 33640 -7410 33760 -7290
rect 33805 -7410 33925 -7290
rect 33970 -7410 34090 -7290
rect 34145 -7410 34265 -7290
rect 34310 -7410 34430 -7290
rect 34475 -7410 34595 -7290
rect 34640 -7410 34760 -7290
rect 34815 -7410 34935 -7290
rect 34980 -7410 35100 -7290
rect 35145 -7410 35265 -7290
rect 35310 -7410 35430 -7290
rect 35485 -7410 35605 -7290
rect 35650 -7410 35770 -7290
rect 35815 -7410 35935 -7290
rect 35980 -7410 36100 -7290
rect 36155 -7410 36275 -7290
rect 30795 -7575 30915 -7455
rect 30960 -7575 31080 -7455
rect 31125 -7575 31245 -7455
rect 31290 -7575 31410 -7455
rect 31465 -7575 31585 -7455
rect 31630 -7575 31750 -7455
rect 31795 -7575 31915 -7455
rect 31960 -7575 32080 -7455
rect 32135 -7575 32255 -7455
rect 32300 -7575 32420 -7455
rect 32465 -7575 32585 -7455
rect 32630 -7575 32750 -7455
rect 32805 -7575 32925 -7455
rect 32970 -7575 33090 -7455
rect 33135 -7575 33255 -7455
rect 33300 -7575 33420 -7455
rect 33475 -7575 33595 -7455
rect 33640 -7575 33760 -7455
rect 33805 -7575 33925 -7455
rect 33970 -7575 34090 -7455
rect 34145 -7575 34265 -7455
rect 34310 -7575 34430 -7455
rect 34475 -7575 34595 -7455
rect 34640 -7575 34760 -7455
rect 34815 -7575 34935 -7455
rect 34980 -7575 35100 -7455
rect 35145 -7575 35265 -7455
rect 35310 -7575 35430 -7455
rect 35485 -7575 35605 -7455
rect 35650 -7575 35770 -7455
rect 35815 -7575 35935 -7455
rect 35980 -7575 36100 -7455
rect 36155 -7575 36275 -7455
rect 30795 -7740 30915 -7620
rect 30960 -7740 31080 -7620
rect 31125 -7740 31245 -7620
rect 31290 -7740 31410 -7620
rect 31465 -7740 31585 -7620
rect 31630 -7740 31750 -7620
rect 31795 -7740 31915 -7620
rect 31960 -7740 32080 -7620
rect 32135 -7740 32255 -7620
rect 32300 -7740 32420 -7620
rect 32465 -7740 32585 -7620
rect 32630 -7740 32750 -7620
rect 32805 -7740 32925 -7620
rect 32970 -7740 33090 -7620
rect 33135 -7740 33255 -7620
rect 33300 -7740 33420 -7620
rect 33475 -7740 33595 -7620
rect 33640 -7740 33760 -7620
rect 33805 -7740 33925 -7620
rect 33970 -7740 34090 -7620
rect 34145 -7740 34265 -7620
rect 34310 -7740 34430 -7620
rect 34475 -7740 34595 -7620
rect 34640 -7740 34760 -7620
rect 34815 -7740 34935 -7620
rect 34980 -7740 35100 -7620
rect 35145 -7740 35265 -7620
rect 35310 -7740 35430 -7620
rect 35485 -7740 35605 -7620
rect 35650 -7740 35770 -7620
rect 35815 -7740 35935 -7620
rect 35980 -7740 36100 -7620
rect 36155 -7740 36275 -7620
rect 30795 -7915 30915 -7795
rect 30960 -7915 31080 -7795
rect 31125 -7915 31245 -7795
rect 31290 -7915 31410 -7795
rect 31465 -7915 31585 -7795
rect 31630 -7915 31750 -7795
rect 31795 -7915 31915 -7795
rect 31960 -7915 32080 -7795
rect 32135 -7915 32255 -7795
rect 32300 -7915 32420 -7795
rect 32465 -7915 32585 -7795
rect 32630 -7915 32750 -7795
rect 32805 -7915 32925 -7795
rect 32970 -7915 33090 -7795
rect 33135 -7915 33255 -7795
rect 33300 -7915 33420 -7795
rect 33475 -7915 33595 -7795
rect 33640 -7915 33760 -7795
rect 33805 -7915 33925 -7795
rect 33970 -7915 34090 -7795
rect 34145 -7915 34265 -7795
rect 34310 -7915 34430 -7795
rect 34475 -7915 34595 -7795
rect 34640 -7915 34760 -7795
rect 34815 -7915 34935 -7795
rect 34980 -7915 35100 -7795
rect 35145 -7915 35265 -7795
rect 35310 -7915 35430 -7795
rect 35485 -7915 35605 -7795
rect 35650 -7915 35770 -7795
rect 35815 -7915 35935 -7795
rect 35980 -7915 36100 -7795
rect 36155 -7915 36275 -7795
rect 30795 -8080 30915 -7960
rect 30960 -8080 31080 -7960
rect 31125 -8080 31245 -7960
rect 31290 -8080 31410 -7960
rect 31465 -8080 31585 -7960
rect 31630 -8080 31750 -7960
rect 31795 -8080 31915 -7960
rect 31960 -8080 32080 -7960
rect 32135 -8080 32255 -7960
rect 32300 -8080 32420 -7960
rect 32465 -8080 32585 -7960
rect 32630 -8080 32750 -7960
rect 32805 -8080 32925 -7960
rect 32970 -8080 33090 -7960
rect 33135 -8080 33255 -7960
rect 33300 -8080 33420 -7960
rect 33475 -8080 33595 -7960
rect 33640 -8080 33760 -7960
rect 33805 -8080 33925 -7960
rect 33970 -8080 34090 -7960
rect 34145 -8080 34265 -7960
rect 34310 -8080 34430 -7960
rect 34475 -8080 34595 -7960
rect 34640 -8080 34760 -7960
rect 34815 -8080 34935 -7960
rect 34980 -8080 35100 -7960
rect 35145 -8080 35265 -7960
rect 35310 -8080 35430 -7960
rect 35485 -8080 35605 -7960
rect 35650 -8080 35770 -7960
rect 35815 -8080 35935 -7960
rect 35980 -8080 36100 -7960
rect 36155 -8080 36275 -7960
rect 30795 -8245 30915 -8125
rect 30960 -8245 31080 -8125
rect 31125 -8245 31245 -8125
rect 31290 -8245 31410 -8125
rect 31465 -8245 31585 -8125
rect 31630 -8245 31750 -8125
rect 31795 -8245 31915 -8125
rect 31960 -8245 32080 -8125
rect 32135 -8245 32255 -8125
rect 32300 -8245 32420 -8125
rect 32465 -8245 32585 -8125
rect 32630 -8245 32750 -8125
rect 32805 -8245 32925 -8125
rect 32970 -8245 33090 -8125
rect 33135 -8245 33255 -8125
rect 33300 -8245 33420 -8125
rect 33475 -8245 33595 -8125
rect 33640 -8245 33760 -8125
rect 33805 -8245 33925 -8125
rect 33970 -8245 34090 -8125
rect 34145 -8245 34265 -8125
rect 34310 -8245 34430 -8125
rect 34475 -8245 34595 -8125
rect 34640 -8245 34760 -8125
rect 34815 -8245 34935 -8125
rect 34980 -8245 35100 -8125
rect 35145 -8245 35265 -8125
rect 35310 -8245 35430 -8125
rect 35485 -8245 35605 -8125
rect 35650 -8245 35770 -8125
rect 35815 -8245 35935 -8125
rect 35980 -8245 36100 -8125
rect 36155 -8245 36275 -8125
rect 30795 -8410 30915 -8290
rect 30960 -8410 31080 -8290
rect 31125 -8410 31245 -8290
rect 31290 -8410 31410 -8290
rect 31465 -8410 31585 -8290
rect 31630 -8410 31750 -8290
rect 31795 -8410 31915 -8290
rect 31960 -8410 32080 -8290
rect 32135 -8410 32255 -8290
rect 32300 -8410 32420 -8290
rect 32465 -8410 32585 -8290
rect 32630 -8410 32750 -8290
rect 32805 -8410 32925 -8290
rect 32970 -8410 33090 -8290
rect 33135 -8410 33255 -8290
rect 33300 -8410 33420 -8290
rect 33475 -8410 33595 -8290
rect 33640 -8410 33760 -8290
rect 33805 -8410 33925 -8290
rect 33970 -8410 34090 -8290
rect 34145 -8410 34265 -8290
rect 34310 -8410 34430 -8290
rect 34475 -8410 34595 -8290
rect 34640 -8410 34760 -8290
rect 34815 -8410 34935 -8290
rect 34980 -8410 35100 -8290
rect 35145 -8410 35265 -8290
rect 35310 -8410 35430 -8290
rect 35485 -8410 35605 -8290
rect 35650 -8410 35770 -8290
rect 35815 -8410 35935 -8290
rect 35980 -8410 36100 -8290
rect 36155 -8410 36275 -8290
rect 30795 -8585 30915 -8465
rect 30960 -8585 31080 -8465
rect 31125 -8585 31245 -8465
rect 31290 -8585 31410 -8465
rect 31465 -8585 31585 -8465
rect 31630 -8585 31750 -8465
rect 31795 -8585 31915 -8465
rect 31960 -8585 32080 -8465
rect 32135 -8585 32255 -8465
rect 32300 -8585 32420 -8465
rect 32465 -8585 32585 -8465
rect 32630 -8585 32750 -8465
rect 32805 -8585 32925 -8465
rect 32970 -8585 33090 -8465
rect 33135 -8585 33255 -8465
rect 33300 -8585 33420 -8465
rect 33475 -8585 33595 -8465
rect 33640 -8585 33760 -8465
rect 33805 -8585 33925 -8465
rect 33970 -8585 34090 -8465
rect 34145 -8585 34265 -8465
rect 34310 -8585 34430 -8465
rect 34475 -8585 34595 -8465
rect 34640 -8585 34760 -8465
rect 34815 -8585 34935 -8465
rect 34980 -8585 35100 -8465
rect 35145 -8585 35265 -8465
rect 35310 -8585 35430 -8465
rect 35485 -8585 35605 -8465
rect 35650 -8585 35770 -8465
rect 35815 -8585 35935 -8465
rect 35980 -8585 36100 -8465
rect 36155 -8585 36275 -8465
rect 30795 -8750 30915 -8630
rect 30960 -8750 31080 -8630
rect 31125 -8750 31245 -8630
rect 31290 -8750 31410 -8630
rect 31465 -8750 31585 -8630
rect 31630 -8750 31750 -8630
rect 31795 -8750 31915 -8630
rect 31960 -8750 32080 -8630
rect 32135 -8750 32255 -8630
rect 32300 -8750 32420 -8630
rect 32465 -8750 32585 -8630
rect 32630 -8750 32750 -8630
rect 32805 -8750 32925 -8630
rect 32970 -8750 33090 -8630
rect 33135 -8750 33255 -8630
rect 33300 -8750 33420 -8630
rect 33475 -8750 33595 -8630
rect 33640 -8750 33760 -8630
rect 33805 -8750 33925 -8630
rect 33970 -8750 34090 -8630
rect 34145 -8750 34265 -8630
rect 34310 -8750 34430 -8630
rect 34475 -8750 34595 -8630
rect 34640 -8750 34760 -8630
rect 34815 -8750 34935 -8630
rect 34980 -8750 35100 -8630
rect 35145 -8750 35265 -8630
rect 35310 -8750 35430 -8630
rect 35485 -8750 35605 -8630
rect 35650 -8750 35770 -8630
rect 35815 -8750 35935 -8630
rect 35980 -8750 36100 -8630
rect 36155 -8750 36275 -8630
rect 30795 -8915 30915 -8795
rect 30960 -8915 31080 -8795
rect 31125 -8915 31245 -8795
rect 31290 -8915 31410 -8795
rect 31465 -8915 31585 -8795
rect 31630 -8915 31750 -8795
rect 31795 -8915 31915 -8795
rect 31960 -8915 32080 -8795
rect 32135 -8915 32255 -8795
rect 32300 -8915 32420 -8795
rect 32465 -8915 32585 -8795
rect 32630 -8915 32750 -8795
rect 32805 -8915 32925 -8795
rect 32970 -8915 33090 -8795
rect 33135 -8915 33255 -8795
rect 33300 -8915 33420 -8795
rect 33475 -8915 33595 -8795
rect 33640 -8915 33760 -8795
rect 33805 -8915 33925 -8795
rect 33970 -8915 34090 -8795
rect 34145 -8915 34265 -8795
rect 34310 -8915 34430 -8795
rect 34475 -8915 34595 -8795
rect 34640 -8915 34760 -8795
rect 34815 -8915 34935 -8795
rect 34980 -8915 35100 -8795
rect 35145 -8915 35265 -8795
rect 35310 -8915 35430 -8795
rect 35485 -8915 35605 -8795
rect 35650 -8915 35770 -8795
rect 35815 -8915 35935 -8795
rect 35980 -8915 36100 -8795
rect 36155 -8915 36275 -8795
rect 30795 -9080 30915 -8960
rect 30960 -9080 31080 -8960
rect 31125 -9080 31245 -8960
rect 31290 -9080 31410 -8960
rect 31465 -9080 31585 -8960
rect 31630 -9080 31750 -8960
rect 31795 -9080 31915 -8960
rect 31960 -9080 32080 -8960
rect 32135 -9080 32255 -8960
rect 32300 -9080 32420 -8960
rect 32465 -9080 32585 -8960
rect 32630 -9080 32750 -8960
rect 32805 -9080 32925 -8960
rect 32970 -9080 33090 -8960
rect 33135 -9080 33255 -8960
rect 33300 -9080 33420 -8960
rect 33475 -9080 33595 -8960
rect 33640 -9080 33760 -8960
rect 33805 -9080 33925 -8960
rect 33970 -9080 34090 -8960
rect 34145 -9080 34265 -8960
rect 34310 -9080 34430 -8960
rect 34475 -9080 34595 -8960
rect 34640 -9080 34760 -8960
rect 34815 -9080 34935 -8960
rect 34980 -9080 35100 -8960
rect 35145 -9080 35265 -8960
rect 35310 -9080 35430 -8960
rect 35485 -9080 35605 -8960
rect 35650 -9080 35770 -8960
rect 35815 -9080 35935 -8960
rect 35980 -9080 36100 -8960
rect 36155 -9080 36275 -8960
rect 30795 -9255 30915 -9135
rect 30960 -9255 31080 -9135
rect 31125 -9255 31245 -9135
rect 31290 -9255 31410 -9135
rect 31465 -9255 31585 -9135
rect 31630 -9255 31750 -9135
rect 31795 -9255 31915 -9135
rect 31960 -9255 32080 -9135
rect 32135 -9255 32255 -9135
rect 32300 -9255 32420 -9135
rect 32465 -9255 32585 -9135
rect 32630 -9255 32750 -9135
rect 32805 -9255 32925 -9135
rect 32970 -9255 33090 -9135
rect 33135 -9255 33255 -9135
rect 33300 -9255 33420 -9135
rect 33475 -9255 33595 -9135
rect 33640 -9255 33760 -9135
rect 33805 -9255 33925 -9135
rect 33970 -9255 34090 -9135
rect 34145 -9255 34265 -9135
rect 34310 -9255 34430 -9135
rect 34475 -9255 34595 -9135
rect 34640 -9255 34760 -9135
rect 34815 -9255 34935 -9135
rect 34980 -9255 35100 -9135
rect 35145 -9255 35265 -9135
rect 35310 -9255 35430 -9135
rect 35485 -9255 35605 -9135
rect 35650 -9255 35770 -9135
rect 35815 -9255 35935 -9135
rect 35980 -9255 36100 -9135
rect 36155 -9255 36275 -9135
rect 30795 -9420 30915 -9300
rect 30960 -9420 31080 -9300
rect 31125 -9420 31245 -9300
rect 31290 -9420 31410 -9300
rect 31465 -9420 31585 -9300
rect 31630 -9420 31750 -9300
rect 31795 -9420 31915 -9300
rect 31960 -9420 32080 -9300
rect 32135 -9420 32255 -9300
rect 32300 -9420 32420 -9300
rect 32465 -9420 32585 -9300
rect 32630 -9420 32750 -9300
rect 32805 -9420 32925 -9300
rect 32970 -9420 33090 -9300
rect 33135 -9420 33255 -9300
rect 33300 -9420 33420 -9300
rect 33475 -9420 33595 -9300
rect 33640 -9420 33760 -9300
rect 33805 -9420 33925 -9300
rect 33970 -9420 34090 -9300
rect 34145 -9420 34265 -9300
rect 34310 -9420 34430 -9300
rect 34475 -9420 34595 -9300
rect 34640 -9420 34760 -9300
rect 34815 -9420 34935 -9300
rect 34980 -9420 35100 -9300
rect 35145 -9420 35265 -9300
rect 35310 -9420 35430 -9300
rect 35485 -9420 35605 -9300
rect 35650 -9420 35770 -9300
rect 35815 -9420 35935 -9300
rect 35980 -9420 36100 -9300
rect 36155 -9420 36275 -9300
rect 30795 -9585 30915 -9465
rect 30960 -9585 31080 -9465
rect 31125 -9585 31245 -9465
rect 31290 -9585 31410 -9465
rect 31465 -9585 31585 -9465
rect 31630 -9585 31750 -9465
rect 31795 -9585 31915 -9465
rect 31960 -9585 32080 -9465
rect 32135 -9585 32255 -9465
rect 32300 -9585 32420 -9465
rect 32465 -9585 32585 -9465
rect 32630 -9585 32750 -9465
rect 32805 -9585 32925 -9465
rect 32970 -9585 33090 -9465
rect 33135 -9585 33255 -9465
rect 33300 -9585 33420 -9465
rect 33475 -9585 33595 -9465
rect 33640 -9585 33760 -9465
rect 33805 -9585 33925 -9465
rect 33970 -9585 34090 -9465
rect 34145 -9585 34265 -9465
rect 34310 -9585 34430 -9465
rect 34475 -9585 34595 -9465
rect 34640 -9585 34760 -9465
rect 34815 -9585 34935 -9465
rect 34980 -9585 35100 -9465
rect 35145 -9585 35265 -9465
rect 35310 -9585 35430 -9465
rect 35485 -9585 35605 -9465
rect 35650 -9585 35770 -9465
rect 35815 -9585 35935 -9465
rect 35980 -9585 36100 -9465
rect 36155 -9585 36275 -9465
rect 30795 -9750 30915 -9630
rect 30960 -9750 31080 -9630
rect 31125 -9750 31245 -9630
rect 31290 -9750 31410 -9630
rect 31465 -9750 31585 -9630
rect 31630 -9750 31750 -9630
rect 31795 -9750 31915 -9630
rect 31960 -9750 32080 -9630
rect 32135 -9750 32255 -9630
rect 32300 -9750 32420 -9630
rect 32465 -9750 32585 -9630
rect 32630 -9750 32750 -9630
rect 32805 -9750 32925 -9630
rect 32970 -9750 33090 -9630
rect 33135 -9750 33255 -9630
rect 33300 -9750 33420 -9630
rect 33475 -9750 33595 -9630
rect 33640 -9750 33760 -9630
rect 33805 -9750 33925 -9630
rect 33970 -9750 34090 -9630
rect 34145 -9750 34265 -9630
rect 34310 -9750 34430 -9630
rect 34475 -9750 34595 -9630
rect 34640 -9750 34760 -9630
rect 34815 -9750 34935 -9630
rect 34980 -9750 35100 -9630
rect 35145 -9750 35265 -9630
rect 35310 -9750 35430 -9630
rect 35485 -9750 35605 -9630
rect 35650 -9750 35770 -9630
rect 35815 -9750 35935 -9630
rect 35980 -9750 36100 -9630
rect 36155 -9750 36275 -9630
rect 36485 -4390 36605 -4270
rect 36650 -4390 36770 -4270
rect 36815 -4390 36935 -4270
rect 36980 -4390 37100 -4270
rect 37155 -4390 37275 -4270
rect 37320 -4390 37440 -4270
rect 37485 -4390 37605 -4270
rect 37650 -4390 37770 -4270
rect 37825 -4390 37945 -4270
rect 37990 -4390 38110 -4270
rect 38155 -4390 38275 -4270
rect 38320 -4390 38440 -4270
rect 38495 -4390 38615 -4270
rect 38660 -4390 38780 -4270
rect 38825 -4390 38945 -4270
rect 38990 -4390 39110 -4270
rect 39165 -4390 39285 -4270
rect 39330 -4390 39450 -4270
rect 39495 -4390 39615 -4270
rect 39660 -4390 39780 -4270
rect 39835 -4390 39955 -4270
rect 40000 -4390 40120 -4270
rect 40165 -4390 40285 -4270
rect 40330 -4390 40450 -4270
rect 40505 -4390 40625 -4270
rect 40670 -4390 40790 -4270
rect 40835 -4390 40955 -4270
rect 41000 -4390 41120 -4270
rect 41175 -4390 41295 -4270
rect 41340 -4390 41460 -4270
rect 41505 -4390 41625 -4270
rect 41670 -4390 41790 -4270
rect 41845 -4390 41965 -4270
rect 36485 -4565 36605 -4445
rect 36650 -4565 36770 -4445
rect 36815 -4565 36935 -4445
rect 36980 -4565 37100 -4445
rect 37155 -4565 37275 -4445
rect 37320 -4565 37440 -4445
rect 37485 -4565 37605 -4445
rect 37650 -4565 37770 -4445
rect 37825 -4565 37945 -4445
rect 37990 -4565 38110 -4445
rect 38155 -4565 38275 -4445
rect 38320 -4565 38440 -4445
rect 38495 -4565 38615 -4445
rect 38660 -4565 38780 -4445
rect 38825 -4565 38945 -4445
rect 38990 -4565 39110 -4445
rect 39165 -4565 39285 -4445
rect 39330 -4565 39450 -4445
rect 39495 -4565 39615 -4445
rect 39660 -4565 39780 -4445
rect 39835 -4565 39955 -4445
rect 40000 -4565 40120 -4445
rect 40165 -4565 40285 -4445
rect 40330 -4565 40450 -4445
rect 40505 -4565 40625 -4445
rect 40670 -4565 40790 -4445
rect 40835 -4565 40955 -4445
rect 41000 -4565 41120 -4445
rect 41175 -4565 41295 -4445
rect 41340 -4565 41460 -4445
rect 41505 -4565 41625 -4445
rect 41670 -4565 41790 -4445
rect 41845 -4565 41965 -4445
rect 36485 -4730 36605 -4610
rect 36650 -4730 36770 -4610
rect 36815 -4730 36935 -4610
rect 36980 -4730 37100 -4610
rect 37155 -4730 37275 -4610
rect 37320 -4730 37440 -4610
rect 37485 -4730 37605 -4610
rect 37650 -4730 37770 -4610
rect 37825 -4730 37945 -4610
rect 37990 -4730 38110 -4610
rect 38155 -4730 38275 -4610
rect 38320 -4730 38440 -4610
rect 38495 -4730 38615 -4610
rect 38660 -4730 38780 -4610
rect 38825 -4730 38945 -4610
rect 38990 -4730 39110 -4610
rect 39165 -4730 39285 -4610
rect 39330 -4730 39450 -4610
rect 39495 -4730 39615 -4610
rect 39660 -4730 39780 -4610
rect 39835 -4730 39955 -4610
rect 40000 -4730 40120 -4610
rect 40165 -4730 40285 -4610
rect 40330 -4730 40450 -4610
rect 40505 -4730 40625 -4610
rect 40670 -4730 40790 -4610
rect 40835 -4730 40955 -4610
rect 41000 -4730 41120 -4610
rect 41175 -4730 41295 -4610
rect 41340 -4730 41460 -4610
rect 41505 -4730 41625 -4610
rect 41670 -4730 41790 -4610
rect 41845 -4730 41965 -4610
rect 36485 -4895 36605 -4775
rect 36650 -4895 36770 -4775
rect 36815 -4895 36935 -4775
rect 36980 -4895 37100 -4775
rect 37155 -4895 37275 -4775
rect 37320 -4895 37440 -4775
rect 37485 -4895 37605 -4775
rect 37650 -4895 37770 -4775
rect 37825 -4895 37945 -4775
rect 37990 -4895 38110 -4775
rect 38155 -4895 38275 -4775
rect 38320 -4895 38440 -4775
rect 38495 -4895 38615 -4775
rect 38660 -4895 38780 -4775
rect 38825 -4895 38945 -4775
rect 38990 -4895 39110 -4775
rect 39165 -4895 39285 -4775
rect 39330 -4895 39450 -4775
rect 39495 -4895 39615 -4775
rect 39660 -4895 39780 -4775
rect 39835 -4895 39955 -4775
rect 40000 -4895 40120 -4775
rect 40165 -4895 40285 -4775
rect 40330 -4895 40450 -4775
rect 40505 -4895 40625 -4775
rect 40670 -4895 40790 -4775
rect 40835 -4895 40955 -4775
rect 41000 -4895 41120 -4775
rect 41175 -4895 41295 -4775
rect 41340 -4895 41460 -4775
rect 41505 -4895 41625 -4775
rect 41670 -4895 41790 -4775
rect 41845 -4895 41965 -4775
rect 36485 -5060 36605 -4940
rect 36650 -5060 36770 -4940
rect 36815 -5060 36935 -4940
rect 36980 -5060 37100 -4940
rect 37155 -5060 37275 -4940
rect 37320 -5060 37440 -4940
rect 37485 -5060 37605 -4940
rect 37650 -5060 37770 -4940
rect 37825 -5060 37945 -4940
rect 37990 -5060 38110 -4940
rect 38155 -5060 38275 -4940
rect 38320 -5060 38440 -4940
rect 38495 -5060 38615 -4940
rect 38660 -5060 38780 -4940
rect 38825 -5060 38945 -4940
rect 38990 -5060 39110 -4940
rect 39165 -5060 39285 -4940
rect 39330 -5060 39450 -4940
rect 39495 -5060 39615 -4940
rect 39660 -5060 39780 -4940
rect 39835 -5060 39955 -4940
rect 40000 -5060 40120 -4940
rect 40165 -5060 40285 -4940
rect 40330 -5060 40450 -4940
rect 40505 -5060 40625 -4940
rect 40670 -5060 40790 -4940
rect 40835 -5060 40955 -4940
rect 41000 -5060 41120 -4940
rect 41175 -5060 41295 -4940
rect 41340 -5060 41460 -4940
rect 41505 -5060 41625 -4940
rect 41670 -5060 41790 -4940
rect 41845 -5060 41965 -4940
rect 36485 -5235 36605 -5115
rect 36650 -5235 36770 -5115
rect 36815 -5235 36935 -5115
rect 36980 -5235 37100 -5115
rect 37155 -5235 37275 -5115
rect 37320 -5235 37440 -5115
rect 37485 -5235 37605 -5115
rect 37650 -5235 37770 -5115
rect 37825 -5235 37945 -5115
rect 37990 -5235 38110 -5115
rect 38155 -5235 38275 -5115
rect 38320 -5235 38440 -5115
rect 38495 -5235 38615 -5115
rect 38660 -5235 38780 -5115
rect 38825 -5235 38945 -5115
rect 38990 -5235 39110 -5115
rect 39165 -5235 39285 -5115
rect 39330 -5235 39450 -5115
rect 39495 -5235 39615 -5115
rect 39660 -5235 39780 -5115
rect 39835 -5235 39955 -5115
rect 40000 -5235 40120 -5115
rect 40165 -5235 40285 -5115
rect 40330 -5235 40450 -5115
rect 40505 -5235 40625 -5115
rect 40670 -5235 40790 -5115
rect 40835 -5235 40955 -5115
rect 41000 -5235 41120 -5115
rect 41175 -5235 41295 -5115
rect 41340 -5235 41460 -5115
rect 41505 -5235 41625 -5115
rect 41670 -5235 41790 -5115
rect 41845 -5235 41965 -5115
rect 36485 -5400 36605 -5280
rect 36650 -5400 36770 -5280
rect 36815 -5400 36935 -5280
rect 36980 -5400 37100 -5280
rect 37155 -5400 37275 -5280
rect 37320 -5400 37440 -5280
rect 37485 -5400 37605 -5280
rect 37650 -5400 37770 -5280
rect 37825 -5400 37945 -5280
rect 37990 -5400 38110 -5280
rect 38155 -5400 38275 -5280
rect 38320 -5400 38440 -5280
rect 38495 -5400 38615 -5280
rect 38660 -5400 38780 -5280
rect 38825 -5400 38945 -5280
rect 38990 -5400 39110 -5280
rect 39165 -5400 39285 -5280
rect 39330 -5400 39450 -5280
rect 39495 -5400 39615 -5280
rect 39660 -5400 39780 -5280
rect 39835 -5400 39955 -5280
rect 40000 -5400 40120 -5280
rect 40165 -5400 40285 -5280
rect 40330 -5400 40450 -5280
rect 40505 -5400 40625 -5280
rect 40670 -5400 40790 -5280
rect 40835 -5400 40955 -5280
rect 41000 -5400 41120 -5280
rect 41175 -5400 41295 -5280
rect 41340 -5400 41460 -5280
rect 41505 -5400 41625 -5280
rect 41670 -5400 41790 -5280
rect 41845 -5400 41965 -5280
rect 36485 -5565 36605 -5445
rect 36650 -5565 36770 -5445
rect 36815 -5565 36935 -5445
rect 36980 -5565 37100 -5445
rect 37155 -5565 37275 -5445
rect 37320 -5565 37440 -5445
rect 37485 -5565 37605 -5445
rect 37650 -5565 37770 -5445
rect 37825 -5565 37945 -5445
rect 37990 -5565 38110 -5445
rect 38155 -5565 38275 -5445
rect 38320 -5565 38440 -5445
rect 38495 -5565 38615 -5445
rect 38660 -5565 38780 -5445
rect 38825 -5565 38945 -5445
rect 38990 -5565 39110 -5445
rect 39165 -5565 39285 -5445
rect 39330 -5565 39450 -5445
rect 39495 -5565 39615 -5445
rect 39660 -5565 39780 -5445
rect 39835 -5565 39955 -5445
rect 40000 -5565 40120 -5445
rect 40165 -5565 40285 -5445
rect 40330 -5565 40450 -5445
rect 40505 -5565 40625 -5445
rect 40670 -5565 40790 -5445
rect 40835 -5565 40955 -5445
rect 41000 -5565 41120 -5445
rect 41175 -5565 41295 -5445
rect 41340 -5565 41460 -5445
rect 41505 -5565 41625 -5445
rect 41670 -5565 41790 -5445
rect 41845 -5565 41965 -5445
rect 36485 -5730 36605 -5610
rect 36650 -5730 36770 -5610
rect 36815 -5730 36935 -5610
rect 36980 -5730 37100 -5610
rect 37155 -5730 37275 -5610
rect 37320 -5730 37440 -5610
rect 37485 -5730 37605 -5610
rect 37650 -5730 37770 -5610
rect 37825 -5730 37945 -5610
rect 37990 -5730 38110 -5610
rect 38155 -5730 38275 -5610
rect 38320 -5730 38440 -5610
rect 38495 -5730 38615 -5610
rect 38660 -5730 38780 -5610
rect 38825 -5730 38945 -5610
rect 38990 -5730 39110 -5610
rect 39165 -5730 39285 -5610
rect 39330 -5730 39450 -5610
rect 39495 -5730 39615 -5610
rect 39660 -5730 39780 -5610
rect 39835 -5730 39955 -5610
rect 40000 -5730 40120 -5610
rect 40165 -5730 40285 -5610
rect 40330 -5730 40450 -5610
rect 40505 -5730 40625 -5610
rect 40670 -5730 40790 -5610
rect 40835 -5730 40955 -5610
rect 41000 -5730 41120 -5610
rect 41175 -5730 41295 -5610
rect 41340 -5730 41460 -5610
rect 41505 -5730 41625 -5610
rect 41670 -5730 41790 -5610
rect 41845 -5730 41965 -5610
rect 36485 -5905 36605 -5785
rect 36650 -5905 36770 -5785
rect 36815 -5905 36935 -5785
rect 36980 -5905 37100 -5785
rect 37155 -5905 37275 -5785
rect 37320 -5905 37440 -5785
rect 37485 -5905 37605 -5785
rect 37650 -5905 37770 -5785
rect 37825 -5905 37945 -5785
rect 37990 -5905 38110 -5785
rect 38155 -5905 38275 -5785
rect 38320 -5905 38440 -5785
rect 38495 -5905 38615 -5785
rect 38660 -5905 38780 -5785
rect 38825 -5905 38945 -5785
rect 38990 -5905 39110 -5785
rect 39165 -5905 39285 -5785
rect 39330 -5905 39450 -5785
rect 39495 -5905 39615 -5785
rect 39660 -5905 39780 -5785
rect 39835 -5905 39955 -5785
rect 40000 -5905 40120 -5785
rect 40165 -5905 40285 -5785
rect 40330 -5905 40450 -5785
rect 40505 -5905 40625 -5785
rect 40670 -5905 40790 -5785
rect 40835 -5905 40955 -5785
rect 41000 -5905 41120 -5785
rect 41175 -5905 41295 -5785
rect 41340 -5905 41460 -5785
rect 41505 -5905 41625 -5785
rect 41670 -5905 41790 -5785
rect 41845 -5905 41965 -5785
rect 36485 -6070 36605 -5950
rect 36650 -6070 36770 -5950
rect 36815 -6070 36935 -5950
rect 36980 -6070 37100 -5950
rect 37155 -6070 37275 -5950
rect 37320 -6070 37440 -5950
rect 37485 -6070 37605 -5950
rect 37650 -6070 37770 -5950
rect 37825 -6070 37945 -5950
rect 37990 -6070 38110 -5950
rect 38155 -6070 38275 -5950
rect 38320 -6070 38440 -5950
rect 38495 -6070 38615 -5950
rect 38660 -6070 38780 -5950
rect 38825 -6070 38945 -5950
rect 38990 -6070 39110 -5950
rect 39165 -6070 39285 -5950
rect 39330 -6070 39450 -5950
rect 39495 -6070 39615 -5950
rect 39660 -6070 39780 -5950
rect 39835 -6070 39955 -5950
rect 40000 -6070 40120 -5950
rect 40165 -6070 40285 -5950
rect 40330 -6070 40450 -5950
rect 40505 -6070 40625 -5950
rect 40670 -6070 40790 -5950
rect 40835 -6070 40955 -5950
rect 41000 -6070 41120 -5950
rect 41175 -6070 41295 -5950
rect 41340 -6070 41460 -5950
rect 41505 -6070 41625 -5950
rect 41670 -6070 41790 -5950
rect 41845 -6070 41965 -5950
rect 36485 -6235 36605 -6115
rect 36650 -6235 36770 -6115
rect 36815 -6235 36935 -6115
rect 36980 -6235 37100 -6115
rect 37155 -6235 37275 -6115
rect 37320 -6235 37440 -6115
rect 37485 -6235 37605 -6115
rect 37650 -6235 37770 -6115
rect 37825 -6235 37945 -6115
rect 37990 -6235 38110 -6115
rect 38155 -6235 38275 -6115
rect 38320 -6235 38440 -6115
rect 38495 -6235 38615 -6115
rect 38660 -6235 38780 -6115
rect 38825 -6235 38945 -6115
rect 38990 -6235 39110 -6115
rect 39165 -6235 39285 -6115
rect 39330 -6235 39450 -6115
rect 39495 -6235 39615 -6115
rect 39660 -6235 39780 -6115
rect 39835 -6235 39955 -6115
rect 40000 -6235 40120 -6115
rect 40165 -6235 40285 -6115
rect 40330 -6235 40450 -6115
rect 40505 -6235 40625 -6115
rect 40670 -6235 40790 -6115
rect 40835 -6235 40955 -6115
rect 41000 -6235 41120 -6115
rect 41175 -6235 41295 -6115
rect 41340 -6235 41460 -6115
rect 41505 -6235 41625 -6115
rect 41670 -6235 41790 -6115
rect 41845 -6235 41965 -6115
rect 36485 -6400 36605 -6280
rect 36650 -6400 36770 -6280
rect 36815 -6400 36935 -6280
rect 36980 -6400 37100 -6280
rect 37155 -6400 37275 -6280
rect 37320 -6400 37440 -6280
rect 37485 -6400 37605 -6280
rect 37650 -6400 37770 -6280
rect 37825 -6400 37945 -6280
rect 37990 -6400 38110 -6280
rect 38155 -6400 38275 -6280
rect 38320 -6400 38440 -6280
rect 38495 -6400 38615 -6280
rect 38660 -6400 38780 -6280
rect 38825 -6400 38945 -6280
rect 38990 -6400 39110 -6280
rect 39165 -6400 39285 -6280
rect 39330 -6400 39450 -6280
rect 39495 -6400 39615 -6280
rect 39660 -6400 39780 -6280
rect 39835 -6400 39955 -6280
rect 40000 -6400 40120 -6280
rect 40165 -6400 40285 -6280
rect 40330 -6400 40450 -6280
rect 40505 -6400 40625 -6280
rect 40670 -6400 40790 -6280
rect 40835 -6400 40955 -6280
rect 41000 -6400 41120 -6280
rect 41175 -6400 41295 -6280
rect 41340 -6400 41460 -6280
rect 41505 -6400 41625 -6280
rect 41670 -6400 41790 -6280
rect 41845 -6400 41965 -6280
rect 36485 -6575 36605 -6455
rect 36650 -6575 36770 -6455
rect 36815 -6575 36935 -6455
rect 36980 -6575 37100 -6455
rect 37155 -6575 37275 -6455
rect 37320 -6575 37440 -6455
rect 37485 -6575 37605 -6455
rect 37650 -6575 37770 -6455
rect 37825 -6575 37945 -6455
rect 37990 -6575 38110 -6455
rect 38155 -6575 38275 -6455
rect 38320 -6575 38440 -6455
rect 38495 -6575 38615 -6455
rect 38660 -6575 38780 -6455
rect 38825 -6575 38945 -6455
rect 38990 -6575 39110 -6455
rect 39165 -6575 39285 -6455
rect 39330 -6575 39450 -6455
rect 39495 -6575 39615 -6455
rect 39660 -6575 39780 -6455
rect 39835 -6575 39955 -6455
rect 40000 -6575 40120 -6455
rect 40165 -6575 40285 -6455
rect 40330 -6575 40450 -6455
rect 40505 -6575 40625 -6455
rect 40670 -6575 40790 -6455
rect 40835 -6575 40955 -6455
rect 41000 -6575 41120 -6455
rect 41175 -6575 41295 -6455
rect 41340 -6575 41460 -6455
rect 41505 -6575 41625 -6455
rect 41670 -6575 41790 -6455
rect 41845 -6575 41965 -6455
rect 36485 -6740 36605 -6620
rect 36650 -6740 36770 -6620
rect 36815 -6740 36935 -6620
rect 36980 -6740 37100 -6620
rect 37155 -6740 37275 -6620
rect 37320 -6740 37440 -6620
rect 37485 -6740 37605 -6620
rect 37650 -6740 37770 -6620
rect 37825 -6740 37945 -6620
rect 37990 -6740 38110 -6620
rect 38155 -6740 38275 -6620
rect 38320 -6740 38440 -6620
rect 38495 -6740 38615 -6620
rect 38660 -6740 38780 -6620
rect 38825 -6740 38945 -6620
rect 38990 -6740 39110 -6620
rect 39165 -6740 39285 -6620
rect 39330 -6740 39450 -6620
rect 39495 -6740 39615 -6620
rect 39660 -6740 39780 -6620
rect 39835 -6740 39955 -6620
rect 40000 -6740 40120 -6620
rect 40165 -6740 40285 -6620
rect 40330 -6740 40450 -6620
rect 40505 -6740 40625 -6620
rect 40670 -6740 40790 -6620
rect 40835 -6740 40955 -6620
rect 41000 -6740 41120 -6620
rect 41175 -6740 41295 -6620
rect 41340 -6740 41460 -6620
rect 41505 -6740 41625 -6620
rect 41670 -6740 41790 -6620
rect 41845 -6740 41965 -6620
rect 36485 -6905 36605 -6785
rect 36650 -6905 36770 -6785
rect 36815 -6905 36935 -6785
rect 36980 -6905 37100 -6785
rect 37155 -6905 37275 -6785
rect 37320 -6905 37440 -6785
rect 37485 -6905 37605 -6785
rect 37650 -6905 37770 -6785
rect 37825 -6905 37945 -6785
rect 37990 -6905 38110 -6785
rect 38155 -6905 38275 -6785
rect 38320 -6905 38440 -6785
rect 38495 -6905 38615 -6785
rect 38660 -6905 38780 -6785
rect 38825 -6905 38945 -6785
rect 38990 -6905 39110 -6785
rect 39165 -6905 39285 -6785
rect 39330 -6905 39450 -6785
rect 39495 -6905 39615 -6785
rect 39660 -6905 39780 -6785
rect 39835 -6905 39955 -6785
rect 40000 -6905 40120 -6785
rect 40165 -6905 40285 -6785
rect 40330 -6905 40450 -6785
rect 40505 -6905 40625 -6785
rect 40670 -6905 40790 -6785
rect 40835 -6905 40955 -6785
rect 41000 -6905 41120 -6785
rect 41175 -6905 41295 -6785
rect 41340 -6905 41460 -6785
rect 41505 -6905 41625 -6785
rect 41670 -6905 41790 -6785
rect 41845 -6905 41965 -6785
rect 36485 -7070 36605 -6950
rect 36650 -7070 36770 -6950
rect 36815 -7070 36935 -6950
rect 36980 -7070 37100 -6950
rect 37155 -7070 37275 -6950
rect 37320 -7070 37440 -6950
rect 37485 -7070 37605 -6950
rect 37650 -7070 37770 -6950
rect 37825 -7070 37945 -6950
rect 37990 -7070 38110 -6950
rect 38155 -7070 38275 -6950
rect 38320 -7070 38440 -6950
rect 38495 -7070 38615 -6950
rect 38660 -7070 38780 -6950
rect 38825 -7070 38945 -6950
rect 38990 -7070 39110 -6950
rect 39165 -7070 39285 -6950
rect 39330 -7070 39450 -6950
rect 39495 -7070 39615 -6950
rect 39660 -7070 39780 -6950
rect 39835 -7070 39955 -6950
rect 40000 -7070 40120 -6950
rect 40165 -7070 40285 -6950
rect 40330 -7070 40450 -6950
rect 40505 -7070 40625 -6950
rect 40670 -7070 40790 -6950
rect 40835 -7070 40955 -6950
rect 41000 -7070 41120 -6950
rect 41175 -7070 41295 -6950
rect 41340 -7070 41460 -6950
rect 41505 -7070 41625 -6950
rect 41670 -7070 41790 -6950
rect 41845 -7070 41965 -6950
rect 36485 -7245 36605 -7125
rect 36650 -7245 36770 -7125
rect 36815 -7245 36935 -7125
rect 36980 -7245 37100 -7125
rect 37155 -7245 37275 -7125
rect 37320 -7245 37440 -7125
rect 37485 -7245 37605 -7125
rect 37650 -7245 37770 -7125
rect 37825 -7245 37945 -7125
rect 37990 -7245 38110 -7125
rect 38155 -7245 38275 -7125
rect 38320 -7245 38440 -7125
rect 38495 -7245 38615 -7125
rect 38660 -7245 38780 -7125
rect 38825 -7245 38945 -7125
rect 38990 -7245 39110 -7125
rect 39165 -7245 39285 -7125
rect 39330 -7245 39450 -7125
rect 39495 -7245 39615 -7125
rect 39660 -7245 39780 -7125
rect 39835 -7245 39955 -7125
rect 40000 -7245 40120 -7125
rect 40165 -7245 40285 -7125
rect 40330 -7245 40450 -7125
rect 40505 -7245 40625 -7125
rect 40670 -7245 40790 -7125
rect 40835 -7245 40955 -7125
rect 41000 -7245 41120 -7125
rect 41175 -7245 41295 -7125
rect 41340 -7245 41460 -7125
rect 41505 -7245 41625 -7125
rect 41670 -7245 41790 -7125
rect 41845 -7245 41965 -7125
rect 36485 -7410 36605 -7290
rect 36650 -7410 36770 -7290
rect 36815 -7410 36935 -7290
rect 36980 -7410 37100 -7290
rect 37155 -7410 37275 -7290
rect 37320 -7410 37440 -7290
rect 37485 -7410 37605 -7290
rect 37650 -7410 37770 -7290
rect 37825 -7410 37945 -7290
rect 37990 -7410 38110 -7290
rect 38155 -7410 38275 -7290
rect 38320 -7410 38440 -7290
rect 38495 -7410 38615 -7290
rect 38660 -7410 38780 -7290
rect 38825 -7410 38945 -7290
rect 38990 -7410 39110 -7290
rect 39165 -7410 39285 -7290
rect 39330 -7410 39450 -7290
rect 39495 -7410 39615 -7290
rect 39660 -7410 39780 -7290
rect 39835 -7410 39955 -7290
rect 40000 -7410 40120 -7290
rect 40165 -7410 40285 -7290
rect 40330 -7410 40450 -7290
rect 40505 -7410 40625 -7290
rect 40670 -7410 40790 -7290
rect 40835 -7410 40955 -7290
rect 41000 -7410 41120 -7290
rect 41175 -7410 41295 -7290
rect 41340 -7410 41460 -7290
rect 41505 -7410 41625 -7290
rect 41670 -7410 41790 -7290
rect 41845 -7410 41965 -7290
rect 36485 -7575 36605 -7455
rect 36650 -7575 36770 -7455
rect 36815 -7575 36935 -7455
rect 36980 -7575 37100 -7455
rect 37155 -7575 37275 -7455
rect 37320 -7575 37440 -7455
rect 37485 -7575 37605 -7455
rect 37650 -7575 37770 -7455
rect 37825 -7575 37945 -7455
rect 37990 -7575 38110 -7455
rect 38155 -7575 38275 -7455
rect 38320 -7575 38440 -7455
rect 38495 -7575 38615 -7455
rect 38660 -7575 38780 -7455
rect 38825 -7575 38945 -7455
rect 38990 -7575 39110 -7455
rect 39165 -7575 39285 -7455
rect 39330 -7575 39450 -7455
rect 39495 -7575 39615 -7455
rect 39660 -7575 39780 -7455
rect 39835 -7575 39955 -7455
rect 40000 -7575 40120 -7455
rect 40165 -7575 40285 -7455
rect 40330 -7575 40450 -7455
rect 40505 -7575 40625 -7455
rect 40670 -7575 40790 -7455
rect 40835 -7575 40955 -7455
rect 41000 -7575 41120 -7455
rect 41175 -7575 41295 -7455
rect 41340 -7575 41460 -7455
rect 41505 -7575 41625 -7455
rect 41670 -7575 41790 -7455
rect 41845 -7575 41965 -7455
rect 36485 -7740 36605 -7620
rect 36650 -7740 36770 -7620
rect 36815 -7740 36935 -7620
rect 36980 -7740 37100 -7620
rect 37155 -7740 37275 -7620
rect 37320 -7740 37440 -7620
rect 37485 -7740 37605 -7620
rect 37650 -7740 37770 -7620
rect 37825 -7740 37945 -7620
rect 37990 -7740 38110 -7620
rect 38155 -7740 38275 -7620
rect 38320 -7740 38440 -7620
rect 38495 -7740 38615 -7620
rect 38660 -7740 38780 -7620
rect 38825 -7740 38945 -7620
rect 38990 -7740 39110 -7620
rect 39165 -7740 39285 -7620
rect 39330 -7740 39450 -7620
rect 39495 -7740 39615 -7620
rect 39660 -7740 39780 -7620
rect 39835 -7740 39955 -7620
rect 40000 -7740 40120 -7620
rect 40165 -7740 40285 -7620
rect 40330 -7740 40450 -7620
rect 40505 -7740 40625 -7620
rect 40670 -7740 40790 -7620
rect 40835 -7740 40955 -7620
rect 41000 -7740 41120 -7620
rect 41175 -7740 41295 -7620
rect 41340 -7740 41460 -7620
rect 41505 -7740 41625 -7620
rect 41670 -7740 41790 -7620
rect 41845 -7740 41965 -7620
rect 36485 -7915 36605 -7795
rect 36650 -7915 36770 -7795
rect 36815 -7915 36935 -7795
rect 36980 -7915 37100 -7795
rect 37155 -7915 37275 -7795
rect 37320 -7915 37440 -7795
rect 37485 -7915 37605 -7795
rect 37650 -7915 37770 -7795
rect 37825 -7915 37945 -7795
rect 37990 -7915 38110 -7795
rect 38155 -7915 38275 -7795
rect 38320 -7915 38440 -7795
rect 38495 -7915 38615 -7795
rect 38660 -7915 38780 -7795
rect 38825 -7915 38945 -7795
rect 38990 -7915 39110 -7795
rect 39165 -7915 39285 -7795
rect 39330 -7915 39450 -7795
rect 39495 -7915 39615 -7795
rect 39660 -7915 39780 -7795
rect 39835 -7915 39955 -7795
rect 40000 -7915 40120 -7795
rect 40165 -7915 40285 -7795
rect 40330 -7915 40450 -7795
rect 40505 -7915 40625 -7795
rect 40670 -7915 40790 -7795
rect 40835 -7915 40955 -7795
rect 41000 -7915 41120 -7795
rect 41175 -7915 41295 -7795
rect 41340 -7915 41460 -7795
rect 41505 -7915 41625 -7795
rect 41670 -7915 41790 -7795
rect 41845 -7915 41965 -7795
rect 36485 -8080 36605 -7960
rect 36650 -8080 36770 -7960
rect 36815 -8080 36935 -7960
rect 36980 -8080 37100 -7960
rect 37155 -8080 37275 -7960
rect 37320 -8080 37440 -7960
rect 37485 -8080 37605 -7960
rect 37650 -8080 37770 -7960
rect 37825 -8080 37945 -7960
rect 37990 -8080 38110 -7960
rect 38155 -8080 38275 -7960
rect 38320 -8080 38440 -7960
rect 38495 -8080 38615 -7960
rect 38660 -8080 38780 -7960
rect 38825 -8080 38945 -7960
rect 38990 -8080 39110 -7960
rect 39165 -8080 39285 -7960
rect 39330 -8080 39450 -7960
rect 39495 -8080 39615 -7960
rect 39660 -8080 39780 -7960
rect 39835 -8080 39955 -7960
rect 40000 -8080 40120 -7960
rect 40165 -8080 40285 -7960
rect 40330 -8080 40450 -7960
rect 40505 -8080 40625 -7960
rect 40670 -8080 40790 -7960
rect 40835 -8080 40955 -7960
rect 41000 -8080 41120 -7960
rect 41175 -8080 41295 -7960
rect 41340 -8080 41460 -7960
rect 41505 -8080 41625 -7960
rect 41670 -8080 41790 -7960
rect 41845 -8080 41965 -7960
rect 36485 -8245 36605 -8125
rect 36650 -8245 36770 -8125
rect 36815 -8245 36935 -8125
rect 36980 -8245 37100 -8125
rect 37155 -8245 37275 -8125
rect 37320 -8245 37440 -8125
rect 37485 -8245 37605 -8125
rect 37650 -8245 37770 -8125
rect 37825 -8245 37945 -8125
rect 37990 -8245 38110 -8125
rect 38155 -8245 38275 -8125
rect 38320 -8245 38440 -8125
rect 38495 -8245 38615 -8125
rect 38660 -8245 38780 -8125
rect 38825 -8245 38945 -8125
rect 38990 -8245 39110 -8125
rect 39165 -8245 39285 -8125
rect 39330 -8245 39450 -8125
rect 39495 -8245 39615 -8125
rect 39660 -8245 39780 -8125
rect 39835 -8245 39955 -8125
rect 40000 -8245 40120 -8125
rect 40165 -8245 40285 -8125
rect 40330 -8245 40450 -8125
rect 40505 -8245 40625 -8125
rect 40670 -8245 40790 -8125
rect 40835 -8245 40955 -8125
rect 41000 -8245 41120 -8125
rect 41175 -8245 41295 -8125
rect 41340 -8245 41460 -8125
rect 41505 -8245 41625 -8125
rect 41670 -8245 41790 -8125
rect 41845 -8245 41965 -8125
rect 36485 -8410 36605 -8290
rect 36650 -8410 36770 -8290
rect 36815 -8410 36935 -8290
rect 36980 -8410 37100 -8290
rect 37155 -8410 37275 -8290
rect 37320 -8410 37440 -8290
rect 37485 -8410 37605 -8290
rect 37650 -8410 37770 -8290
rect 37825 -8410 37945 -8290
rect 37990 -8410 38110 -8290
rect 38155 -8410 38275 -8290
rect 38320 -8410 38440 -8290
rect 38495 -8410 38615 -8290
rect 38660 -8410 38780 -8290
rect 38825 -8410 38945 -8290
rect 38990 -8410 39110 -8290
rect 39165 -8410 39285 -8290
rect 39330 -8410 39450 -8290
rect 39495 -8410 39615 -8290
rect 39660 -8410 39780 -8290
rect 39835 -8410 39955 -8290
rect 40000 -8410 40120 -8290
rect 40165 -8410 40285 -8290
rect 40330 -8410 40450 -8290
rect 40505 -8410 40625 -8290
rect 40670 -8410 40790 -8290
rect 40835 -8410 40955 -8290
rect 41000 -8410 41120 -8290
rect 41175 -8410 41295 -8290
rect 41340 -8410 41460 -8290
rect 41505 -8410 41625 -8290
rect 41670 -8410 41790 -8290
rect 41845 -8410 41965 -8290
rect 36485 -8585 36605 -8465
rect 36650 -8585 36770 -8465
rect 36815 -8585 36935 -8465
rect 36980 -8585 37100 -8465
rect 37155 -8585 37275 -8465
rect 37320 -8585 37440 -8465
rect 37485 -8585 37605 -8465
rect 37650 -8585 37770 -8465
rect 37825 -8585 37945 -8465
rect 37990 -8585 38110 -8465
rect 38155 -8585 38275 -8465
rect 38320 -8585 38440 -8465
rect 38495 -8585 38615 -8465
rect 38660 -8585 38780 -8465
rect 38825 -8585 38945 -8465
rect 38990 -8585 39110 -8465
rect 39165 -8585 39285 -8465
rect 39330 -8585 39450 -8465
rect 39495 -8585 39615 -8465
rect 39660 -8585 39780 -8465
rect 39835 -8585 39955 -8465
rect 40000 -8585 40120 -8465
rect 40165 -8585 40285 -8465
rect 40330 -8585 40450 -8465
rect 40505 -8585 40625 -8465
rect 40670 -8585 40790 -8465
rect 40835 -8585 40955 -8465
rect 41000 -8585 41120 -8465
rect 41175 -8585 41295 -8465
rect 41340 -8585 41460 -8465
rect 41505 -8585 41625 -8465
rect 41670 -8585 41790 -8465
rect 41845 -8585 41965 -8465
rect 36485 -8750 36605 -8630
rect 36650 -8750 36770 -8630
rect 36815 -8750 36935 -8630
rect 36980 -8750 37100 -8630
rect 37155 -8750 37275 -8630
rect 37320 -8750 37440 -8630
rect 37485 -8750 37605 -8630
rect 37650 -8750 37770 -8630
rect 37825 -8750 37945 -8630
rect 37990 -8750 38110 -8630
rect 38155 -8750 38275 -8630
rect 38320 -8750 38440 -8630
rect 38495 -8750 38615 -8630
rect 38660 -8750 38780 -8630
rect 38825 -8750 38945 -8630
rect 38990 -8750 39110 -8630
rect 39165 -8750 39285 -8630
rect 39330 -8750 39450 -8630
rect 39495 -8750 39615 -8630
rect 39660 -8750 39780 -8630
rect 39835 -8750 39955 -8630
rect 40000 -8750 40120 -8630
rect 40165 -8750 40285 -8630
rect 40330 -8750 40450 -8630
rect 40505 -8750 40625 -8630
rect 40670 -8750 40790 -8630
rect 40835 -8750 40955 -8630
rect 41000 -8750 41120 -8630
rect 41175 -8750 41295 -8630
rect 41340 -8750 41460 -8630
rect 41505 -8750 41625 -8630
rect 41670 -8750 41790 -8630
rect 41845 -8750 41965 -8630
rect 36485 -8915 36605 -8795
rect 36650 -8915 36770 -8795
rect 36815 -8915 36935 -8795
rect 36980 -8915 37100 -8795
rect 37155 -8915 37275 -8795
rect 37320 -8915 37440 -8795
rect 37485 -8915 37605 -8795
rect 37650 -8915 37770 -8795
rect 37825 -8915 37945 -8795
rect 37990 -8915 38110 -8795
rect 38155 -8915 38275 -8795
rect 38320 -8915 38440 -8795
rect 38495 -8915 38615 -8795
rect 38660 -8915 38780 -8795
rect 38825 -8915 38945 -8795
rect 38990 -8915 39110 -8795
rect 39165 -8915 39285 -8795
rect 39330 -8915 39450 -8795
rect 39495 -8915 39615 -8795
rect 39660 -8915 39780 -8795
rect 39835 -8915 39955 -8795
rect 40000 -8915 40120 -8795
rect 40165 -8915 40285 -8795
rect 40330 -8915 40450 -8795
rect 40505 -8915 40625 -8795
rect 40670 -8915 40790 -8795
rect 40835 -8915 40955 -8795
rect 41000 -8915 41120 -8795
rect 41175 -8915 41295 -8795
rect 41340 -8915 41460 -8795
rect 41505 -8915 41625 -8795
rect 41670 -8915 41790 -8795
rect 41845 -8915 41965 -8795
rect 36485 -9080 36605 -8960
rect 36650 -9080 36770 -8960
rect 36815 -9080 36935 -8960
rect 36980 -9080 37100 -8960
rect 37155 -9080 37275 -8960
rect 37320 -9080 37440 -8960
rect 37485 -9080 37605 -8960
rect 37650 -9080 37770 -8960
rect 37825 -9080 37945 -8960
rect 37990 -9080 38110 -8960
rect 38155 -9080 38275 -8960
rect 38320 -9080 38440 -8960
rect 38495 -9080 38615 -8960
rect 38660 -9080 38780 -8960
rect 38825 -9080 38945 -8960
rect 38990 -9080 39110 -8960
rect 39165 -9080 39285 -8960
rect 39330 -9080 39450 -8960
rect 39495 -9080 39615 -8960
rect 39660 -9080 39780 -8960
rect 39835 -9080 39955 -8960
rect 40000 -9080 40120 -8960
rect 40165 -9080 40285 -8960
rect 40330 -9080 40450 -8960
rect 40505 -9080 40625 -8960
rect 40670 -9080 40790 -8960
rect 40835 -9080 40955 -8960
rect 41000 -9080 41120 -8960
rect 41175 -9080 41295 -8960
rect 41340 -9080 41460 -8960
rect 41505 -9080 41625 -8960
rect 41670 -9080 41790 -8960
rect 41845 -9080 41965 -8960
rect 36485 -9255 36605 -9135
rect 36650 -9255 36770 -9135
rect 36815 -9255 36935 -9135
rect 36980 -9255 37100 -9135
rect 37155 -9255 37275 -9135
rect 37320 -9255 37440 -9135
rect 37485 -9255 37605 -9135
rect 37650 -9255 37770 -9135
rect 37825 -9255 37945 -9135
rect 37990 -9255 38110 -9135
rect 38155 -9255 38275 -9135
rect 38320 -9255 38440 -9135
rect 38495 -9255 38615 -9135
rect 38660 -9255 38780 -9135
rect 38825 -9255 38945 -9135
rect 38990 -9255 39110 -9135
rect 39165 -9255 39285 -9135
rect 39330 -9255 39450 -9135
rect 39495 -9255 39615 -9135
rect 39660 -9255 39780 -9135
rect 39835 -9255 39955 -9135
rect 40000 -9255 40120 -9135
rect 40165 -9255 40285 -9135
rect 40330 -9255 40450 -9135
rect 40505 -9255 40625 -9135
rect 40670 -9255 40790 -9135
rect 40835 -9255 40955 -9135
rect 41000 -9255 41120 -9135
rect 41175 -9255 41295 -9135
rect 41340 -9255 41460 -9135
rect 41505 -9255 41625 -9135
rect 41670 -9255 41790 -9135
rect 41845 -9255 41965 -9135
rect 36485 -9420 36605 -9300
rect 36650 -9420 36770 -9300
rect 36815 -9420 36935 -9300
rect 36980 -9420 37100 -9300
rect 37155 -9420 37275 -9300
rect 37320 -9420 37440 -9300
rect 37485 -9420 37605 -9300
rect 37650 -9420 37770 -9300
rect 37825 -9420 37945 -9300
rect 37990 -9420 38110 -9300
rect 38155 -9420 38275 -9300
rect 38320 -9420 38440 -9300
rect 38495 -9420 38615 -9300
rect 38660 -9420 38780 -9300
rect 38825 -9420 38945 -9300
rect 38990 -9420 39110 -9300
rect 39165 -9420 39285 -9300
rect 39330 -9420 39450 -9300
rect 39495 -9420 39615 -9300
rect 39660 -9420 39780 -9300
rect 39835 -9420 39955 -9300
rect 40000 -9420 40120 -9300
rect 40165 -9420 40285 -9300
rect 40330 -9420 40450 -9300
rect 40505 -9420 40625 -9300
rect 40670 -9420 40790 -9300
rect 40835 -9420 40955 -9300
rect 41000 -9420 41120 -9300
rect 41175 -9420 41295 -9300
rect 41340 -9420 41460 -9300
rect 41505 -9420 41625 -9300
rect 41670 -9420 41790 -9300
rect 41845 -9420 41965 -9300
rect 36485 -9585 36605 -9465
rect 36650 -9585 36770 -9465
rect 36815 -9585 36935 -9465
rect 36980 -9585 37100 -9465
rect 37155 -9585 37275 -9465
rect 37320 -9585 37440 -9465
rect 37485 -9585 37605 -9465
rect 37650 -9585 37770 -9465
rect 37825 -9585 37945 -9465
rect 37990 -9585 38110 -9465
rect 38155 -9585 38275 -9465
rect 38320 -9585 38440 -9465
rect 38495 -9585 38615 -9465
rect 38660 -9585 38780 -9465
rect 38825 -9585 38945 -9465
rect 38990 -9585 39110 -9465
rect 39165 -9585 39285 -9465
rect 39330 -9585 39450 -9465
rect 39495 -9585 39615 -9465
rect 39660 -9585 39780 -9465
rect 39835 -9585 39955 -9465
rect 40000 -9585 40120 -9465
rect 40165 -9585 40285 -9465
rect 40330 -9585 40450 -9465
rect 40505 -9585 40625 -9465
rect 40670 -9585 40790 -9465
rect 40835 -9585 40955 -9465
rect 41000 -9585 41120 -9465
rect 41175 -9585 41295 -9465
rect 41340 -9585 41460 -9465
rect 41505 -9585 41625 -9465
rect 41670 -9585 41790 -9465
rect 41845 -9585 41965 -9465
rect 36485 -9750 36605 -9630
rect 36650 -9750 36770 -9630
rect 36815 -9750 36935 -9630
rect 36980 -9750 37100 -9630
rect 37155 -9750 37275 -9630
rect 37320 -9750 37440 -9630
rect 37485 -9750 37605 -9630
rect 37650 -9750 37770 -9630
rect 37825 -9750 37945 -9630
rect 37990 -9750 38110 -9630
rect 38155 -9750 38275 -9630
rect 38320 -9750 38440 -9630
rect 38495 -9750 38615 -9630
rect 38660 -9750 38780 -9630
rect 38825 -9750 38945 -9630
rect 38990 -9750 39110 -9630
rect 39165 -9750 39285 -9630
rect 39330 -9750 39450 -9630
rect 39495 -9750 39615 -9630
rect 39660 -9750 39780 -9630
rect 39835 -9750 39955 -9630
rect 40000 -9750 40120 -9630
rect 40165 -9750 40285 -9630
rect 40330 -9750 40450 -9630
rect 40505 -9750 40625 -9630
rect 40670 -9750 40790 -9630
rect 40835 -9750 40955 -9630
rect 41000 -9750 41120 -9630
rect 41175 -9750 41295 -9630
rect 41340 -9750 41460 -9630
rect 41505 -9750 41625 -9630
rect 41670 -9750 41790 -9630
rect 41845 -9750 41965 -9630
rect 42175 -4390 42295 -4270
rect 42340 -4390 42460 -4270
rect 42505 -4390 42625 -4270
rect 42670 -4390 42790 -4270
rect 42845 -4390 42965 -4270
rect 43010 -4390 43130 -4270
rect 43175 -4390 43295 -4270
rect 43340 -4390 43460 -4270
rect 43515 -4390 43635 -4270
rect 43680 -4390 43800 -4270
rect 43845 -4390 43965 -4270
rect 44010 -4390 44130 -4270
rect 44185 -4390 44305 -4270
rect 44350 -4390 44470 -4270
rect 44515 -4390 44635 -4270
rect 44680 -4390 44800 -4270
rect 44855 -4390 44975 -4270
rect 45020 -4390 45140 -4270
rect 45185 -4390 45305 -4270
rect 45350 -4390 45470 -4270
rect 45525 -4390 45645 -4270
rect 45690 -4390 45810 -4270
rect 45855 -4390 45975 -4270
rect 46020 -4390 46140 -4270
rect 46195 -4390 46315 -4270
rect 46360 -4390 46480 -4270
rect 46525 -4390 46645 -4270
rect 46690 -4390 46810 -4270
rect 46865 -4390 46985 -4270
rect 47030 -4390 47150 -4270
rect 47195 -4390 47315 -4270
rect 47360 -4390 47480 -4270
rect 47535 -4390 47655 -4270
rect 42175 -4565 42295 -4445
rect 42340 -4565 42460 -4445
rect 42505 -4565 42625 -4445
rect 42670 -4565 42790 -4445
rect 42845 -4565 42965 -4445
rect 43010 -4565 43130 -4445
rect 43175 -4565 43295 -4445
rect 43340 -4565 43460 -4445
rect 43515 -4565 43635 -4445
rect 43680 -4565 43800 -4445
rect 43845 -4565 43965 -4445
rect 44010 -4565 44130 -4445
rect 44185 -4565 44305 -4445
rect 44350 -4565 44470 -4445
rect 44515 -4565 44635 -4445
rect 44680 -4565 44800 -4445
rect 44855 -4565 44975 -4445
rect 45020 -4565 45140 -4445
rect 45185 -4565 45305 -4445
rect 45350 -4565 45470 -4445
rect 45525 -4565 45645 -4445
rect 45690 -4565 45810 -4445
rect 45855 -4565 45975 -4445
rect 46020 -4565 46140 -4445
rect 46195 -4565 46315 -4445
rect 46360 -4565 46480 -4445
rect 46525 -4565 46645 -4445
rect 46690 -4565 46810 -4445
rect 46865 -4565 46985 -4445
rect 47030 -4565 47150 -4445
rect 47195 -4565 47315 -4445
rect 47360 -4565 47480 -4445
rect 47535 -4565 47655 -4445
rect 42175 -4730 42295 -4610
rect 42340 -4730 42460 -4610
rect 42505 -4730 42625 -4610
rect 42670 -4730 42790 -4610
rect 42845 -4730 42965 -4610
rect 43010 -4730 43130 -4610
rect 43175 -4730 43295 -4610
rect 43340 -4730 43460 -4610
rect 43515 -4730 43635 -4610
rect 43680 -4730 43800 -4610
rect 43845 -4730 43965 -4610
rect 44010 -4730 44130 -4610
rect 44185 -4730 44305 -4610
rect 44350 -4730 44470 -4610
rect 44515 -4730 44635 -4610
rect 44680 -4730 44800 -4610
rect 44855 -4730 44975 -4610
rect 45020 -4730 45140 -4610
rect 45185 -4730 45305 -4610
rect 45350 -4730 45470 -4610
rect 45525 -4730 45645 -4610
rect 45690 -4730 45810 -4610
rect 45855 -4730 45975 -4610
rect 46020 -4730 46140 -4610
rect 46195 -4730 46315 -4610
rect 46360 -4730 46480 -4610
rect 46525 -4730 46645 -4610
rect 46690 -4730 46810 -4610
rect 46865 -4730 46985 -4610
rect 47030 -4730 47150 -4610
rect 47195 -4730 47315 -4610
rect 47360 -4730 47480 -4610
rect 47535 -4730 47655 -4610
rect 42175 -4895 42295 -4775
rect 42340 -4895 42460 -4775
rect 42505 -4895 42625 -4775
rect 42670 -4895 42790 -4775
rect 42845 -4895 42965 -4775
rect 43010 -4895 43130 -4775
rect 43175 -4895 43295 -4775
rect 43340 -4895 43460 -4775
rect 43515 -4895 43635 -4775
rect 43680 -4895 43800 -4775
rect 43845 -4895 43965 -4775
rect 44010 -4895 44130 -4775
rect 44185 -4895 44305 -4775
rect 44350 -4895 44470 -4775
rect 44515 -4895 44635 -4775
rect 44680 -4895 44800 -4775
rect 44855 -4895 44975 -4775
rect 45020 -4895 45140 -4775
rect 45185 -4895 45305 -4775
rect 45350 -4895 45470 -4775
rect 45525 -4895 45645 -4775
rect 45690 -4895 45810 -4775
rect 45855 -4895 45975 -4775
rect 46020 -4895 46140 -4775
rect 46195 -4895 46315 -4775
rect 46360 -4895 46480 -4775
rect 46525 -4895 46645 -4775
rect 46690 -4895 46810 -4775
rect 46865 -4895 46985 -4775
rect 47030 -4895 47150 -4775
rect 47195 -4895 47315 -4775
rect 47360 -4895 47480 -4775
rect 47535 -4895 47655 -4775
rect 42175 -5060 42295 -4940
rect 42340 -5060 42460 -4940
rect 42505 -5060 42625 -4940
rect 42670 -5060 42790 -4940
rect 42845 -5060 42965 -4940
rect 43010 -5060 43130 -4940
rect 43175 -5060 43295 -4940
rect 43340 -5060 43460 -4940
rect 43515 -5060 43635 -4940
rect 43680 -5060 43800 -4940
rect 43845 -5060 43965 -4940
rect 44010 -5060 44130 -4940
rect 44185 -5060 44305 -4940
rect 44350 -5060 44470 -4940
rect 44515 -5060 44635 -4940
rect 44680 -5060 44800 -4940
rect 44855 -5060 44975 -4940
rect 45020 -5060 45140 -4940
rect 45185 -5060 45305 -4940
rect 45350 -5060 45470 -4940
rect 45525 -5060 45645 -4940
rect 45690 -5060 45810 -4940
rect 45855 -5060 45975 -4940
rect 46020 -5060 46140 -4940
rect 46195 -5060 46315 -4940
rect 46360 -5060 46480 -4940
rect 46525 -5060 46645 -4940
rect 46690 -5060 46810 -4940
rect 46865 -5060 46985 -4940
rect 47030 -5060 47150 -4940
rect 47195 -5060 47315 -4940
rect 47360 -5060 47480 -4940
rect 47535 -5060 47655 -4940
rect 42175 -5235 42295 -5115
rect 42340 -5235 42460 -5115
rect 42505 -5235 42625 -5115
rect 42670 -5235 42790 -5115
rect 42845 -5235 42965 -5115
rect 43010 -5235 43130 -5115
rect 43175 -5235 43295 -5115
rect 43340 -5235 43460 -5115
rect 43515 -5235 43635 -5115
rect 43680 -5235 43800 -5115
rect 43845 -5235 43965 -5115
rect 44010 -5235 44130 -5115
rect 44185 -5235 44305 -5115
rect 44350 -5235 44470 -5115
rect 44515 -5235 44635 -5115
rect 44680 -5235 44800 -5115
rect 44855 -5235 44975 -5115
rect 45020 -5235 45140 -5115
rect 45185 -5235 45305 -5115
rect 45350 -5235 45470 -5115
rect 45525 -5235 45645 -5115
rect 45690 -5235 45810 -5115
rect 45855 -5235 45975 -5115
rect 46020 -5235 46140 -5115
rect 46195 -5235 46315 -5115
rect 46360 -5235 46480 -5115
rect 46525 -5235 46645 -5115
rect 46690 -5235 46810 -5115
rect 46865 -5235 46985 -5115
rect 47030 -5235 47150 -5115
rect 47195 -5235 47315 -5115
rect 47360 -5235 47480 -5115
rect 47535 -5235 47655 -5115
rect 42175 -5400 42295 -5280
rect 42340 -5400 42460 -5280
rect 42505 -5400 42625 -5280
rect 42670 -5400 42790 -5280
rect 42845 -5400 42965 -5280
rect 43010 -5400 43130 -5280
rect 43175 -5400 43295 -5280
rect 43340 -5400 43460 -5280
rect 43515 -5400 43635 -5280
rect 43680 -5400 43800 -5280
rect 43845 -5400 43965 -5280
rect 44010 -5400 44130 -5280
rect 44185 -5400 44305 -5280
rect 44350 -5400 44470 -5280
rect 44515 -5400 44635 -5280
rect 44680 -5400 44800 -5280
rect 44855 -5400 44975 -5280
rect 45020 -5400 45140 -5280
rect 45185 -5400 45305 -5280
rect 45350 -5400 45470 -5280
rect 45525 -5400 45645 -5280
rect 45690 -5400 45810 -5280
rect 45855 -5400 45975 -5280
rect 46020 -5400 46140 -5280
rect 46195 -5400 46315 -5280
rect 46360 -5400 46480 -5280
rect 46525 -5400 46645 -5280
rect 46690 -5400 46810 -5280
rect 46865 -5400 46985 -5280
rect 47030 -5400 47150 -5280
rect 47195 -5400 47315 -5280
rect 47360 -5400 47480 -5280
rect 47535 -5400 47655 -5280
rect 42175 -5565 42295 -5445
rect 42340 -5565 42460 -5445
rect 42505 -5565 42625 -5445
rect 42670 -5565 42790 -5445
rect 42845 -5565 42965 -5445
rect 43010 -5565 43130 -5445
rect 43175 -5565 43295 -5445
rect 43340 -5565 43460 -5445
rect 43515 -5565 43635 -5445
rect 43680 -5565 43800 -5445
rect 43845 -5565 43965 -5445
rect 44010 -5565 44130 -5445
rect 44185 -5565 44305 -5445
rect 44350 -5565 44470 -5445
rect 44515 -5565 44635 -5445
rect 44680 -5565 44800 -5445
rect 44855 -5565 44975 -5445
rect 45020 -5565 45140 -5445
rect 45185 -5565 45305 -5445
rect 45350 -5565 45470 -5445
rect 45525 -5565 45645 -5445
rect 45690 -5565 45810 -5445
rect 45855 -5565 45975 -5445
rect 46020 -5565 46140 -5445
rect 46195 -5565 46315 -5445
rect 46360 -5565 46480 -5445
rect 46525 -5565 46645 -5445
rect 46690 -5565 46810 -5445
rect 46865 -5565 46985 -5445
rect 47030 -5565 47150 -5445
rect 47195 -5565 47315 -5445
rect 47360 -5565 47480 -5445
rect 47535 -5565 47655 -5445
rect 42175 -5730 42295 -5610
rect 42340 -5730 42460 -5610
rect 42505 -5730 42625 -5610
rect 42670 -5730 42790 -5610
rect 42845 -5730 42965 -5610
rect 43010 -5730 43130 -5610
rect 43175 -5730 43295 -5610
rect 43340 -5730 43460 -5610
rect 43515 -5730 43635 -5610
rect 43680 -5730 43800 -5610
rect 43845 -5730 43965 -5610
rect 44010 -5730 44130 -5610
rect 44185 -5730 44305 -5610
rect 44350 -5730 44470 -5610
rect 44515 -5730 44635 -5610
rect 44680 -5730 44800 -5610
rect 44855 -5730 44975 -5610
rect 45020 -5730 45140 -5610
rect 45185 -5730 45305 -5610
rect 45350 -5730 45470 -5610
rect 45525 -5730 45645 -5610
rect 45690 -5730 45810 -5610
rect 45855 -5730 45975 -5610
rect 46020 -5730 46140 -5610
rect 46195 -5730 46315 -5610
rect 46360 -5730 46480 -5610
rect 46525 -5730 46645 -5610
rect 46690 -5730 46810 -5610
rect 46865 -5730 46985 -5610
rect 47030 -5730 47150 -5610
rect 47195 -5730 47315 -5610
rect 47360 -5730 47480 -5610
rect 47535 -5730 47655 -5610
rect 42175 -5905 42295 -5785
rect 42340 -5905 42460 -5785
rect 42505 -5905 42625 -5785
rect 42670 -5905 42790 -5785
rect 42845 -5905 42965 -5785
rect 43010 -5905 43130 -5785
rect 43175 -5905 43295 -5785
rect 43340 -5905 43460 -5785
rect 43515 -5905 43635 -5785
rect 43680 -5905 43800 -5785
rect 43845 -5905 43965 -5785
rect 44010 -5905 44130 -5785
rect 44185 -5905 44305 -5785
rect 44350 -5905 44470 -5785
rect 44515 -5905 44635 -5785
rect 44680 -5905 44800 -5785
rect 44855 -5905 44975 -5785
rect 45020 -5905 45140 -5785
rect 45185 -5905 45305 -5785
rect 45350 -5905 45470 -5785
rect 45525 -5905 45645 -5785
rect 45690 -5905 45810 -5785
rect 45855 -5905 45975 -5785
rect 46020 -5905 46140 -5785
rect 46195 -5905 46315 -5785
rect 46360 -5905 46480 -5785
rect 46525 -5905 46645 -5785
rect 46690 -5905 46810 -5785
rect 46865 -5905 46985 -5785
rect 47030 -5905 47150 -5785
rect 47195 -5905 47315 -5785
rect 47360 -5905 47480 -5785
rect 47535 -5905 47655 -5785
rect 42175 -6070 42295 -5950
rect 42340 -6070 42460 -5950
rect 42505 -6070 42625 -5950
rect 42670 -6070 42790 -5950
rect 42845 -6070 42965 -5950
rect 43010 -6070 43130 -5950
rect 43175 -6070 43295 -5950
rect 43340 -6070 43460 -5950
rect 43515 -6070 43635 -5950
rect 43680 -6070 43800 -5950
rect 43845 -6070 43965 -5950
rect 44010 -6070 44130 -5950
rect 44185 -6070 44305 -5950
rect 44350 -6070 44470 -5950
rect 44515 -6070 44635 -5950
rect 44680 -6070 44800 -5950
rect 44855 -6070 44975 -5950
rect 45020 -6070 45140 -5950
rect 45185 -6070 45305 -5950
rect 45350 -6070 45470 -5950
rect 45525 -6070 45645 -5950
rect 45690 -6070 45810 -5950
rect 45855 -6070 45975 -5950
rect 46020 -6070 46140 -5950
rect 46195 -6070 46315 -5950
rect 46360 -6070 46480 -5950
rect 46525 -6070 46645 -5950
rect 46690 -6070 46810 -5950
rect 46865 -6070 46985 -5950
rect 47030 -6070 47150 -5950
rect 47195 -6070 47315 -5950
rect 47360 -6070 47480 -5950
rect 47535 -6070 47655 -5950
rect 42175 -6235 42295 -6115
rect 42340 -6235 42460 -6115
rect 42505 -6235 42625 -6115
rect 42670 -6235 42790 -6115
rect 42845 -6235 42965 -6115
rect 43010 -6235 43130 -6115
rect 43175 -6235 43295 -6115
rect 43340 -6235 43460 -6115
rect 43515 -6235 43635 -6115
rect 43680 -6235 43800 -6115
rect 43845 -6235 43965 -6115
rect 44010 -6235 44130 -6115
rect 44185 -6235 44305 -6115
rect 44350 -6235 44470 -6115
rect 44515 -6235 44635 -6115
rect 44680 -6235 44800 -6115
rect 44855 -6235 44975 -6115
rect 45020 -6235 45140 -6115
rect 45185 -6235 45305 -6115
rect 45350 -6235 45470 -6115
rect 45525 -6235 45645 -6115
rect 45690 -6235 45810 -6115
rect 45855 -6235 45975 -6115
rect 46020 -6235 46140 -6115
rect 46195 -6235 46315 -6115
rect 46360 -6235 46480 -6115
rect 46525 -6235 46645 -6115
rect 46690 -6235 46810 -6115
rect 46865 -6235 46985 -6115
rect 47030 -6235 47150 -6115
rect 47195 -6235 47315 -6115
rect 47360 -6235 47480 -6115
rect 47535 -6235 47655 -6115
rect 42175 -6400 42295 -6280
rect 42340 -6400 42460 -6280
rect 42505 -6400 42625 -6280
rect 42670 -6400 42790 -6280
rect 42845 -6400 42965 -6280
rect 43010 -6400 43130 -6280
rect 43175 -6400 43295 -6280
rect 43340 -6400 43460 -6280
rect 43515 -6400 43635 -6280
rect 43680 -6400 43800 -6280
rect 43845 -6400 43965 -6280
rect 44010 -6400 44130 -6280
rect 44185 -6400 44305 -6280
rect 44350 -6400 44470 -6280
rect 44515 -6400 44635 -6280
rect 44680 -6400 44800 -6280
rect 44855 -6400 44975 -6280
rect 45020 -6400 45140 -6280
rect 45185 -6400 45305 -6280
rect 45350 -6400 45470 -6280
rect 45525 -6400 45645 -6280
rect 45690 -6400 45810 -6280
rect 45855 -6400 45975 -6280
rect 46020 -6400 46140 -6280
rect 46195 -6400 46315 -6280
rect 46360 -6400 46480 -6280
rect 46525 -6400 46645 -6280
rect 46690 -6400 46810 -6280
rect 46865 -6400 46985 -6280
rect 47030 -6400 47150 -6280
rect 47195 -6400 47315 -6280
rect 47360 -6400 47480 -6280
rect 47535 -6400 47655 -6280
rect 42175 -6575 42295 -6455
rect 42340 -6575 42460 -6455
rect 42505 -6575 42625 -6455
rect 42670 -6575 42790 -6455
rect 42845 -6575 42965 -6455
rect 43010 -6575 43130 -6455
rect 43175 -6575 43295 -6455
rect 43340 -6575 43460 -6455
rect 43515 -6575 43635 -6455
rect 43680 -6575 43800 -6455
rect 43845 -6575 43965 -6455
rect 44010 -6575 44130 -6455
rect 44185 -6575 44305 -6455
rect 44350 -6575 44470 -6455
rect 44515 -6575 44635 -6455
rect 44680 -6575 44800 -6455
rect 44855 -6575 44975 -6455
rect 45020 -6575 45140 -6455
rect 45185 -6575 45305 -6455
rect 45350 -6575 45470 -6455
rect 45525 -6575 45645 -6455
rect 45690 -6575 45810 -6455
rect 45855 -6575 45975 -6455
rect 46020 -6575 46140 -6455
rect 46195 -6575 46315 -6455
rect 46360 -6575 46480 -6455
rect 46525 -6575 46645 -6455
rect 46690 -6575 46810 -6455
rect 46865 -6575 46985 -6455
rect 47030 -6575 47150 -6455
rect 47195 -6575 47315 -6455
rect 47360 -6575 47480 -6455
rect 47535 -6575 47655 -6455
rect 42175 -6740 42295 -6620
rect 42340 -6740 42460 -6620
rect 42505 -6740 42625 -6620
rect 42670 -6740 42790 -6620
rect 42845 -6740 42965 -6620
rect 43010 -6740 43130 -6620
rect 43175 -6740 43295 -6620
rect 43340 -6740 43460 -6620
rect 43515 -6740 43635 -6620
rect 43680 -6740 43800 -6620
rect 43845 -6740 43965 -6620
rect 44010 -6740 44130 -6620
rect 44185 -6740 44305 -6620
rect 44350 -6740 44470 -6620
rect 44515 -6740 44635 -6620
rect 44680 -6740 44800 -6620
rect 44855 -6740 44975 -6620
rect 45020 -6740 45140 -6620
rect 45185 -6740 45305 -6620
rect 45350 -6740 45470 -6620
rect 45525 -6740 45645 -6620
rect 45690 -6740 45810 -6620
rect 45855 -6740 45975 -6620
rect 46020 -6740 46140 -6620
rect 46195 -6740 46315 -6620
rect 46360 -6740 46480 -6620
rect 46525 -6740 46645 -6620
rect 46690 -6740 46810 -6620
rect 46865 -6740 46985 -6620
rect 47030 -6740 47150 -6620
rect 47195 -6740 47315 -6620
rect 47360 -6740 47480 -6620
rect 47535 -6740 47655 -6620
rect 42175 -6905 42295 -6785
rect 42340 -6905 42460 -6785
rect 42505 -6905 42625 -6785
rect 42670 -6905 42790 -6785
rect 42845 -6905 42965 -6785
rect 43010 -6905 43130 -6785
rect 43175 -6905 43295 -6785
rect 43340 -6905 43460 -6785
rect 43515 -6905 43635 -6785
rect 43680 -6905 43800 -6785
rect 43845 -6905 43965 -6785
rect 44010 -6905 44130 -6785
rect 44185 -6905 44305 -6785
rect 44350 -6905 44470 -6785
rect 44515 -6905 44635 -6785
rect 44680 -6905 44800 -6785
rect 44855 -6905 44975 -6785
rect 45020 -6905 45140 -6785
rect 45185 -6905 45305 -6785
rect 45350 -6905 45470 -6785
rect 45525 -6905 45645 -6785
rect 45690 -6905 45810 -6785
rect 45855 -6905 45975 -6785
rect 46020 -6905 46140 -6785
rect 46195 -6905 46315 -6785
rect 46360 -6905 46480 -6785
rect 46525 -6905 46645 -6785
rect 46690 -6905 46810 -6785
rect 46865 -6905 46985 -6785
rect 47030 -6905 47150 -6785
rect 47195 -6905 47315 -6785
rect 47360 -6905 47480 -6785
rect 47535 -6905 47655 -6785
rect 42175 -7070 42295 -6950
rect 42340 -7070 42460 -6950
rect 42505 -7070 42625 -6950
rect 42670 -7070 42790 -6950
rect 42845 -7070 42965 -6950
rect 43010 -7070 43130 -6950
rect 43175 -7070 43295 -6950
rect 43340 -7070 43460 -6950
rect 43515 -7070 43635 -6950
rect 43680 -7070 43800 -6950
rect 43845 -7070 43965 -6950
rect 44010 -7070 44130 -6950
rect 44185 -7070 44305 -6950
rect 44350 -7070 44470 -6950
rect 44515 -7070 44635 -6950
rect 44680 -7070 44800 -6950
rect 44855 -7070 44975 -6950
rect 45020 -7070 45140 -6950
rect 45185 -7070 45305 -6950
rect 45350 -7070 45470 -6950
rect 45525 -7070 45645 -6950
rect 45690 -7070 45810 -6950
rect 45855 -7070 45975 -6950
rect 46020 -7070 46140 -6950
rect 46195 -7070 46315 -6950
rect 46360 -7070 46480 -6950
rect 46525 -7070 46645 -6950
rect 46690 -7070 46810 -6950
rect 46865 -7070 46985 -6950
rect 47030 -7070 47150 -6950
rect 47195 -7070 47315 -6950
rect 47360 -7070 47480 -6950
rect 47535 -7070 47655 -6950
rect 42175 -7245 42295 -7125
rect 42340 -7245 42460 -7125
rect 42505 -7245 42625 -7125
rect 42670 -7245 42790 -7125
rect 42845 -7245 42965 -7125
rect 43010 -7245 43130 -7125
rect 43175 -7245 43295 -7125
rect 43340 -7245 43460 -7125
rect 43515 -7245 43635 -7125
rect 43680 -7245 43800 -7125
rect 43845 -7245 43965 -7125
rect 44010 -7245 44130 -7125
rect 44185 -7245 44305 -7125
rect 44350 -7245 44470 -7125
rect 44515 -7245 44635 -7125
rect 44680 -7245 44800 -7125
rect 44855 -7245 44975 -7125
rect 45020 -7245 45140 -7125
rect 45185 -7245 45305 -7125
rect 45350 -7245 45470 -7125
rect 45525 -7245 45645 -7125
rect 45690 -7245 45810 -7125
rect 45855 -7245 45975 -7125
rect 46020 -7245 46140 -7125
rect 46195 -7245 46315 -7125
rect 46360 -7245 46480 -7125
rect 46525 -7245 46645 -7125
rect 46690 -7245 46810 -7125
rect 46865 -7245 46985 -7125
rect 47030 -7245 47150 -7125
rect 47195 -7245 47315 -7125
rect 47360 -7245 47480 -7125
rect 47535 -7245 47655 -7125
rect 42175 -7410 42295 -7290
rect 42340 -7410 42460 -7290
rect 42505 -7410 42625 -7290
rect 42670 -7410 42790 -7290
rect 42845 -7410 42965 -7290
rect 43010 -7410 43130 -7290
rect 43175 -7410 43295 -7290
rect 43340 -7410 43460 -7290
rect 43515 -7410 43635 -7290
rect 43680 -7410 43800 -7290
rect 43845 -7410 43965 -7290
rect 44010 -7410 44130 -7290
rect 44185 -7410 44305 -7290
rect 44350 -7410 44470 -7290
rect 44515 -7410 44635 -7290
rect 44680 -7410 44800 -7290
rect 44855 -7410 44975 -7290
rect 45020 -7410 45140 -7290
rect 45185 -7410 45305 -7290
rect 45350 -7410 45470 -7290
rect 45525 -7410 45645 -7290
rect 45690 -7410 45810 -7290
rect 45855 -7410 45975 -7290
rect 46020 -7410 46140 -7290
rect 46195 -7410 46315 -7290
rect 46360 -7410 46480 -7290
rect 46525 -7410 46645 -7290
rect 46690 -7410 46810 -7290
rect 46865 -7410 46985 -7290
rect 47030 -7410 47150 -7290
rect 47195 -7410 47315 -7290
rect 47360 -7410 47480 -7290
rect 47535 -7410 47655 -7290
rect 42175 -7575 42295 -7455
rect 42340 -7575 42460 -7455
rect 42505 -7575 42625 -7455
rect 42670 -7575 42790 -7455
rect 42845 -7575 42965 -7455
rect 43010 -7575 43130 -7455
rect 43175 -7575 43295 -7455
rect 43340 -7575 43460 -7455
rect 43515 -7575 43635 -7455
rect 43680 -7575 43800 -7455
rect 43845 -7575 43965 -7455
rect 44010 -7575 44130 -7455
rect 44185 -7575 44305 -7455
rect 44350 -7575 44470 -7455
rect 44515 -7575 44635 -7455
rect 44680 -7575 44800 -7455
rect 44855 -7575 44975 -7455
rect 45020 -7575 45140 -7455
rect 45185 -7575 45305 -7455
rect 45350 -7575 45470 -7455
rect 45525 -7575 45645 -7455
rect 45690 -7575 45810 -7455
rect 45855 -7575 45975 -7455
rect 46020 -7575 46140 -7455
rect 46195 -7575 46315 -7455
rect 46360 -7575 46480 -7455
rect 46525 -7575 46645 -7455
rect 46690 -7575 46810 -7455
rect 46865 -7575 46985 -7455
rect 47030 -7575 47150 -7455
rect 47195 -7575 47315 -7455
rect 47360 -7575 47480 -7455
rect 47535 -7575 47655 -7455
rect 42175 -7740 42295 -7620
rect 42340 -7740 42460 -7620
rect 42505 -7740 42625 -7620
rect 42670 -7740 42790 -7620
rect 42845 -7740 42965 -7620
rect 43010 -7740 43130 -7620
rect 43175 -7740 43295 -7620
rect 43340 -7740 43460 -7620
rect 43515 -7740 43635 -7620
rect 43680 -7740 43800 -7620
rect 43845 -7740 43965 -7620
rect 44010 -7740 44130 -7620
rect 44185 -7740 44305 -7620
rect 44350 -7740 44470 -7620
rect 44515 -7740 44635 -7620
rect 44680 -7740 44800 -7620
rect 44855 -7740 44975 -7620
rect 45020 -7740 45140 -7620
rect 45185 -7740 45305 -7620
rect 45350 -7740 45470 -7620
rect 45525 -7740 45645 -7620
rect 45690 -7740 45810 -7620
rect 45855 -7740 45975 -7620
rect 46020 -7740 46140 -7620
rect 46195 -7740 46315 -7620
rect 46360 -7740 46480 -7620
rect 46525 -7740 46645 -7620
rect 46690 -7740 46810 -7620
rect 46865 -7740 46985 -7620
rect 47030 -7740 47150 -7620
rect 47195 -7740 47315 -7620
rect 47360 -7740 47480 -7620
rect 47535 -7740 47655 -7620
rect 42175 -7915 42295 -7795
rect 42340 -7915 42460 -7795
rect 42505 -7915 42625 -7795
rect 42670 -7915 42790 -7795
rect 42845 -7915 42965 -7795
rect 43010 -7915 43130 -7795
rect 43175 -7915 43295 -7795
rect 43340 -7915 43460 -7795
rect 43515 -7915 43635 -7795
rect 43680 -7915 43800 -7795
rect 43845 -7915 43965 -7795
rect 44010 -7915 44130 -7795
rect 44185 -7915 44305 -7795
rect 44350 -7915 44470 -7795
rect 44515 -7915 44635 -7795
rect 44680 -7915 44800 -7795
rect 44855 -7915 44975 -7795
rect 45020 -7915 45140 -7795
rect 45185 -7915 45305 -7795
rect 45350 -7915 45470 -7795
rect 45525 -7915 45645 -7795
rect 45690 -7915 45810 -7795
rect 45855 -7915 45975 -7795
rect 46020 -7915 46140 -7795
rect 46195 -7915 46315 -7795
rect 46360 -7915 46480 -7795
rect 46525 -7915 46645 -7795
rect 46690 -7915 46810 -7795
rect 46865 -7915 46985 -7795
rect 47030 -7915 47150 -7795
rect 47195 -7915 47315 -7795
rect 47360 -7915 47480 -7795
rect 47535 -7915 47655 -7795
rect 42175 -8080 42295 -7960
rect 42340 -8080 42460 -7960
rect 42505 -8080 42625 -7960
rect 42670 -8080 42790 -7960
rect 42845 -8080 42965 -7960
rect 43010 -8080 43130 -7960
rect 43175 -8080 43295 -7960
rect 43340 -8080 43460 -7960
rect 43515 -8080 43635 -7960
rect 43680 -8080 43800 -7960
rect 43845 -8080 43965 -7960
rect 44010 -8080 44130 -7960
rect 44185 -8080 44305 -7960
rect 44350 -8080 44470 -7960
rect 44515 -8080 44635 -7960
rect 44680 -8080 44800 -7960
rect 44855 -8080 44975 -7960
rect 45020 -8080 45140 -7960
rect 45185 -8080 45305 -7960
rect 45350 -8080 45470 -7960
rect 45525 -8080 45645 -7960
rect 45690 -8080 45810 -7960
rect 45855 -8080 45975 -7960
rect 46020 -8080 46140 -7960
rect 46195 -8080 46315 -7960
rect 46360 -8080 46480 -7960
rect 46525 -8080 46645 -7960
rect 46690 -8080 46810 -7960
rect 46865 -8080 46985 -7960
rect 47030 -8080 47150 -7960
rect 47195 -8080 47315 -7960
rect 47360 -8080 47480 -7960
rect 47535 -8080 47655 -7960
rect 42175 -8245 42295 -8125
rect 42340 -8245 42460 -8125
rect 42505 -8245 42625 -8125
rect 42670 -8245 42790 -8125
rect 42845 -8245 42965 -8125
rect 43010 -8245 43130 -8125
rect 43175 -8245 43295 -8125
rect 43340 -8245 43460 -8125
rect 43515 -8245 43635 -8125
rect 43680 -8245 43800 -8125
rect 43845 -8245 43965 -8125
rect 44010 -8245 44130 -8125
rect 44185 -8245 44305 -8125
rect 44350 -8245 44470 -8125
rect 44515 -8245 44635 -8125
rect 44680 -8245 44800 -8125
rect 44855 -8245 44975 -8125
rect 45020 -8245 45140 -8125
rect 45185 -8245 45305 -8125
rect 45350 -8245 45470 -8125
rect 45525 -8245 45645 -8125
rect 45690 -8245 45810 -8125
rect 45855 -8245 45975 -8125
rect 46020 -8245 46140 -8125
rect 46195 -8245 46315 -8125
rect 46360 -8245 46480 -8125
rect 46525 -8245 46645 -8125
rect 46690 -8245 46810 -8125
rect 46865 -8245 46985 -8125
rect 47030 -8245 47150 -8125
rect 47195 -8245 47315 -8125
rect 47360 -8245 47480 -8125
rect 47535 -8245 47655 -8125
rect 42175 -8410 42295 -8290
rect 42340 -8410 42460 -8290
rect 42505 -8410 42625 -8290
rect 42670 -8410 42790 -8290
rect 42845 -8410 42965 -8290
rect 43010 -8410 43130 -8290
rect 43175 -8410 43295 -8290
rect 43340 -8410 43460 -8290
rect 43515 -8410 43635 -8290
rect 43680 -8410 43800 -8290
rect 43845 -8410 43965 -8290
rect 44010 -8410 44130 -8290
rect 44185 -8410 44305 -8290
rect 44350 -8410 44470 -8290
rect 44515 -8410 44635 -8290
rect 44680 -8410 44800 -8290
rect 44855 -8410 44975 -8290
rect 45020 -8410 45140 -8290
rect 45185 -8410 45305 -8290
rect 45350 -8410 45470 -8290
rect 45525 -8410 45645 -8290
rect 45690 -8410 45810 -8290
rect 45855 -8410 45975 -8290
rect 46020 -8410 46140 -8290
rect 46195 -8410 46315 -8290
rect 46360 -8410 46480 -8290
rect 46525 -8410 46645 -8290
rect 46690 -8410 46810 -8290
rect 46865 -8410 46985 -8290
rect 47030 -8410 47150 -8290
rect 47195 -8410 47315 -8290
rect 47360 -8410 47480 -8290
rect 47535 -8410 47655 -8290
rect 42175 -8585 42295 -8465
rect 42340 -8585 42460 -8465
rect 42505 -8585 42625 -8465
rect 42670 -8585 42790 -8465
rect 42845 -8585 42965 -8465
rect 43010 -8585 43130 -8465
rect 43175 -8585 43295 -8465
rect 43340 -8585 43460 -8465
rect 43515 -8585 43635 -8465
rect 43680 -8585 43800 -8465
rect 43845 -8585 43965 -8465
rect 44010 -8585 44130 -8465
rect 44185 -8585 44305 -8465
rect 44350 -8585 44470 -8465
rect 44515 -8585 44635 -8465
rect 44680 -8585 44800 -8465
rect 44855 -8585 44975 -8465
rect 45020 -8585 45140 -8465
rect 45185 -8585 45305 -8465
rect 45350 -8585 45470 -8465
rect 45525 -8585 45645 -8465
rect 45690 -8585 45810 -8465
rect 45855 -8585 45975 -8465
rect 46020 -8585 46140 -8465
rect 46195 -8585 46315 -8465
rect 46360 -8585 46480 -8465
rect 46525 -8585 46645 -8465
rect 46690 -8585 46810 -8465
rect 46865 -8585 46985 -8465
rect 47030 -8585 47150 -8465
rect 47195 -8585 47315 -8465
rect 47360 -8585 47480 -8465
rect 47535 -8585 47655 -8465
rect 42175 -8750 42295 -8630
rect 42340 -8750 42460 -8630
rect 42505 -8750 42625 -8630
rect 42670 -8750 42790 -8630
rect 42845 -8750 42965 -8630
rect 43010 -8750 43130 -8630
rect 43175 -8750 43295 -8630
rect 43340 -8750 43460 -8630
rect 43515 -8750 43635 -8630
rect 43680 -8750 43800 -8630
rect 43845 -8750 43965 -8630
rect 44010 -8750 44130 -8630
rect 44185 -8750 44305 -8630
rect 44350 -8750 44470 -8630
rect 44515 -8750 44635 -8630
rect 44680 -8750 44800 -8630
rect 44855 -8750 44975 -8630
rect 45020 -8750 45140 -8630
rect 45185 -8750 45305 -8630
rect 45350 -8750 45470 -8630
rect 45525 -8750 45645 -8630
rect 45690 -8750 45810 -8630
rect 45855 -8750 45975 -8630
rect 46020 -8750 46140 -8630
rect 46195 -8750 46315 -8630
rect 46360 -8750 46480 -8630
rect 46525 -8750 46645 -8630
rect 46690 -8750 46810 -8630
rect 46865 -8750 46985 -8630
rect 47030 -8750 47150 -8630
rect 47195 -8750 47315 -8630
rect 47360 -8750 47480 -8630
rect 47535 -8750 47655 -8630
rect 42175 -8915 42295 -8795
rect 42340 -8915 42460 -8795
rect 42505 -8915 42625 -8795
rect 42670 -8915 42790 -8795
rect 42845 -8915 42965 -8795
rect 43010 -8915 43130 -8795
rect 43175 -8915 43295 -8795
rect 43340 -8915 43460 -8795
rect 43515 -8915 43635 -8795
rect 43680 -8915 43800 -8795
rect 43845 -8915 43965 -8795
rect 44010 -8915 44130 -8795
rect 44185 -8915 44305 -8795
rect 44350 -8915 44470 -8795
rect 44515 -8915 44635 -8795
rect 44680 -8915 44800 -8795
rect 44855 -8915 44975 -8795
rect 45020 -8915 45140 -8795
rect 45185 -8915 45305 -8795
rect 45350 -8915 45470 -8795
rect 45525 -8915 45645 -8795
rect 45690 -8915 45810 -8795
rect 45855 -8915 45975 -8795
rect 46020 -8915 46140 -8795
rect 46195 -8915 46315 -8795
rect 46360 -8915 46480 -8795
rect 46525 -8915 46645 -8795
rect 46690 -8915 46810 -8795
rect 46865 -8915 46985 -8795
rect 47030 -8915 47150 -8795
rect 47195 -8915 47315 -8795
rect 47360 -8915 47480 -8795
rect 47535 -8915 47655 -8795
rect 42175 -9080 42295 -8960
rect 42340 -9080 42460 -8960
rect 42505 -9080 42625 -8960
rect 42670 -9080 42790 -8960
rect 42845 -9080 42965 -8960
rect 43010 -9080 43130 -8960
rect 43175 -9080 43295 -8960
rect 43340 -9080 43460 -8960
rect 43515 -9080 43635 -8960
rect 43680 -9080 43800 -8960
rect 43845 -9080 43965 -8960
rect 44010 -9080 44130 -8960
rect 44185 -9080 44305 -8960
rect 44350 -9080 44470 -8960
rect 44515 -9080 44635 -8960
rect 44680 -9080 44800 -8960
rect 44855 -9080 44975 -8960
rect 45020 -9080 45140 -8960
rect 45185 -9080 45305 -8960
rect 45350 -9080 45470 -8960
rect 45525 -9080 45645 -8960
rect 45690 -9080 45810 -8960
rect 45855 -9080 45975 -8960
rect 46020 -9080 46140 -8960
rect 46195 -9080 46315 -8960
rect 46360 -9080 46480 -8960
rect 46525 -9080 46645 -8960
rect 46690 -9080 46810 -8960
rect 46865 -9080 46985 -8960
rect 47030 -9080 47150 -8960
rect 47195 -9080 47315 -8960
rect 47360 -9080 47480 -8960
rect 47535 -9080 47655 -8960
rect 42175 -9255 42295 -9135
rect 42340 -9255 42460 -9135
rect 42505 -9255 42625 -9135
rect 42670 -9255 42790 -9135
rect 42845 -9255 42965 -9135
rect 43010 -9255 43130 -9135
rect 43175 -9255 43295 -9135
rect 43340 -9255 43460 -9135
rect 43515 -9255 43635 -9135
rect 43680 -9255 43800 -9135
rect 43845 -9255 43965 -9135
rect 44010 -9255 44130 -9135
rect 44185 -9255 44305 -9135
rect 44350 -9255 44470 -9135
rect 44515 -9255 44635 -9135
rect 44680 -9255 44800 -9135
rect 44855 -9255 44975 -9135
rect 45020 -9255 45140 -9135
rect 45185 -9255 45305 -9135
rect 45350 -9255 45470 -9135
rect 45525 -9255 45645 -9135
rect 45690 -9255 45810 -9135
rect 45855 -9255 45975 -9135
rect 46020 -9255 46140 -9135
rect 46195 -9255 46315 -9135
rect 46360 -9255 46480 -9135
rect 46525 -9255 46645 -9135
rect 46690 -9255 46810 -9135
rect 46865 -9255 46985 -9135
rect 47030 -9255 47150 -9135
rect 47195 -9255 47315 -9135
rect 47360 -9255 47480 -9135
rect 47535 -9255 47655 -9135
rect 42175 -9420 42295 -9300
rect 42340 -9420 42460 -9300
rect 42505 -9420 42625 -9300
rect 42670 -9420 42790 -9300
rect 42845 -9420 42965 -9300
rect 43010 -9420 43130 -9300
rect 43175 -9420 43295 -9300
rect 43340 -9420 43460 -9300
rect 43515 -9420 43635 -9300
rect 43680 -9420 43800 -9300
rect 43845 -9420 43965 -9300
rect 44010 -9420 44130 -9300
rect 44185 -9420 44305 -9300
rect 44350 -9420 44470 -9300
rect 44515 -9420 44635 -9300
rect 44680 -9420 44800 -9300
rect 44855 -9420 44975 -9300
rect 45020 -9420 45140 -9300
rect 45185 -9420 45305 -9300
rect 45350 -9420 45470 -9300
rect 45525 -9420 45645 -9300
rect 45690 -9420 45810 -9300
rect 45855 -9420 45975 -9300
rect 46020 -9420 46140 -9300
rect 46195 -9420 46315 -9300
rect 46360 -9420 46480 -9300
rect 46525 -9420 46645 -9300
rect 46690 -9420 46810 -9300
rect 46865 -9420 46985 -9300
rect 47030 -9420 47150 -9300
rect 47195 -9420 47315 -9300
rect 47360 -9420 47480 -9300
rect 47535 -9420 47655 -9300
rect 42175 -9585 42295 -9465
rect 42340 -9585 42460 -9465
rect 42505 -9585 42625 -9465
rect 42670 -9585 42790 -9465
rect 42845 -9585 42965 -9465
rect 43010 -9585 43130 -9465
rect 43175 -9585 43295 -9465
rect 43340 -9585 43460 -9465
rect 43515 -9585 43635 -9465
rect 43680 -9585 43800 -9465
rect 43845 -9585 43965 -9465
rect 44010 -9585 44130 -9465
rect 44185 -9585 44305 -9465
rect 44350 -9585 44470 -9465
rect 44515 -9585 44635 -9465
rect 44680 -9585 44800 -9465
rect 44855 -9585 44975 -9465
rect 45020 -9585 45140 -9465
rect 45185 -9585 45305 -9465
rect 45350 -9585 45470 -9465
rect 45525 -9585 45645 -9465
rect 45690 -9585 45810 -9465
rect 45855 -9585 45975 -9465
rect 46020 -9585 46140 -9465
rect 46195 -9585 46315 -9465
rect 46360 -9585 46480 -9465
rect 46525 -9585 46645 -9465
rect 46690 -9585 46810 -9465
rect 46865 -9585 46985 -9465
rect 47030 -9585 47150 -9465
rect 47195 -9585 47315 -9465
rect 47360 -9585 47480 -9465
rect 47535 -9585 47655 -9465
rect 42175 -9750 42295 -9630
rect 42340 -9750 42460 -9630
rect 42505 -9750 42625 -9630
rect 42670 -9750 42790 -9630
rect 42845 -9750 42965 -9630
rect 43010 -9750 43130 -9630
rect 43175 -9750 43295 -9630
rect 43340 -9750 43460 -9630
rect 43515 -9750 43635 -9630
rect 43680 -9750 43800 -9630
rect 43845 -9750 43965 -9630
rect 44010 -9750 44130 -9630
rect 44185 -9750 44305 -9630
rect 44350 -9750 44470 -9630
rect 44515 -9750 44635 -9630
rect 44680 -9750 44800 -9630
rect 44855 -9750 44975 -9630
rect 45020 -9750 45140 -9630
rect 45185 -9750 45305 -9630
rect 45350 -9750 45470 -9630
rect 45525 -9750 45645 -9630
rect 45690 -9750 45810 -9630
rect 45855 -9750 45975 -9630
rect 46020 -9750 46140 -9630
rect 46195 -9750 46315 -9630
rect 46360 -9750 46480 -9630
rect 46525 -9750 46645 -9630
rect 46690 -9750 46810 -9630
rect 46865 -9750 46985 -9630
rect 47030 -9750 47150 -9630
rect 47195 -9750 47315 -9630
rect 47360 -9750 47480 -9630
rect 47535 -9750 47655 -9630
rect 47865 -4390 47985 -4270
rect 48030 -4390 48150 -4270
rect 48195 -4390 48315 -4270
rect 48360 -4390 48480 -4270
rect 48535 -4390 48655 -4270
rect 48700 -4390 48820 -4270
rect 48865 -4390 48985 -4270
rect 49030 -4390 49150 -4270
rect 49205 -4390 49325 -4270
rect 49370 -4390 49490 -4270
rect 49535 -4390 49655 -4270
rect 49700 -4390 49820 -4270
rect 49875 -4390 49995 -4270
rect 50040 -4390 50160 -4270
rect 50205 -4390 50325 -4270
rect 50370 -4390 50490 -4270
rect 50545 -4390 50665 -4270
rect 50710 -4390 50830 -4270
rect 50875 -4390 50995 -4270
rect 51040 -4390 51160 -4270
rect 51215 -4390 51335 -4270
rect 51380 -4390 51500 -4270
rect 51545 -4390 51665 -4270
rect 51710 -4390 51830 -4270
rect 51885 -4390 52005 -4270
rect 52050 -4390 52170 -4270
rect 52215 -4390 52335 -4270
rect 52380 -4390 52500 -4270
rect 52555 -4390 52675 -4270
rect 52720 -4390 52840 -4270
rect 52885 -4390 53005 -4270
rect 53050 -4390 53170 -4270
rect 53225 -4390 53345 -4270
rect 47865 -4565 47985 -4445
rect 48030 -4565 48150 -4445
rect 48195 -4565 48315 -4445
rect 48360 -4565 48480 -4445
rect 48535 -4565 48655 -4445
rect 48700 -4565 48820 -4445
rect 48865 -4565 48985 -4445
rect 49030 -4565 49150 -4445
rect 49205 -4565 49325 -4445
rect 49370 -4565 49490 -4445
rect 49535 -4565 49655 -4445
rect 49700 -4565 49820 -4445
rect 49875 -4565 49995 -4445
rect 50040 -4565 50160 -4445
rect 50205 -4565 50325 -4445
rect 50370 -4565 50490 -4445
rect 50545 -4565 50665 -4445
rect 50710 -4565 50830 -4445
rect 50875 -4565 50995 -4445
rect 51040 -4565 51160 -4445
rect 51215 -4565 51335 -4445
rect 51380 -4565 51500 -4445
rect 51545 -4565 51665 -4445
rect 51710 -4565 51830 -4445
rect 51885 -4565 52005 -4445
rect 52050 -4565 52170 -4445
rect 52215 -4565 52335 -4445
rect 52380 -4565 52500 -4445
rect 52555 -4565 52675 -4445
rect 52720 -4565 52840 -4445
rect 52885 -4565 53005 -4445
rect 53050 -4565 53170 -4445
rect 53225 -4565 53345 -4445
rect 47865 -4730 47985 -4610
rect 48030 -4730 48150 -4610
rect 48195 -4730 48315 -4610
rect 48360 -4730 48480 -4610
rect 48535 -4730 48655 -4610
rect 48700 -4730 48820 -4610
rect 48865 -4730 48985 -4610
rect 49030 -4730 49150 -4610
rect 49205 -4730 49325 -4610
rect 49370 -4730 49490 -4610
rect 49535 -4730 49655 -4610
rect 49700 -4730 49820 -4610
rect 49875 -4730 49995 -4610
rect 50040 -4730 50160 -4610
rect 50205 -4730 50325 -4610
rect 50370 -4730 50490 -4610
rect 50545 -4730 50665 -4610
rect 50710 -4730 50830 -4610
rect 50875 -4730 50995 -4610
rect 51040 -4730 51160 -4610
rect 51215 -4730 51335 -4610
rect 51380 -4730 51500 -4610
rect 51545 -4730 51665 -4610
rect 51710 -4730 51830 -4610
rect 51885 -4730 52005 -4610
rect 52050 -4730 52170 -4610
rect 52215 -4730 52335 -4610
rect 52380 -4730 52500 -4610
rect 52555 -4730 52675 -4610
rect 52720 -4730 52840 -4610
rect 52885 -4730 53005 -4610
rect 53050 -4730 53170 -4610
rect 53225 -4730 53345 -4610
rect 47865 -4895 47985 -4775
rect 48030 -4895 48150 -4775
rect 48195 -4895 48315 -4775
rect 48360 -4895 48480 -4775
rect 48535 -4895 48655 -4775
rect 48700 -4895 48820 -4775
rect 48865 -4895 48985 -4775
rect 49030 -4895 49150 -4775
rect 49205 -4895 49325 -4775
rect 49370 -4895 49490 -4775
rect 49535 -4895 49655 -4775
rect 49700 -4895 49820 -4775
rect 49875 -4895 49995 -4775
rect 50040 -4895 50160 -4775
rect 50205 -4895 50325 -4775
rect 50370 -4895 50490 -4775
rect 50545 -4895 50665 -4775
rect 50710 -4895 50830 -4775
rect 50875 -4895 50995 -4775
rect 51040 -4895 51160 -4775
rect 51215 -4895 51335 -4775
rect 51380 -4895 51500 -4775
rect 51545 -4895 51665 -4775
rect 51710 -4895 51830 -4775
rect 51885 -4895 52005 -4775
rect 52050 -4895 52170 -4775
rect 52215 -4895 52335 -4775
rect 52380 -4895 52500 -4775
rect 52555 -4895 52675 -4775
rect 52720 -4895 52840 -4775
rect 52885 -4895 53005 -4775
rect 53050 -4895 53170 -4775
rect 53225 -4895 53345 -4775
rect 47865 -5060 47985 -4940
rect 48030 -5060 48150 -4940
rect 48195 -5060 48315 -4940
rect 48360 -5060 48480 -4940
rect 48535 -5060 48655 -4940
rect 48700 -5060 48820 -4940
rect 48865 -5060 48985 -4940
rect 49030 -5060 49150 -4940
rect 49205 -5060 49325 -4940
rect 49370 -5060 49490 -4940
rect 49535 -5060 49655 -4940
rect 49700 -5060 49820 -4940
rect 49875 -5060 49995 -4940
rect 50040 -5060 50160 -4940
rect 50205 -5060 50325 -4940
rect 50370 -5060 50490 -4940
rect 50545 -5060 50665 -4940
rect 50710 -5060 50830 -4940
rect 50875 -5060 50995 -4940
rect 51040 -5060 51160 -4940
rect 51215 -5060 51335 -4940
rect 51380 -5060 51500 -4940
rect 51545 -5060 51665 -4940
rect 51710 -5060 51830 -4940
rect 51885 -5060 52005 -4940
rect 52050 -5060 52170 -4940
rect 52215 -5060 52335 -4940
rect 52380 -5060 52500 -4940
rect 52555 -5060 52675 -4940
rect 52720 -5060 52840 -4940
rect 52885 -5060 53005 -4940
rect 53050 -5060 53170 -4940
rect 53225 -5060 53345 -4940
rect 47865 -5235 47985 -5115
rect 48030 -5235 48150 -5115
rect 48195 -5235 48315 -5115
rect 48360 -5235 48480 -5115
rect 48535 -5235 48655 -5115
rect 48700 -5235 48820 -5115
rect 48865 -5235 48985 -5115
rect 49030 -5235 49150 -5115
rect 49205 -5235 49325 -5115
rect 49370 -5235 49490 -5115
rect 49535 -5235 49655 -5115
rect 49700 -5235 49820 -5115
rect 49875 -5235 49995 -5115
rect 50040 -5235 50160 -5115
rect 50205 -5235 50325 -5115
rect 50370 -5235 50490 -5115
rect 50545 -5235 50665 -5115
rect 50710 -5235 50830 -5115
rect 50875 -5235 50995 -5115
rect 51040 -5235 51160 -5115
rect 51215 -5235 51335 -5115
rect 51380 -5235 51500 -5115
rect 51545 -5235 51665 -5115
rect 51710 -5235 51830 -5115
rect 51885 -5235 52005 -5115
rect 52050 -5235 52170 -5115
rect 52215 -5235 52335 -5115
rect 52380 -5235 52500 -5115
rect 52555 -5235 52675 -5115
rect 52720 -5235 52840 -5115
rect 52885 -5235 53005 -5115
rect 53050 -5235 53170 -5115
rect 53225 -5235 53345 -5115
rect 47865 -5400 47985 -5280
rect 48030 -5400 48150 -5280
rect 48195 -5400 48315 -5280
rect 48360 -5400 48480 -5280
rect 48535 -5400 48655 -5280
rect 48700 -5400 48820 -5280
rect 48865 -5400 48985 -5280
rect 49030 -5400 49150 -5280
rect 49205 -5400 49325 -5280
rect 49370 -5400 49490 -5280
rect 49535 -5400 49655 -5280
rect 49700 -5400 49820 -5280
rect 49875 -5400 49995 -5280
rect 50040 -5400 50160 -5280
rect 50205 -5400 50325 -5280
rect 50370 -5400 50490 -5280
rect 50545 -5400 50665 -5280
rect 50710 -5400 50830 -5280
rect 50875 -5400 50995 -5280
rect 51040 -5400 51160 -5280
rect 51215 -5400 51335 -5280
rect 51380 -5400 51500 -5280
rect 51545 -5400 51665 -5280
rect 51710 -5400 51830 -5280
rect 51885 -5400 52005 -5280
rect 52050 -5400 52170 -5280
rect 52215 -5400 52335 -5280
rect 52380 -5400 52500 -5280
rect 52555 -5400 52675 -5280
rect 52720 -5400 52840 -5280
rect 52885 -5400 53005 -5280
rect 53050 -5400 53170 -5280
rect 53225 -5400 53345 -5280
rect 47865 -5565 47985 -5445
rect 48030 -5565 48150 -5445
rect 48195 -5565 48315 -5445
rect 48360 -5565 48480 -5445
rect 48535 -5565 48655 -5445
rect 48700 -5565 48820 -5445
rect 48865 -5565 48985 -5445
rect 49030 -5565 49150 -5445
rect 49205 -5565 49325 -5445
rect 49370 -5565 49490 -5445
rect 49535 -5565 49655 -5445
rect 49700 -5565 49820 -5445
rect 49875 -5565 49995 -5445
rect 50040 -5565 50160 -5445
rect 50205 -5565 50325 -5445
rect 50370 -5565 50490 -5445
rect 50545 -5565 50665 -5445
rect 50710 -5565 50830 -5445
rect 50875 -5565 50995 -5445
rect 51040 -5565 51160 -5445
rect 51215 -5565 51335 -5445
rect 51380 -5565 51500 -5445
rect 51545 -5565 51665 -5445
rect 51710 -5565 51830 -5445
rect 51885 -5565 52005 -5445
rect 52050 -5565 52170 -5445
rect 52215 -5565 52335 -5445
rect 52380 -5565 52500 -5445
rect 52555 -5565 52675 -5445
rect 52720 -5565 52840 -5445
rect 52885 -5565 53005 -5445
rect 53050 -5565 53170 -5445
rect 53225 -5565 53345 -5445
rect 47865 -5730 47985 -5610
rect 48030 -5730 48150 -5610
rect 48195 -5730 48315 -5610
rect 48360 -5730 48480 -5610
rect 48535 -5730 48655 -5610
rect 48700 -5730 48820 -5610
rect 48865 -5730 48985 -5610
rect 49030 -5730 49150 -5610
rect 49205 -5730 49325 -5610
rect 49370 -5730 49490 -5610
rect 49535 -5730 49655 -5610
rect 49700 -5730 49820 -5610
rect 49875 -5730 49995 -5610
rect 50040 -5730 50160 -5610
rect 50205 -5730 50325 -5610
rect 50370 -5730 50490 -5610
rect 50545 -5730 50665 -5610
rect 50710 -5730 50830 -5610
rect 50875 -5730 50995 -5610
rect 51040 -5730 51160 -5610
rect 51215 -5730 51335 -5610
rect 51380 -5730 51500 -5610
rect 51545 -5730 51665 -5610
rect 51710 -5730 51830 -5610
rect 51885 -5730 52005 -5610
rect 52050 -5730 52170 -5610
rect 52215 -5730 52335 -5610
rect 52380 -5730 52500 -5610
rect 52555 -5730 52675 -5610
rect 52720 -5730 52840 -5610
rect 52885 -5730 53005 -5610
rect 53050 -5730 53170 -5610
rect 53225 -5730 53345 -5610
rect 47865 -5905 47985 -5785
rect 48030 -5905 48150 -5785
rect 48195 -5905 48315 -5785
rect 48360 -5905 48480 -5785
rect 48535 -5905 48655 -5785
rect 48700 -5905 48820 -5785
rect 48865 -5905 48985 -5785
rect 49030 -5905 49150 -5785
rect 49205 -5905 49325 -5785
rect 49370 -5905 49490 -5785
rect 49535 -5905 49655 -5785
rect 49700 -5905 49820 -5785
rect 49875 -5905 49995 -5785
rect 50040 -5905 50160 -5785
rect 50205 -5905 50325 -5785
rect 50370 -5905 50490 -5785
rect 50545 -5905 50665 -5785
rect 50710 -5905 50830 -5785
rect 50875 -5905 50995 -5785
rect 51040 -5905 51160 -5785
rect 51215 -5905 51335 -5785
rect 51380 -5905 51500 -5785
rect 51545 -5905 51665 -5785
rect 51710 -5905 51830 -5785
rect 51885 -5905 52005 -5785
rect 52050 -5905 52170 -5785
rect 52215 -5905 52335 -5785
rect 52380 -5905 52500 -5785
rect 52555 -5905 52675 -5785
rect 52720 -5905 52840 -5785
rect 52885 -5905 53005 -5785
rect 53050 -5905 53170 -5785
rect 53225 -5905 53345 -5785
rect 47865 -6070 47985 -5950
rect 48030 -6070 48150 -5950
rect 48195 -6070 48315 -5950
rect 48360 -6070 48480 -5950
rect 48535 -6070 48655 -5950
rect 48700 -6070 48820 -5950
rect 48865 -6070 48985 -5950
rect 49030 -6070 49150 -5950
rect 49205 -6070 49325 -5950
rect 49370 -6070 49490 -5950
rect 49535 -6070 49655 -5950
rect 49700 -6070 49820 -5950
rect 49875 -6070 49995 -5950
rect 50040 -6070 50160 -5950
rect 50205 -6070 50325 -5950
rect 50370 -6070 50490 -5950
rect 50545 -6070 50665 -5950
rect 50710 -6070 50830 -5950
rect 50875 -6070 50995 -5950
rect 51040 -6070 51160 -5950
rect 51215 -6070 51335 -5950
rect 51380 -6070 51500 -5950
rect 51545 -6070 51665 -5950
rect 51710 -6070 51830 -5950
rect 51885 -6070 52005 -5950
rect 52050 -6070 52170 -5950
rect 52215 -6070 52335 -5950
rect 52380 -6070 52500 -5950
rect 52555 -6070 52675 -5950
rect 52720 -6070 52840 -5950
rect 52885 -6070 53005 -5950
rect 53050 -6070 53170 -5950
rect 53225 -6070 53345 -5950
rect 47865 -6235 47985 -6115
rect 48030 -6235 48150 -6115
rect 48195 -6235 48315 -6115
rect 48360 -6235 48480 -6115
rect 48535 -6235 48655 -6115
rect 48700 -6235 48820 -6115
rect 48865 -6235 48985 -6115
rect 49030 -6235 49150 -6115
rect 49205 -6235 49325 -6115
rect 49370 -6235 49490 -6115
rect 49535 -6235 49655 -6115
rect 49700 -6235 49820 -6115
rect 49875 -6235 49995 -6115
rect 50040 -6235 50160 -6115
rect 50205 -6235 50325 -6115
rect 50370 -6235 50490 -6115
rect 50545 -6235 50665 -6115
rect 50710 -6235 50830 -6115
rect 50875 -6235 50995 -6115
rect 51040 -6235 51160 -6115
rect 51215 -6235 51335 -6115
rect 51380 -6235 51500 -6115
rect 51545 -6235 51665 -6115
rect 51710 -6235 51830 -6115
rect 51885 -6235 52005 -6115
rect 52050 -6235 52170 -6115
rect 52215 -6235 52335 -6115
rect 52380 -6235 52500 -6115
rect 52555 -6235 52675 -6115
rect 52720 -6235 52840 -6115
rect 52885 -6235 53005 -6115
rect 53050 -6235 53170 -6115
rect 53225 -6235 53345 -6115
rect 47865 -6400 47985 -6280
rect 48030 -6400 48150 -6280
rect 48195 -6400 48315 -6280
rect 48360 -6400 48480 -6280
rect 48535 -6400 48655 -6280
rect 48700 -6400 48820 -6280
rect 48865 -6400 48985 -6280
rect 49030 -6400 49150 -6280
rect 49205 -6400 49325 -6280
rect 49370 -6400 49490 -6280
rect 49535 -6400 49655 -6280
rect 49700 -6400 49820 -6280
rect 49875 -6400 49995 -6280
rect 50040 -6400 50160 -6280
rect 50205 -6400 50325 -6280
rect 50370 -6400 50490 -6280
rect 50545 -6400 50665 -6280
rect 50710 -6400 50830 -6280
rect 50875 -6400 50995 -6280
rect 51040 -6400 51160 -6280
rect 51215 -6400 51335 -6280
rect 51380 -6400 51500 -6280
rect 51545 -6400 51665 -6280
rect 51710 -6400 51830 -6280
rect 51885 -6400 52005 -6280
rect 52050 -6400 52170 -6280
rect 52215 -6400 52335 -6280
rect 52380 -6400 52500 -6280
rect 52555 -6400 52675 -6280
rect 52720 -6400 52840 -6280
rect 52885 -6400 53005 -6280
rect 53050 -6400 53170 -6280
rect 53225 -6400 53345 -6280
rect 47865 -6575 47985 -6455
rect 48030 -6575 48150 -6455
rect 48195 -6575 48315 -6455
rect 48360 -6575 48480 -6455
rect 48535 -6575 48655 -6455
rect 48700 -6575 48820 -6455
rect 48865 -6575 48985 -6455
rect 49030 -6575 49150 -6455
rect 49205 -6575 49325 -6455
rect 49370 -6575 49490 -6455
rect 49535 -6575 49655 -6455
rect 49700 -6575 49820 -6455
rect 49875 -6575 49995 -6455
rect 50040 -6575 50160 -6455
rect 50205 -6575 50325 -6455
rect 50370 -6575 50490 -6455
rect 50545 -6575 50665 -6455
rect 50710 -6575 50830 -6455
rect 50875 -6575 50995 -6455
rect 51040 -6575 51160 -6455
rect 51215 -6575 51335 -6455
rect 51380 -6575 51500 -6455
rect 51545 -6575 51665 -6455
rect 51710 -6575 51830 -6455
rect 51885 -6575 52005 -6455
rect 52050 -6575 52170 -6455
rect 52215 -6575 52335 -6455
rect 52380 -6575 52500 -6455
rect 52555 -6575 52675 -6455
rect 52720 -6575 52840 -6455
rect 52885 -6575 53005 -6455
rect 53050 -6575 53170 -6455
rect 53225 -6575 53345 -6455
rect 47865 -6740 47985 -6620
rect 48030 -6740 48150 -6620
rect 48195 -6740 48315 -6620
rect 48360 -6740 48480 -6620
rect 48535 -6740 48655 -6620
rect 48700 -6740 48820 -6620
rect 48865 -6740 48985 -6620
rect 49030 -6740 49150 -6620
rect 49205 -6740 49325 -6620
rect 49370 -6740 49490 -6620
rect 49535 -6740 49655 -6620
rect 49700 -6740 49820 -6620
rect 49875 -6740 49995 -6620
rect 50040 -6740 50160 -6620
rect 50205 -6740 50325 -6620
rect 50370 -6740 50490 -6620
rect 50545 -6740 50665 -6620
rect 50710 -6740 50830 -6620
rect 50875 -6740 50995 -6620
rect 51040 -6740 51160 -6620
rect 51215 -6740 51335 -6620
rect 51380 -6740 51500 -6620
rect 51545 -6740 51665 -6620
rect 51710 -6740 51830 -6620
rect 51885 -6740 52005 -6620
rect 52050 -6740 52170 -6620
rect 52215 -6740 52335 -6620
rect 52380 -6740 52500 -6620
rect 52555 -6740 52675 -6620
rect 52720 -6740 52840 -6620
rect 52885 -6740 53005 -6620
rect 53050 -6740 53170 -6620
rect 53225 -6740 53345 -6620
rect 47865 -6905 47985 -6785
rect 48030 -6905 48150 -6785
rect 48195 -6905 48315 -6785
rect 48360 -6905 48480 -6785
rect 48535 -6905 48655 -6785
rect 48700 -6905 48820 -6785
rect 48865 -6905 48985 -6785
rect 49030 -6905 49150 -6785
rect 49205 -6905 49325 -6785
rect 49370 -6905 49490 -6785
rect 49535 -6905 49655 -6785
rect 49700 -6905 49820 -6785
rect 49875 -6905 49995 -6785
rect 50040 -6905 50160 -6785
rect 50205 -6905 50325 -6785
rect 50370 -6905 50490 -6785
rect 50545 -6905 50665 -6785
rect 50710 -6905 50830 -6785
rect 50875 -6905 50995 -6785
rect 51040 -6905 51160 -6785
rect 51215 -6905 51335 -6785
rect 51380 -6905 51500 -6785
rect 51545 -6905 51665 -6785
rect 51710 -6905 51830 -6785
rect 51885 -6905 52005 -6785
rect 52050 -6905 52170 -6785
rect 52215 -6905 52335 -6785
rect 52380 -6905 52500 -6785
rect 52555 -6905 52675 -6785
rect 52720 -6905 52840 -6785
rect 52885 -6905 53005 -6785
rect 53050 -6905 53170 -6785
rect 53225 -6905 53345 -6785
rect 47865 -7070 47985 -6950
rect 48030 -7070 48150 -6950
rect 48195 -7070 48315 -6950
rect 48360 -7070 48480 -6950
rect 48535 -7070 48655 -6950
rect 48700 -7070 48820 -6950
rect 48865 -7070 48985 -6950
rect 49030 -7070 49150 -6950
rect 49205 -7070 49325 -6950
rect 49370 -7070 49490 -6950
rect 49535 -7070 49655 -6950
rect 49700 -7070 49820 -6950
rect 49875 -7070 49995 -6950
rect 50040 -7070 50160 -6950
rect 50205 -7070 50325 -6950
rect 50370 -7070 50490 -6950
rect 50545 -7070 50665 -6950
rect 50710 -7070 50830 -6950
rect 50875 -7070 50995 -6950
rect 51040 -7070 51160 -6950
rect 51215 -7070 51335 -6950
rect 51380 -7070 51500 -6950
rect 51545 -7070 51665 -6950
rect 51710 -7070 51830 -6950
rect 51885 -7070 52005 -6950
rect 52050 -7070 52170 -6950
rect 52215 -7070 52335 -6950
rect 52380 -7070 52500 -6950
rect 52555 -7070 52675 -6950
rect 52720 -7070 52840 -6950
rect 52885 -7070 53005 -6950
rect 53050 -7070 53170 -6950
rect 53225 -7070 53345 -6950
rect 47865 -7245 47985 -7125
rect 48030 -7245 48150 -7125
rect 48195 -7245 48315 -7125
rect 48360 -7245 48480 -7125
rect 48535 -7245 48655 -7125
rect 48700 -7245 48820 -7125
rect 48865 -7245 48985 -7125
rect 49030 -7245 49150 -7125
rect 49205 -7245 49325 -7125
rect 49370 -7245 49490 -7125
rect 49535 -7245 49655 -7125
rect 49700 -7245 49820 -7125
rect 49875 -7245 49995 -7125
rect 50040 -7245 50160 -7125
rect 50205 -7245 50325 -7125
rect 50370 -7245 50490 -7125
rect 50545 -7245 50665 -7125
rect 50710 -7245 50830 -7125
rect 50875 -7245 50995 -7125
rect 51040 -7245 51160 -7125
rect 51215 -7245 51335 -7125
rect 51380 -7245 51500 -7125
rect 51545 -7245 51665 -7125
rect 51710 -7245 51830 -7125
rect 51885 -7245 52005 -7125
rect 52050 -7245 52170 -7125
rect 52215 -7245 52335 -7125
rect 52380 -7245 52500 -7125
rect 52555 -7245 52675 -7125
rect 52720 -7245 52840 -7125
rect 52885 -7245 53005 -7125
rect 53050 -7245 53170 -7125
rect 53225 -7245 53345 -7125
rect 47865 -7410 47985 -7290
rect 48030 -7410 48150 -7290
rect 48195 -7410 48315 -7290
rect 48360 -7410 48480 -7290
rect 48535 -7410 48655 -7290
rect 48700 -7410 48820 -7290
rect 48865 -7410 48985 -7290
rect 49030 -7410 49150 -7290
rect 49205 -7410 49325 -7290
rect 49370 -7410 49490 -7290
rect 49535 -7410 49655 -7290
rect 49700 -7410 49820 -7290
rect 49875 -7410 49995 -7290
rect 50040 -7410 50160 -7290
rect 50205 -7410 50325 -7290
rect 50370 -7410 50490 -7290
rect 50545 -7410 50665 -7290
rect 50710 -7410 50830 -7290
rect 50875 -7410 50995 -7290
rect 51040 -7410 51160 -7290
rect 51215 -7410 51335 -7290
rect 51380 -7410 51500 -7290
rect 51545 -7410 51665 -7290
rect 51710 -7410 51830 -7290
rect 51885 -7410 52005 -7290
rect 52050 -7410 52170 -7290
rect 52215 -7410 52335 -7290
rect 52380 -7410 52500 -7290
rect 52555 -7410 52675 -7290
rect 52720 -7410 52840 -7290
rect 52885 -7410 53005 -7290
rect 53050 -7410 53170 -7290
rect 53225 -7410 53345 -7290
rect 47865 -7575 47985 -7455
rect 48030 -7575 48150 -7455
rect 48195 -7575 48315 -7455
rect 48360 -7575 48480 -7455
rect 48535 -7575 48655 -7455
rect 48700 -7575 48820 -7455
rect 48865 -7575 48985 -7455
rect 49030 -7575 49150 -7455
rect 49205 -7575 49325 -7455
rect 49370 -7575 49490 -7455
rect 49535 -7575 49655 -7455
rect 49700 -7575 49820 -7455
rect 49875 -7575 49995 -7455
rect 50040 -7575 50160 -7455
rect 50205 -7575 50325 -7455
rect 50370 -7575 50490 -7455
rect 50545 -7575 50665 -7455
rect 50710 -7575 50830 -7455
rect 50875 -7575 50995 -7455
rect 51040 -7575 51160 -7455
rect 51215 -7575 51335 -7455
rect 51380 -7575 51500 -7455
rect 51545 -7575 51665 -7455
rect 51710 -7575 51830 -7455
rect 51885 -7575 52005 -7455
rect 52050 -7575 52170 -7455
rect 52215 -7575 52335 -7455
rect 52380 -7575 52500 -7455
rect 52555 -7575 52675 -7455
rect 52720 -7575 52840 -7455
rect 52885 -7575 53005 -7455
rect 53050 -7575 53170 -7455
rect 53225 -7575 53345 -7455
rect 47865 -7740 47985 -7620
rect 48030 -7740 48150 -7620
rect 48195 -7740 48315 -7620
rect 48360 -7740 48480 -7620
rect 48535 -7740 48655 -7620
rect 48700 -7740 48820 -7620
rect 48865 -7740 48985 -7620
rect 49030 -7740 49150 -7620
rect 49205 -7740 49325 -7620
rect 49370 -7740 49490 -7620
rect 49535 -7740 49655 -7620
rect 49700 -7740 49820 -7620
rect 49875 -7740 49995 -7620
rect 50040 -7740 50160 -7620
rect 50205 -7740 50325 -7620
rect 50370 -7740 50490 -7620
rect 50545 -7740 50665 -7620
rect 50710 -7740 50830 -7620
rect 50875 -7740 50995 -7620
rect 51040 -7740 51160 -7620
rect 51215 -7740 51335 -7620
rect 51380 -7740 51500 -7620
rect 51545 -7740 51665 -7620
rect 51710 -7740 51830 -7620
rect 51885 -7740 52005 -7620
rect 52050 -7740 52170 -7620
rect 52215 -7740 52335 -7620
rect 52380 -7740 52500 -7620
rect 52555 -7740 52675 -7620
rect 52720 -7740 52840 -7620
rect 52885 -7740 53005 -7620
rect 53050 -7740 53170 -7620
rect 53225 -7740 53345 -7620
rect 47865 -7915 47985 -7795
rect 48030 -7915 48150 -7795
rect 48195 -7915 48315 -7795
rect 48360 -7915 48480 -7795
rect 48535 -7915 48655 -7795
rect 48700 -7915 48820 -7795
rect 48865 -7915 48985 -7795
rect 49030 -7915 49150 -7795
rect 49205 -7915 49325 -7795
rect 49370 -7915 49490 -7795
rect 49535 -7915 49655 -7795
rect 49700 -7915 49820 -7795
rect 49875 -7915 49995 -7795
rect 50040 -7915 50160 -7795
rect 50205 -7915 50325 -7795
rect 50370 -7915 50490 -7795
rect 50545 -7915 50665 -7795
rect 50710 -7915 50830 -7795
rect 50875 -7915 50995 -7795
rect 51040 -7915 51160 -7795
rect 51215 -7915 51335 -7795
rect 51380 -7915 51500 -7795
rect 51545 -7915 51665 -7795
rect 51710 -7915 51830 -7795
rect 51885 -7915 52005 -7795
rect 52050 -7915 52170 -7795
rect 52215 -7915 52335 -7795
rect 52380 -7915 52500 -7795
rect 52555 -7915 52675 -7795
rect 52720 -7915 52840 -7795
rect 52885 -7915 53005 -7795
rect 53050 -7915 53170 -7795
rect 53225 -7915 53345 -7795
rect 47865 -8080 47985 -7960
rect 48030 -8080 48150 -7960
rect 48195 -8080 48315 -7960
rect 48360 -8080 48480 -7960
rect 48535 -8080 48655 -7960
rect 48700 -8080 48820 -7960
rect 48865 -8080 48985 -7960
rect 49030 -8080 49150 -7960
rect 49205 -8080 49325 -7960
rect 49370 -8080 49490 -7960
rect 49535 -8080 49655 -7960
rect 49700 -8080 49820 -7960
rect 49875 -8080 49995 -7960
rect 50040 -8080 50160 -7960
rect 50205 -8080 50325 -7960
rect 50370 -8080 50490 -7960
rect 50545 -8080 50665 -7960
rect 50710 -8080 50830 -7960
rect 50875 -8080 50995 -7960
rect 51040 -8080 51160 -7960
rect 51215 -8080 51335 -7960
rect 51380 -8080 51500 -7960
rect 51545 -8080 51665 -7960
rect 51710 -8080 51830 -7960
rect 51885 -8080 52005 -7960
rect 52050 -8080 52170 -7960
rect 52215 -8080 52335 -7960
rect 52380 -8080 52500 -7960
rect 52555 -8080 52675 -7960
rect 52720 -8080 52840 -7960
rect 52885 -8080 53005 -7960
rect 53050 -8080 53170 -7960
rect 53225 -8080 53345 -7960
rect 47865 -8245 47985 -8125
rect 48030 -8245 48150 -8125
rect 48195 -8245 48315 -8125
rect 48360 -8245 48480 -8125
rect 48535 -8245 48655 -8125
rect 48700 -8245 48820 -8125
rect 48865 -8245 48985 -8125
rect 49030 -8245 49150 -8125
rect 49205 -8245 49325 -8125
rect 49370 -8245 49490 -8125
rect 49535 -8245 49655 -8125
rect 49700 -8245 49820 -8125
rect 49875 -8245 49995 -8125
rect 50040 -8245 50160 -8125
rect 50205 -8245 50325 -8125
rect 50370 -8245 50490 -8125
rect 50545 -8245 50665 -8125
rect 50710 -8245 50830 -8125
rect 50875 -8245 50995 -8125
rect 51040 -8245 51160 -8125
rect 51215 -8245 51335 -8125
rect 51380 -8245 51500 -8125
rect 51545 -8245 51665 -8125
rect 51710 -8245 51830 -8125
rect 51885 -8245 52005 -8125
rect 52050 -8245 52170 -8125
rect 52215 -8245 52335 -8125
rect 52380 -8245 52500 -8125
rect 52555 -8245 52675 -8125
rect 52720 -8245 52840 -8125
rect 52885 -8245 53005 -8125
rect 53050 -8245 53170 -8125
rect 53225 -8245 53345 -8125
rect 47865 -8410 47985 -8290
rect 48030 -8410 48150 -8290
rect 48195 -8410 48315 -8290
rect 48360 -8410 48480 -8290
rect 48535 -8410 48655 -8290
rect 48700 -8410 48820 -8290
rect 48865 -8410 48985 -8290
rect 49030 -8410 49150 -8290
rect 49205 -8410 49325 -8290
rect 49370 -8410 49490 -8290
rect 49535 -8410 49655 -8290
rect 49700 -8410 49820 -8290
rect 49875 -8410 49995 -8290
rect 50040 -8410 50160 -8290
rect 50205 -8410 50325 -8290
rect 50370 -8410 50490 -8290
rect 50545 -8410 50665 -8290
rect 50710 -8410 50830 -8290
rect 50875 -8410 50995 -8290
rect 51040 -8410 51160 -8290
rect 51215 -8410 51335 -8290
rect 51380 -8410 51500 -8290
rect 51545 -8410 51665 -8290
rect 51710 -8410 51830 -8290
rect 51885 -8410 52005 -8290
rect 52050 -8410 52170 -8290
rect 52215 -8410 52335 -8290
rect 52380 -8410 52500 -8290
rect 52555 -8410 52675 -8290
rect 52720 -8410 52840 -8290
rect 52885 -8410 53005 -8290
rect 53050 -8410 53170 -8290
rect 53225 -8410 53345 -8290
rect 47865 -8585 47985 -8465
rect 48030 -8585 48150 -8465
rect 48195 -8585 48315 -8465
rect 48360 -8585 48480 -8465
rect 48535 -8585 48655 -8465
rect 48700 -8585 48820 -8465
rect 48865 -8585 48985 -8465
rect 49030 -8585 49150 -8465
rect 49205 -8585 49325 -8465
rect 49370 -8585 49490 -8465
rect 49535 -8585 49655 -8465
rect 49700 -8585 49820 -8465
rect 49875 -8585 49995 -8465
rect 50040 -8585 50160 -8465
rect 50205 -8585 50325 -8465
rect 50370 -8585 50490 -8465
rect 50545 -8585 50665 -8465
rect 50710 -8585 50830 -8465
rect 50875 -8585 50995 -8465
rect 51040 -8585 51160 -8465
rect 51215 -8585 51335 -8465
rect 51380 -8585 51500 -8465
rect 51545 -8585 51665 -8465
rect 51710 -8585 51830 -8465
rect 51885 -8585 52005 -8465
rect 52050 -8585 52170 -8465
rect 52215 -8585 52335 -8465
rect 52380 -8585 52500 -8465
rect 52555 -8585 52675 -8465
rect 52720 -8585 52840 -8465
rect 52885 -8585 53005 -8465
rect 53050 -8585 53170 -8465
rect 53225 -8585 53345 -8465
rect 47865 -8750 47985 -8630
rect 48030 -8750 48150 -8630
rect 48195 -8750 48315 -8630
rect 48360 -8750 48480 -8630
rect 48535 -8750 48655 -8630
rect 48700 -8750 48820 -8630
rect 48865 -8750 48985 -8630
rect 49030 -8750 49150 -8630
rect 49205 -8750 49325 -8630
rect 49370 -8750 49490 -8630
rect 49535 -8750 49655 -8630
rect 49700 -8750 49820 -8630
rect 49875 -8750 49995 -8630
rect 50040 -8750 50160 -8630
rect 50205 -8750 50325 -8630
rect 50370 -8750 50490 -8630
rect 50545 -8750 50665 -8630
rect 50710 -8750 50830 -8630
rect 50875 -8750 50995 -8630
rect 51040 -8750 51160 -8630
rect 51215 -8750 51335 -8630
rect 51380 -8750 51500 -8630
rect 51545 -8750 51665 -8630
rect 51710 -8750 51830 -8630
rect 51885 -8750 52005 -8630
rect 52050 -8750 52170 -8630
rect 52215 -8750 52335 -8630
rect 52380 -8750 52500 -8630
rect 52555 -8750 52675 -8630
rect 52720 -8750 52840 -8630
rect 52885 -8750 53005 -8630
rect 53050 -8750 53170 -8630
rect 53225 -8750 53345 -8630
rect 47865 -8915 47985 -8795
rect 48030 -8915 48150 -8795
rect 48195 -8915 48315 -8795
rect 48360 -8915 48480 -8795
rect 48535 -8915 48655 -8795
rect 48700 -8915 48820 -8795
rect 48865 -8915 48985 -8795
rect 49030 -8915 49150 -8795
rect 49205 -8915 49325 -8795
rect 49370 -8915 49490 -8795
rect 49535 -8915 49655 -8795
rect 49700 -8915 49820 -8795
rect 49875 -8915 49995 -8795
rect 50040 -8915 50160 -8795
rect 50205 -8915 50325 -8795
rect 50370 -8915 50490 -8795
rect 50545 -8915 50665 -8795
rect 50710 -8915 50830 -8795
rect 50875 -8915 50995 -8795
rect 51040 -8915 51160 -8795
rect 51215 -8915 51335 -8795
rect 51380 -8915 51500 -8795
rect 51545 -8915 51665 -8795
rect 51710 -8915 51830 -8795
rect 51885 -8915 52005 -8795
rect 52050 -8915 52170 -8795
rect 52215 -8915 52335 -8795
rect 52380 -8915 52500 -8795
rect 52555 -8915 52675 -8795
rect 52720 -8915 52840 -8795
rect 52885 -8915 53005 -8795
rect 53050 -8915 53170 -8795
rect 53225 -8915 53345 -8795
rect 47865 -9080 47985 -8960
rect 48030 -9080 48150 -8960
rect 48195 -9080 48315 -8960
rect 48360 -9080 48480 -8960
rect 48535 -9080 48655 -8960
rect 48700 -9080 48820 -8960
rect 48865 -9080 48985 -8960
rect 49030 -9080 49150 -8960
rect 49205 -9080 49325 -8960
rect 49370 -9080 49490 -8960
rect 49535 -9080 49655 -8960
rect 49700 -9080 49820 -8960
rect 49875 -9080 49995 -8960
rect 50040 -9080 50160 -8960
rect 50205 -9080 50325 -8960
rect 50370 -9080 50490 -8960
rect 50545 -9080 50665 -8960
rect 50710 -9080 50830 -8960
rect 50875 -9080 50995 -8960
rect 51040 -9080 51160 -8960
rect 51215 -9080 51335 -8960
rect 51380 -9080 51500 -8960
rect 51545 -9080 51665 -8960
rect 51710 -9080 51830 -8960
rect 51885 -9080 52005 -8960
rect 52050 -9080 52170 -8960
rect 52215 -9080 52335 -8960
rect 52380 -9080 52500 -8960
rect 52555 -9080 52675 -8960
rect 52720 -9080 52840 -8960
rect 52885 -9080 53005 -8960
rect 53050 -9080 53170 -8960
rect 53225 -9080 53345 -8960
rect 47865 -9255 47985 -9135
rect 48030 -9255 48150 -9135
rect 48195 -9255 48315 -9135
rect 48360 -9255 48480 -9135
rect 48535 -9255 48655 -9135
rect 48700 -9255 48820 -9135
rect 48865 -9255 48985 -9135
rect 49030 -9255 49150 -9135
rect 49205 -9255 49325 -9135
rect 49370 -9255 49490 -9135
rect 49535 -9255 49655 -9135
rect 49700 -9255 49820 -9135
rect 49875 -9255 49995 -9135
rect 50040 -9255 50160 -9135
rect 50205 -9255 50325 -9135
rect 50370 -9255 50490 -9135
rect 50545 -9255 50665 -9135
rect 50710 -9255 50830 -9135
rect 50875 -9255 50995 -9135
rect 51040 -9255 51160 -9135
rect 51215 -9255 51335 -9135
rect 51380 -9255 51500 -9135
rect 51545 -9255 51665 -9135
rect 51710 -9255 51830 -9135
rect 51885 -9255 52005 -9135
rect 52050 -9255 52170 -9135
rect 52215 -9255 52335 -9135
rect 52380 -9255 52500 -9135
rect 52555 -9255 52675 -9135
rect 52720 -9255 52840 -9135
rect 52885 -9255 53005 -9135
rect 53050 -9255 53170 -9135
rect 53225 -9255 53345 -9135
rect 47865 -9420 47985 -9300
rect 48030 -9420 48150 -9300
rect 48195 -9420 48315 -9300
rect 48360 -9420 48480 -9300
rect 48535 -9420 48655 -9300
rect 48700 -9420 48820 -9300
rect 48865 -9420 48985 -9300
rect 49030 -9420 49150 -9300
rect 49205 -9420 49325 -9300
rect 49370 -9420 49490 -9300
rect 49535 -9420 49655 -9300
rect 49700 -9420 49820 -9300
rect 49875 -9420 49995 -9300
rect 50040 -9420 50160 -9300
rect 50205 -9420 50325 -9300
rect 50370 -9420 50490 -9300
rect 50545 -9420 50665 -9300
rect 50710 -9420 50830 -9300
rect 50875 -9420 50995 -9300
rect 51040 -9420 51160 -9300
rect 51215 -9420 51335 -9300
rect 51380 -9420 51500 -9300
rect 51545 -9420 51665 -9300
rect 51710 -9420 51830 -9300
rect 51885 -9420 52005 -9300
rect 52050 -9420 52170 -9300
rect 52215 -9420 52335 -9300
rect 52380 -9420 52500 -9300
rect 52555 -9420 52675 -9300
rect 52720 -9420 52840 -9300
rect 52885 -9420 53005 -9300
rect 53050 -9420 53170 -9300
rect 53225 -9420 53345 -9300
rect 47865 -9585 47985 -9465
rect 48030 -9585 48150 -9465
rect 48195 -9585 48315 -9465
rect 48360 -9585 48480 -9465
rect 48535 -9585 48655 -9465
rect 48700 -9585 48820 -9465
rect 48865 -9585 48985 -9465
rect 49030 -9585 49150 -9465
rect 49205 -9585 49325 -9465
rect 49370 -9585 49490 -9465
rect 49535 -9585 49655 -9465
rect 49700 -9585 49820 -9465
rect 49875 -9585 49995 -9465
rect 50040 -9585 50160 -9465
rect 50205 -9585 50325 -9465
rect 50370 -9585 50490 -9465
rect 50545 -9585 50665 -9465
rect 50710 -9585 50830 -9465
rect 50875 -9585 50995 -9465
rect 51040 -9585 51160 -9465
rect 51215 -9585 51335 -9465
rect 51380 -9585 51500 -9465
rect 51545 -9585 51665 -9465
rect 51710 -9585 51830 -9465
rect 51885 -9585 52005 -9465
rect 52050 -9585 52170 -9465
rect 52215 -9585 52335 -9465
rect 52380 -9585 52500 -9465
rect 52555 -9585 52675 -9465
rect 52720 -9585 52840 -9465
rect 52885 -9585 53005 -9465
rect 53050 -9585 53170 -9465
rect 53225 -9585 53345 -9465
rect 47865 -9750 47985 -9630
rect 48030 -9750 48150 -9630
rect 48195 -9750 48315 -9630
rect 48360 -9750 48480 -9630
rect 48535 -9750 48655 -9630
rect 48700 -9750 48820 -9630
rect 48865 -9750 48985 -9630
rect 49030 -9750 49150 -9630
rect 49205 -9750 49325 -9630
rect 49370 -9750 49490 -9630
rect 49535 -9750 49655 -9630
rect 49700 -9750 49820 -9630
rect 49875 -9750 49995 -9630
rect 50040 -9750 50160 -9630
rect 50205 -9750 50325 -9630
rect 50370 -9750 50490 -9630
rect 50545 -9750 50665 -9630
rect 50710 -9750 50830 -9630
rect 50875 -9750 50995 -9630
rect 51040 -9750 51160 -9630
rect 51215 -9750 51335 -9630
rect 51380 -9750 51500 -9630
rect 51545 -9750 51665 -9630
rect 51710 -9750 51830 -9630
rect 51885 -9750 52005 -9630
rect 52050 -9750 52170 -9630
rect 52215 -9750 52335 -9630
rect 52380 -9750 52500 -9630
rect 52555 -9750 52675 -9630
rect 52720 -9750 52840 -9630
rect 52885 -9750 53005 -9630
rect 53050 -9750 53170 -9630
rect 53225 -9750 53345 -9630
rect 30795 -10170 30915 -10050
rect 30970 -10170 31090 -10050
rect 31135 -10170 31255 -10050
rect 31300 -10170 31420 -10050
rect 31465 -10170 31585 -10050
rect 31640 -10170 31760 -10050
rect 31805 -10170 31925 -10050
rect 31970 -10170 32090 -10050
rect 32135 -10170 32255 -10050
rect 32310 -10170 32430 -10050
rect 32475 -10170 32595 -10050
rect 32640 -10170 32760 -10050
rect 32805 -10170 32925 -10050
rect 32980 -10170 33100 -10050
rect 33145 -10170 33265 -10050
rect 33310 -10170 33430 -10050
rect 33475 -10170 33595 -10050
rect 33650 -10170 33770 -10050
rect 33815 -10170 33935 -10050
rect 33980 -10170 34100 -10050
rect 34145 -10170 34265 -10050
rect 34320 -10170 34440 -10050
rect 34485 -10170 34605 -10050
rect 34650 -10170 34770 -10050
rect 34815 -10170 34935 -10050
rect 34990 -10170 35110 -10050
rect 35155 -10170 35275 -10050
rect 35320 -10170 35440 -10050
rect 35485 -10170 35605 -10050
rect 35660 -10170 35780 -10050
rect 35825 -10170 35945 -10050
rect 35990 -10170 36110 -10050
rect 36155 -10170 36275 -10050
rect 30795 -10335 30915 -10215
rect 30970 -10335 31090 -10215
rect 31135 -10335 31255 -10215
rect 31300 -10335 31420 -10215
rect 31465 -10335 31585 -10215
rect 31640 -10335 31760 -10215
rect 31805 -10335 31925 -10215
rect 31970 -10335 32090 -10215
rect 32135 -10335 32255 -10215
rect 32310 -10335 32430 -10215
rect 32475 -10335 32595 -10215
rect 32640 -10335 32760 -10215
rect 32805 -10335 32925 -10215
rect 32980 -10335 33100 -10215
rect 33145 -10335 33265 -10215
rect 33310 -10335 33430 -10215
rect 33475 -10335 33595 -10215
rect 33650 -10335 33770 -10215
rect 33815 -10335 33935 -10215
rect 33980 -10335 34100 -10215
rect 34145 -10335 34265 -10215
rect 34320 -10335 34440 -10215
rect 34485 -10335 34605 -10215
rect 34650 -10335 34770 -10215
rect 34815 -10335 34935 -10215
rect 34990 -10335 35110 -10215
rect 35155 -10335 35275 -10215
rect 35320 -10335 35440 -10215
rect 35485 -10335 35605 -10215
rect 35660 -10335 35780 -10215
rect 35825 -10335 35945 -10215
rect 35990 -10335 36110 -10215
rect 36155 -10335 36275 -10215
rect 30795 -10500 30915 -10380
rect 30970 -10500 31090 -10380
rect 31135 -10500 31255 -10380
rect 31300 -10500 31420 -10380
rect 31465 -10500 31585 -10380
rect 31640 -10500 31760 -10380
rect 31805 -10500 31925 -10380
rect 31970 -10500 32090 -10380
rect 32135 -10500 32255 -10380
rect 32310 -10500 32430 -10380
rect 32475 -10500 32595 -10380
rect 32640 -10500 32760 -10380
rect 32805 -10500 32925 -10380
rect 32980 -10500 33100 -10380
rect 33145 -10500 33265 -10380
rect 33310 -10500 33430 -10380
rect 33475 -10500 33595 -10380
rect 33650 -10500 33770 -10380
rect 33815 -10500 33935 -10380
rect 33980 -10500 34100 -10380
rect 34145 -10500 34265 -10380
rect 34320 -10500 34440 -10380
rect 34485 -10500 34605 -10380
rect 34650 -10500 34770 -10380
rect 34815 -10500 34935 -10380
rect 34990 -10500 35110 -10380
rect 35155 -10500 35275 -10380
rect 35320 -10500 35440 -10380
rect 35485 -10500 35605 -10380
rect 35660 -10500 35780 -10380
rect 35825 -10500 35945 -10380
rect 35990 -10500 36110 -10380
rect 36155 -10500 36275 -10380
rect 30795 -10665 30915 -10545
rect 30970 -10665 31090 -10545
rect 31135 -10665 31255 -10545
rect 31300 -10665 31420 -10545
rect 31465 -10665 31585 -10545
rect 31640 -10665 31760 -10545
rect 31805 -10665 31925 -10545
rect 31970 -10665 32090 -10545
rect 32135 -10665 32255 -10545
rect 32310 -10665 32430 -10545
rect 32475 -10665 32595 -10545
rect 32640 -10665 32760 -10545
rect 32805 -10665 32925 -10545
rect 32980 -10665 33100 -10545
rect 33145 -10665 33265 -10545
rect 33310 -10665 33430 -10545
rect 33475 -10665 33595 -10545
rect 33650 -10665 33770 -10545
rect 33815 -10665 33935 -10545
rect 33980 -10665 34100 -10545
rect 34145 -10665 34265 -10545
rect 34320 -10665 34440 -10545
rect 34485 -10665 34605 -10545
rect 34650 -10665 34770 -10545
rect 34815 -10665 34935 -10545
rect 34990 -10665 35110 -10545
rect 35155 -10665 35275 -10545
rect 35320 -10665 35440 -10545
rect 35485 -10665 35605 -10545
rect 35660 -10665 35780 -10545
rect 35825 -10665 35945 -10545
rect 35990 -10665 36110 -10545
rect 36155 -10665 36275 -10545
rect 30795 -10840 30915 -10720
rect 30970 -10840 31090 -10720
rect 31135 -10840 31255 -10720
rect 31300 -10840 31420 -10720
rect 31465 -10840 31585 -10720
rect 31640 -10840 31760 -10720
rect 31805 -10840 31925 -10720
rect 31970 -10840 32090 -10720
rect 32135 -10840 32255 -10720
rect 32310 -10840 32430 -10720
rect 32475 -10840 32595 -10720
rect 32640 -10840 32760 -10720
rect 32805 -10840 32925 -10720
rect 32980 -10840 33100 -10720
rect 33145 -10840 33265 -10720
rect 33310 -10840 33430 -10720
rect 33475 -10840 33595 -10720
rect 33650 -10840 33770 -10720
rect 33815 -10840 33935 -10720
rect 33980 -10840 34100 -10720
rect 34145 -10840 34265 -10720
rect 34320 -10840 34440 -10720
rect 34485 -10840 34605 -10720
rect 34650 -10840 34770 -10720
rect 34815 -10840 34935 -10720
rect 34990 -10840 35110 -10720
rect 35155 -10840 35275 -10720
rect 35320 -10840 35440 -10720
rect 35485 -10840 35605 -10720
rect 35660 -10840 35780 -10720
rect 35825 -10840 35945 -10720
rect 35990 -10840 36110 -10720
rect 36155 -10840 36275 -10720
rect 30795 -11005 30915 -10885
rect 30970 -11005 31090 -10885
rect 31135 -11005 31255 -10885
rect 31300 -11005 31420 -10885
rect 31465 -11005 31585 -10885
rect 31640 -11005 31760 -10885
rect 31805 -11005 31925 -10885
rect 31970 -11005 32090 -10885
rect 32135 -11005 32255 -10885
rect 32310 -11005 32430 -10885
rect 32475 -11005 32595 -10885
rect 32640 -11005 32760 -10885
rect 32805 -11005 32925 -10885
rect 32980 -11005 33100 -10885
rect 33145 -11005 33265 -10885
rect 33310 -11005 33430 -10885
rect 33475 -11005 33595 -10885
rect 33650 -11005 33770 -10885
rect 33815 -11005 33935 -10885
rect 33980 -11005 34100 -10885
rect 34145 -11005 34265 -10885
rect 34320 -11005 34440 -10885
rect 34485 -11005 34605 -10885
rect 34650 -11005 34770 -10885
rect 34815 -11005 34935 -10885
rect 34990 -11005 35110 -10885
rect 35155 -11005 35275 -10885
rect 35320 -11005 35440 -10885
rect 35485 -11005 35605 -10885
rect 35660 -11005 35780 -10885
rect 35825 -11005 35945 -10885
rect 35990 -11005 36110 -10885
rect 36155 -11005 36275 -10885
rect 30795 -11170 30915 -11050
rect 30970 -11170 31090 -11050
rect 31135 -11170 31255 -11050
rect 31300 -11170 31420 -11050
rect 31465 -11170 31585 -11050
rect 31640 -11170 31760 -11050
rect 31805 -11170 31925 -11050
rect 31970 -11170 32090 -11050
rect 32135 -11170 32255 -11050
rect 32310 -11170 32430 -11050
rect 32475 -11170 32595 -11050
rect 32640 -11170 32760 -11050
rect 32805 -11170 32925 -11050
rect 32980 -11170 33100 -11050
rect 33145 -11170 33265 -11050
rect 33310 -11170 33430 -11050
rect 33475 -11170 33595 -11050
rect 33650 -11170 33770 -11050
rect 33815 -11170 33935 -11050
rect 33980 -11170 34100 -11050
rect 34145 -11170 34265 -11050
rect 34320 -11170 34440 -11050
rect 34485 -11170 34605 -11050
rect 34650 -11170 34770 -11050
rect 34815 -11170 34935 -11050
rect 34990 -11170 35110 -11050
rect 35155 -11170 35275 -11050
rect 35320 -11170 35440 -11050
rect 35485 -11170 35605 -11050
rect 35660 -11170 35780 -11050
rect 35825 -11170 35945 -11050
rect 35990 -11170 36110 -11050
rect 36155 -11170 36275 -11050
rect 30795 -11335 30915 -11215
rect 30970 -11335 31090 -11215
rect 31135 -11335 31255 -11215
rect 31300 -11335 31420 -11215
rect 31465 -11335 31585 -11215
rect 31640 -11335 31760 -11215
rect 31805 -11335 31925 -11215
rect 31970 -11335 32090 -11215
rect 32135 -11335 32255 -11215
rect 32310 -11335 32430 -11215
rect 32475 -11335 32595 -11215
rect 32640 -11335 32760 -11215
rect 32805 -11335 32925 -11215
rect 32980 -11335 33100 -11215
rect 33145 -11335 33265 -11215
rect 33310 -11335 33430 -11215
rect 33475 -11335 33595 -11215
rect 33650 -11335 33770 -11215
rect 33815 -11335 33935 -11215
rect 33980 -11335 34100 -11215
rect 34145 -11335 34265 -11215
rect 34320 -11335 34440 -11215
rect 34485 -11335 34605 -11215
rect 34650 -11335 34770 -11215
rect 34815 -11335 34935 -11215
rect 34990 -11335 35110 -11215
rect 35155 -11335 35275 -11215
rect 35320 -11335 35440 -11215
rect 35485 -11335 35605 -11215
rect 35660 -11335 35780 -11215
rect 35825 -11335 35945 -11215
rect 35990 -11335 36110 -11215
rect 36155 -11335 36275 -11215
rect 30795 -11510 30915 -11390
rect 30970 -11510 31090 -11390
rect 31135 -11510 31255 -11390
rect 31300 -11510 31420 -11390
rect 31465 -11510 31585 -11390
rect 31640 -11510 31760 -11390
rect 31805 -11510 31925 -11390
rect 31970 -11510 32090 -11390
rect 32135 -11510 32255 -11390
rect 32310 -11510 32430 -11390
rect 32475 -11510 32595 -11390
rect 32640 -11510 32760 -11390
rect 32805 -11510 32925 -11390
rect 32980 -11510 33100 -11390
rect 33145 -11510 33265 -11390
rect 33310 -11510 33430 -11390
rect 33475 -11510 33595 -11390
rect 33650 -11510 33770 -11390
rect 33815 -11510 33935 -11390
rect 33980 -11510 34100 -11390
rect 34145 -11510 34265 -11390
rect 34320 -11510 34440 -11390
rect 34485 -11510 34605 -11390
rect 34650 -11510 34770 -11390
rect 34815 -11510 34935 -11390
rect 34990 -11510 35110 -11390
rect 35155 -11510 35275 -11390
rect 35320 -11510 35440 -11390
rect 35485 -11510 35605 -11390
rect 35660 -11510 35780 -11390
rect 35825 -11510 35945 -11390
rect 35990 -11510 36110 -11390
rect 36155 -11510 36275 -11390
rect 30795 -11675 30915 -11555
rect 30970 -11675 31090 -11555
rect 31135 -11675 31255 -11555
rect 31300 -11675 31420 -11555
rect 31465 -11675 31585 -11555
rect 31640 -11675 31760 -11555
rect 31805 -11675 31925 -11555
rect 31970 -11675 32090 -11555
rect 32135 -11675 32255 -11555
rect 32310 -11675 32430 -11555
rect 32475 -11675 32595 -11555
rect 32640 -11675 32760 -11555
rect 32805 -11675 32925 -11555
rect 32980 -11675 33100 -11555
rect 33145 -11675 33265 -11555
rect 33310 -11675 33430 -11555
rect 33475 -11675 33595 -11555
rect 33650 -11675 33770 -11555
rect 33815 -11675 33935 -11555
rect 33980 -11675 34100 -11555
rect 34145 -11675 34265 -11555
rect 34320 -11675 34440 -11555
rect 34485 -11675 34605 -11555
rect 34650 -11675 34770 -11555
rect 34815 -11675 34935 -11555
rect 34990 -11675 35110 -11555
rect 35155 -11675 35275 -11555
rect 35320 -11675 35440 -11555
rect 35485 -11675 35605 -11555
rect 35660 -11675 35780 -11555
rect 35825 -11675 35945 -11555
rect 35990 -11675 36110 -11555
rect 36155 -11675 36275 -11555
rect 30795 -11840 30915 -11720
rect 30970 -11840 31090 -11720
rect 31135 -11840 31255 -11720
rect 31300 -11840 31420 -11720
rect 31465 -11840 31585 -11720
rect 31640 -11840 31760 -11720
rect 31805 -11840 31925 -11720
rect 31970 -11840 32090 -11720
rect 32135 -11840 32255 -11720
rect 32310 -11840 32430 -11720
rect 32475 -11840 32595 -11720
rect 32640 -11840 32760 -11720
rect 32805 -11840 32925 -11720
rect 32980 -11840 33100 -11720
rect 33145 -11840 33265 -11720
rect 33310 -11840 33430 -11720
rect 33475 -11840 33595 -11720
rect 33650 -11840 33770 -11720
rect 33815 -11840 33935 -11720
rect 33980 -11840 34100 -11720
rect 34145 -11840 34265 -11720
rect 34320 -11840 34440 -11720
rect 34485 -11840 34605 -11720
rect 34650 -11840 34770 -11720
rect 34815 -11840 34935 -11720
rect 34990 -11840 35110 -11720
rect 35155 -11840 35275 -11720
rect 35320 -11840 35440 -11720
rect 35485 -11840 35605 -11720
rect 35660 -11840 35780 -11720
rect 35825 -11840 35945 -11720
rect 35990 -11840 36110 -11720
rect 36155 -11840 36275 -11720
rect 30795 -12005 30915 -11885
rect 30970 -12005 31090 -11885
rect 31135 -12005 31255 -11885
rect 31300 -12005 31420 -11885
rect 31465 -12005 31585 -11885
rect 31640 -12005 31760 -11885
rect 31805 -12005 31925 -11885
rect 31970 -12005 32090 -11885
rect 32135 -12005 32255 -11885
rect 32310 -12005 32430 -11885
rect 32475 -12005 32595 -11885
rect 32640 -12005 32760 -11885
rect 32805 -12005 32925 -11885
rect 32980 -12005 33100 -11885
rect 33145 -12005 33265 -11885
rect 33310 -12005 33430 -11885
rect 33475 -12005 33595 -11885
rect 33650 -12005 33770 -11885
rect 33815 -12005 33935 -11885
rect 33980 -12005 34100 -11885
rect 34145 -12005 34265 -11885
rect 34320 -12005 34440 -11885
rect 34485 -12005 34605 -11885
rect 34650 -12005 34770 -11885
rect 34815 -12005 34935 -11885
rect 34990 -12005 35110 -11885
rect 35155 -12005 35275 -11885
rect 35320 -12005 35440 -11885
rect 35485 -12005 35605 -11885
rect 35660 -12005 35780 -11885
rect 35825 -12005 35945 -11885
rect 35990 -12005 36110 -11885
rect 36155 -12005 36275 -11885
rect 30795 -12180 30915 -12060
rect 30970 -12180 31090 -12060
rect 31135 -12180 31255 -12060
rect 31300 -12180 31420 -12060
rect 31465 -12180 31585 -12060
rect 31640 -12180 31760 -12060
rect 31805 -12180 31925 -12060
rect 31970 -12180 32090 -12060
rect 32135 -12180 32255 -12060
rect 32310 -12180 32430 -12060
rect 32475 -12180 32595 -12060
rect 32640 -12180 32760 -12060
rect 32805 -12180 32925 -12060
rect 32980 -12180 33100 -12060
rect 33145 -12180 33265 -12060
rect 33310 -12180 33430 -12060
rect 33475 -12180 33595 -12060
rect 33650 -12180 33770 -12060
rect 33815 -12180 33935 -12060
rect 33980 -12180 34100 -12060
rect 34145 -12180 34265 -12060
rect 34320 -12180 34440 -12060
rect 34485 -12180 34605 -12060
rect 34650 -12180 34770 -12060
rect 34815 -12180 34935 -12060
rect 34990 -12180 35110 -12060
rect 35155 -12180 35275 -12060
rect 35320 -12180 35440 -12060
rect 35485 -12180 35605 -12060
rect 35660 -12180 35780 -12060
rect 35825 -12180 35945 -12060
rect 35990 -12180 36110 -12060
rect 36155 -12180 36275 -12060
rect 30795 -12345 30915 -12225
rect 30970 -12345 31090 -12225
rect 31135 -12345 31255 -12225
rect 31300 -12345 31420 -12225
rect 31465 -12345 31585 -12225
rect 31640 -12345 31760 -12225
rect 31805 -12345 31925 -12225
rect 31970 -12345 32090 -12225
rect 32135 -12345 32255 -12225
rect 32310 -12345 32430 -12225
rect 32475 -12345 32595 -12225
rect 32640 -12345 32760 -12225
rect 32805 -12345 32925 -12225
rect 32980 -12345 33100 -12225
rect 33145 -12345 33265 -12225
rect 33310 -12345 33430 -12225
rect 33475 -12345 33595 -12225
rect 33650 -12345 33770 -12225
rect 33815 -12345 33935 -12225
rect 33980 -12345 34100 -12225
rect 34145 -12345 34265 -12225
rect 34320 -12345 34440 -12225
rect 34485 -12345 34605 -12225
rect 34650 -12345 34770 -12225
rect 34815 -12345 34935 -12225
rect 34990 -12345 35110 -12225
rect 35155 -12345 35275 -12225
rect 35320 -12345 35440 -12225
rect 35485 -12345 35605 -12225
rect 35660 -12345 35780 -12225
rect 35825 -12345 35945 -12225
rect 35990 -12345 36110 -12225
rect 36155 -12345 36275 -12225
rect 30795 -12510 30915 -12390
rect 30970 -12510 31090 -12390
rect 31135 -12510 31255 -12390
rect 31300 -12510 31420 -12390
rect 31465 -12510 31585 -12390
rect 31640 -12510 31760 -12390
rect 31805 -12510 31925 -12390
rect 31970 -12510 32090 -12390
rect 32135 -12510 32255 -12390
rect 32310 -12510 32430 -12390
rect 32475 -12510 32595 -12390
rect 32640 -12510 32760 -12390
rect 32805 -12510 32925 -12390
rect 32980 -12510 33100 -12390
rect 33145 -12510 33265 -12390
rect 33310 -12510 33430 -12390
rect 33475 -12510 33595 -12390
rect 33650 -12510 33770 -12390
rect 33815 -12510 33935 -12390
rect 33980 -12510 34100 -12390
rect 34145 -12510 34265 -12390
rect 34320 -12510 34440 -12390
rect 34485 -12510 34605 -12390
rect 34650 -12510 34770 -12390
rect 34815 -12510 34935 -12390
rect 34990 -12510 35110 -12390
rect 35155 -12510 35275 -12390
rect 35320 -12510 35440 -12390
rect 35485 -12510 35605 -12390
rect 35660 -12510 35780 -12390
rect 35825 -12510 35945 -12390
rect 35990 -12510 36110 -12390
rect 36155 -12510 36275 -12390
rect 30795 -12675 30915 -12555
rect 30970 -12675 31090 -12555
rect 31135 -12675 31255 -12555
rect 31300 -12675 31420 -12555
rect 31465 -12675 31585 -12555
rect 31640 -12675 31760 -12555
rect 31805 -12675 31925 -12555
rect 31970 -12675 32090 -12555
rect 32135 -12675 32255 -12555
rect 32310 -12675 32430 -12555
rect 32475 -12675 32595 -12555
rect 32640 -12675 32760 -12555
rect 32805 -12675 32925 -12555
rect 32980 -12675 33100 -12555
rect 33145 -12675 33265 -12555
rect 33310 -12675 33430 -12555
rect 33475 -12675 33595 -12555
rect 33650 -12675 33770 -12555
rect 33815 -12675 33935 -12555
rect 33980 -12675 34100 -12555
rect 34145 -12675 34265 -12555
rect 34320 -12675 34440 -12555
rect 34485 -12675 34605 -12555
rect 34650 -12675 34770 -12555
rect 34815 -12675 34935 -12555
rect 34990 -12675 35110 -12555
rect 35155 -12675 35275 -12555
rect 35320 -12675 35440 -12555
rect 35485 -12675 35605 -12555
rect 35660 -12675 35780 -12555
rect 35825 -12675 35945 -12555
rect 35990 -12675 36110 -12555
rect 36155 -12675 36275 -12555
rect 30795 -12850 30915 -12730
rect 30970 -12850 31090 -12730
rect 31135 -12850 31255 -12730
rect 31300 -12850 31420 -12730
rect 31465 -12850 31585 -12730
rect 31640 -12850 31760 -12730
rect 31805 -12850 31925 -12730
rect 31970 -12850 32090 -12730
rect 32135 -12850 32255 -12730
rect 32310 -12850 32430 -12730
rect 32475 -12850 32595 -12730
rect 32640 -12850 32760 -12730
rect 32805 -12850 32925 -12730
rect 32980 -12850 33100 -12730
rect 33145 -12850 33265 -12730
rect 33310 -12850 33430 -12730
rect 33475 -12850 33595 -12730
rect 33650 -12850 33770 -12730
rect 33815 -12850 33935 -12730
rect 33980 -12850 34100 -12730
rect 34145 -12850 34265 -12730
rect 34320 -12850 34440 -12730
rect 34485 -12850 34605 -12730
rect 34650 -12850 34770 -12730
rect 34815 -12850 34935 -12730
rect 34990 -12850 35110 -12730
rect 35155 -12850 35275 -12730
rect 35320 -12850 35440 -12730
rect 35485 -12850 35605 -12730
rect 35660 -12850 35780 -12730
rect 35825 -12850 35945 -12730
rect 35990 -12850 36110 -12730
rect 36155 -12850 36275 -12730
rect 30795 -13015 30915 -12895
rect 30970 -13015 31090 -12895
rect 31135 -13015 31255 -12895
rect 31300 -13015 31420 -12895
rect 31465 -13015 31585 -12895
rect 31640 -13015 31760 -12895
rect 31805 -13015 31925 -12895
rect 31970 -13015 32090 -12895
rect 32135 -13015 32255 -12895
rect 32310 -13015 32430 -12895
rect 32475 -13015 32595 -12895
rect 32640 -13015 32760 -12895
rect 32805 -13015 32925 -12895
rect 32980 -13015 33100 -12895
rect 33145 -13015 33265 -12895
rect 33310 -13015 33430 -12895
rect 33475 -13015 33595 -12895
rect 33650 -13015 33770 -12895
rect 33815 -13015 33935 -12895
rect 33980 -13015 34100 -12895
rect 34145 -13015 34265 -12895
rect 34320 -13015 34440 -12895
rect 34485 -13015 34605 -12895
rect 34650 -13015 34770 -12895
rect 34815 -13015 34935 -12895
rect 34990 -13015 35110 -12895
rect 35155 -13015 35275 -12895
rect 35320 -13015 35440 -12895
rect 35485 -13015 35605 -12895
rect 35660 -13015 35780 -12895
rect 35825 -13015 35945 -12895
rect 35990 -13015 36110 -12895
rect 36155 -13015 36275 -12895
rect 30795 -13180 30915 -13060
rect 30970 -13180 31090 -13060
rect 31135 -13180 31255 -13060
rect 31300 -13180 31420 -13060
rect 31465 -13180 31585 -13060
rect 31640 -13180 31760 -13060
rect 31805 -13180 31925 -13060
rect 31970 -13180 32090 -13060
rect 32135 -13180 32255 -13060
rect 32310 -13180 32430 -13060
rect 32475 -13180 32595 -13060
rect 32640 -13180 32760 -13060
rect 32805 -13180 32925 -13060
rect 32980 -13180 33100 -13060
rect 33145 -13180 33265 -13060
rect 33310 -13180 33430 -13060
rect 33475 -13180 33595 -13060
rect 33650 -13180 33770 -13060
rect 33815 -13180 33935 -13060
rect 33980 -13180 34100 -13060
rect 34145 -13180 34265 -13060
rect 34320 -13180 34440 -13060
rect 34485 -13180 34605 -13060
rect 34650 -13180 34770 -13060
rect 34815 -13180 34935 -13060
rect 34990 -13180 35110 -13060
rect 35155 -13180 35275 -13060
rect 35320 -13180 35440 -13060
rect 35485 -13180 35605 -13060
rect 35660 -13180 35780 -13060
rect 35825 -13180 35945 -13060
rect 35990 -13180 36110 -13060
rect 36155 -13180 36275 -13060
rect 30795 -13345 30915 -13225
rect 30970 -13345 31090 -13225
rect 31135 -13345 31255 -13225
rect 31300 -13345 31420 -13225
rect 31465 -13345 31585 -13225
rect 31640 -13345 31760 -13225
rect 31805 -13345 31925 -13225
rect 31970 -13345 32090 -13225
rect 32135 -13345 32255 -13225
rect 32310 -13345 32430 -13225
rect 32475 -13345 32595 -13225
rect 32640 -13345 32760 -13225
rect 32805 -13345 32925 -13225
rect 32980 -13345 33100 -13225
rect 33145 -13345 33265 -13225
rect 33310 -13345 33430 -13225
rect 33475 -13345 33595 -13225
rect 33650 -13345 33770 -13225
rect 33815 -13345 33935 -13225
rect 33980 -13345 34100 -13225
rect 34145 -13345 34265 -13225
rect 34320 -13345 34440 -13225
rect 34485 -13345 34605 -13225
rect 34650 -13345 34770 -13225
rect 34815 -13345 34935 -13225
rect 34990 -13345 35110 -13225
rect 35155 -13345 35275 -13225
rect 35320 -13345 35440 -13225
rect 35485 -13345 35605 -13225
rect 35660 -13345 35780 -13225
rect 35825 -13345 35945 -13225
rect 35990 -13345 36110 -13225
rect 36155 -13345 36275 -13225
rect 30795 -13520 30915 -13400
rect 30970 -13520 31090 -13400
rect 31135 -13520 31255 -13400
rect 31300 -13520 31420 -13400
rect 31465 -13520 31585 -13400
rect 31640 -13520 31760 -13400
rect 31805 -13520 31925 -13400
rect 31970 -13520 32090 -13400
rect 32135 -13520 32255 -13400
rect 32310 -13520 32430 -13400
rect 32475 -13520 32595 -13400
rect 32640 -13520 32760 -13400
rect 32805 -13520 32925 -13400
rect 32980 -13520 33100 -13400
rect 33145 -13520 33265 -13400
rect 33310 -13520 33430 -13400
rect 33475 -13520 33595 -13400
rect 33650 -13520 33770 -13400
rect 33815 -13520 33935 -13400
rect 33980 -13520 34100 -13400
rect 34145 -13520 34265 -13400
rect 34320 -13520 34440 -13400
rect 34485 -13520 34605 -13400
rect 34650 -13520 34770 -13400
rect 34815 -13520 34935 -13400
rect 34990 -13520 35110 -13400
rect 35155 -13520 35275 -13400
rect 35320 -13520 35440 -13400
rect 35485 -13520 35605 -13400
rect 35660 -13520 35780 -13400
rect 35825 -13520 35945 -13400
rect 35990 -13520 36110 -13400
rect 36155 -13520 36275 -13400
rect 30795 -13685 30915 -13565
rect 30970 -13685 31090 -13565
rect 31135 -13685 31255 -13565
rect 31300 -13685 31420 -13565
rect 31465 -13685 31585 -13565
rect 31640 -13685 31760 -13565
rect 31805 -13685 31925 -13565
rect 31970 -13685 32090 -13565
rect 32135 -13685 32255 -13565
rect 32310 -13685 32430 -13565
rect 32475 -13685 32595 -13565
rect 32640 -13685 32760 -13565
rect 32805 -13685 32925 -13565
rect 32980 -13685 33100 -13565
rect 33145 -13685 33265 -13565
rect 33310 -13685 33430 -13565
rect 33475 -13685 33595 -13565
rect 33650 -13685 33770 -13565
rect 33815 -13685 33935 -13565
rect 33980 -13685 34100 -13565
rect 34145 -13685 34265 -13565
rect 34320 -13685 34440 -13565
rect 34485 -13685 34605 -13565
rect 34650 -13685 34770 -13565
rect 34815 -13685 34935 -13565
rect 34990 -13685 35110 -13565
rect 35155 -13685 35275 -13565
rect 35320 -13685 35440 -13565
rect 35485 -13685 35605 -13565
rect 35660 -13685 35780 -13565
rect 35825 -13685 35945 -13565
rect 35990 -13685 36110 -13565
rect 36155 -13685 36275 -13565
rect 30795 -13850 30915 -13730
rect 30970 -13850 31090 -13730
rect 31135 -13850 31255 -13730
rect 31300 -13850 31420 -13730
rect 31465 -13850 31585 -13730
rect 31640 -13850 31760 -13730
rect 31805 -13850 31925 -13730
rect 31970 -13850 32090 -13730
rect 32135 -13850 32255 -13730
rect 32310 -13850 32430 -13730
rect 32475 -13850 32595 -13730
rect 32640 -13850 32760 -13730
rect 32805 -13850 32925 -13730
rect 32980 -13850 33100 -13730
rect 33145 -13850 33265 -13730
rect 33310 -13850 33430 -13730
rect 33475 -13850 33595 -13730
rect 33650 -13850 33770 -13730
rect 33815 -13850 33935 -13730
rect 33980 -13850 34100 -13730
rect 34145 -13850 34265 -13730
rect 34320 -13850 34440 -13730
rect 34485 -13850 34605 -13730
rect 34650 -13850 34770 -13730
rect 34815 -13850 34935 -13730
rect 34990 -13850 35110 -13730
rect 35155 -13850 35275 -13730
rect 35320 -13850 35440 -13730
rect 35485 -13850 35605 -13730
rect 35660 -13850 35780 -13730
rect 35825 -13850 35945 -13730
rect 35990 -13850 36110 -13730
rect 36155 -13850 36275 -13730
rect 30795 -14015 30915 -13895
rect 30970 -14015 31090 -13895
rect 31135 -14015 31255 -13895
rect 31300 -14015 31420 -13895
rect 31465 -14015 31585 -13895
rect 31640 -14015 31760 -13895
rect 31805 -14015 31925 -13895
rect 31970 -14015 32090 -13895
rect 32135 -14015 32255 -13895
rect 32310 -14015 32430 -13895
rect 32475 -14015 32595 -13895
rect 32640 -14015 32760 -13895
rect 32805 -14015 32925 -13895
rect 32980 -14015 33100 -13895
rect 33145 -14015 33265 -13895
rect 33310 -14015 33430 -13895
rect 33475 -14015 33595 -13895
rect 33650 -14015 33770 -13895
rect 33815 -14015 33935 -13895
rect 33980 -14015 34100 -13895
rect 34145 -14015 34265 -13895
rect 34320 -14015 34440 -13895
rect 34485 -14015 34605 -13895
rect 34650 -14015 34770 -13895
rect 34815 -14015 34935 -13895
rect 34990 -14015 35110 -13895
rect 35155 -14015 35275 -13895
rect 35320 -14015 35440 -13895
rect 35485 -14015 35605 -13895
rect 35660 -14015 35780 -13895
rect 35825 -14015 35945 -13895
rect 35990 -14015 36110 -13895
rect 36155 -14015 36275 -13895
rect 30795 -14190 30915 -14070
rect 30970 -14190 31090 -14070
rect 31135 -14190 31255 -14070
rect 31300 -14190 31420 -14070
rect 31465 -14190 31585 -14070
rect 31640 -14190 31760 -14070
rect 31805 -14190 31925 -14070
rect 31970 -14190 32090 -14070
rect 32135 -14190 32255 -14070
rect 32310 -14190 32430 -14070
rect 32475 -14190 32595 -14070
rect 32640 -14190 32760 -14070
rect 32805 -14190 32925 -14070
rect 32980 -14190 33100 -14070
rect 33145 -14190 33265 -14070
rect 33310 -14190 33430 -14070
rect 33475 -14190 33595 -14070
rect 33650 -14190 33770 -14070
rect 33815 -14190 33935 -14070
rect 33980 -14190 34100 -14070
rect 34145 -14190 34265 -14070
rect 34320 -14190 34440 -14070
rect 34485 -14190 34605 -14070
rect 34650 -14190 34770 -14070
rect 34815 -14190 34935 -14070
rect 34990 -14190 35110 -14070
rect 35155 -14190 35275 -14070
rect 35320 -14190 35440 -14070
rect 35485 -14190 35605 -14070
rect 35660 -14190 35780 -14070
rect 35825 -14190 35945 -14070
rect 35990 -14190 36110 -14070
rect 36155 -14190 36275 -14070
rect 30795 -14355 30915 -14235
rect 30970 -14355 31090 -14235
rect 31135 -14355 31255 -14235
rect 31300 -14355 31420 -14235
rect 31465 -14355 31585 -14235
rect 31640 -14355 31760 -14235
rect 31805 -14355 31925 -14235
rect 31970 -14355 32090 -14235
rect 32135 -14355 32255 -14235
rect 32310 -14355 32430 -14235
rect 32475 -14355 32595 -14235
rect 32640 -14355 32760 -14235
rect 32805 -14355 32925 -14235
rect 32980 -14355 33100 -14235
rect 33145 -14355 33265 -14235
rect 33310 -14355 33430 -14235
rect 33475 -14355 33595 -14235
rect 33650 -14355 33770 -14235
rect 33815 -14355 33935 -14235
rect 33980 -14355 34100 -14235
rect 34145 -14355 34265 -14235
rect 34320 -14355 34440 -14235
rect 34485 -14355 34605 -14235
rect 34650 -14355 34770 -14235
rect 34815 -14355 34935 -14235
rect 34990 -14355 35110 -14235
rect 35155 -14355 35275 -14235
rect 35320 -14355 35440 -14235
rect 35485 -14355 35605 -14235
rect 35660 -14355 35780 -14235
rect 35825 -14355 35945 -14235
rect 35990 -14355 36110 -14235
rect 36155 -14355 36275 -14235
rect 30795 -14520 30915 -14400
rect 30970 -14520 31090 -14400
rect 31135 -14520 31255 -14400
rect 31300 -14520 31420 -14400
rect 31465 -14520 31585 -14400
rect 31640 -14520 31760 -14400
rect 31805 -14520 31925 -14400
rect 31970 -14520 32090 -14400
rect 32135 -14520 32255 -14400
rect 32310 -14520 32430 -14400
rect 32475 -14520 32595 -14400
rect 32640 -14520 32760 -14400
rect 32805 -14520 32925 -14400
rect 32980 -14520 33100 -14400
rect 33145 -14520 33265 -14400
rect 33310 -14520 33430 -14400
rect 33475 -14520 33595 -14400
rect 33650 -14520 33770 -14400
rect 33815 -14520 33935 -14400
rect 33980 -14520 34100 -14400
rect 34145 -14520 34265 -14400
rect 34320 -14520 34440 -14400
rect 34485 -14520 34605 -14400
rect 34650 -14520 34770 -14400
rect 34815 -14520 34935 -14400
rect 34990 -14520 35110 -14400
rect 35155 -14520 35275 -14400
rect 35320 -14520 35440 -14400
rect 35485 -14520 35605 -14400
rect 35660 -14520 35780 -14400
rect 35825 -14520 35945 -14400
rect 35990 -14520 36110 -14400
rect 36155 -14520 36275 -14400
rect 30795 -14685 30915 -14565
rect 30970 -14685 31090 -14565
rect 31135 -14685 31255 -14565
rect 31300 -14685 31420 -14565
rect 31465 -14685 31585 -14565
rect 31640 -14685 31760 -14565
rect 31805 -14685 31925 -14565
rect 31970 -14685 32090 -14565
rect 32135 -14685 32255 -14565
rect 32310 -14685 32430 -14565
rect 32475 -14685 32595 -14565
rect 32640 -14685 32760 -14565
rect 32805 -14685 32925 -14565
rect 32980 -14685 33100 -14565
rect 33145 -14685 33265 -14565
rect 33310 -14685 33430 -14565
rect 33475 -14685 33595 -14565
rect 33650 -14685 33770 -14565
rect 33815 -14685 33935 -14565
rect 33980 -14685 34100 -14565
rect 34145 -14685 34265 -14565
rect 34320 -14685 34440 -14565
rect 34485 -14685 34605 -14565
rect 34650 -14685 34770 -14565
rect 34815 -14685 34935 -14565
rect 34990 -14685 35110 -14565
rect 35155 -14685 35275 -14565
rect 35320 -14685 35440 -14565
rect 35485 -14685 35605 -14565
rect 35660 -14685 35780 -14565
rect 35825 -14685 35945 -14565
rect 35990 -14685 36110 -14565
rect 36155 -14685 36275 -14565
rect 30795 -14860 30915 -14740
rect 30970 -14860 31090 -14740
rect 31135 -14860 31255 -14740
rect 31300 -14860 31420 -14740
rect 31465 -14860 31585 -14740
rect 31640 -14860 31760 -14740
rect 31805 -14860 31925 -14740
rect 31970 -14860 32090 -14740
rect 32135 -14860 32255 -14740
rect 32310 -14860 32430 -14740
rect 32475 -14860 32595 -14740
rect 32640 -14860 32760 -14740
rect 32805 -14860 32925 -14740
rect 32980 -14860 33100 -14740
rect 33145 -14860 33265 -14740
rect 33310 -14860 33430 -14740
rect 33475 -14860 33595 -14740
rect 33650 -14860 33770 -14740
rect 33815 -14860 33935 -14740
rect 33980 -14860 34100 -14740
rect 34145 -14860 34265 -14740
rect 34320 -14860 34440 -14740
rect 34485 -14860 34605 -14740
rect 34650 -14860 34770 -14740
rect 34815 -14860 34935 -14740
rect 34990 -14860 35110 -14740
rect 35155 -14860 35275 -14740
rect 35320 -14860 35440 -14740
rect 35485 -14860 35605 -14740
rect 35660 -14860 35780 -14740
rect 35825 -14860 35945 -14740
rect 35990 -14860 36110 -14740
rect 36155 -14860 36275 -14740
rect 30795 -15025 30915 -14905
rect 30970 -15025 31090 -14905
rect 31135 -15025 31255 -14905
rect 31300 -15025 31420 -14905
rect 31465 -15025 31585 -14905
rect 31640 -15025 31760 -14905
rect 31805 -15025 31925 -14905
rect 31970 -15025 32090 -14905
rect 32135 -15025 32255 -14905
rect 32310 -15025 32430 -14905
rect 32475 -15025 32595 -14905
rect 32640 -15025 32760 -14905
rect 32805 -15025 32925 -14905
rect 32980 -15025 33100 -14905
rect 33145 -15025 33265 -14905
rect 33310 -15025 33430 -14905
rect 33475 -15025 33595 -14905
rect 33650 -15025 33770 -14905
rect 33815 -15025 33935 -14905
rect 33980 -15025 34100 -14905
rect 34145 -15025 34265 -14905
rect 34320 -15025 34440 -14905
rect 34485 -15025 34605 -14905
rect 34650 -15025 34770 -14905
rect 34815 -15025 34935 -14905
rect 34990 -15025 35110 -14905
rect 35155 -15025 35275 -14905
rect 35320 -15025 35440 -14905
rect 35485 -15025 35605 -14905
rect 35660 -15025 35780 -14905
rect 35825 -15025 35945 -14905
rect 35990 -15025 36110 -14905
rect 36155 -15025 36275 -14905
rect 30795 -15190 30915 -15070
rect 30970 -15190 31090 -15070
rect 31135 -15190 31255 -15070
rect 31300 -15190 31420 -15070
rect 31465 -15190 31585 -15070
rect 31640 -15190 31760 -15070
rect 31805 -15190 31925 -15070
rect 31970 -15190 32090 -15070
rect 32135 -15190 32255 -15070
rect 32310 -15190 32430 -15070
rect 32475 -15190 32595 -15070
rect 32640 -15190 32760 -15070
rect 32805 -15190 32925 -15070
rect 32980 -15190 33100 -15070
rect 33145 -15190 33265 -15070
rect 33310 -15190 33430 -15070
rect 33475 -15190 33595 -15070
rect 33650 -15190 33770 -15070
rect 33815 -15190 33935 -15070
rect 33980 -15190 34100 -15070
rect 34145 -15190 34265 -15070
rect 34320 -15190 34440 -15070
rect 34485 -15190 34605 -15070
rect 34650 -15190 34770 -15070
rect 34815 -15190 34935 -15070
rect 34990 -15190 35110 -15070
rect 35155 -15190 35275 -15070
rect 35320 -15190 35440 -15070
rect 35485 -15190 35605 -15070
rect 35660 -15190 35780 -15070
rect 35825 -15190 35945 -15070
rect 35990 -15190 36110 -15070
rect 36155 -15190 36275 -15070
rect 30795 -15355 30915 -15235
rect 30970 -15355 31090 -15235
rect 31135 -15355 31255 -15235
rect 31300 -15355 31420 -15235
rect 31465 -15355 31585 -15235
rect 31640 -15355 31760 -15235
rect 31805 -15355 31925 -15235
rect 31970 -15355 32090 -15235
rect 32135 -15355 32255 -15235
rect 32310 -15355 32430 -15235
rect 32475 -15355 32595 -15235
rect 32640 -15355 32760 -15235
rect 32805 -15355 32925 -15235
rect 32980 -15355 33100 -15235
rect 33145 -15355 33265 -15235
rect 33310 -15355 33430 -15235
rect 33475 -15355 33595 -15235
rect 33650 -15355 33770 -15235
rect 33815 -15355 33935 -15235
rect 33980 -15355 34100 -15235
rect 34145 -15355 34265 -15235
rect 34320 -15355 34440 -15235
rect 34485 -15355 34605 -15235
rect 34650 -15355 34770 -15235
rect 34815 -15355 34935 -15235
rect 34990 -15355 35110 -15235
rect 35155 -15355 35275 -15235
rect 35320 -15355 35440 -15235
rect 35485 -15355 35605 -15235
rect 35660 -15355 35780 -15235
rect 35825 -15355 35945 -15235
rect 35990 -15355 36110 -15235
rect 36155 -15355 36275 -15235
rect 30795 -15530 30915 -15410
rect 30970 -15530 31090 -15410
rect 31135 -15530 31255 -15410
rect 31300 -15530 31420 -15410
rect 31465 -15530 31585 -15410
rect 31640 -15530 31760 -15410
rect 31805 -15530 31925 -15410
rect 31970 -15530 32090 -15410
rect 32135 -15530 32255 -15410
rect 32310 -15530 32430 -15410
rect 32475 -15530 32595 -15410
rect 32640 -15530 32760 -15410
rect 32805 -15530 32925 -15410
rect 32980 -15530 33100 -15410
rect 33145 -15530 33265 -15410
rect 33310 -15530 33430 -15410
rect 33475 -15530 33595 -15410
rect 33650 -15530 33770 -15410
rect 33815 -15530 33935 -15410
rect 33980 -15530 34100 -15410
rect 34145 -15530 34265 -15410
rect 34320 -15530 34440 -15410
rect 34485 -15530 34605 -15410
rect 34650 -15530 34770 -15410
rect 34815 -15530 34935 -15410
rect 34990 -15530 35110 -15410
rect 35155 -15530 35275 -15410
rect 35320 -15530 35440 -15410
rect 35485 -15530 35605 -15410
rect 35660 -15530 35780 -15410
rect 35825 -15530 35945 -15410
rect 35990 -15530 36110 -15410
rect 36155 -15530 36275 -15410
rect 36485 -10170 36605 -10050
rect 36660 -10170 36780 -10050
rect 36825 -10170 36945 -10050
rect 36990 -10170 37110 -10050
rect 37155 -10170 37275 -10050
rect 37330 -10170 37450 -10050
rect 37495 -10170 37615 -10050
rect 37660 -10170 37780 -10050
rect 37825 -10170 37945 -10050
rect 38000 -10170 38120 -10050
rect 38165 -10170 38285 -10050
rect 38330 -10170 38450 -10050
rect 38495 -10170 38615 -10050
rect 38670 -10170 38790 -10050
rect 38835 -10170 38955 -10050
rect 39000 -10170 39120 -10050
rect 39165 -10170 39285 -10050
rect 39340 -10170 39460 -10050
rect 39505 -10170 39625 -10050
rect 39670 -10170 39790 -10050
rect 39835 -10170 39955 -10050
rect 40010 -10170 40130 -10050
rect 40175 -10170 40295 -10050
rect 40340 -10170 40460 -10050
rect 40505 -10170 40625 -10050
rect 40680 -10170 40800 -10050
rect 40845 -10170 40965 -10050
rect 41010 -10170 41130 -10050
rect 41175 -10170 41295 -10050
rect 41350 -10170 41470 -10050
rect 41515 -10170 41635 -10050
rect 41680 -10170 41800 -10050
rect 41845 -10170 41965 -10050
rect 36485 -10335 36605 -10215
rect 36660 -10335 36780 -10215
rect 36825 -10335 36945 -10215
rect 36990 -10335 37110 -10215
rect 37155 -10335 37275 -10215
rect 37330 -10335 37450 -10215
rect 37495 -10335 37615 -10215
rect 37660 -10335 37780 -10215
rect 37825 -10335 37945 -10215
rect 38000 -10335 38120 -10215
rect 38165 -10335 38285 -10215
rect 38330 -10335 38450 -10215
rect 38495 -10335 38615 -10215
rect 38670 -10335 38790 -10215
rect 38835 -10335 38955 -10215
rect 39000 -10335 39120 -10215
rect 39165 -10335 39285 -10215
rect 39340 -10335 39460 -10215
rect 39505 -10335 39625 -10215
rect 39670 -10335 39790 -10215
rect 39835 -10335 39955 -10215
rect 40010 -10335 40130 -10215
rect 40175 -10335 40295 -10215
rect 40340 -10335 40460 -10215
rect 40505 -10335 40625 -10215
rect 40680 -10335 40800 -10215
rect 40845 -10335 40965 -10215
rect 41010 -10335 41130 -10215
rect 41175 -10335 41295 -10215
rect 41350 -10335 41470 -10215
rect 41515 -10335 41635 -10215
rect 41680 -10335 41800 -10215
rect 41845 -10335 41965 -10215
rect 36485 -10500 36605 -10380
rect 36660 -10500 36780 -10380
rect 36825 -10500 36945 -10380
rect 36990 -10500 37110 -10380
rect 37155 -10500 37275 -10380
rect 37330 -10500 37450 -10380
rect 37495 -10500 37615 -10380
rect 37660 -10500 37780 -10380
rect 37825 -10500 37945 -10380
rect 38000 -10500 38120 -10380
rect 38165 -10500 38285 -10380
rect 38330 -10500 38450 -10380
rect 38495 -10500 38615 -10380
rect 38670 -10500 38790 -10380
rect 38835 -10500 38955 -10380
rect 39000 -10500 39120 -10380
rect 39165 -10500 39285 -10380
rect 39340 -10500 39460 -10380
rect 39505 -10500 39625 -10380
rect 39670 -10500 39790 -10380
rect 39835 -10500 39955 -10380
rect 40010 -10500 40130 -10380
rect 40175 -10500 40295 -10380
rect 40340 -10500 40460 -10380
rect 40505 -10500 40625 -10380
rect 40680 -10500 40800 -10380
rect 40845 -10500 40965 -10380
rect 41010 -10500 41130 -10380
rect 41175 -10500 41295 -10380
rect 41350 -10500 41470 -10380
rect 41515 -10500 41635 -10380
rect 41680 -10500 41800 -10380
rect 41845 -10500 41965 -10380
rect 36485 -10665 36605 -10545
rect 36660 -10665 36780 -10545
rect 36825 -10665 36945 -10545
rect 36990 -10665 37110 -10545
rect 37155 -10665 37275 -10545
rect 37330 -10665 37450 -10545
rect 37495 -10665 37615 -10545
rect 37660 -10665 37780 -10545
rect 37825 -10665 37945 -10545
rect 38000 -10665 38120 -10545
rect 38165 -10665 38285 -10545
rect 38330 -10665 38450 -10545
rect 38495 -10665 38615 -10545
rect 38670 -10665 38790 -10545
rect 38835 -10665 38955 -10545
rect 39000 -10665 39120 -10545
rect 39165 -10665 39285 -10545
rect 39340 -10665 39460 -10545
rect 39505 -10665 39625 -10545
rect 39670 -10665 39790 -10545
rect 39835 -10665 39955 -10545
rect 40010 -10665 40130 -10545
rect 40175 -10665 40295 -10545
rect 40340 -10665 40460 -10545
rect 40505 -10665 40625 -10545
rect 40680 -10665 40800 -10545
rect 40845 -10665 40965 -10545
rect 41010 -10665 41130 -10545
rect 41175 -10665 41295 -10545
rect 41350 -10665 41470 -10545
rect 41515 -10665 41635 -10545
rect 41680 -10665 41800 -10545
rect 41845 -10665 41965 -10545
rect 36485 -10840 36605 -10720
rect 36660 -10840 36780 -10720
rect 36825 -10840 36945 -10720
rect 36990 -10840 37110 -10720
rect 37155 -10840 37275 -10720
rect 37330 -10840 37450 -10720
rect 37495 -10840 37615 -10720
rect 37660 -10840 37780 -10720
rect 37825 -10840 37945 -10720
rect 38000 -10840 38120 -10720
rect 38165 -10840 38285 -10720
rect 38330 -10840 38450 -10720
rect 38495 -10840 38615 -10720
rect 38670 -10840 38790 -10720
rect 38835 -10840 38955 -10720
rect 39000 -10840 39120 -10720
rect 39165 -10840 39285 -10720
rect 39340 -10840 39460 -10720
rect 39505 -10840 39625 -10720
rect 39670 -10840 39790 -10720
rect 39835 -10840 39955 -10720
rect 40010 -10840 40130 -10720
rect 40175 -10840 40295 -10720
rect 40340 -10840 40460 -10720
rect 40505 -10840 40625 -10720
rect 40680 -10840 40800 -10720
rect 40845 -10840 40965 -10720
rect 41010 -10840 41130 -10720
rect 41175 -10840 41295 -10720
rect 41350 -10840 41470 -10720
rect 41515 -10840 41635 -10720
rect 41680 -10840 41800 -10720
rect 41845 -10840 41965 -10720
rect 36485 -11005 36605 -10885
rect 36660 -11005 36780 -10885
rect 36825 -11005 36945 -10885
rect 36990 -11005 37110 -10885
rect 37155 -11005 37275 -10885
rect 37330 -11005 37450 -10885
rect 37495 -11005 37615 -10885
rect 37660 -11005 37780 -10885
rect 37825 -11005 37945 -10885
rect 38000 -11005 38120 -10885
rect 38165 -11005 38285 -10885
rect 38330 -11005 38450 -10885
rect 38495 -11005 38615 -10885
rect 38670 -11005 38790 -10885
rect 38835 -11005 38955 -10885
rect 39000 -11005 39120 -10885
rect 39165 -11005 39285 -10885
rect 39340 -11005 39460 -10885
rect 39505 -11005 39625 -10885
rect 39670 -11005 39790 -10885
rect 39835 -11005 39955 -10885
rect 40010 -11005 40130 -10885
rect 40175 -11005 40295 -10885
rect 40340 -11005 40460 -10885
rect 40505 -11005 40625 -10885
rect 40680 -11005 40800 -10885
rect 40845 -11005 40965 -10885
rect 41010 -11005 41130 -10885
rect 41175 -11005 41295 -10885
rect 41350 -11005 41470 -10885
rect 41515 -11005 41635 -10885
rect 41680 -11005 41800 -10885
rect 41845 -11005 41965 -10885
rect 36485 -11170 36605 -11050
rect 36660 -11170 36780 -11050
rect 36825 -11170 36945 -11050
rect 36990 -11170 37110 -11050
rect 37155 -11170 37275 -11050
rect 37330 -11170 37450 -11050
rect 37495 -11170 37615 -11050
rect 37660 -11170 37780 -11050
rect 37825 -11170 37945 -11050
rect 38000 -11170 38120 -11050
rect 38165 -11170 38285 -11050
rect 38330 -11170 38450 -11050
rect 38495 -11170 38615 -11050
rect 38670 -11170 38790 -11050
rect 38835 -11170 38955 -11050
rect 39000 -11170 39120 -11050
rect 39165 -11170 39285 -11050
rect 39340 -11170 39460 -11050
rect 39505 -11170 39625 -11050
rect 39670 -11170 39790 -11050
rect 39835 -11170 39955 -11050
rect 40010 -11170 40130 -11050
rect 40175 -11170 40295 -11050
rect 40340 -11170 40460 -11050
rect 40505 -11170 40625 -11050
rect 40680 -11170 40800 -11050
rect 40845 -11170 40965 -11050
rect 41010 -11170 41130 -11050
rect 41175 -11170 41295 -11050
rect 41350 -11170 41470 -11050
rect 41515 -11170 41635 -11050
rect 41680 -11170 41800 -11050
rect 41845 -11170 41965 -11050
rect 36485 -11335 36605 -11215
rect 36660 -11335 36780 -11215
rect 36825 -11335 36945 -11215
rect 36990 -11335 37110 -11215
rect 37155 -11335 37275 -11215
rect 37330 -11335 37450 -11215
rect 37495 -11335 37615 -11215
rect 37660 -11335 37780 -11215
rect 37825 -11335 37945 -11215
rect 38000 -11335 38120 -11215
rect 38165 -11335 38285 -11215
rect 38330 -11335 38450 -11215
rect 38495 -11335 38615 -11215
rect 38670 -11335 38790 -11215
rect 38835 -11335 38955 -11215
rect 39000 -11335 39120 -11215
rect 39165 -11335 39285 -11215
rect 39340 -11335 39460 -11215
rect 39505 -11335 39625 -11215
rect 39670 -11335 39790 -11215
rect 39835 -11335 39955 -11215
rect 40010 -11335 40130 -11215
rect 40175 -11335 40295 -11215
rect 40340 -11335 40460 -11215
rect 40505 -11335 40625 -11215
rect 40680 -11335 40800 -11215
rect 40845 -11335 40965 -11215
rect 41010 -11335 41130 -11215
rect 41175 -11335 41295 -11215
rect 41350 -11335 41470 -11215
rect 41515 -11335 41635 -11215
rect 41680 -11335 41800 -11215
rect 41845 -11335 41965 -11215
rect 36485 -11510 36605 -11390
rect 36660 -11510 36780 -11390
rect 36825 -11510 36945 -11390
rect 36990 -11510 37110 -11390
rect 37155 -11510 37275 -11390
rect 37330 -11510 37450 -11390
rect 37495 -11510 37615 -11390
rect 37660 -11510 37780 -11390
rect 37825 -11510 37945 -11390
rect 38000 -11510 38120 -11390
rect 38165 -11510 38285 -11390
rect 38330 -11510 38450 -11390
rect 38495 -11510 38615 -11390
rect 38670 -11510 38790 -11390
rect 38835 -11510 38955 -11390
rect 39000 -11510 39120 -11390
rect 39165 -11510 39285 -11390
rect 39340 -11510 39460 -11390
rect 39505 -11510 39625 -11390
rect 39670 -11510 39790 -11390
rect 39835 -11510 39955 -11390
rect 40010 -11510 40130 -11390
rect 40175 -11510 40295 -11390
rect 40340 -11510 40460 -11390
rect 40505 -11510 40625 -11390
rect 40680 -11510 40800 -11390
rect 40845 -11510 40965 -11390
rect 41010 -11510 41130 -11390
rect 41175 -11510 41295 -11390
rect 41350 -11510 41470 -11390
rect 41515 -11510 41635 -11390
rect 41680 -11510 41800 -11390
rect 41845 -11510 41965 -11390
rect 36485 -11675 36605 -11555
rect 36660 -11675 36780 -11555
rect 36825 -11675 36945 -11555
rect 36990 -11675 37110 -11555
rect 37155 -11675 37275 -11555
rect 37330 -11675 37450 -11555
rect 37495 -11675 37615 -11555
rect 37660 -11675 37780 -11555
rect 37825 -11675 37945 -11555
rect 38000 -11675 38120 -11555
rect 38165 -11675 38285 -11555
rect 38330 -11675 38450 -11555
rect 38495 -11675 38615 -11555
rect 38670 -11675 38790 -11555
rect 38835 -11675 38955 -11555
rect 39000 -11675 39120 -11555
rect 39165 -11675 39285 -11555
rect 39340 -11675 39460 -11555
rect 39505 -11675 39625 -11555
rect 39670 -11675 39790 -11555
rect 39835 -11675 39955 -11555
rect 40010 -11675 40130 -11555
rect 40175 -11675 40295 -11555
rect 40340 -11675 40460 -11555
rect 40505 -11675 40625 -11555
rect 40680 -11675 40800 -11555
rect 40845 -11675 40965 -11555
rect 41010 -11675 41130 -11555
rect 41175 -11675 41295 -11555
rect 41350 -11675 41470 -11555
rect 41515 -11675 41635 -11555
rect 41680 -11675 41800 -11555
rect 41845 -11675 41965 -11555
rect 36485 -11840 36605 -11720
rect 36660 -11840 36780 -11720
rect 36825 -11840 36945 -11720
rect 36990 -11840 37110 -11720
rect 37155 -11840 37275 -11720
rect 37330 -11840 37450 -11720
rect 37495 -11840 37615 -11720
rect 37660 -11840 37780 -11720
rect 37825 -11840 37945 -11720
rect 38000 -11840 38120 -11720
rect 38165 -11840 38285 -11720
rect 38330 -11840 38450 -11720
rect 38495 -11840 38615 -11720
rect 38670 -11840 38790 -11720
rect 38835 -11840 38955 -11720
rect 39000 -11840 39120 -11720
rect 39165 -11840 39285 -11720
rect 39340 -11840 39460 -11720
rect 39505 -11840 39625 -11720
rect 39670 -11840 39790 -11720
rect 39835 -11840 39955 -11720
rect 40010 -11840 40130 -11720
rect 40175 -11840 40295 -11720
rect 40340 -11840 40460 -11720
rect 40505 -11840 40625 -11720
rect 40680 -11840 40800 -11720
rect 40845 -11840 40965 -11720
rect 41010 -11840 41130 -11720
rect 41175 -11840 41295 -11720
rect 41350 -11840 41470 -11720
rect 41515 -11840 41635 -11720
rect 41680 -11840 41800 -11720
rect 41845 -11840 41965 -11720
rect 36485 -12005 36605 -11885
rect 36660 -12005 36780 -11885
rect 36825 -12005 36945 -11885
rect 36990 -12005 37110 -11885
rect 37155 -12005 37275 -11885
rect 37330 -12005 37450 -11885
rect 37495 -12005 37615 -11885
rect 37660 -12005 37780 -11885
rect 37825 -12005 37945 -11885
rect 38000 -12005 38120 -11885
rect 38165 -12005 38285 -11885
rect 38330 -12005 38450 -11885
rect 38495 -12005 38615 -11885
rect 38670 -12005 38790 -11885
rect 38835 -12005 38955 -11885
rect 39000 -12005 39120 -11885
rect 39165 -12005 39285 -11885
rect 39340 -12005 39460 -11885
rect 39505 -12005 39625 -11885
rect 39670 -12005 39790 -11885
rect 39835 -12005 39955 -11885
rect 40010 -12005 40130 -11885
rect 40175 -12005 40295 -11885
rect 40340 -12005 40460 -11885
rect 40505 -12005 40625 -11885
rect 40680 -12005 40800 -11885
rect 40845 -12005 40965 -11885
rect 41010 -12005 41130 -11885
rect 41175 -12005 41295 -11885
rect 41350 -12005 41470 -11885
rect 41515 -12005 41635 -11885
rect 41680 -12005 41800 -11885
rect 41845 -12005 41965 -11885
rect 36485 -12180 36605 -12060
rect 36660 -12180 36780 -12060
rect 36825 -12180 36945 -12060
rect 36990 -12180 37110 -12060
rect 37155 -12180 37275 -12060
rect 37330 -12180 37450 -12060
rect 37495 -12180 37615 -12060
rect 37660 -12180 37780 -12060
rect 37825 -12180 37945 -12060
rect 38000 -12180 38120 -12060
rect 38165 -12180 38285 -12060
rect 38330 -12180 38450 -12060
rect 38495 -12180 38615 -12060
rect 38670 -12180 38790 -12060
rect 38835 -12180 38955 -12060
rect 39000 -12180 39120 -12060
rect 39165 -12180 39285 -12060
rect 39340 -12180 39460 -12060
rect 39505 -12180 39625 -12060
rect 39670 -12180 39790 -12060
rect 39835 -12180 39955 -12060
rect 40010 -12180 40130 -12060
rect 40175 -12180 40295 -12060
rect 40340 -12180 40460 -12060
rect 40505 -12180 40625 -12060
rect 40680 -12180 40800 -12060
rect 40845 -12180 40965 -12060
rect 41010 -12180 41130 -12060
rect 41175 -12180 41295 -12060
rect 41350 -12180 41470 -12060
rect 41515 -12180 41635 -12060
rect 41680 -12180 41800 -12060
rect 41845 -12180 41965 -12060
rect 36485 -12345 36605 -12225
rect 36660 -12345 36780 -12225
rect 36825 -12345 36945 -12225
rect 36990 -12345 37110 -12225
rect 37155 -12345 37275 -12225
rect 37330 -12345 37450 -12225
rect 37495 -12345 37615 -12225
rect 37660 -12345 37780 -12225
rect 37825 -12345 37945 -12225
rect 38000 -12345 38120 -12225
rect 38165 -12345 38285 -12225
rect 38330 -12345 38450 -12225
rect 38495 -12345 38615 -12225
rect 38670 -12345 38790 -12225
rect 38835 -12345 38955 -12225
rect 39000 -12345 39120 -12225
rect 39165 -12345 39285 -12225
rect 39340 -12345 39460 -12225
rect 39505 -12345 39625 -12225
rect 39670 -12345 39790 -12225
rect 39835 -12345 39955 -12225
rect 40010 -12345 40130 -12225
rect 40175 -12345 40295 -12225
rect 40340 -12345 40460 -12225
rect 40505 -12345 40625 -12225
rect 40680 -12345 40800 -12225
rect 40845 -12345 40965 -12225
rect 41010 -12345 41130 -12225
rect 41175 -12345 41295 -12225
rect 41350 -12345 41470 -12225
rect 41515 -12345 41635 -12225
rect 41680 -12345 41800 -12225
rect 41845 -12345 41965 -12225
rect 36485 -12510 36605 -12390
rect 36660 -12510 36780 -12390
rect 36825 -12510 36945 -12390
rect 36990 -12510 37110 -12390
rect 37155 -12510 37275 -12390
rect 37330 -12510 37450 -12390
rect 37495 -12510 37615 -12390
rect 37660 -12510 37780 -12390
rect 37825 -12510 37945 -12390
rect 38000 -12510 38120 -12390
rect 38165 -12510 38285 -12390
rect 38330 -12510 38450 -12390
rect 38495 -12510 38615 -12390
rect 38670 -12510 38790 -12390
rect 38835 -12510 38955 -12390
rect 39000 -12510 39120 -12390
rect 39165 -12510 39285 -12390
rect 39340 -12510 39460 -12390
rect 39505 -12510 39625 -12390
rect 39670 -12510 39790 -12390
rect 39835 -12510 39955 -12390
rect 40010 -12510 40130 -12390
rect 40175 -12510 40295 -12390
rect 40340 -12510 40460 -12390
rect 40505 -12510 40625 -12390
rect 40680 -12510 40800 -12390
rect 40845 -12510 40965 -12390
rect 41010 -12510 41130 -12390
rect 41175 -12510 41295 -12390
rect 41350 -12510 41470 -12390
rect 41515 -12510 41635 -12390
rect 41680 -12510 41800 -12390
rect 41845 -12510 41965 -12390
rect 36485 -12675 36605 -12555
rect 36660 -12675 36780 -12555
rect 36825 -12675 36945 -12555
rect 36990 -12675 37110 -12555
rect 37155 -12675 37275 -12555
rect 37330 -12675 37450 -12555
rect 37495 -12675 37615 -12555
rect 37660 -12675 37780 -12555
rect 37825 -12675 37945 -12555
rect 38000 -12675 38120 -12555
rect 38165 -12675 38285 -12555
rect 38330 -12675 38450 -12555
rect 38495 -12675 38615 -12555
rect 38670 -12675 38790 -12555
rect 38835 -12675 38955 -12555
rect 39000 -12675 39120 -12555
rect 39165 -12675 39285 -12555
rect 39340 -12675 39460 -12555
rect 39505 -12675 39625 -12555
rect 39670 -12675 39790 -12555
rect 39835 -12675 39955 -12555
rect 40010 -12675 40130 -12555
rect 40175 -12675 40295 -12555
rect 40340 -12675 40460 -12555
rect 40505 -12675 40625 -12555
rect 40680 -12675 40800 -12555
rect 40845 -12675 40965 -12555
rect 41010 -12675 41130 -12555
rect 41175 -12675 41295 -12555
rect 41350 -12675 41470 -12555
rect 41515 -12675 41635 -12555
rect 41680 -12675 41800 -12555
rect 41845 -12675 41965 -12555
rect 36485 -12850 36605 -12730
rect 36660 -12850 36780 -12730
rect 36825 -12850 36945 -12730
rect 36990 -12850 37110 -12730
rect 37155 -12850 37275 -12730
rect 37330 -12850 37450 -12730
rect 37495 -12850 37615 -12730
rect 37660 -12850 37780 -12730
rect 37825 -12850 37945 -12730
rect 38000 -12850 38120 -12730
rect 38165 -12850 38285 -12730
rect 38330 -12850 38450 -12730
rect 38495 -12850 38615 -12730
rect 38670 -12850 38790 -12730
rect 38835 -12850 38955 -12730
rect 39000 -12850 39120 -12730
rect 39165 -12850 39285 -12730
rect 39340 -12850 39460 -12730
rect 39505 -12850 39625 -12730
rect 39670 -12850 39790 -12730
rect 39835 -12850 39955 -12730
rect 40010 -12850 40130 -12730
rect 40175 -12850 40295 -12730
rect 40340 -12850 40460 -12730
rect 40505 -12850 40625 -12730
rect 40680 -12850 40800 -12730
rect 40845 -12850 40965 -12730
rect 41010 -12850 41130 -12730
rect 41175 -12850 41295 -12730
rect 41350 -12850 41470 -12730
rect 41515 -12850 41635 -12730
rect 41680 -12850 41800 -12730
rect 41845 -12850 41965 -12730
rect 36485 -13015 36605 -12895
rect 36660 -13015 36780 -12895
rect 36825 -13015 36945 -12895
rect 36990 -13015 37110 -12895
rect 37155 -13015 37275 -12895
rect 37330 -13015 37450 -12895
rect 37495 -13015 37615 -12895
rect 37660 -13015 37780 -12895
rect 37825 -13015 37945 -12895
rect 38000 -13015 38120 -12895
rect 38165 -13015 38285 -12895
rect 38330 -13015 38450 -12895
rect 38495 -13015 38615 -12895
rect 38670 -13015 38790 -12895
rect 38835 -13015 38955 -12895
rect 39000 -13015 39120 -12895
rect 39165 -13015 39285 -12895
rect 39340 -13015 39460 -12895
rect 39505 -13015 39625 -12895
rect 39670 -13015 39790 -12895
rect 39835 -13015 39955 -12895
rect 40010 -13015 40130 -12895
rect 40175 -13015 40295 -12895
rect 40340 -13015 40460 -12895
rect 40505 -13015 40625 -12895
rect 40680 -13015 40800 -12895
rect 40845 -13015 40965 -12895
rect 41010 -13015 41130 -12895
rect 41175 -13015 41295 -12895
rect 41350 -13015 41470 -12895
rect 41515 -13015 41635 -12895
rect 41680 -13015 41800 -12895
rect 41845 -13015 41965 -12895
rect 36485 -13180 36605 -13060
rect 36660 -13180 36780 -13060
rect 36825 -13180 36945 -13060
rect 36990 -13180 37110 -13060
rect 37155 -13180 37275 -13060
rect 37330 -13180 37450 -13060
rect 37495 -13180 37615 -13060
rect 37660 -13180 37780 -13060
rect 37825 -13180 37945 -13060
rect 38000 -13180 38120 -13060
rect 38165 -13180 38285 -13060
rect 38330 -13180 38450 -13060
rect 38495 -13180 38615 -13060
rect 38670 -13180 38790 -13060
rect 38835 -13180 38955 -13060
rect 39000 -13180 39120 -13060
rect 39165 -13180 39285 -13060
rect 39340 -13180 39460 -13060
rect 39505 -13180 39625 -13060
rect 39670 -13180 39790 -13060
rect 39835 -13180 39955 -13060
rect 40010 -13180 40130 -13060
rect 40175 -13180 40295 -13060
rect 40340 -13180 40460 -13060
rect 40505 -13180 40625 -13060
rect 40680 -13180 40800 -13060
rect 40845 -13180 40965 -13060
rect 41010 -13180 41130 -13060
rect 41175 -13180 41295 -13060
rect 41350 -13180 41470 -13060
rect 41515 -13180 41635 -13060
rect 41680 -13180 41800 -13060
rect 41845 -13180 41965 -13060
rect 36485 -13345 36605 -13225
rect 36660 -13345 36780 -13225
rect 36825 -13345 36945 -13225
rect 36990 -13345 37110 -13225
rect 37155 -13345 37275 -13225
rect 37330 -13345 37450 -13225
rect 37495 -13345 37615 -13225
rect 37660 -13345 37780 -13225
rect 37825 -13345 37945 -13225
rect 38000 -13345 38120 -13225
rect 38165 -13345 38285 -13225
rect 38330 -13345 38450 -13225
rect 38495 -13345 38615 -13225
rect 38670 -13345 38790 -13225
rect 38835 -13345 38955 -13225
rect 39000 -13345 39120 -13225
rect 39165 -13345 39285 -13225
rect 39340 -13345 39460 -13225
rect 39505 -13345 39625 -13225
rect 39670 -13345 39790 -13225
rect 39835 -13345 39955 -13225
rect 40010 -13345 40130 -13225
rect 40175 -13345 40295 -13225
rect 40340 -13345 40460 -13225
rect 40505 -13345 40625 -13225
rect 40680 -13345 40800 -13225
rect 40845 -13345 40965 -13225
rect 41010 -13345 41130 -13225
rect 41175 -13345 41295 -13225
rect 41350 -13345 41470 -13225
rect 41515 -13345 41635 -13225
rect 41680 -13345 41800 -13225
rect 41845 -13345 41965 -13225
rect 36485 -13520 36605 -13400
rect 36660 -13520 36780 -13400
rect 36825 -13520 36945 -13400
rect 36990 -13520 37110 -13400
rect 37155 -13520 37275 -13400
rect 37330 -13520 37450 -13400
rect 37495 -13520 37615 -13400
rect 37660 -13520 37780 -13400
rect 37825 -13520 37945 -13400
rect 38000 -13520 38120 -13400
rect 38165 -13520 38285 -13400
rect 38330 -13520 38450 -13400
rect 38495 -13520 38615 -13400
rect 38670 -13520 38790 -13400
rect 38835 -13520 38955 -13400
rect 39000 -13520 39120 -13400
rect 39165 -13520 39285 -13400
rect 39340 -13520 39460 -13400
rect 39505 -13520 39625 -13400
rect 39670 -13520 39790 -13400
rect 39835 -13520 39955 -13400
rect 40010 -13520 40130 -13400
rect 40175 -13520 40295 -13400
rect 40340 -13520 40460 -13400
rect 40505 -13520 40625 -13400
rect 40680 -13520 40800 -13400
rect 40845 -13520 40965 -13400
rect 41010 -13520 41130 -13400
rect 41175 -13520 41295 -13400
rect 41350 -13520 41470 -13400
rect 41515 -13520 41635 -13400
rect 41680 -13520 41800 -13400
rect 41845 -13520 41965 -13400
rect 36485 -13685 36605 -13565
rect 36660 -13685 36780 -13565
rect 36825 -13685 36945 -13565
rect 36990 -13685 37110 -13565
rect 37155 -13685 37275 -13565
rect 37330 -13685 37450 -13565
rect 37495 -13685 37615 -13565
rect 37660 -13685 37780 -13565
rect 37825 -13685 37945 -13565
rect 38000 -13685 38120 -13565
rect 38165 -13685 38285 -13565
rect 38330 -13685 38450 -13565
rect 38495 -13685 38615 -13565
rect 38670 -13685 38790 -13565
rect 38835 -13685 38955 -13565
rect 39000 -13685 39120 -13565
rect 39165 -13685 39285 -13565
rect 39340 -13685 39460 -13565
rect 39505 -13685 39625 -13565
rect 39670 -13685 39790 -13565
rect 39835 -13685 39955 -13565
rect 40010 -13685 40130 -13565
rect 40175 -13685 40295 -13565
rect 40340 -13685 40460 -13565
rect 40505 -13685 40625 -13565
rect 40680 -13685 40800 -13565
rect 40845 -13685 40965 -13565
rect 41010 -13685 41130 -13565
rect 41175 -13685 41295 -13565
rect 41350 -13685 41470 -13565
rect 41515 -13685 41635 -13565
rect 41680 -13685 41800 -13565
rect 41845 -13685 41965 -13565
rect 36485 -13850 36605 -13730
rect 36660 -13850 36780 -13730
rect 36825 -13850 36945 -13730
rect 36990 -13850 37110 -13730
rect 37155 -13850 37275 -13730
rect 37330 -13850 37450 -13730
rect 37495 -13850 37615 -13730
rect 37660 -13850 37780 -13730
rect 37825 -13850 37945 -13730
rect 38000 -13850 38120 -13730
rect 38165 -13850 38285 -13730
rect 38330 -13850 38450 -13730
rect 38495 -13850 38615 -13730
rect 38670 -13850 38790 -13730
rect 38835 -13850 38955 -13730
rect 39000 -13850 39120 -13730
rect 39165 -13850 39285 -13730
rect 39340 -13850 39460 -13730
rect 39505 -13850 39625 -13730
rect 39670 -13850 39790 -13730
rect 39835 -13850 39955 -13730
rect 40010 -13850 40130 -13730
rect 40175 -13850 40295 -13730
rect 40340 -13850 40460 -13730
rect 40505 -13850 40625 -13730
rect 40680 -13850 40800 -13730
rect 40845 -13850 40965 -13730
rect 41010 -13850 41130 -13730
rect 41175 -13850 41295 -13730
rect 41350 -13850 41470 -13730
rect 41515 -13850 41635 -13730
rect 41680 -13850 41800 -13730
rect 41845 -13850 41965 -13730
rect 36485 -14015 36605 -13895
rect 36660 -14015 36780 -13895
rect 36825 -14015 36945 -13895
rect 36990 -14015 37110 -13895
rect 37155 -14015 37275 -13895
rect 37330 -14015 37450 -13895
rect 37495 -14015 37615 -13895
rect 37660 -14015 37780 -13895
rect 37825 -14015 37945 -13895
rect 38000 -14015 38120 -13895
rect 38165 -14015 38285 -13895
rect 38330 -14015 38450 -13895
rect 38495 -14015 38615 -13895
rect 38670 -14015 38790 -13895
rect 38835 -14015 38955 -13895
rect 39000 -14015 39120 -13895
rect 39165 -14015 39285 -13895
rect 39340 -14015 39460 -13895
rect 39505 -14015 39625 -13895
rect 39670 -14015 39790 -13895
rect 39835 -14015 39955 -13895
rect 40010 -14015 40130 -13895
rect 40175 -14015 40295 -13895
rect 40340 -14015 40460 -13895
rect 40505 -14015 40625 -13895
rect 40680 -14015 40800 -13895
rect 40845 -14015 40965 -13895
rect 41010 -14015 41130 -13895
rect 41175 -14015 41295 -13895
rect 41350 -14015 41470 -13895
rect 41515 -14015 41635 -13895
rect 41680 -14015 41800 -13895
rect 41845 -14015 41965 -13895
rect 36485 -14190 36605 -14070
rect 36660 -14190 36780 -14070
rect 36825 -14190 36945 -14070
rect 36990 -14190 37110 -14070
rect 37155 -14190 37275 -14070
rect 37330 -14190 37450 -14070
rect 37495 -14190 37615 -14070
rect 37660 -14190 37780 -14070
rect 37825 -14190 37945 -14070
rect 38000 -14190 38120 -14070
rect 38165 -14190 38285 -14070
rect 38330 -14190 38450 -14070
rect 38495 -14190 38615 -14070
rect 38670 -14190 38790 -14070
rect 38835 -14190 38955 -14070
rect 39000 -14190 39120 -14070
rect 39165 -14190 39285 -14070
rect 39340 -14190 39460 -14070
rect 39505 -14190 39625 -14070
rect 39670 -14190 39790 -14070
rect 39835 -14190 39955 -14070
rect 40010 -14190 40130 -14070
rect 40175 -14190 40295 -14070
rect 40340 -14190 40460 -14070
rect 40505 -14190 40625 -14070
rect 40680 -14190 40800 -14070
rect 40845 -14190 40965 -14070
rect 41010 -14190 41130 -14070
rect 41175 -14190 41295 -14070
rect 41350 -14190 41470 -14070
rect 41515 -14190 41635 -14070
rect 41680 -14190 41800 -14070
rect 41845 -14190 41965 -14070
rect 36485 -14355 36605 -14235
rect 36660 -14355 36780 -14235
rect 36825 -14355 36945 -14235
rect 36990 -14355 37110 -14235
rect 37155 -14355 37275 -14235
rect 37330 -14355 37450 -14235
rect 37495 -14355 37615 -14235
rect 37660 -14355 37780 -14235
rect 37825 -14355 37945 -14235
rect 38000 -14355 38120 -14235
rect 38165 -14355 38285 -14235
rect 38330 -14355 38450 -14235
rect 38495 -14355 38615 -14235
rect 38670 -14355 38790 -14235
rect 38835 -14355 38955 -14235
rect 39000 -14355 39120 -14235
rect 39165 -14355 39285 -14235
rect 39340 -14355 39460 -14235
rect 39505 -14355 39625 -14235
rect 39670 -14355 39790 -14235
rect 39835 -14355 39955 -14235
rect 40010 -14355 40130 -14235
rect 40175 -14355 40295 -14235
rect 40340 -14355 40460 -14235
rect 40505 -14355 40625 -14235
rect 40680 -14355 40800 -14235
rect 40845 -14355 40965 -14235
rect 41010 -14355 41130 -14235
rect 41175 -14355 41295 -14235
rect 41350 -14355 41470 -14235
rect 41515 -14355 41635 -14235
rect 41680 -14355 41800 -14235
rect 41845 -14355 41965 -14235
rect 36485 -14520 36605 -14400
rect 36660 -14520 36780 -14400
rect 36825 -14520 36945 -14400
rect 36990 -14520 37110 -14400
rect 37155 -14520 37275 -14400
rect 37330 -14520 37450 -14400
rect 37495 -14520 37615 -14400
rect 37660 -14520 37780 -14400
rect 37825 -14520 37945 -14400
rect 38000 -14520 38120 -14400
rect 38165 -14520 38285 -14400
rect 38330 -14520 38450 -14400
rect 38495 -14520 38615 -14400
rect 38670 -14520 38790 -14400
rect 38835 -14520 38955 -14400
rect 39000 -14520 39120 -14400
rect 39165 -14520 39285 -14400
rect 39340 -14520 39460 -14400
rect 39505 -14520 39625 -14400
rect 39670 -14520 39790 -14400
rect 39835 -14520 39955 -14400
rect 40010 -14520 40130 -14400
rect 40175 -14520 40295 -14400
rect 40340 -14520 40460 -14400
rect 40505 -14520 40625 -14400
rect 40680 -14520 40800 -14400
rect 40845 -14520 40965 -14400
rect 41010 -14520 41130 -14400
rect 41175 -14520 41295 -14400
rect 41350 -14520 41470 -14400
rect 41515 -14520 41635 -14400
rect 41680 -14520 41800 -14400
rect 41845 -14520 41965 -14400
rect 36485 -14685 36605 -14565
rect 36660 -14685 36780 -14565
rect 36825 -14685 36945 -14565
rect 36990 -14685 37110 -14565
rect 37155 -14685 37275 -14565
rect 37330 -14685 37450 -14565
rect 37495 -14685 37615 -14565
rect 37660 -14685 37780 -14565
rect 37825 -14685 37945 -14565
rect 38000 -14685 38120 -14565
rect 38165 -14685 38285 -14565
rect 38330 -14685 38450 -14565
rect 38495 -14685 38615 -14565
rect 38670 -14685 38790 -14565
rect 38835 -14685 38955 -14565
rect 39000 -14685 39120 -14565
rect 39165 -14685 39285 -14565
rect 39340 -14685 39460 -14565
rect 39505 -14685 39625 -14565
rect 39670 -14685 39790 -14565
rect 39835 -14685 39955 -14565
rect 40010 -14685 40130 -14565
rect 40175 -14685 40295 -14565
rect 40340 -14685 40460 -14565
rect 40505 -14685 40625 -14565
rect 40680 -14685 40800 -14565
rect 40845 -14685 40965 -14565
rect 41010 -14685 41130 -14565
rect 41175 -14685 41295 -14565
rect 41350 -14685 41470 -14565
rect 41515 -14685 41635 -14565
rect 41680 -14685 41800 -14565
rect 41845 -14685 41965 -14565
rect 36485 -14860 36605 -14740
rect 36660 -14860 36780 -14740
rect 36825 -14860 36945 -14740
rect 36990 -14860 37110 -14740
rect 37155 -14860 37275 -14740
rect 37330 -14860 37450 -14740
rect 37495 -14860 37615 -14740
rect 37660 -14860 37780 -14740
rect 37825 -14860 37945 -14740
rect 38000 -14860 38120 -14740
rect 38165 -14860 38285 -14740
rect 38330 -14860 38450 -14740
rect 38495 -14860 38615 -14740
rect 38670 -14860 38790 -14740
rect 38835 -14860 38955 -14740
rect 39000 -14860 39120 -14740
rect 39165 -14860 39285 -14740
rect 39340 -14860 39460 -14740
rect 39505 -14860 39625 -14740
rect 39670 -14860 39790 -14740
rect 39835 -14860 39955 -14740
rect 40010 -14860 40130 -14740
rect 40175 -14860 40295 -14740
rect 40340 -14860 40460 -14740
rect 40505 -14860 40625 -14740
rect 40680 -14860 40800 -14740
rect 40845 -14860 40965 -14740
rect 41010 -14860 41130 -14740
rect 41175 -14860 41295 -14740
rect 41350 -14860 41470 -14740
rect 41515 -14860 41635 -14740
rect 41680 -14860 41800 -14740
rect 41845 -14860 41965 -14740
rect 36485 -15025 36605 -14905
rect 36660 -15025 36780 -14905
rect 36825 -15025 36945 -14905
rect 36990 -15025 37110 -14905
rect 37155 -15025 37275 -14905
rect 37330 -15025 37450 -14905
rect 37495 -15025 37615 -14905
rect 37660 -15025 37780 -14905
rect 37825 -15025 37945 -14905
rect 38000 -15025 38120 -14905
rect 38165 -15025 38285 -14905
rect 38330 -15025 38450 -14905
rect 38495 -15025 38615 -14905
rect 38670 -15025 38790 -14905
rect 38835 -15025 38955 -14905
rect 39000 -15025 39120 -14905
rect 39165 -15025 39285 -14905
rect 39340 -15025 39460 -14905
rect 39505 -15025 39625 -14905
rect 39670 -15025 39790 -14905
rect 39835 -15025 39955 -14905
rect 40010 -15025 40130 -14905
rect 40175 -15025 40295 -14905
rect 40340 -15025 40460 -14905
rect 40505 -15025 40625 -14905
rect 40680 -15025 40800 -14905
rect 40845 -15025 40965 -14905
rect 41010 -15025 41130 -14905
rect 41175 -15025 41295 -14905
rect 41350 -15025 41470 -14905
rect 41515 -15025 41635 -14905
rect 41680 -15025 41800 -14905
rect 41845 -15025 41965 -14905
rect 36485 -15190 36605 -15070
rect 36660 -15190 36780 -15070
rect 36825 -15190 36945 -15070
rect 36990 -15190 37110 -15070
rect 37155 -15190 37275 -15070
rect 37330 -15190 37450 -15070
rect 37495 -15190 37615 -15070
rect 37660 -15190 37780 -15070
rect 37825 -15190 37945 -15070
rect 38000 -15190 38120 -15070
rect 38165 -15190 38285 -15070
rect 38330 -15190 38450 -15070
rect 38495 -15190 38615 -15070
rect 38670 -15190 38790 -15070
rect 38835 -15190 38955 -15070
rect 39000 -15190 39120 -15070
rect 39165 -15190 39285 -15070
rect 39340 -15190 39460 -15070
rect 39505 -15190 39625 -15070
rect 39670 -15190 39790 -15070
rect 39835 -15190 39955 -15070
rect 40010 -15190 40130 -15070
rect 40175 -15190 40295 -15070
rect 40340 -15190 40460 -15070
rect 40505 -15190 40625 -15070
rect 40680 -15190 40800 -15070
rect 40845 -15190 40965 -15070
rect 41010 -15190 41130 -15070
rect 41175 -15190 41295 -15070
rect 41350 -15190 41470 -15070
rect 41515 -15190 41635 -15070
rect 41680 -15190 41800 -15070
rect 41845 -15190 41965 -15070
rect 36485 -15355 36605 -15235
rect 36660 -15355 36780 -15235
rect 36825 -15355 36945 -15235
rect 36990 -15355 37110 -15235
rect 37155 -15355 37275 -15235
rect 37330 -15355 37450 -15235
rect 37495 -15355 37615 -15235
rect 37660 -15355 37780 -15235
rect 37825 -15355 37945 -15235
rect 38000 -15355 38120 -15235
rect 38165 -15355 38285 -15235
rect 38330 -15355 38450 -15235
rect 38495 -15355 38615 -15235
rect 38670 -15355 38790 -15235
rect 38835 -15355 38955 -15235
rect 39000 -15355 39120 -15235
rect 39165 -15355 39285 -15235
rect 39340 -15355 39460 -15235
rect 39505 -15355 39625 -15235
rect 39670 -15355 39790 -15235
rect 39835 -15355 39955 -15235
rect 40010 -15355 40130 -15235
rect 40175 -15355 40295 -15235
rect 40340 -15355 40460 -15235
rect 40505 -15355 40625 -15235
rect 40680 -15355 40800 -15235
rect 40845 -15355 40965 -15235
rect 41010 -15355 41130 -15235
rect 41175 -15355 41295 -15235
rect 41350 -15355 41470 -15235
rect 41515 -15355 41635 -15235
rect 41680 -15355 41800 -15235
rect 41845 -15355 41965 -15235
rect 36485 -15530 36605 -15410
rect 36660 -15530 36780 -15410
rect 36825 -15530 36945 -15410
rect 36990 -15530 37110 -15410
rect 37155 -15530 37275 -15410
rect 37330 -15530 37450 -15410
rect 37495 -15530 37615 -15410
rect 37660 -15530 37780 -15410
rect 37825 -15530 37945 -15410
rect 38000 -15530 38120 -15410
rect 38165 -15530 38285 -15410
rect 38330 -15530 38450 -15410
rect 38495 -15530 38615 -15410
rect 38670 -15530 38790 -15410
rect 38835 -15530 38955 -15410
rect 39000 -15530 39120 -15410
rect 39165 -15530 39285 -15410
rect 39340 -15530 39460 -15410
rect 39505 -15530 39625 -15410
rect 39670 -15530 39790 -15410
rect 39835 -15530 39955 -15410
rect 40010 -15530 40130 -15410
rect 40175 -15530 40295 -15410
rect 40340 -15530 40460 -15410
rect 40505 -15530 40625 -15410
rect 40680 -15530 40800 -15410
rect 40845 -15530 40965 -15410
rect 41010 -15530 41130 -15410
rect 41175 -15530 41295 -15410
rect 41350 -15530 41470 -15410
rect 41515 -15530 41635 -15410
rect 41680 -15530 41800 -15410
rect 41845 -15530 41965 -15410
rect 42175 -10170 42295 -10050
rect 42350 -10170 42470 -10050
rect 42515 -10170 42635 -10050
rect 42680 -10170 42800 -10050
rect 42845 -10170 42965 -10050
rect 43020 -10170 43140 -10050
rect 43185 -10170 43305 -10050
rect 43350 -10170 43470 -10050
rect 43515 -10170 43635 -10050
rect 43690 -10170 43810 -10050
rect 43855 -10170 43975 -10050
rect 44020 -10170 44140 -10050
rect 44185 -10170 44305 -10050
rect 44360 -10170 44480 -10050
rect 44525 -10170 44645 -10050
rect 44690 -10170 44810 -10050
rect 44855 -10170 44975 -10050
rect 45030 -10170 45150 -10050
rect 45195 -10170 45315 -10050
rect 45360 -10170 45480 -10050
rect 45525 -10170 45645 -10050
rect 45700 -10170 45820 -10050
rect 45865 -10170 45985 -10050
rect 46030 -10170 46150 -10050
rect 46195 -10170 46315 -10050
rect 46370 -10170 46490 -10050
rect 46535 -10170 46655 -10050
rect 46700 -10170 46820 -10050
rect 46865 -10170 46985 -10050
rect 47040 -10170 47160 -10050
rect 47205 -10170 47325 -10050
rect 47370 -10170 47490 -10050
rect 47535 -10170 47655 -10050
rect 42175 -10335 42295 -10215
rect 42350 -10335 42470 -10215
rect 42515 -10335 42635 -10215
rect 42680 -10335 42800 -10215
rect 42845 -10335 42965 -10215
rect 43020 -10335 43140 -10215
rect 43185 -10335 43305 -10215
rect 43350 -10335 43470 -10215
rect 43515 -10335 43635 -10215
rect 43690 -10335 43810 -10215
rect 43855 -10335 43975 -10215
rect 44020 -10335 44140 -10215
rect 44185 -10335 44305 -10215
rect 44360 -10335 44480 -10215
rect 44525 -10335 44645 -10215
rect 44690 -10335 44810 -10215
rect 44855 -10335 44975 -10215
rect 45030 -10335 45150 -10215
rect 45195 -10335 45315 -10215
rect 45360 -10335 45480 -10215
rect 45525 -10335 45645 -10215
rect 45700 -10335 45820 -10215
rect 45865 -10335 45985 -10215
rect 46030 -10335 46150 -10215
rect 46195 -10335 46315 -10215
rect 46370 -10335 46490 -10215
rect 46535 -10335 46655 -10215
rect 46700 -10335 46820 -10215
rect 46865 -10335 46985 -10215
rect 47040 -10335 47160 -10215
rect 47205 -10335 47325 -10215
rect 47370 -10335 47490 -10215
rect 47535 -10335 47655 -10215
rect 42175 -10500 42295 -10380
rect 42350 -10500 42470 -10380
rect 42515 -10500 42635 -10380
rect 42680 -10500 42800 -10380
rect 42845 -10500 42965 -10380
rect 43020 -10500 43140 -10380
rect 43185 -10500 43305 -10380
rect 43350 -10500 43470 -10380
rect 43515 -10500 43635 -10380
rect 43690 -10500 43810 -10380
rect 43855 -10500 43975 -10380
rect 44020 -10500 44140 -10380
rect 44185 -10500 44305 -10380
rect 44360 -10500 44480 -10380
rect 44525 -10500 44645 -10380
rect 44690 -10500 44810 -10380
rect 44855 -10500 44975 -10380
rect 45030 -10500 45150 -10380
rect 45195 -10500 45315 -10380
rect 45360 -10500 45480 -10380
rect 45525 -10500 45645 -10380
rect 45700 -10500 45820 -10380
rect 45865 -10500 45985 -10380
rect 46030 -10500 46150 -10380
rect 46195 -10500 46315 -10380
rect 46370 -10500 46490 -10380
rect 46535 -10500 46655 -10380
rect 46700 -10500 46820 -10380
rect 46865 -10500 46985 -10380
rect 47040 -10500 47160 -10380
rect 47205 -10500 47325 -10380
rect 47370 -10500 47490 -10380
rect 47535 -10500 47655 -10380
rect 42175 -10665 42295 -10545
rect 42350 -10665 42470 -10545
rect 42515 -10665 42635 -10545
rect 42680 -10665 42800 -10545
rect 42845 -10665 42965 -10545
rect 43020 -10665 43140 -10545
rect 43185 -10665 43305 -10545
rect 43350 -10665 43470 -10545
rect 43515 -10665 43635 -10545
rect 43690 -10665 43810 -10545
rect 43855 -10665 43975 -10545
rect 44020 -10665 44140 -10545
rect 44185 -10665 44305 -10545
rect 44360 -10665 44480 -10545
rect 44525 -10665 44645 -10545
rect 44690 -10665 44810 -10545
rect 44855 -10665 44975 -10545
rect 45030 -10665 45150 -10545
rect 45195 -10665 45315 -10545
rect 45360 -10665 45480 -10545
rect 45525 -10665 45645 -10545
rect 45700 -10665 45820 -10545
rect 45865 -10665 45985 -10545
rect 46030 -10665 46150 -10545
rect 46195 -10665 46315 -10545
rect 46370 -10665 46490 -10545
rect 46535 -10665 46655 -10545
rect 46700 -10665 46820 -10545
rect 46865 -10665 46985 -10545
rect 47040 -10665 47160 -10545
rect 47205 -10665 47325 -10545
rect 47370 -10665 47490 -10545
rect 47535 -10665 47655 -10545
rect 42175 -10840 42295 -10720
rect 42350 -10840 42470 -10720
rect 42515 -10840 42635 -10720
rect 42680 -10840 42800 -10720
rect 42845 -10840 42965 -10720
rect 43020 -10840 43140 -10720
rect 43185 -10840 43305 -10720
rect 43350 -10840 43470 -10720
rect 43515 -10840 43635 -10720
rect 43690 -10840 43810 -10720
rect 43855 -10840 43975 -10720
rect 44020 -10840 44140 -10720
rect 44185 -10840 44305 -10720
rect 44360 -10840 44480 -10720
rect 44525 -10840 44645 -10720
rect 44690 -10840 44810 -10720
rect 44855 -10840 44975 -10720
rect 45030 -10840 45150 -10720
rect 45195 -10840 45315 -10720
rect 45360 -10840 45480 -10720
rect 45525 -10840 45645 -10720
rect 45700 -10840 45820 -10720
rect 45865 -10840 45985 -10720
rect 46030 -10840 46150 -10720
rect 46195 -10840 46315 -10720
rect 46370 -10840 46490 -10720
rect 46535 -10840 46655 -10720
rect 46700 -10840 46820 -10720
rect 46865 -10840 46985 -10720
rect 47040 -10840 47160 -10720
rect 47205 -10840 47325 -10720
rect 47370 -10840 47490 -10720
rect 47535 -10840 47655 -10720
rect 42175 -11005 42295 -10885
rect 42350 -11005 42470 -10885
rect 42515 -11005 42635 -10885
rect 42680 -11005 42800 -10885
rect 42845 -11005 42965 -10885
rect 43020 -11005 43140 -10885
rect 43185 -11005 43305 -10885
rect 43350 -11005 43470 -10885
rect 43515 -11005 43635 -10885
rect 43690 -11005 43810 -10885
rect 43855 -11005 43975 -10885
rect 44020 -11005 44140 -10885
rect 44185 -11005 44305 -10885
rect 44360 -11005 44480 -10885
rect 44525 -11005 44645 -10885
rect 44690 -11005 44810 -10885
rect 44855 -11005 44975 -10885
rect 45030 -11005 45150 -10885
rect 45195 -11005 45315 -10885
rect 45360 -11005 45480 -10885
rect 45525 -11005 45645 -10885
rect 45700 -11005 45820 -10885
rect 45865 -11005 45985 -10885
rect 46030 -11005 46150 -10885
rect 46195 -11005 46315 -10885
rect 46370 -11005 46490 -10885
rect 46535 -11005 46655 -10885
rect 46700 -11005 46820 -10885
rect 46865 -11005 46985 -10885
rect 47040 -11005 47160 -10885
rect 47205 -11005 47325 -10885
rect 47370 -11005 47490 -10885
rect 47535 -11005 47655 -10885
rect 42175 -11170 42295 -11050
rect 42350 -11170 42470 -11050
rect 42515 -11170 42635 -11050
rect 42680 -11170 42800 -11050
rect 42845 -11170 42965 -11050
rect 43020 -11170 43140 -11050
rect 43185 -11170 43305 -11050
rect 43350 -11170 43470 -11050
rect 43515 -11170 43635 -11050
rect 43690 -11170 43810 -11050
rect 43855 -11170 43975 -11050
rect 44020 -11170 44140 -11050
rect 44185 -11170 44305 -11050
rect 44360 -11170 44480 -11050
rect 44525 -11170 44645 -11050
rect 44690 -11170 44810 -11050
rect 44855 -11170 44975 -11050
rect 45030 -11170 45150 -11050
rect 45195 -11170 45315 -11050
rect 45360 -11170 45480 -11050
rect 45525 -11170 45645 -11050
rect 45700 -11170 45820 -11050
rect 45865 -11170 45985 -11050
rect 46030 -11170 46150 -11050
rect 46195 -11170 46315 -11050
rect 46370 -11170 46490 -11050
rect 46535 -11170 46655 -11050
rect 46700 -11170 46820 -11050
rect 46865 -11170 46985 -11050
rect 47040 -11170 47160 -11050
rect 47205 -11170 47325 -11050
rect 47370 -11170 47490 -11050
rect 47535 -11170 47655 -11050
rect 42175 -11335 42295 -11215
rect 42350 -11335 42470 -11215
rect 42515 -11335 42635 -11215
rect 42680 -11335 42800 -11215
rect 42845 -11335 42965 -11215
rect 43020 -11335 43140 -11215
rect 43185 -11335 43305 -11215
rect 43350 -11335 43470 -11215
rect 43515 -11335 43635 -11215
rect 43690 -11335 43810 -11215
rect 43855 -11335 43975 -11215
rect 44020 -11335 44140 -11215
rect 44185 -11335 44305 -11215
rect 44360 -11335 44480 -11215
rect 44525 -11335 44645 -11215
rect 44690 -11335 44810 -11215
rect 44855 -11335 44975 -11215
rect 45030 -11335 45150 -11215
rect 45195 -11335 45315 -11215
rect 45360 -11335 45480 -11215
rect 45525 -11335 45645 -11215
rect 45700 -11335 45820 -11215
rect 45865 -11335 45985 -11215
rect 46030 -11335 46150 -11215
rect 46195 -11335 46315 -11215
rect 46370 -11335 46490 -11215
rect 46535 -11335 46655 -11215
rect 46700 -11335 46820 -11215
rect 46865 -11335 46985 -11215
rect 47040 -11335 47160 -11215
rect 47205 -11335 47325 -11215
rect 47370 -11335 47490 -11215
rect 47535 -11335 47655 -11215
rect 42175 -11510 42295 -11390
rect 42350 -11510 42470 -11390
rect 42515 -11510 42635 -11390
rect 42680 -11510 42800 -11390
rect 42845 -11510 42965 -11390
rect 43020 -11510 43140 -11390
rect 43185 -11510 43305 -11390
rect 43350 -11510 43470 -11390
rect 43515 -11510 43635 -11390
rect 43690 -11510 43810 -11390
rect 43855 -11510 43975 -11390
rect 44020 -11510 44140 -11390
rect 44185 -11510 44305 -11390
rect 44360 -11510 44480 -11390
rect 44525 -11510 44645 -11390
rect 44690 -11510 44810 -11390
rect 44855 -11510 44975 -11390
rect 45030 -11510 45150 -11390
rect 45195 -11510 45315 -11390
rect 45360 -11510 45480 -11390
rect 45525 -11510 45645 -11390
rect 45700 -11510 45820 -11390
rect 45865 -11510 45985 -11390
rect 46030 -11510 46150 -11390
rect 46195 -11510 46315 -11390
rect 46370 -11510 46490 -11390
rect 46535 -11510 46655 -11390
rect 46700 -11510 46820 -11390
rect 46865 -11510 46985 -11390
rect 47040 -11510 47160 -11390
rect 47205 -11510 47325 -11390
rect 47370 -11510 47490 -11390
rect 47535 -11510 47655 -11390
rect 42175 -11675 42295 -11555
rect 42350 -11675 42470 -11555
rect 42515 -11675 42635 -11555
rect 42680 -11675 42800 -11555
rect 42845 -11675 42965 -11555
rect 43020 -11675 43140 -11555
rect 43185 -11675 43305 -11555
rect 43350 -11675 43470 -11555
rect 43515 -11675 43635 -11555
rect 43690 -11675 43810 -11555
rect 43855 -11675 43975 -11555
rect 44020 -11675 44140 -11555
rect 44185 -11675 44305 -11555
rect 44360 -11675 44480 -11555
rect 44525 -11675 44645 -11555
rect 44690 -11675 44810 -11555
rect 44855 -11675 44975 -11555
rect 45030 -11675 45150 -11555
rect 45195 -11675 45315 -11555
rect 45360 -11675 45480 -11555
rect 45525 -11675 45645 -11555
rect 45700 -11675 45820 -11555
rect 45865 -11675 45985 -11555
rect 46030 -11675 46150 -11555
rect 46195 -11675 46315 -11555
rect 46370 -11675 46490 -11555
rect 46535 -11675 46655 -11555
rect 46700 -11675 46820 -11555
rect 46865 -11675 46985 -11555
rect 47040 -11675 47160 -11555
rect 47205 -11675 47325 -11555
rect 47370 -11675 47490 -11555
rect 47535 -11675 47655 -11555
rect 42175 -11840 42295 -11720
rect 42350 -11840 42470 -11720
rect 42515 -11840 42635 -11720
rect 42680 -11840 42800 -11720
rect 42845 -11840 42965 -11720
rect 43020 -11840 43140 -11720
rect 43185 -11840 43305 -11720
rect 43350 -11840 43470 -11720
rect 43515 -11840 43635 -11720
rect 43690 -11840 43810 -11720
rect 43855 -11840 43975 -11720
rect 44020 -11840 44140 -11720
rect 44185 -11840 44305 -11720
rect 44360 -11840 44480 -11720
rect 44525 -11840 44645 -11720
rect 44690 -11840 44810 -11720
rect 44855 -11840 44975 -11720
rect 45030 -11840 45150 -11720
rect 45195 -11840 45315 -11720
rect 45360 -11840 45480 -11720
rect 45525 -11840 45645 -11720
rect 45700 -11840 45820 -11720
rect 45865 -11840 45985 -11720
rect 46030 -11840 46150 -11720
rect 46195 -11840 46315 -11720
rect 46370 -11840 46490 -11720
rect 46535 -11840 46655 -11720
rect 46700 -11840 46820 -11720
rect 46865 -11840 46985 -11720
rect 47040 -11840 47160 -11720
rect 47205 -11840 47325 -11720
rect 47370 -11840 47490 -11720
rect 47535 -11840 47655 -11720
rect 42175 -12005 42295 -11885
rect 42350 -12005 42470 -11885
rect 42515 -12005 42635 -11885
rect 42680 -12005 42800 -11885
rect 42845 -12005 42965 -11885
rect 43020 -12005 43140 -11885
rect 43185 -12005 43305 -11885
rect 43350 -12005 43470 -11885
rect 43515 -12005 43635 -11885
rect 43690 -12005 43810 -11885
rect 43855 -12005 43975 -11885
rect 44020 -12005 44140 -11885
rect 44185 -12005 44305 -11885
rect 44360 -12005 44480 -11885
rect 44525 -12005 44645 -11885
rect 44690 -12005 44810 -11885
rect 44855 -12005 44975 -11885
rect 45030 -12005 45150 -11885
rect 45195 -12005 45315 -11885
rect 45360 -12005 45480 -11885
rect 45525 -12005 45645 -11885
rect 45700 -12005 45820 -11885
rect 45865 -12005 45985 -11885
rect 46030 -12005 46150 -11885
rect 46195 -12005 46315 -11885
rect 46370 -12005 46490 -11885
rect 46535 -12005 46655 -11885
rect 46700 -12005 46820 -11885
rect 46865 -12005 46985 -11885
rect 47040 -12005 47160 -11885
rect 47205 -12005 47325 -11885
rect 47370 -12005 47490 -11885
rect 47535 -12005 47655 -11885
rect 42175 -12180 42295 -12060
rect 42350 -12180 42470 -12060
rect 42515 -12180 42635 -12060
rect 42680 -12180 42800 -12060
rect 42845 -12180 42965 -12060
rect 43020 -12180 43140 -12060
rect 43185 -12180 43305 -12060
rect 43350 -12180 43470 -12060
rect 43515 -12180 43635 -12060
rect 43690 -12180 43810 -12060
rect 43855 -12180 43975 -12060
rect 44020 -12180 44140 -12060
rect 44185 -12180 44305 -12060
rect 44360 -12180 44480 -12060
rect 44525 -12180 44645 -12060
rect 44690 -12180 44810 -12060
rect 44855 -12180 44975 -12060
rect 45030 -12180 45150 -12060
rect 45195 -12180 45315 -12060
rect 45360 -12180 45480 -12060
rect 45525 -12180 45645 -12060
rect 45700 -12180 45820 -12060
rect 45865 -12180 45985 -12060
rect 46030 -12180 46150 -12060
rect 46195 -12180 46315 -12060
rect 46370 -12180 46490 -12060
rect 46535 -12180 46655 -12060
rect 46700 -12180 46820 -12060
rect 46865 -12180 46985 -12060
rect 47040 -12180 47160 -12060
rect 47205 -12180 47325 -12060
rect 47370 -12180 47490 -12060
rect 47535 -12180 47655 -12060
rect 42175 -12345 42295 -12225
rect 42350 -12345 42470 -12225
rect 42515 -12345 42635 -12225
rect 42680 -12345 42800 -12225
rect 42845 -12345 42965 -12225
rect 43020 -12345 43140 -12225
rect 43185 -12345 43305 -12225
rect 43350 -12345 43470 -12225
rect 43515 -12345 43635 -12225
rect 43690 -12345 43810 -12225
rect 43855 -12345 43975 -12225
rect 44020 -12345 44140 -12225
rect 44185 -12345 44305 -12225
rect 44360 -12345 44480 -12225
rect 44525 -12345 44645 -12225
rect 44690 -12345 44810 -12225
rect 44855 -12345 44975 -12225
rect 45030 -12345 45150 -12225
rect 45195 -12345 45315 -12225
rect 45360 -12345 45480 -12225
rect 45525 -12345 45645 -12225
rect 45700 -12345 45820 -12225
rect 45865 -12345 45985 -12225
rect 46030 -12345 46150 -12225
rect 46195 -12345 46315 -12225
rect 46370 -12345 46490 -12225
rect 46535 -12345 46655 -12225
rect 46700 -12345 46820 -12225
rect 46865 -12345 46985 -12225
rect 47040 -12345 47160 -12225
rect 47205 -12345 47325 -12225
rect 47370 -12345 47490 -12225
rect 47535 -12345 47655 -12225
rect 42175 -12510 42295 -12390
rect 42350 -12510 42470 -12390
rect 42515 -12510 42635 -12390
rect 42680 -12510 42800 -12390
rect 42845 -12510 42965 -12390
rect 43020 -12510 43140 -12390
rect 43185 -12510 43305 -12390
rect 43350 -12510 43470 -12390
rect 43515 -12510 43635 -12390
rect 43690 -12510 43810 -12390
rect 43855 -12510 43975 -12390
rect 44020 -12510 44140 -12390
rect 44185 -12510 44305 -12390
rect 44360 -12510 44480 -12390
rect 44525 -12510 44645 -12390
rect 44690 -12510 44810 -12390
rect 44855 -12510 44975 -12390
rect 45030 -12510 45150 -12390
rect 45195 -12510 45315 -12390
rect 45360 -12510 45480 -12390
rect 45525 -12510 45645 -12390
rect 45700 -12510 45820 -12390
rect 45865 -12510 45985 -12390
rect 46030 -12510 46150 -12390
rect 46195 -12510 46315 -12390
rect 46370 -12510 46490 -12390
rect 46535 -12510 46655 -12390
rect 46700 -12510 46820 -12390
rect 46865 -12510 46985 -12390
rect 47040 -12510 47160 -12390
rect 47205 -12510 47325 -12390
rect 47370 -12510 47490 -12390
rect 47535 -12510 47655 -12390
rect 42175 -12675 42295 -12555
rect 42350 -12675 42470 -12555
rect 42515 -12675 42635 -12555
rect 42680 -12675 42800 -12555
rect 42845 -12675 42965 -12555
rect 43020 -12675 43140 -12555
rect 43185 -12675 43305 -12555
rect 43350 -12675 43470 -12555
rect 43515 -12675 43635 -12555
rect 43690 -12675 43810 -12555
rect 43855 -12675 43975 -12555
rect 44020 -12675 44140 -12555
rect 44185 -12675 44305 -12555
rect 44360 -12675 44480 -12555
rect 44525 -12675 44645 -12555
rect 44690 -12675 44810 -12555
rect 44855 -12675 44975 -12555
rect 45030 -12675 45150 -12555
rect 45195 -12675 45315 -12555
rect 45360 -12675 45480 -12555
rect 45525 -12675 45645 -12555
rect 45700 -12675 45820 -12555
rect 45865 -12675 45985 -12555
rect 46030 -12675 46150 -12555
rect 46195 -12675 46315 -12555
rect 46370 -12675 46490 -12555
rect 46535 -12675 46655 -12555
rect 46700 -12675 46820 -12555
rect 46865 -12675 46985 -12555
rect 47040 -12675 47160 -12555
rect 47205 -12675 47325 -12555
rect 47370 -12675 47490 -12555
rect 47535 -12675 47655 -12555
rect 42175 -12850 42295 -12730
rect 42350 -12850 42470 -12730
rect 42515 -12850 42635 -12730
rect 42680 -12850 42800 -12730
rect 42845 -12850 42965 -12730
rect 43020 -12850 43140 -12730
rect 43185 -12850 43305 -12730
rect 43350 -12850 43470 -12730
rect 43515 -12850 43635 -12730
rect 43690 -12850 43810 -12730
rect 43855 -12850 43975 -12730
rect 44020 -12850 44140 -12730
rect 44185 -12850 44305 -12730
rect 44360 -12850 44480 -12730
rect 44525 -12850 44645 -12730
rect 44690 -12850 44810 -12730
rect 44855 -12850 44975 -12730
rect 45030 -12850 45150 -12730
rect 45195 -12850 45315 -12730
rect 45360 -12850 45480 -12730
rect 45525 -12850 45645 -12730
rect 45700 -12850 45820 -12730
rect 45865 -12850 45985 -12730
rect 46030 -12850 46150 -12730
rect 46195 -12850 46315 -12730
rect 46370 -12850 46490 -12730
rect 46535 -12850 46655 -12730
rect 46700 -12850 46820 -12730
rect 46865 -12850 46985 -12730
rect 47040 -12850 47160 -12730
rect 47205 -12850 47325 -12730
rect 47370 -12850 47490 -12730
rect 47535 -12850 47655 -12730
rect 42175 -13015 42295 -12895
rect 42350 -13015 42470 -12895
rect 42515 -13015 42635 -12895
rect 42680 -13015 42800 -12895
rect 42845 -13015 42965 -12895
rect 43020 -13015 43140 -12895
rect 43185 -13015 43305 -12895
rect 43350 -13015 43470 -12895
rect 43515 -13015 43635 -12895
rect 43690 -13015 43810 -12895
rect 43855 -13015 43975 -12895
rect 44020 -13015 44140 -12895
rect 44185 -13015 44305 -12895
rect 44360 -13015 44480 -12895
rect 44525 -13015 44645 -12895
rect 44690 -13015 44810 -12895
rect 44855 -13015 44975 -12895
rect 45030 -13015 45150 -12895
rect 45195 -13015 45315 -12895
rect 45360 -13015 45480 -12895
rect 45525 -13015 45645 -12895
rect 45700 -13015 45820 -12895
rect 45865 -13015 45985 -12895
rect 46030 -13015 46150 -12895
rect 46195 -13015 46315 -12895
rect 46370 -13015 46490 -12895
rect 46535 -13015 46655 -12895
rect 46700 -13015 46820 -12895
rect 46865 -13015 46985 -12895
rect 47040 -13015 47160 -12895
rect 47205 -13015 47325 -12895
rect 47370 -13015 47490 -12895
rect 47535 -13015 47655 -12895
rect 42175 -13180 42295 -13060
rect 42350 -13180 42470 -13060
rect 42515 -13180 42635 -13060
rect 42680 -13180 42800 -13060
rect 42845 -13180 42965 -13060
rect 43020 -13180 43140 -13060
rect 43185 -13180 43305 -13060
rect 43350 -13180 43470 -13060
rect 43515 -13180 43635 -13060
rect 43690 -13180 43810 -13060
rect 43855 -13180 43975 -13060
rect 44020 -13180 44140 -13060
rect 44185 -13180 44305 -13060
rect 44360 -13180 44480 -13060
rect 44525 -13180 44645 -13060
rect 44690 -13180 44810 -13060
rect 44855 -13180 44975 -13060
rect 45030 -13180 45150 -13060
rect 45195 -13180 45315 -13060
rect 45360 -13180 45480 -13060
rect 45525 -13180 45645 -13060
rect 45700 -13180 45820 -13060
rect 45865 -13180 45985 -13060
rect 46030 -13180 46150 -13060
rect 46195 -13180 46315 -13060
rect 46370 -13180 46490 -13060
rect 46535 -13180 46655 -13060
rect 46700 -13180 46820 -13060
rect 46865 -13180 46985 -13060
rect 47040 -13180 47160 -13060
rect 47205 -13180 47325 -13060
rect 47370 -13180 47490 -13060
rect 47535 -13180 47655 -13060
rect 42175 -13345 42295 -13225
rect 42350 -13345 42470 -13225
rect 42515 -13345 42635 -13225
rect 42680 -13345 42800 -13225
rect 42845 -13345 42965 -13225
rect 43020 -13345 43140 -13225
rect 43185 -13345 43305 -13225
rect 43350 -13345 43470 -13225
rect 43515 -13345 43635 -13225
rect 43690 -13345 43810 -13225
rect 43855 -13345 43975 -13225
rect 44020 -13345 44140 -13225
rect 44185 -13345 44305 -13225
rect 44360 -13345 44480 -13225
rect 44525 -13345 44645 -13225
rect 44690 -13345 44810 -13225
rect 44855 -13345 44975 -13225
rect 45030 -13345 45150 -13225
rect 45195 -13345 45315 -13225
rect 45360 -13345 45480 -13225
rect 45525 -13345 45645 -13225
rect 45700 -13345 45820 -13225
rect 45865 -13345 45985 -13225
rect 46030 -13345 46150 -13225
rect 46195 -13345 46315 -13225
rect 46370 -13345 46490 -13225
rect 46535 -13345 46655 -13225
rect 46700 -13345 46820 -13225
rect 46865 -13345 46985 -13225
rect 47040 -13345 47160 -13225
rect 47205 -13345 47325 -13225
rect 47370 -13345 47490 -13225
rect 47535 -13345 47655 -13225
rect 42175 -13520 42295 -13400
rect 42350 -13520 42470 -13400
rect 42515 -13520 42635 -13400
rect 42680 -13520 42800 -13400
rect 42845 -13520 42965 -13400
rect 43020 -13520 43140 -13400
rect 43185 -13520 43305 -13400
rect 43350 -13520 43470 -13400
rect 43515 -13520 43635 -13400
rect 43690 -13520 43810 -13400
rect 43855 -13520 43975 -13400
rect 44020 -13520 44140 -13400
rect 44185 -13520 44305 -13400
rect 44360 -13520 44480 -13400
rect 44525 -13520 44645 -13400
rect 44690 -13520 44810 -13400
rect 44855 -13520 44975 -13400
rect 45030 -13520 45150 -13400
rect 45195 -13520 45315 -13400
rect 45360 -13520 45480 -13400
rect 45525 -13520 45645 -13400
rect 45700 -13520 45820 -13400
rect 45865 -13520 45985 -13400
rect 46030 -13520 46150 -13400
rect 46195 -13520 46315 -13400
rect 46370 -13520 46490 -13400
rect 46535 -13520 46655 -13400
rect 46700 -13520 46820 -13400
rect 46865 -13520 46985 -13400
rect 47040 -13520 47160 -13400
rect 47205 -13520 47325 -13400
rect 47370 -13520 47490 -13400
rect 47535 -13520 47655 -13400
rect 42175 -13685 42295 -13565
rect 42350 -13685 42470 -13565
rect 42515 -13685 42635 -13565
rect 42680 -13685 42800 -13565
rect 42845 -13685 42965 -13565
rect 43020 -13685 43140 -13565
rect 43185 -13685 43305 -13565
rect 43350 -13685 43470 -13565
rect 43515 -13685 43635 -13565
rect 43690 -13685 43810 -13565
rect 43855 -13685 43975 -13565
rect 44020 -13685 44140 -13565
rect 44185 -13685 44305 -13565
rect 44360 -13685 44480 -13565
rect 44525 -13685 44645 -13565
rect 44690 -13685 44810 -13565
rect 44855 -13685 44975 -13565
rect 45030 -13685 45150 -13565
rect 45195 -13685 45315 -13565
rect 45360 -13685 45480 -13565
rect 45525 -13685 45645 -13565
rect 45700 -13685 45820 -13565
rect 45865 -13685 45985 -13565
rect 46030 -13685 46150 -13565
rect 46195 -13685 46315 -13565
rect 46370 -13685 46490 -13565
rect 46535 -13685 46655 -13565
rect 46700 -13685 46820 -13565
rect 46865 -13685 46985 -13565
rect 47040 -13685 47160 -13565
rect 47205 -13685 47325 -13565
rect 47370 -13685 47490 -13565
rect 47535 -13685 47655 -13565
rect 42175 -13850 42295 -13730
rect 42350 -13850 42470 -13730
rect 42515 -13850 42635 -13730
rect 42680 -13850 42800 -13730
rect 42845 -13850 42965 -13730
rect 43020 -13850 43140 -13730
rect 43185 -13850 43305 -13730
rect 43350 -13850 43470 -13730
rect 43515 -13850 43635 -13730
rect 43690 -13850 43810 -13730
rect 43855 -13850 43975 -13730
rect 44020 -13850 44140 -13730
rect 44185 -13850 44305 -13730
rect 44360 -13850 44480 -13730
rect 44525 -13850 44645 -13730
rect 44690 -13850 44810 -13730
rect 44855 -13850 44975 -13730
rect 45030 -13850 45150 -13730
rect 45195 -13850 45315 -13730
rect 45360 -13850 45480 -13730
rect 45525 -13850 45645 -13730
rect 45700 -13850 45820 -13730
rect 45865 -13850 45985 -13730
rect 46030 -13850 46150 -13730
rect 46195 -13850 46315 -13730
rect 46370 -13850 46490 -13730
rect 46535 -13850 46655 -13730
rect 46700 -13850 46820 -13730
rect 46865 -13850 46985 -13730
rect 47040 -13850 47160 -13730
rect 47205 -13850 47325 -13730
rect 47370 -13850 47490 -13730
rect 47535 -13850 47655 -13730
rect 42175 -14015 42295 -13895
rect 42350 -14015 42470 -13895
rect 42515 -14015 42635 -13895
rect 42680 -14015 42800 -13895
rect 42845 -14015 42965 -13895
rect 43020 -14015 43140 -13895
rect 43185 -14015 43305 -13895
rect 43350 -14015 43470 -13895
rect 43515 -14015 43635 -13895
rect 43690 -14015 43810 -13895
rect 43855 -14015 43975 -13895
rect 44020 -14015 44140 -13895
rect 44185 -14015 44305 -13895
rect 44360 -14015 44480 -13895
rect 44525 -14015 44645 -13895
rect 44690 -14015 44810 -13895
rect 44855 -14015 44975 -13895
rect 45030 -14015 45150 -13895
rect 45195 -14015 45315 -13895
rect 45360 -14015 45480 -13895
rect 45525 -14015 45645 -13895
rect 45700 -14015 45820 -13895
rect 45865 -14015 45985 -13895
rect 46030 -14015 46150 -13895
rect 46195 -14015 46315 -13895
rect 46370 -14015 46490 -13895
rect 46535 -14015 46655 -13895
rect 46700 -14015 46820 -13895
rect 46865 -14015 46985 -13895
rect 47040 -14015 47160 -13895
rect 47205 -14015 47325 -13895
rect 47370 -14015 47490 -13895
rect 47535 -14015 47655 -13895
rect 42175 -14190 42295 -14070
rect 42350 -14190 42470 -14070
rect 42515 -14190 42635 -14070
rect 42680 -14190 42800 -14070
rect 42845 -14190 42965 -14070
rect 43020 -14190 43140 -14070
rect 43185 -14190 43305 -14070
rect 43350 -14190 43470 -14070
rect 43515 -14190 43635 -14070
rect 43690 -14190 43810 -14070
rect 43855 -14190 43975 -14070
rect 44020 -14190 44140 -14070
rect 44185 -14190 44305 -14070
rect 44360 -14190 44480 -14070
rect 44525 -14190 44645 -14070
rect 44690 -14190 44810 -14070
rect 44855 -14190 44975 -14070
rect 45030 -14190 45150 -14070
rect 45195 -14190 45315 -14070
rect 45360 -14190 45480 -14070
rect 45525 -14190 45645 -14070
rect 45700 -14190 45820 -14070
rect 45865 -14190 45985 -14070
rect 46030 -14190 46150 -14070
rect 46195 -14190 46315 -14070
rect 46370 -14190 46490 -14070
rect 46535 -14190 46655 -14070
rect 46700 -14190 46820 -14070
rect 46865 -14190 46985 -14070
rect 47040 -14190 47160 -14070
rect 47205 -14190 47325 -14070
rect 47370 -14190 47490 -14070
rect 47535 -14190 47655 -14070
rect 42175 -14355 42295 -14235
rect 42350 -14355 42470 -14235
rect 42515 -14355 42635 -14235
rect 42680 -14355 42800 -14235
rect 42845 -14355 42965 -14235
rect 43020 -14355 43140 -14235
rect 43185 -14355 43305 -14235
rect 43350 -14355 43470 -14235
rect 43515 -14355 43635 -14235
rect 43690 -14355 43810 -14235
rect 43855 -14355 43975 -14235
rect 44020 -14355 44140 -14235
rect 44185 -14355 44305 -14235
rect 44360 -14355 44480 -14235
rect 44525 -14355 44645 -14235
rect 44690 -14355 44810 -14235
rect 44855 -14355 44975 -14235
rect 45030 -14355 45150 -14235
rect 45195 -14355 45315 -14235
rect 45360 -14355 45480 -14235
rect 45525 -14355 45645 -14235
rect 45700 -14355 45820 -14235
rect 45865 -14355 45985 -14235
rect 46030 -14355 46150 -14235
rect 46195 -14355 46315 -14235
rect 46370 -14355 46490 -14235
rect 46535 -14355 46655 -14235
rect 46700 -14355 46820 -14235
rect 46865 -14355 46985 -14235
rect 47040 -14355 47160 -14235
rect 47205 -14355 47325 -14235
rect 47370 -14355 47490 -14235
rect 47535 -14355 47655 -14235
rect 42175 -14520 42295 -14400
rect 42350 -14520 42470 -14400
rect 42515 -14520 42635 -14400
rect 42680 -14520 42800 -14400
rect 42845 -14520 42965 -14400
rect 43020 -14520 43140 -14400
rect 43185 -14520 43305 -14400
rect 43350 -14520 43470 -14400
rect 43515 -14520 43635 -14400
rect 43690 -14520 43810 -14400
rect 43855 -14520 43975 -14400
rect 44020 -14520 44140 -14400
rect 44185 -14520 44305 -14400
rect 44360 -14520 44480 -14400
rect 44525 -14520 44645 -14400
rect 44690 -14520 44810 -14400
rect 44855 -14520 44975 -14400
rect 45030 -14520 45150 -14400
rect 45195 -14520 45315 -14400
rect 45360 -14520 45480 -14400
rect 45525 -14520 45645 -14400
rect 45700 -14520 45820 -14400
rect 45865 -14520 45985 -14400
rect 46030 -14520 46150 -14400
rect 46195 -14520 46315 -14400
rect 46370 -14520 46490 -14400
rect 46535 -14520 46655 -14400
rect 46700 -14520 46820 -14400
rect 46865 -14520 46985 -14400
rect 47040 -14520 47160 -14400
rect 47205 -14520 47325 -14400
rect 47370 -14520 47490 -14400
rect 47535 -14520 47655 -14400
rect 42175 -14685 42295 -14565
rect 42350 -14685 42470 -14565
rect 42515 -14685 42635 -14565
rect 42680 -14685 42800 -14565
rect 42845 -14685 42965 -14565
rect 43020 -14685 43140 -14565
rect 43185 -14685 43305 -14565
rect 43350 -14685 43470 -14565
rect 43515 -14685 43635 -14565
rect 43690 -14685 43810 -14565
rect 43855 -14685 43975 -14565
rect 44020 -14685 44140 -14565
rect 44185 -14685 44305 -14565
rect 44360 -14685 44480 -14565
rect 44525 -14685 44645 -14565
rect 44690 -14685 44810 -14565
rect 44855 -14685 44975 -14565
rect 45030 -14685 45150 -14565
rect 45195 -14685 45315 -14565
rect 45360 -14685 45480 -14565
rect 45525 -14685 45645 -14565
rect 45700 -14685 45820 -14565
rect 45865 -14685 45985 -14565
rect 46030 -14685 46150 -14565
rect 46195 -14685 46315 -14565
rect 46370 -14685 46490 -14565
rect 46535 -14685 46655 -14565
rect 46700 -14685 46820 -14565
rect 46865 -14685 46985 -14565
rect 47040 -14685 47160 -14565
rect 47205 -14685 47325 -14565
rect 47370 -14685 47490 -14565
rect 47535 -14685 47655 -14565
rect 42175 -14860 42295 -14740
rect 42350 -14860 42470 -14740
rect 42515 -14860 42635 -14740
rect 42680 -14860 42800 -14740
rect 42845 -14860 42965 -14740
rect 43020 -14860 43140 -14740
rect 43185 -14860 43305 -14740
rect 43350 -14860 43470 -14740
rect 43515 -14860 43635 -14740
rect 43690 -14860 43810 -14740
rect 43855 -14860 43975 -14740
rect 44020 -14860 44140 -14740
rect 44185 -14860 44305 -14740
rect 44360 -14860 44480 -14740
rect 44525 -14860 44645 -14740
rect 44690 -14860 44810 -14740
rect 44855 -14860 44975 -14740
rect 45030 -14860 45150 -14740
rect 45195 -14860 45315 -14740
rect 45360 -14860 45480 -14740
rect 45525 -14860 45645 -14740
rect 45700 -14860 45820 -14740
rect 45865 -14860 45985 -14740
rect 46030 -14860 46150 -14740
rect 46195 -14860 46315 -14740
rect 46370 -14860 46490 -14740
rect 46535 -14860 46655 -14740
rect 46700 -14860 46820 -14740
rect 46865 -14860 46985 -14740
rect 47040 -14860 47160 -14740
rect 47205 -14860 47325 -14740
rect 47370 -14860 47490 -14740
rect 47535 -14860 47655 -14740
rect 42175 -15025 42295 -14905
rect 42350 -15025 42470 -14905
rect 42515 -15025 42635 -14905
rect 42680 -15025 42800 -14905
rect 42845 -15025 42965 -14905
rect 43020 -15025 43140 -14905
rect 43185 -15025 43305 -14905
rect 43350 -15025 43470 -14905
rect 43515 -15025 43635 -14905
rect 43690 -15025 43810 -14905
rect 43855 -15025 43975 -14905
rect 44020 -15025 44140 -14905
rect 44185 -15025 44305 -14905
rect 44360 -15025 44480 -14905
rect 44525 -15025 44645 -14905
rect 44690 -15025 44810 -14905
rect 44855 -15025 44975 -14905
rect 45030 -15025 45150 -14905
rect 45195 -15025 45315 -14905
rect 45360 -15025 45480 -14905
rect 45525 -15025 45645 -14905
rect 45700 -15025 45820 -14905
rect 45865 -15025 45985 -14905
rect 46030 -15025 46150 -14905
rect 46195 -15025 46315 -14905
rect 46370 -15025 46490 -14905
rect 46535 -15025 46655 -14905
rect 46700 -15025 46820 -14905
rect 46865 -15025 46985 -14905
rect 47040 -15025 47160 -14905
rect 47205 -15025 47325 -14905
rect 47370 -15025 47490 -14905
rect 47535 -15025 47655 -14905
rect 42175 -15190 42295 -15070
rect 42350 -15190 42470 -15070
rect 42515 -15190 42635 -15070
rect 42680 -15190 42800 -15070
rect 42845 -15190 42965 -15070
rect 43020 -15190 43140 -15070
rect 43185 -15190 43305 -15070
rect 43350 -15190 43470 -15070
rect 43515 -15190 43635 -15070
rect 43690 -15190 43810 -15070
rect 43855 -15190 43975 -15070
rect 44020 -15190 44140 -15070
rect 44185 -15190 44305 -15070
rect 44360 -15190 44480 -15070
rect 44525 -15190 44645 -15070
rect 44690 -15190 44810 -15070
rect 44855 -15190 44975 -15070
rect 45030 -15190 45150 -15070
rect 45195 -15190 45315 -15070
rect 45360 -15190 45480 -15070
rect 45525 -15190 45645 -15070
rect 45700 -15190 45820 -15070
rect 45865 -15190 45985 -15070
rect 46030 -15190 46150 -15070
rect 46195 -15190 46315 -15070
rect 46370 -15190 46490 -15070
rect 46535 -15190 46655 -15070
rect 46700 -15190 46820 -15070
rect 46865 -15190 46985 -15070
rect 47040 -15190 47160 -15070
rect 47205 -15190 47325 -15070
rect 47370 -15190 47490 -15070
rect 47535 -15190 47655 -15070
rect 42175 -15355 42295 -15235
rect 42350 -15355 42470 -15235
rect 42515 -15355 42635 -15235
rect 42680 -15355 42800 -15235
rect 42845 -15355 42965 -15235
rect 43020 -15355 43140 -15235
rect 43185 -15355 43305 -15235
rect 43350 -15355 43470 -15235
rect 43515 -15355 43635 -15235
rect 43690 -15355 43810 -15235
rect 43855 -15355 43975 -15235
rect 44020 -15355 44140 -15235
rect 44185 -15355 44305 -15235
rect 44360 -15355 44480 -15235
rect 44525 -15355 44645 -15235
rect 44690 -15355 44810 -15235
rect 44855 -15355 44975 -15235
rect 45030 -15355 45150 -15235
rect 45195 -15355 45315 -15235
rect 45360 -15355 45480 -15235
rect 45525 -15355 45645 -15235
rect 45700 -15355 45820 -15235
rect 45865 -15355 45985 -15235
rect 46030 -15355 46150 -15235
rect 46195 -15355 46315 -15235
rect 46370 -15355 46490 -15235
rect 46535 -15355 46655 -15235
rect 46700 -15355 46820 -15235
rect 46865 -15355 46985 -15235
rect 47040 -15355 47160 -15235
rect 47205 -15355 47325 -15235
rect 47370 -15355 47490 -15235
rect 47535 -15355 47655 -15235
rect 42175 -15530 42295 -15410
rect 42350 -15530 42470 -15410
rect 42515 -15530 42635 -15410
rect 42680 -15530 42800 -15410
rect 42845 -15530 42965 -15410
rect 43020 -15530 43140 -15410
rect 43185 -15530 43305 -15410
rect 43350 -15530 43470 -15410
rect 43515 -15530 43635 -15410
rect 43690 -15530 43810 -15410
rect 43855 -15530 43975 -15410
rect 44020 -15530 44140 -15410
rect 44185 -15530 44305 -15410
rect 44360 -15530 44480 -15410
rect 44525 -15530 44645 -15410
rect 44690 -15530 44810 -15410
rect 44855 -15530 44975 -15410
rect 45030 -15530 45150 -15410
rect 45195 -15530 45315 -15410
rect 45360 -15530 45480 -15410
rect 45525 -15530 45645 -15410
rect 45700 -15530 45820 -15410
rect 45865 -15530 45985 -15410
rect 46030 -15530 46150 -15410
rect 46195 -15530 46315 -15410
rect 46370 -15530 46490 -15410
rect 46535 -15530 46655 -15410
rect 46700 -15530 46820 -15410
rect 46865 -15530 46985 -15410
rect 47040 -15530 47160 -15410
rect 47205 -15530 47325 -15410
rect 47370 -15530 47490 -15410
rect 47535 -15530 47655 -15410
rect 47865 -10170 47985 -10050
rect 48040 -10170 48160 -10050
rect 48205 -10170 48325 -10050
rect 48370 -10170 48490 -10050
rect 48535 -10170 48655 -10050
rect 48710 -10170 48830 -10050
rect 48875 -10170 48995 -10050
rect 49040 -10170 49160 -10050
rect 49205 -10170 49325 -10050
rect 49380 -10170 49500 -10050
rect 49545 -10170 49665 -10050
rect 49710 -10170 49830 -10050
rect 49875 -10170 49995 -10050
rect 50050 -10170 50170 -10050
rect 50215 -10170 50335 -10050
rect 50380 -10170 50500 -10050
rect 50545 -10170 50665 -10050
rect 50720 -10170 50840 -10050
rect 50885 -10170 51005 -10050
rect 51050 -10170 51170 -10050
rect 51215 -10170 51335 -10050
rect 51390 -10170 51510 -10050
rect 51555 -10170 51675 -10050
rect 51720 -10170 51840 -10050
rect 51885 -10170 52005 -10050
rect 52060 -10170 52180 -10050
rect 52225 -10170 52345 -10050
rect 52390 -10170 52510 -10050
rect 52555 -10170 52675 -10050
rect 52730 -10170 52850 -10050
rect 52895 -10170 53015 -10050
rect 53060 -10170 53180 -10050
rect 53225 -10170 53345 -10050
rect 47865 -10335 47985 -10215
rect 48040 -10335 48160 -10215
rect 48205 -10335 48325 -10215
rect 48370 -10335 48490 -10215
rect 48535 -10335 48655 -10215
rect 48710 -10335 48830 -10215
rect 48875 -10335 48995 -10215
rect 49040 -10335 49160 -10215
rect 49205 -10335 49325 -10215
rect 49380 -10335 49500 -10215
rect 49545 -10335 49665 -10215
rect 49710 -10335 49830 -10215
rect 49875 -10335 49995 -10215
rect 50050 -10335 50170 -10215
rect 50215 -10335 50335 -10215
rect 50380 -10335 50500 -10215
rect 50545 -10335 50665 -10215
rect 50720 -10335 50840 -10215
rect 50885 -10335 51005 -10215
rect 51050 -10335 51170 -10215
rect 51215 -10335 51335 -10215
rect 51390 -10335 51510 -10215
rect 51555 -10335 51675 -10215
rect 51720 -10335 51840 -10215
rect 51885 -10335 52005 -10215
rect 52060 -10335 52180 -10215
rect 52225 -10335 52345 -10215
rect 52390 -10335 52510 -10215
rect 52555 -10335 52675 -10215
rect 52730 -10335 52850 -10215
rect 52895 -10335 53015 -10215
rect 53060 -10335 53180 -10215
rect 53225 -10335 53345 -10215
rect 47865 -10500 47985 -10380
rect 48040 -10500 48160 -10380
rect 48205 -10500 48325 -10380
rect 48370 -10500 48490 -10380
rect 48535 -10500 48655 -10380
rect 48710 -10500 48830 -10380
rect 48875 -10500 48995 -10380
rect 49040 -10500 49160 -10380
rect 49205 -10500 49325 -10380
rect 49380 -10500 49500 -10380
rect 49545 -10500 49665 -10380
rect 49710 -10500 49830 -10380
rect 49875 -10500 49995 -10380
rect 50050 -10500 50170 -10380
rect 50215 -10500 50335 -10380
rect 50380 -10500 50500 -10380
rect 50545 -10500 50665 -10380
rect 50720 -10500 50840 -10380
rect 50885 -10500 51005 -10380
rect 51050 -10500 51170 -10380
rect 51215 -10500 51335 -10380
rect 51390 -10500 51510 -10380
rect 51555 -10500 51675 -10380
rect 51720 -10500 51840 -10380
rect 51885 -10500 52005 -10380
rect 52060 -10500 52180 -10380
rect 52225 -10500 52345 -10380
rect 52390 -10500 52510 -10380
rect 52555 -10500 52675 -10380
rect 52730 -10500 52850 -10380
rect 52895 -10500 53015 -10380
rect 53060 -10500 53180 -10380
rect 53225 -10500 53345 -10380
rect 47865 -10665 47985 -10545
rect 48040 -10665 48160 -10545
rect 48205 -10665 48325 -10545
rect 48370 -10665 48490 -10545
rect 48535 -10665 48655 -10545
rect 48710 -10665 48830 -10545
rect 48875 -10665 48995 -10545
rect 49040 -10665 49160 -10545
rect 49205 -10665 49325 -10545
rect 49380 -10665 49500 -10545
rect 49545 -10665 49665 -10545
rect 49710 -10665 49830 -10545
rect 49875 -10665 49995 -10545
rect 50050 -10665 50170 -10545
rect 50215 -10665 50335 -10545
rect 50380 -10665 50500 -10545
rect 50545 -10665 50665 -10545
rect 50720 -10665 50840 -10545
rect 50885 -10665 51005 -10545
rect 51050 -10665 51170 -10545
rect 51215 -10665 51335 -10545
rect 51390 -10665 51510 -10545
rect 51555 -10665 51675 -10545
rect 51720 -10665 51840 -10545
rect 51885 -10665 52005 -10545
rect 52060 -10665 52180 -10545
rect 52225 -10665 52345 -10545
rect 52390 -10665 52510 -10545
rect 52555 -10665 52675 -10545
rect 52730 -10665 52850 -10545
rect 52895 -10665 53015 -10545
rect 53060 -10665 53180 -10545
rect 53225 -10665 53345 -10545
rect 47865 -10840 47985 -10720
rect 48040 -10840 48160 -10720
rect 48205 -10840 48325 -10720
rect 48370 -10840 48490 -10720
rect 48535 -10840 48655 -10720
rect 48710 -10840 48830 -10720
rect 48875 -10840 48995 -10720
rect 49040 -10840 49160 -10720
rect 49205 -10840 49325 -10720
rect 49380 -10840 49500 -10720
rect 49545 -10840 49665 -10720
rect 49710 -10840 49830 -10720
rect 49875 -10840 49995 -10720
rect 50050 -10840 50170 -10720
rect 50215 -10840 50335 -10720
rect 50380 -10840 50500 -10720
rect 50545 -10840 50665 -10720
rect 50720 -10840 50840 -10720
rect 50885 -10840 51005 -10720
rect 51050 -10840 51170 -10720
rect 51215 -10840 51335 -10720
rect 51390 -10840 51510 -10720
rect 51555 -10840 51675 -10720
rect 51720 -10840 51840 -10720
rect 51885 -10840 52005 -10720
rect 52060 -10840 52180 -10720
rect 52225 -10840 52345 -10720
rect 52390 -10840 52510 -10720
rect 52555 -10840 52675 -10720
rect 52730 -10840 52850 -10720
rect 52895 -10840 53015 -10720
rect 53060 -10840 53180 -10720
rect 53225 -10840 53345 -10720
rect 47865 -11005 47985 -10885
rect 48040 -11005 48160 -10885
rect 48205 -11005 48325 -10885
rect 48370 -11005 48490 -10885
rect 48535 -11005 48655 -10885
rect 48710 -11005 48830 -10885
rect 48875 -11005 48995 -10885
rect 49040 -11005 49160 -10885
rect 49205 -11005 49325 -10885
rect 49380 -11005 49500 -10885
rect 49545 -11005 49665 -10885
rect 49710 -11005 49830 -10885
rect 49875 -11005 49995 -10885
rect 50050 -11005 50170 -10885
rect 50215 -11005 50335 -10885
rect 50380 -11005 50500 -10885
rect 50545 -11005 50665 -10885
rect 50720 -11005 50840 -10885
rect 50885 -11005 51005 -10885
rect 51050 -11005 51170 -10885
rect 51215 -11005 51335 -10885
rect 51390 -11005 51510 -10885
rect 51555 -11005 51675 -10885
rect 51720 -11005 51840 -10885
rect 51885 -11005 52005 -10885
rect 52060 -11005 52180 -10885
rect 52225 -11005 52345 -10885
rect 52390 -11005 52510 -10885
rect 52555 -11005 52675 -10885
rect 52730 -11005 52850 -10885
rect 52895 -11005 53015 -10885
rect 53060 -11005 53180 -10885
rect 53225 -11005 53345 -10885
rect 47865 -11170 47985 -11050
rect 48040 -11170 48160 -11050
rect 48205 -11170 48325 -11050
rect 48370 -11170 48490 -11050
rect 48535 -11170 48655 -11050
rect 48710 -11170 48830 -11050
rect 48875 -11170 48995 -11050
rect 49040 -11170 49160 -11050
rect 49205 -11170 49325 -11050
rect 49380 -11170 49500 -11050
rect 49545 -11170 49665 -11050
rect 49710 -11170 49830 -11050
rect 49875 -11170 49995 -11050
rect 50050 -11170 50170 -11050
rect 50215 -11170 50335 -11050
rect 50380 -11170 50500 -11050
rect 50545 -11170 50665 -11050
rect 50720 -11170 50840 -11050
rect 50885 -11170 51005 -11050
rect 51050 -11170 51170 -11050
rect 51215 -11170 51335 -11050
rect 51390 -11170 51510 -11050
rect 51555 -11170 51675 -11050
rect 51720 -11170 51840 -11050
rect 51885 -11170 52005 -11050
rect 52060 -11170 52180 -11050
rect 52225 -11170 52345 -11050
rect 52390 -11170 52510 -11050
rect 52555 -11170 52675 -11050
rect 52730 -11170 52850 -11050
rect 52895 -11170 53015 -11050
rect 53060 -11170 53180 -11050
rect 53225 -11170 53345 -11050
rect 47865 -11335 47985 -11215
rect 48040 -11335 48160 -11215
rect 48205 -11335 48325 -11215
rect 48370 -11335 48490 -11215
rect 48535 -11335 48655 -11215
rect 48710 -11335 48830 -11215
rect 48875 -11335 48995 -11215
rect 49040 -11335 49160 -11215
rect 49205 -11335 49325 -11215
rect 49380 -11335 49500 -11215
rect 49545 -11335 49665 -11215
rect 49710 -11335 49830 -11215
rect 49875 -11335 49995 -11215
rect 50050 -11335 50170 -11215
rect 50215 -11335 50335 -11215
rect 50380 -11335 50500 -11215
rect 50545 -11335 50665 -11215
rect 50720 -11335 50840 -11215
rect 50885 -11335 51005 -11215
rect 51050 -11335 51170 -11215
rect 51215 -11335 51335 -11215
rect 51390 -11335 51510 -11215
rect 51555 -11335 51675 -11215
rect 51720 -11335 51840 -11215
rect 51885 -11335 52005 -11215
rect 52060 -11335 52180 -11215
rect 52225 -11335 52345 -11215
rect 52390 -11335 52510 -11215
rect 52555 -11335 52675 -11215
rect 52730 -11335 52850 -11215
rect 52895 -11335 53015 -11215
rect 53060 -11335 53180 -11215
rect 53225 -11335 53345 -11215
rect 47865 -11510 47985 -11390
rect 48040 -11510 48160 -11390
rect 48205 -11510 48325 -11390
rect 48370 -11510 48490 -11390
rect 48535 -11510 48655 -11390
rect 48710 -11510 48830 -11390
rect 48875 -11510 48995 -11390
rect 49040 -11510 49160 -11390
rect 49205 -11510 49325 -11390
rect 49380 -11510 49500 -11390
rect 49545 -11510 49665 -11390
rect 49710 -11510 49830 -11390
rect 49875 -11510 49995 -11390
rect 50050 -11510 50170 -11390
rect 50215 -11510 50335 -11390
rect 50380 -11510 50500 -11390
rect 50545 -11510 50665 -11390
rect 50720 -11510 50840 -11390
rect 50885 -11510 51005 -11390
rect 51050 -11510 51170 -11390
rect 51215 -11510 51335 -11390
rect 51390 -11510 51510 -11390
rect 51555 -11510 51675 -11390
rect 51720 -11510 51840 -11390
rect 51885 -11510 52005 -11390
rect 52060 -11510 52180 -11390
rect 52225 -11510 52345 -11390
rect 52390 -11510 52510 -11390
rect 52555 -11510 52675 -11390
rect 52730 -11510 52850 -11390
rect 52895 -11510 53015 -11390
rect 53060 -11510 53180 -11390
rect 53225 -11510 53345 -11390
rect 47865 -11675 47985 -11555
rect 48040 -11675 48160 -11555
rect 48205 -11675 48325 -11555
rect 48370 -11675 48490 -11555
rect 48535 -11675 48655 -11555
rect 48710 -11675 48830 -11555
rect 48875 -11675 48995 -11555
rect 49040 -11675 49160 -11555
rect 49205 -11675 49325 -11555
rect 49380 -11675 49500 -11555
rect 49545 -11675 49665 -11555
rect 49710 -11675 49830 -11555
rect 49875 -11675 49995 -11555
rect 50050 -11675 50170 -11555
rect 50215 -11675 50335 -11555
rect 50380 -11675 50500 -11555
rect 50545 -11675 50665 -11555
rect 50720 -11675 50840 -11555
rect 50885 -11675 51005 -11555
rect 51050 -11675 51170 -11555
rect 51215 -11675 51335 -11555
rect 51390 -11675 51510 -11555
rect 51555 -11675 51675 -11555
rect 51720 -11675 51840 -11555
rect 51885 -11675 52005 -11555
rect 52060 -11675 52180 -11555
rect 52225 -11675 52345 -11555
rect 52390 -11675 52510 -11555
rect 52555 -11675 52675 -11555
rect 52730 -11675 52850 -11555
rect 52895 -11675 53015 -11555
rect 53060 -11675 53180 -11555
rect 53225 -11675 53345 -11555
rect 47865 -11840 47985 -11720
rect 48040 -11840 48160 -11720
rect 48205 -11840 48325 -11720
rect 48370 -11840 48490 -11720
rect 48535 -11840 48655 -11720
rect 48710 -11840 48830 -11720
rect 48875 -11840 48995 -11720
rect 49040 -11840 49160 -11720
rect 49205 -11840 49325 -11720
rect 49380 -11840 49500 -11720
rect 49545 -11840 49665 -11720
rect 49710 -11840 49830 -11720
rect 49875 -11840 49995 -11720
rect 50050 -11840 50170 -11720
rect 50215 -11840 50335 -11720
rect 50380 -11840 50500 -11720
rect 50545 -11840 50665 -11720
rect 50720 -11840 50840 -11720
rect 50885 -11840 51005 -11720
rect 51050 -11840 51170 -11720
rect 51215 -11840 51335 -11720
rect 51390 -11840 51510 -11720
rect 51555 -11840 51675 -11720
rect 51720 -11840 51840 -11720
rect 51885 -11840 52005 -11720
rect 52060 -11840 52180 -11720
rect 52225 -11840 52345 -11720
rect 52390 -11840 52510 -11720
rect 52555 -11840 52675 -11720
rect 52730 -11840 52850 -11720
rect 52895 -11840 53015 -11720
rect 53060 -11840 53180 -11720
rect 53225 -11840 53345 -11720
rect 47865 -12005 47985 -11885
rect 48040 -12005 48160 -11885
rect 48205 -12005 48325 -11885
rect 48370 -12005 48490 -11885
rect 48535 -12005 48655 -11885
rect 48710 -12005 48830 -11885
rect 48875 -12005 48995 -11885
rect 49040 -12005 49160 -11885
rect 49205 -12005 49325 -11885
rect 49380 -12005 49500 -11885
rect 49545 -12005 49665 -11885
rect 49710 -12005 49830 -11885
rect 49875 -12005 49995 -11885
rect 50050 -12005 50170 -11885
rect 50215 -12005 50335 -11885
rect 50380 -12005 50500 -11885
rect 50545 -12005 50665 -11885
rect 50720 -12005 50840 -11885
rect 50885 -12005 51005 -11885
rect 51050 -12005 51170 -11885
rect 51215 -12005 51335 -11885
rect 51390 -12005 51510 -11885
rect 51555 -12005 51675 -11885
rect 51720 -12005 51840 -11885
rect 51885 -12005 52005 -11885
rect 52060 -12005 52180 -11885
rect 52225 -12005 52345 -11885
rect 52390 -12005 52510 -11885
rect 52555 -12005 52675 -11885
rect 52730 -12005 52850 -11885
rect 52895 -12005 53015 -11885
rect 53060 -12005 53180 -11885
rect 53225 -12005 53345 -11885
rect 47865 -12180 47985 -12060
rect 48040 -12180 48160 -12060
rect 48205 -12180 48325 -12060
rect 48370 -12180 48490 -12060
rect 48535 -12180 48655 -12060
rect 48710 -12180 48830 -12060
rect 48875 -12180 48995 -12060
rect 49040 -12180 49160 -12060
rect 49205 -12180 49325 -12060
rect 49380 -12180 49500 -12060
rect 49545 -12180 49665 -12060
rect 49710 -12180 49830 -12060
rect 49875 -12180 49995 -12060
rect 50050 -12180 50170 -12060
rect 50215 -12180 50335 -12060
rect 50380 -12180 50500 -12060
rect 50545 -12180 50665 -12060
rect 50720 -12180 50840 -12060
rect 50885 -12180 51005 -12060
rect 51050 -12180 51170 -12060
rect 51215 -12180 51335 -12060
rect 51390 -12180 51510 -12060
rect 51555 -12180 51675 -12060
rect 51720 -12180 51840 -12060
rect 51885 -12180 52005 -12060
rect 52060 -12180 52180 -12060
rect 52225 -12180 52345 -12060
rect 52390 -12180 52510 -12060
rect 52555 -12180 52675 -12060
rect 52730 -12180 52850 -12060
rect 52895 -12180 53015 -12060
rect 53060 -12180 53180 -12060
rect 53225 -12180 53345 -12060
rect 47865 -12345 47985 -12225
rect 48040 -12345 48160 -12225
rect 48205 -12345 48325 -12225
rect 48370 -12345 48490 -12225
rect 48535 -12345 48655 -12225
rect 48710 -12345 48830 -12225
rect 48875 -12345 48995 -12225
rect 49040 -12345 49160 -12225
rect 49205 -12345 49325 -12225
rect 49380 -12345 49500 -12225
rect 49545 -12345 49665 -12225
rect 49710 -12345 49830 -12225
rect 49875 -12345 49995 -12225
rect 50050 -12345 50170 -12225
rect 50215 -12345 50335 -12225
rect 50380 -12345 50500 -12225
rect 50545 -12345 50665 -12225
rect 50720 -12345 50840 -12225
rect 50885 -12345 51005 -12225
rect 51050 -12345 51170 -12225
rect 51215 -12345 51335 -12225
rect 51390 -12345 51510 -12225
rect 51555 -12345 51675 -12225
rect 51720 -12345 51840 -12225
rect 51885 -12345 52005 -12225
rect 52060 -12345 52180 -12225
rect 52225 -12345 52345 -12225
rect 52390 -12345 52510 -12225
rect 52555 -12345 52675 -12225
rect 52730 -12345 52850 -12225
rect 52895 -12345 53015 -12225
rect 53060 -12345 53180 -12225
rect 53225 -12345 53345 -12225
rect 47865 -12510 47985 -12390
rect 48040 -12510 48160 -12390
rect 48205 -12510 48325 -12390
rect 48370 -12510 48490 -12390
rect 48535 -12510 48655 -12390
rect 48710 -12510 48830 -12390
rect 48875 -12510 48995 -12390
rect 49040 -12510 49160 -12390
rect 49205 -12510 49325 -12390
rect 49380 -12510 49500 -12390
rect 49545 -12510 49665 -12390
rect 49710 -12510 49830 -12390
rect 49875 -12510 49995 -12390
rect 50050 -12510 50170 -12390
rect 50215 -12510 50335 -12390
rect 50380 -12510 50500 -12390
rect 50545 -12510 50665 -12390
rect 50720 -12510 50840 -12390
rect 50885 -12510 51005 -12390
rect 51050 -12510 51170 -12390
rect 51215 -12510 51335 -12390
rect 51390 -12510 51510 -12390
rect 51555 -12510 51675 -12390
rect 51720 -12510 51840 -12390
rect 51885 -12510 52005 -12390
rect 52060 -12510 52180 -12390
rect 52225 -12510 52345 -12390
rect 52390 -12510 52510 -12390
rect 52555 -12510 52675 -12390
rect 52730 -12510 52850 -12390
rect 52895 -12510 53015 -12390
rect 53060 -12510 53180 -12390
rect 53225 -12510 53345 -12390
rect 47865 -12675 47985 -12555
rect 48040 -12675 48160 -12555
rect 48205 -12675 48325 -12555
rect 48370 -12675 48490 -12555
rect 48535 -12675 48655 -12555
rect 48710 -12675 48830 -12555
rect 48875 -12675 48995 -12555
rect 49040 -12675 49160 -12555
rect 49205 -12675 49325 -12555
rect 49380 -12675 49500 -12555
rect 49545 -12675 49665 -12555
rect 49710 -12675 49830 -12555
rect 49875 -12675 49995 -12555
rect 50050 -12675 50170 -12555
rect 50215 -12675 50335 -12555
rect 50380 -12675 50500 -12555
rect 50545 -12675 50665 -12555
rect 50720 -12675 50840 -12555
rect 50885 -12675 51005 -12555
rect 51050 -12675 51170 -12555
rect 51215 -12675 51335 -12555
rect 51390 -12675 51510 -12555
rect 51555 -12675 51675 -12555
rect 51720 -12675 51840 -12555
rect 51885 -12675 52005 -12555
rect 52060 -12675 52180 -12555
rect 52225 -12675 52345 -12555
rect 52390 -12675 52510 -12555
rect 52555 -12675 52675 -12555
rect 52730 -12675 52850 -12555
rect 52895 -12675 53015 -12555
rect 53060 -12675 53180 -12555
rect 53225 -12675 53345 -12555
rect 47865 -12850 47985 -12730
rect 48040 -12850 48160 -12730
rect 48205 -12850 48325 -12730
rect 48370 -12850 48490 -12730
rect 48535 -12850 48655 -12730
rect 48710 -12850 48830 -12730
rect 48875 -12850 48995 -12730
rect 49040 -12850 49160 -12730
rect 49205 -12850 49325 -12730
rect 49380 -12850 49500 -12730
rect 49545 -12850 49665 -12730
rect 49710 -12850 49830 -12730
rect 49875 -12850 49995 -12730
rect 50050 -12850 50170 -12730
rect 50215 -12850 50335 -12730
rect 50380 -12850 50500 -12730
rect 50545 -12850 50665 -12730
rect 50720 -12850 50840 -12730
rect 50885 -12850 51005 -12730
rect 51050 -12850 51170 -12730
rect 51215 -12850 51335 -12730
rect 51390 -12850 51510 -12730
rect 51555 -12850 51675 -12730
rect 51720 -12850 51840 -12730
rect 51885 -12850 52005 -12730
rect 52060 -12850 52180 -12730
rect 52225 -12850 52345 -12730
rect 52390 -12850 52510 -12730
rect 52555 -12850 52675 -12730
rect 52730 -12850 52850 -12730
rect 52895 -12850 53015 -12730
rect 53060 -12850 53180 -12730
rect 53225 -12850 53345 -12730
rect 47865 -13015 47985 -12895
rect 48040 -13015 48160 -12895
rect 48205 -13015 48325 -12895
rect 48370 -13015 48490 -12895
rect 48535 -13015 48655 -12895
rect 48710 -13015 48830 -12895
rect 48875 -13015 48995 -12895
rect 49040 -13015 49160 -12895
rect 49205 -13015 49325 -12895
rect 49380 -13015 49500 -12895
rect 49545 -13015 49665 -12895
rect 49710 -13015 49830 -12895
rect 49875 -13015 49995 -12895
rect 50050 -13015 50170 -12895
rect 50215 -13015 50335 -12895
rect 50380 -13015 50500 -12895
rect 50545 -13015 50665 -12895
rect 50720 -13015 50840 -12895
rect 50885 -13015 51005 -12895
rect 51050 -13015 51170 -12895
rect 51215 -13015 51335 -12895
rect 51390 -13015 51510 -12895
rect 51555 -13015 51675 -12895
rect 51720 -13015 51840 -12895
rect 51885 -13015 52005 -12895
rect 52060 -13015 52180 -12895
rect 52225 -13015 52345 -12895
rect 52390 -13015 52510 -12895
rect 52555 -13015 52675 -12895
rect 52730 -13015 52850 -12895
rect 52895 -13015 53015 -12895
rect 53060 -13015 53180 -12895
rect 53225 -13015 53345 -12895
rect 47865 -13180 47985 -13060
rect 48040 -13180 48160 -13060
rect 48205 -13180 48325 -13060
rect 48370 -13180 48490 -13060
rect 48535 -13180 48655 -13060
rect 48710 -13180 48830 -13060
rect 48875 -13180 48995 -13060
rect 49040 -13180 49160 -13060
rect 49205 -13180 49325 -13060
rect 49380 -13180 49500 -13060
rect 49545 -13180 49665 -13060
rect 49710 -13180 49830 -13060
rect 49875 -13180 49995 -13060
rect 50050 -13180 50170 -13060
rect 50215 -13180 50335 -13060
rect 50380 -13180 50500 -13060
rect 50545 -13180 50665 -13060
rect 50720 -13180 50840 -13060
rect 50885 -13180 51005 -13060
rect 51050 -13180 51170 -13060
rect 51215 -13180 51335 -13060
rect 51390 -13180 51510 -13060
rect 51555 -13180 51675 -13060
rect 51720 -13180 51840 -13060
rect 51885 -13180 52005 -13060
rect 52060 -13180 52180 -13060
rect 52225 -13180 52345 -13060
rect 52390 -13180 52510 -13060
rect 52555 -13180 52675 -13060
rect 52730 -13180 52850 -13060
rect 52895 -13180 53015 -13060
rect 53060 -13180 53180 -13060
rect 53225 -13180 53345 -13060
rect 47865 -13345 47985 -13225
rect 48040 -13345 48160 -13225
rect 48205 -13345 48325 -13225
rect 48370 -13345 48490 -13225
rect 48535 -13345 48655 -13225
rect 48710 -13345 48830 -13225
rect 48875 -13345 48995 -13225
rect 49040 -13345 49160 -13225
rect 49205 -13345 49325 -13225
rect 49380 -13345 49500 -13225
rect 49545 -13345 49665 -13225
rect 49710 -13345 49830 -13225
rect 49875 -13345 49995 -13225
rect 50050 -13345 50170 -13225
rect 50215 -13345 50335 -13225
rect 50380 -13345 50500 -13225
rect 50545 -13345 50665 -13225
rect 50720 -13345 50840 -13225
rect 50885 -13345 51005 -13225
rect 51050 -13345 51170 -13225
rect 51215 -13345 51335 -13225
rect 51390 -13345 51510 -13225
rect 51555 -13345 51675 -13225
rect 51720 -13345 51840 -13225
rect 51885 -13345 52005 -13225
rect 52060 -13345 52180 -13225
rect 52225 -13345 52345 -13225
rect 52390 -13345 52510 -13225
rect 52555 -13345 52675 -13225
rect 52730 -13345 52850 -13225
rect 52895 -13345 53015 -13225
rect 53060 -13345 53180 -13225
rect 53225 -13345 53345 -13225
rect 47865 -13520 47985 -13400
rect 48040 -13520 48160 -13400
rect 48205 -13520 48325 -13400
rect 48370 -13520 48490 -13400
rect 48535 -13520 48655 -13400
rect 48710 -13520 48830 -13400
rect 48875 -13520 48995 -13400
rect 49040 -13520 49160 -13400
rect 49205 -13520 49325 -13400
rect 49380 -13520 49500 -13400
rect 49545 -13520 49665 -13400
rect 49710 -13520 49830 -13400
rect 49875 -13520 49995 -13400
rect 50050 -13520 50170 -13400
rect 50215 -13520 50335 -13400
rect 50380 -13520 50500 -13400
rect 50545 -13520 50665 -13400
rect 50720 -13520 50840 -13400
rect 50885 -13520 51005 -13400
rect 51050 -13520 51170 -13400
rect 51215 -13520 51335 -13400
rect 51390 -13520 51510 -13400
rect 51555 -13520 51675 -13400
rect 51720 -13520 51840 -13400
rect 51885 -13520 52005 -13400
rect 52060 -13520 52180 -13400
rect 52225 -13520 52345 -13400
rect 52390 -13520 52510 -13400
rect 52555 -13520 52675 -13400
rect 52730 -13520 52850 -13400
rect 52895 -13520 53015 -13400
rect 53060 -13520 53180 -13400
rect 53225 -13520 53345 -13400
rect 47865 -13685 47985 -13565
rect 48040 -13685 48160 -13565
rect 48205 -13685 48325 -13565
rect 48370 -13685 48490 -13565
rect 48535 -13685 48655 -13565
rect 48710 -13685 48830 -13565
rect 48875 -13685 48995 -13565
rect 49040 -13685 49160 -13565
rect 49205 -13685 49325 -13565
rect 49380 -13685 49500 -13565
rect 49545 -13685 49665 -13565
rect 49710 -13685 49830 -13565
rect 49875 -13685 49995 -13565
rect 50050 -13685 50170 -13565
rect 50215 -13685 50335 -13565
rect 50380 -13685 50500 -13565
rect 50545 -13685 50665 -13565
rect 50720 -13685 50840 -13565
rect 50885 -13685 51005 -13565
rect 51050 -13685 51170 -13565
rect 51215 -13685 51335 -13565
rect 51390 -13685 51510 -13565
rect 51555 -13685 51675 -13565
rect 51720 -13685 51840 -13565
rect 51885 -13685 52005 -13565
rect 52060 -13685 52180 -13565
rect 52225 -13685 52345 -13565
rect 52390 -13685 52510 -13565
rect 52555 -13685 52675 -13565
rect 52730 -13685 52850 -13565
rect 52895 -13685 53015 -13565
rect 53060 -13685 53180 -13565
rect 53225 -13685 53345 -13565
rect 47865 -13850 47985 -13730
rect 48040 -13850 48160 -13730
rect 48205 -13850 48325 -13730
rect 48370 -13850 48490 -13730
rect 48535 -13850 48655 -13730
rect 48710 -13850 48830 -13730
rect 48875 -13850 48995 -13730
rect 49040 -13850 49160 -13730
rect 49205 -13850 49325 -13730
rect 49380 -13850 49500 -13730
rect 49545 -13850 49665 -13730
rect 49710 -13850 49830 -13730
rect 49875 -13850 49995 -13730
rect 50050 -13850 50170 -13730
rect 50215 -13850 50335 -13730
rect 50380 -13850 50500 -13730
rect 50545 -13850 50665 -13730
rect 50720 -13850 50840 -13730
rect 50885 -13850 51005 -13730
rect 51050 -13850 51170 -13730
rect 51215 -13850 51335 -13730
rect 51390 -13850 51510 -13730
rect 51555 -13850 51675 -13730
rect 51720 -13850 51840 -13730
rect 51885 -13850 52005 -13730
rect 52060 -13850 52180 -13730
rect 52225 -13850 52345 -13730
rect 52390 -13850 52510 -13730
rect 52555 -13850 52675 -13730
rect 52730 -13850 52850 -13730
rect 52895 -13850 53015 -13730
rect 53060 -13850 53180 -13730
rect 53225 -13850 53345 -13730
rect 47865 -14015 47985 -13895
rect 48040 -14015 48160 -13895
rect 48205 -14015 48325 -13895
rect 48370 -14015 48490 -13895
rect 48535 -14015 48655 -13895
rect 48710 -14015 48830 -13895
rect 48875 -14015 48995 -13895
rect 49040 -14015 49160 -13895
rect 49205 -14015 49325 -13895
rect 49380 -14015 49500 -13895
rect 49545 -14015 49665 -13895
rect 49710 -14015 49830 -13895
rect 49875 -14015 49995 -13895
rect 50050 -14015 50170 -13895
rect 50215 -14015 50335 -13895
rect 50380 -14015 50500 -13895
rect 50545 -14015 50665 -13895
rect 50720 -14015 50840 -13895
rect 50885 -14015 51005 -13895
rect 51050 -14015 51170 -13895
rect 51215 -14015 51335 -13895
rect 51390 -14015 51510 -13895
rect 51555 -14015 51675 -13895
rect 51720 -14015 51840 -13895
rect 51885 -14015 52005 -13895
rect 52060 -14015 52180 -13895
rect 52225 -14015 52345 -13895
rect 52390 -14015 52510 -13895
rect 52555 -14015 52675 -13895
rect 52730 -14015 52850 -13895
rect 52895 -14015 53015 -13895
rect 53060 -14015 53180 -13895
rect 53225 -14015 53345 -13895
rect 47865 -14190 47985 -14070
rect 48040 -14190 48160 -14070
rect 48205 -14190 48325 -14070
rect 48370 -14190 48490 -14070
rect 48535 -14190 48655 -14070
rect 48710 -14190 48830 -14070
rect 48875 -14190 48995 -14070
rect 49040 -14190 49160 -14070
rect 49205 -14190 49325 -14070
rect 49380 -14190 49500 -14070
rect 49545 -14190 49665 -14070
rect 49710 -14190 49830 -14070
rect 49875 -14190 49995 -14070
rect 50050 -14190 50170 -14070
rect 50215 -14190 50335 -14070
rect 50380 -14190 50500 -14070
rect 50545 -14190 50665 -14070
rect 50720 -14190 50840 -14070
rect 50885 -14190 51005 -14070
rect 51050 -14190 51170 -14070
rect 51215 -14190 51335 -14070
rect 51390 -14190 51510 -14070
rect 51555 -14190 51675 -14070
rect 51720 -14190 51840 -14070
rect 51885 -14190 52005 -14070
rect 52060 -14190 52180 -14070
rect 52225 -14190 52345 -14070
rect 52390 -14190 52510 -14070
rect 52555 -14190 52675 -14070
rect 52730 -14190 52850 -14070
rect 52895 -14190 53015 -14070
rect 53060 -14190 53180 -14070
rect 53225 -14190 53345 -14070
rect 47865 -14355 47985 -14235
rect 48040 -14355 48160 -14235
rect 48205 -14355 48325 -14235
rect 48370 -14355 48490 -14235
rect 48535 -14355 48655 -14235
rect 48710 -14355 48830 -14235
rect 48875 -14355 48995 -14235
rect 49040 -14355 49160 -14235
rect 49205 -14355 49325 -14235
rect 49380 -14355 49500 -14235
rect 49545 -14355 49665 -14235
rect 49710 -14355 49830 -14235
rect 49875 -14355 49995 -14235
rect 50050 -14355 50170 -14235
rect 50215 -14355 50335 -14235
rect 50380 -14355 50500 -14235
rect 50545 -14355 50665 -14235
rect 50720 -14355 50840 -14235
rect 50885 -14355 51005 -14235
rect 51050 -14355 51170 -14235
rect 51215 -14355 51335 -14235
rect 51390 -14355 51510 -14235
rect 51555 -14355 51675 -14235
rect 51720 -14355 51840 -14235
rect 51885 -14355 52005 -14235
rect 52060 -14355 52180 -14235
rect 52225 -14355 52345 -14235
rect 52390 -14355 52510 -14235
rect 52555 -14355 52675 -14235
rect 52730 -14355 52850 -14235
rect 52895 -14355 53015 -14235
rect 53060 -14355 53180 -14235
rect 53225 -14355 53345 -14235
rect 47865 -14520 47985 -14400
rect 48040 -14520 48160 -14400
rect 48205 -14520 48325 -14400
rect 48370 -14520 48490 -14400
rect 48535 -14520 48655 -14400
rect 48710 -14520 48830 -14400
rect 48875 -14520 48995 -14400
rect 49040 -14520 49160 -14400
rect 49205 -14520 49325 -14400
rect 49380 -14520 49500 -14400
rect 49545 -14520 49665 -14400
rect 49710 -14520 49830 -14400
rect 49875 -14520 49995 -14400
rect 50050 -14520 50170 -14400
rect 50215 -14520 50335 -14400
rect 50380 -14520 50500 -14400
rect 50545 -14520 50665 -14400
rect 50720 -14520 50840 -14400
rect 50885 -14520 51005 -14400
rect 51050 -14520 51170 -14400
rect 51215 -14520 51335 -14400
rect 51390 -14520 51510 -14400
rect 51555 -14520 51675 -14400
rect 51720 -14520 51840 -14400
rect 51885 -14520 52005 -14400
rect 52060 -14520 52180 -14400
rect 52225 -14520 52345 -14400
rect 52390 -14520 52510 -14400
rect 52555 -14520 52675 -14400
rect 52730 -14520 52850 -14400
rect 52895 -14520 53015 -14400
rect 53060 -14520 53180 -14400
rect 53225 -14520 53345 -14400
rect 47865 -14685 47985 -14565
rect 48040 -14685 48160 -14565
rect 48205 -14685 48325 -14565
rect 48370 -14685 48490 -14565
rect 48535 -14685 48655 -14565
rect 48710 -14685 48830 -14565
rect 48875 -14685 48995 -14565
rect 49040 -14685 49160 -14565
rect 49205 -14685 49325 -14565
rect 49380 -14685 49500 -14565
rect 49545 -14685 49665 -14565
rect 49710 -14685 49830 -14565
rect 49875 -14685 49995 -14565
rect 50050 -14685 50170 -14565
rect 50215 -14685 50335 -14565
rect 50380 -14685 50500 -14565
rect 50545 -14685 50665 -14565
rect 50720 -14685 50840 -14565
rect 50885 -14685 51005 -14565
rect 51050 -14685 51170 -14565
rect 51215 -14685 51335 -14565
rect 51390 -14685 51510 -14565
rect 51555 -14685 51675 -14565
rect 51720 -14685 51840 -14565
rect 51885 -14685 52005 -14565
rect 52060 -14685 52180 -14565
rect 52225 -14685 52345 -14565
rect 52390 -14685 52510 -14565
rect 52555 -14685 52675 -14565
rect 52730 -14685 52850 -14565
rect 52895 -14685 53015 -14565
rect 53060 -14685 53180 -14565
rect 53225 -14685 53345 -14565
rect 47865 -14860 47985 -14740
rect 48040 -14860 48160 -14740
rect 48205 -14860 48325 -14740
rect 48370 -14860 48490 -14740
rect 48535 -14860 48655 -14740
rect 48710 -14860 48830 -14740
rect 48875 -14860 48995 -14740
rect 49040 -14860 49160 -14740
rect 49205 -14860 49325 -14740
rect 49380 -14860 49500 -14740
rect 49545 -14860 49665 -14740
rect 49710 -14860 49830 -14740
rect 49875 -14860 49995 -14740
rect 50050 -14860 50170 -14740
rect 50215 -14860 50335 -14740
rect 50380 -14860 50500 -14740
rect 50545 -14860 50665 -14740
rect 50720 -14860 50840 -14740
rect 50885 -14860 51005 -14740
rect 51050 -14860 51170 -14740
rect 51215 -14860 51335 -14740
rect 51390 -14860 51510 -14740
rect 51555 -14860 51675 -14740
rect 51720 -14860 51840 -14740
rect 51885 -14860 52005 -14740
rect 52060 -14860 52180 -14740
rect 52225 -14860 52345 -14740
rect 52390 -14860 52510 -14740
rect 52555 -14860 52675 -14740
rect 52730 -14860 52850 -14740
rect 52895 -14860 53015 -14740
rect 53060 -14860 53180 -14740
rect 53225 -14860 53345 -14740
rect 47865 -15025 47985 -14905
rect 48040 -15025 48160 -14905
rect 48205 -15025 48325 -14905
rect 48370 -15025 48490 -14905
rect 48535 -15025 48655 -14905
rect 48710 -15025 48830 -14905
rect 48875 -15025 48995 -14905
rect 49040 -15025 49160 -14905
rect 49205 -15025 49325 -14905
rect 49380 -15025 49500 -14905
rect 49545 -15025 49665 -14905
rect 49710 -15025 49830 -14905
rect 49875 -15025 49995 -14905
rect 50050 -15025 50170 -14905
rect 50215 -15025 50335 -14905
rect 50380 -15025 50500 -14905
rect 50545 -15025 50665 -14905
rect 50720 -15025 50840 -14905
rect 50885 -15025 51005 -14905
rect 51050 -15025 51170 -14905
rect 51215 -15025 51335 -14905
rect 51390 -15025 51510 -14905
rect 51555 -15025 51675 -14905
rect 51720 -15025 51840 -14905
rect 51885 -15025 52005 -14905
rect 52060 -15025 52180 -14905
rect 52225 -15025 52345 -14905
rect 52390 -15025 52510 -14905
rect 52555 -15025 52675 -14905
rect 52730 -15025 52850 -14905
rect 52895 -15025 53015 -14905
rect 53060 -15025 53180 -14905
rect 53225 -15025 53345 -14905
rect 47865 -15190 47985 -15070
rect 48040 -15190 48160 -15070
rect 48205 -15190 48325 -15070
rect 48370 -15190 48490 -15070
rect 48535 -15190 48655 -15070
rect 48710 -15190 48830 -15070
rect 48875 -15190 48995 -15070
rect 49040 -15190 49160 -15070
rect 49205 -15190 49325 -15070
rect 49380 -15190 49500 -15070
rect 49545 -15190 49665 -15070
rect 49710 -15190 49830 -15070
rect 49875 -15190 49995 -15070
rect 50050 -15190 50170 -15070
rect 50215 -15190 50335 -15070
rect 50380 -15190 50500 -15070
rect 50545 -15190 50665 -15070
rect 50720 -15190 50840 -15070
rect 50885 -15190 51005 -15070
rect 51050 -15190 51170 -15070
rect 51215 -15190 51335 -15070
rect 51390 -15190 51510 -15070
rect 51555 -15190 51675 -15070
rect 51720 -15190 51840 -15070
rect 51885 -15190 52005 -15070
rect 52060 -15190 52180 -15070
rect 52225 -15190 52345 -15070
rect 52390 -15190 52510 -15070
rect 52555 -15190 52675 -15070
rect 52730 -15190 52850 -15070
rect 52895 -15190 53015 -15070
rect 53060 -15190 53180 -15070
rect 53225 -15190 53345 -15070
rect 47865 -15355 47985 -15235
rect 48040 -15355 48160 -15235
rect 48205 -15355 48325 -15235
rect 48370 -15355 48490 -15235
rect 48535 -15355 48655 -15235
rect 48710 -15355 48830 -15235
rect 48875 -15355 48995 -15235
rect 49040 -15355 49160 -15235
rect 49205 -15355 49325 -15235
rect 49380 -15355 49500 -15235
rect 49545 -15355 49665 -15235
rect 49710 -15355 49830 -15235
rect 49875 -15355 49995 -15235
rect 50050 -15355 50170 -15235
rect 50215 -15355 50335 -15235
rect 50380 -15355 50500 -15235
rect 50545 -15355 50665 -15235
rect 50720 -15355 50840 -15235
rect 50885 -15355 51005 -15235
rect 51050 -15355 51170 -15235
rect 51215 -15355 51335 -15235
rect 51390 -15355 51510 -15235
rect 51555 -15355 51675 -15235
rect 51720 -15355 51840 -15235
rect 51885 -15355 52005 -15235
rect 52060 -15355 52180 -15235
rect 52225 -15355 52345 -15235
rect 52390 -15355 52510 -15235
rect 52555 -15355 52675 -15235
rect 52730 -15355 52850 -15235
rect 52895 -15355 53015 -15235
rect 53060 -15355 53180 -15235
rect 53225 -15355 53345 -15235
rect 47865 -15530 47985 -15410
rect 48040 -15530 48160 -15410
rect 48205 -15530 48325 -15410
rect 48370 -15530 48490 -15410
rect 48535 -15530 48655 -15410
rect 48710 -15530 48830 -15410
rect 48875 -15530 48995 -15410
rect 49040 -15530 49160 -15410
rect 49205 -15530 49325 -15410
rect 49380 -15530 49500 -15410
rect 49545 -15530 49665 -15410
rect 49710 -15530 49830 -15410
rect 49875 -15530 49995 -15410
rect 50050 -15530 50170 -15410
rect 50215 -15530 50335 -15410
rect 50380 -15530 50500 -15410
rect 50545 -15530 50665 -15410
rect 50720 -15530 50840 -15410
rect 50885 -15530 51005 -15410
rect 51050 -15530 51170 -15410
rect 51215 -15530 51335 -15410
rect 51390 -15530 51510 -15410
rect 51555 -15530 51675 -15410
rect 51720 -15530 51840 -15410
rect 51885 -15530 52005 -15410
rect 52060 -15530 52180 -15410
rect 52225 -15530 52345 -15410
rect 52390 -15530 52510 -15410
rect 52555 -15530 52675 -15410
rect 52730 -15530 52850 -15410
rect 52895 -15530 53015 -15410
rect 53060 -15530 53180 -15410
rect 53225 -15530 53345 -15410
<< metal4 >>
rect 30770 7200 53370 7225
rect 30770 7080 30795 7200
rect 30915 7080 30960 7200
rect 31080 7080 31125 7200
rect 31245 7080 31290 7200
rect 31410 7080 31465 7200
rect 31585 7080 31630 7200
rect 31750 7080 31795 7200
rect 31915 7080 31960 7200
rect 32080 7080 32135 7200
rect 32255 7080 32300 7200
rect 32420 7080 32465 7200
rect 32585 7080 32630 7200
rect 32750 7080 32805 7200
rect 32925 7080 32970 7200
rect 33090 7080 33135 7200
rect 33255 7080 33300 7200
rect 33420 7080 33475 7200
rect 33595 7080 33640 7200
rect 33760 7080 33805 7200
rect 33925 7080 33970 7200
rect 34090 7080 34145 7200
rect 34265 7080 34310 7200
rect 34430 7080 34475 7200
rect 34595 7080 34640 7200
rect 34760 7080 34815 7200
rect 34935 7080 34980 7200
rect 35100 7080 35145 7200
rect 35265 7080 35310 7200
rect 35430 7080 35485 7200
rect 35605 7080 35650 7200
rect 35770 7080 35815 7200
rect 35935 7080 35980 7200
rect 36100 7080 36155 7200
rect 36275 7080 36485 7200
rect 36605 7080 36650 7200
rect 36770 7080 36815 7200
rect 36935 7080 36980 7200
rect 37100 7080 37155 7200
rect 37275 7080 37320 7200
rect 37440 7080 37485 7200
rect 37605 7080 37650 7200
rect 37770 7080 37825 7200
rect 37945 7080 37990 7200
rect 38110 7080 38155 7200
rect 38275 7080 38320 7200
rect 38440 7080 38495 7200
rect 38615 7080 38660 7200
rect 38780 7080 38825 7200
rect 38945 7080 38990 7200
rect 39110 7080 39165 7200
rect 39285 7080 39330 7200
rect 39450 7080 39495 7200
rect 39615 7080 39660 7200
rect 39780 7080 39835 7200
rect 39955 7080 40000 7200
rect 40120 7080 40165 7200
rect 40285 7080 40330 7200
rect 40450 7080 40505 7200
rect 40625 7080 40670 7200
rect 40790 7080 40835 7200
rect 40955 7080 41000 7200
rect 41120 7080 41175 7200
rect 41295 7080 41340 7200
rect 41460 7080 41505 7200
rect 41625 7080 41670 7200
rect 41790 7080 41845 7200
rect 41965 7080 42175 7200
rect 42295 7080 42340 7200
rect 42460 7080 42505 7200
rect 42625 7080 42670 7200
rect 42790 7080 42845 7200
rect 42965 7080 43010 7200
rect 43130 7080 43175 7200
rect 43295 7080 43340 7200
rect 43460 7080 43515 7200
rect 43635 7080 43680 7200
rect 43800 7080 43845 7200
rect 43965 7080 44010 7200
rect 44130 7080 44185 7200
rect 44305 7080 44350 7200
rect 44470 7080 44515 7200
rect 44635 7080 44680 7200
rect 44800 7080 44855 7200
rect 44975 7080 45020 7200
rect 45140 7080 45185 7200
rect 45305 7080 45350 7200
rect 45470 7080 45525 7200
rect 45645 7080 45690 7200
rect 45810 7080 45855 7200
rect 45975 7080 46020 7200
rect 46140 7080 46195 7200
rect 46315 7080 46360 7200
rect 46480 7080 46525 7200
rect 46645 7080 46690 7200
rect 46810 7080 46865 7200
rect 46985 7080 47030 7200
rect 47150 7080 47195 7200
rect 47315 7080 47360 7200
rect 47480 7080 47535 7200
rect 47655 7080 47865 7200
rect 47985 7080 48030 7200
rect 48150 7080 48195 7200
rect 48315 7080 48360 7200
rect 48480 7080 48535 7200
rect 48655 7080 48700 7200
rect 48820 7080 48865 7200
rect 48985 7080 49030 7200
rect 49150 7080 49205 7200
rect 49325 7080 49370 7200
rect 49490 7080 49535 7200
rect 49655 7080 49700 7200
rect 49820 7080 49875 7200
rect 49995 7080 50040 7200
rect 50160 7080 50205 7200
rect 50325 7080 50370 7200
rect 50490 7080 50545 7200
rect 50665 7080 50710 7200
rect 50830 7080 50875 7200
rect 50995 7080 51040 7200
rect 51160 7080 51215 7200
rect 51335 7080 51380 7200
rect 51500 7080 51545 7200
rect 51665 7080 51710 7200
rect 51830 7080 51885 7200
rect 52005 7080 52050 7200
rect 52170 7080 52215 7200
rect 52335 7080 52380 7200
rect 52500 7080 52555 7200
rect 52675 7080 52720 7200
rect 52840 7080 52885 7200
rect 53005 7080 53050 7200
rect 53170 7080 53225 7200
rect 53345 7080 53370 7200
rect 30770 7025 53370 7080
rect 30770 6905 30795 7025
rect 30915 6905 30960 7025
rect 31080 6905 31125 7025
rect 31245 6905 31290 7025
rect 31410 6905 31465 7025
rect 31585 6905 31630 7025
rect 31750 6905 31795 7025
rect 31915 6905 31960 7025
rect 32080 6905 32135 7025
rect 32255 6905 32300 7025
rect 32420 6905 32465 7025
rect 32585 6905 32630 7025
rect 32750 6905 32805 7025
rect 32925 6905 32970 7025
rect 33090 6905 33135 7025
rect 33255 6905 33300 7025
rect 33420 6905 33475 7025
rect 33595 6905 33640 7025
rect 33760 6905 33805 7025
rect 33925 6905 33970 7025
rect 34090 6905 34145 7025
rect 34265 6905 34310 7025
rect 34430 6905 34475 7025
rect 34595 6905 34640 7025
rect 34760 6905 34815 7025
rect 34935 6905 34980 7025
rect 35100 6905 35145 7025
rect 35265 6905 35310 7025
rect 35430 6905 35485 7025
rect 35605 6905 35650 7025
rect 35770 6905 35815 7025
rect 35935 6905 35980 7025
rect 36100 6905 36155 7025
rect 36275 6905 36485 7025
rect 36605 6905 36650 7025
rect 36770 6905 36815 7025
rect 36935 6905 36980 7025
rect 37100 6905 37155 7025
rect 37275 6905 37320 7025
rect 37440 6905 37485 7025
rect 37605 6905 37650 7025
rect 37770 6905 37825 7025
rect 37945 6905 37990 7025
rect 38110 6905 38155 7025
rect 38275 6905 38320 7025
rect 38440 6905 38495 7025
rect 38615 6905 38660 7025
rect 38780 6905 38825 7025
rect 38945 6905 38990 7025
rect 39110 6905 39165 7025
rect 39285 6905 39330 7025
rect 39450 6905 39495 7025
rect 39615 6905 39660 7025
rect 39780 6905 39835 7025
rect 39955 6905 40000 7025
rect 40120 6905 40165 7025
rect 40285 6905 40330 7025
rect 40450 6905 40505 7025
rect 40625 6905 40670 7025
rect 40790 6905 40835 7025
rect 40955 6905 41000 7025
rect 41120 6905 41175 7025
rect 41295 6905 41340 7025
rect 41460 6905 41505 7025
rect 41625 6905 41670 7025
rect 41790 6905 41845 7025
rect 41965 6905 42175 7025
rect 42295 6905 42340 7025
rect 42460 6905 42505 7025
rect 42625 6905 42670 7025
rect 42790 6905 42845 7025
rect 42965 6905 43010 7025
rect 43130 6905 43175 7025
rect 43295 6905 43340 7025
rect 43460 6905 43515 7025
rect 43635 6905 43680 7025
rect 43800 6905 43845 7025
rect 43965 6905 44010 7025
rect 44130 6905 44185 7025
rect 44305 6905 44350 7025
rect 44470 6905 44515 7025
rect 44635 6905 44680 7025
rect 44800 6905 44855 7025
rect 44975 6905 45020 7025
rect 45140 6905 45185 7025
rect 45305 6905 45350 7025
rect 45470 6905 45525 7025
rect 45645 6905 45690 7025
rect 45810 6905 45855 7025
rect 45975 6905 46020 7025
rect 46140 6905 46195 7025
rect 46315 6905 46360 7025
rect 46480 6905 46525 7025
rect 46645 6905 46690 7025
rect 46810 6905 46865 7025
rect 46985 6905 47030 7025
rect 47150 6905 47195 7025
rect 47315 6905 47360 7025
rect 47480 6905 47535 7025
rect 47655 6905 47865 7025
rect 47985 6905 48030 7025
rect 48150 6905 48195 7025
rect 48315 6905 48360 7025
rect 48480 6905 48535 7025
rect 48655 6905 48700 7025
rect 48820 6905 48865 7025
rect 48985 6905 49030 7025
rect 49150 6905 49205 7025
rect 49325 6905 49370 7025
rect 49490 6905 49535 7025
rect 49655 6905 49700 7025
rect 49820 6905 49875 7025
rect 49995 6905 50040 7025
rect 50160 6905 50205 7025
rect 50325 6905 50370 7025
rect 50490 6905 50545 7025
rect 50665 6905 50710 7025
rect 50830 6905 50875 7025
rect 50995 6905 51040 7025
rect 51160 6905 51215 7025
rect 51335 6905 51380 7025
rect 51500 6905 51545 7025
rect 51665 6905 51710 7025
rect 51830 6905 51885 7025
rect 52005 6905 52050 7025
rect 52170 6905 52215 7025
rect 52335 6905 52380 7025
rect 52500 6905 52555 7025
rect 52675 6905 52720 7025
rect 52840 6905 52885 7025
rect 53005 6905 53050 7025
rect 53170 6905 53225 7025
rect 53345 6905 53370 7025
rect 30770 6860 53370 6905
rect 30770 6740 30795 6860
rect 30915 6740 30960 6860
rect 31080 6740 31125 6860
rect 31245 6740 31290 6860
rect 31410 6740 31465 6860
rect 31585 6740 31630 6860
rect 31750 6740 31795 6860
rect 31915 6740 31960 6860
rect 32080 6740 32135 6860
rect 32255 6740 32300 6860
rect 32420 6740 32465 6860
rect 32585 6740 32630 6860
rect 32750 6740 32805 6860
rect 32925 6740 32970 6860
rect 33090 6740 33135 6860
rect 33255 6740 33300 6860
rect 33420 6740 33475 6860
rect 33595 6740 33640 6860
rect 33760 6740 33805 6860
rect 33925 6740 33970 6860
rect 34090 6740 34145 6860
rect 34265 6740 34310 6860
rect 34430 6740 34475 6860
rect 34595 6740 34640 6860
rect 34760 6740 34815 6860
rect 34935 6740 34980 6860
rect 35100 6740 35145 6860
rect 35265 6740 35310 6860
rect 35430 6740 35485 6860
rect 35605 6740 35650 6860
rect 35770 6740 35815 6860
rect 35935 6740 35980 6860
rect 36100 6740 36155 6860
rect 36275 6740 36485 6860
rect 36605 6740 36650 6860
rect 36770 6740 36815 6860
rect 36935 6740 36980 6860
rect 37100 6740 37155 6860
rect 37275 6740 37320 6860
rect 37440 6740 37485 6860
rect 37605 6740 37650 6860
rect 37770 6740 37825 6860
rect 37945 6740 37990 6860
rect 38110 6740 38155 6860
rect 38275 6740 38320 6860
rect 38440 6740 38495 6860
rect 38615 6740 38660 6860
rect 38780 6740 38825 6860
rect 38945 6740 38990 6860
rect 39110 6740 39165 6860
rect 39285 6740 39330 6860
rect 39450 6740 39495 6860
rect 39615 6740 39660 6860
rect 39780 6740 39835 6860
rect 39955 6740 40000 6860
rect 40120 6740 40165 6860
rect 40285 6740 40330 6860
rect 40450 6740 40505 6860
rect 40625 6740 40670 6860
rect 40790 6740 40835 6860
rect 40955 6740 41000 6860
rect 41120 6740 41175 6860
rect 41295 6740 41340 6860
rect 41460 6740 41505 6860
rect 41625 6740 41670 6860
rect 41790 6740 41845 6860
rect 41965 6740 42175 6860
rect 42295 6740 42340 6860
rect 42460 6740 42505 6860
rect 42625 6740 42670 6860
rect 42790 6740 42845 6860
rect 42965 6740 43010 6860
rect 43130 6740 43175 6860
rect 43295 6740 43340 6860
rect 43460 6740 43515 6860
rect 43635 6740 43680 6860
rect 43800 6740 43845 6860
rect 43965 6740 44010 6860
rect 44130 6740 44185 6860
rect 44305 6740 44350 6860
rect 44470 6740 44515 6860
rect 44635 6740 44680 6860
rect 44800 6740 44855 6860
rect 44975 6740 45020 6860
rect 45140 6740 45185 6860
rect 45305 6740 45350 6860
rect 45470 6740 45525 6860
rect 45645 6740 45690 6860
rect 45810 6740 45855 6860
rect 45975 6740 46020 6860
rect 46140 6740 46195 6860
rect 46315 6740 46360 6860
rect 46480 6740 46525 6860
rect 46645 6740 46690 6860
rect 46810 6740 46865 6860
rect 46985 6740 47030 6860
rect 47150 6740 47195 6860
rect 47315 6740 47360 6860
rect 47480 6740 47535 6860
rect 47655 6740 47865 6860
rect 47985 6740 48030 6860
rect 48150 6740 48195 6860
rect 48315 6740 48360 6860
rect 48480 6740 48535 6860
rect 48655 6740 48700 6860
rect 48820 6740 48865 6860
rect 48985 6740 49030 6860
rect 49150 6740 49205 6860
rect 49325 6740 49370 6860
rect 49490 6740 49535 6860
rect 49655 6740 49700 6860
rect 49820 6740 49875 6860
rect 49995 6740 50040 6860
rect 50160 6740 50205 6860
rect 50325 6740 50370 6860
rect 50490 6740 50545 6860
rect 50665 6740 50710 6860
rect 50830 6740 50875 6860
rect 50995 6740 51040 6860
rect 51160 6740 51215 6860
rect 51335 6740 51380 6860
rect 51500 6740 51545 6860
rect 51665 6740 51710 6860
rect 51830 6740 51885 6860
rect 52005 6740 52050 6860
rect 52170 6740 52215 6860
rect 52335 6740 52380 6860
rect 52500 6740 52555 6860
rect 52675 6740 52720 6860
rect 52840 6740 52885 6860
rect 53005 6740 53050 6860
rect 53170 6740 53225 6860
rect 53345 6740 53370 6860
rect 30770 6695 53370 6740
rect 30770 6575 30795 6695
rect 30915 6575 30960 6695
rect 31080 6575 31125 6695
rect 31245 6575 31290 6695
rect 31410 6575 31465 6695
rect 31585 6575 31630 6695
rect 31750 6575 31795 6695
rect 31915 6575 31960 6695
rect 32080 6575 32135 6695
rect 32255 6575 32300 6695
rect 32420 6575 32465 6695
rect 32585 6575 32630 6695
rect 32750 6575 32805 6695
rect 32925 6575 32970 6695
rect 33090 6575 33135 6695
rect 33255 6575 33300 6695
rect 33420 6575 33475 6695
rect 33595 6575 33640 6695
rect 33760 6575 33805 6695
rect 33925 6575 33970 6695
rect 34090 6575 34145 6695
rect 34265 6575 34310 6695
rect 34430 6575 34475 6695
rect 34595 6575 34640 6695
rect 34760 6575 34815 6695
rect 34935 6575 34980 6695
rect 35100 6575 35145 6695
rect 35265 6575 35310 6695
rect 35430 6575 35485 6695
rect 35605 6575 35650 6695
rect 35770 6575 35815 6695
rect 35935 6575 35980 6695
rect 36100 6575 36155 6695
rect 36275 6575 36485 6695
rect 36605 6575 36650 6695
rect 36770 6575 36815 6695
rect 36935 6575 36980 6695
rect 37100 6575 37155 6695
rect 37275 6575 37320 6695
rect 37440 6575 37485 6695
rect 37605 6575 37650 6695
rect 37770 6575 37825 6695
rect 37945 6575 37990 6695
rect 38110 6575 38155 6695
rect 38275 6575 38320 6695
rect 38440 6575 38495 6695
rect 38615 6575 38660 6695
rect 38780 6575 38825 6695
rect 38945 6575 38990 6695
rect 39110 6575 39165 6695
rect 39285 6575 39330 6695
rect 39450 6575 39495 6695
rect 39615 6575 39660 6695
rect 39780 6575 39835 6695
rect 39955 6575 40000 6695
rect 40120 6575 40165 6695
rect 40285 6575 40330 6695
rect 40450 6575 40505 6695
rect 40625 6575 40670 6695
rect 40790 6575 40835 6695
rect 40955 6575 41000 6695
rect 41120 6575 41175 6695
rect 41295 6575 41340 6695
rect 41460 6575 41505 6695
rect 41625 6575 41670 6695
rect 41790 6575 41845 6695
rect 41965 6575 42175 6695
rect 42295 6575 42340 6695
rect 42460 6575 42505 6695
rect 42625 6575 42670 6695
rect 42790 6575 42845 6695
rect 42965 6575 43010 6695
rect 43130 6575 43175 6695
rect 43295 6575 43340 6695
rect 43460 6575 43515 6695
rect 43635 6575 43680 6695
rect 43800 6575 43845 6695
rect 43965 6575 44010 6695
rect 44130 6575 44185 6695
rect 44305 6575 44350 6695
rect 44470 6575 44515 6695
rect 44635 6575 44680 6695
rect 44800 6575 44855 6695
rect 44975 6575 45020 6695
rect 45140 6575 45185 6695
rect 45305 6575 45350 6695
rect 45470 6575 45525 6695
rect 45645 6575 45690 6695
rect 45810 6575 45855 6695
rect 45975 6575 46020 6695
rect 46140 6575 46195 6695
rect 46315 6575 46360 6695
rect 46480 6575 46525 6695
rect 46645 6575 46690 6695
rect 46810 6575 46865 6695
rect 46985 6575 47030 6695
rect 47150 6575 47195 6695
rect 47315 6575 47360 6695
rect 47480 6575 47535 6695
rect 47655 6575 47865 6695
rect 47985 6575 48030 6695
rect 48150 6575 48195 6695
rect 48315 6575 48360 6695
rect 48480 6575 48535 6695
rect 48655 6575 48700 6695
rect 48820 6575 48865 6695
rect 48985 6575 49030 6695
rect 49150 6575 49205 6695
rect 49325 6575 49370 6695
rect 49490 6575 49535 6695
rect 49655 6575 49700 6695
rect 49820 6575 49875 6695
rect 49995 6575 50040 6695
rect 50160 6575 50205 6695
rect 50325 6575 50370 6695
rect 50490 6575 50545 6695
rect 50665 6575 50710 6695
rect 50830 6575 50875 6695
rect 50995 6575 51040 6695
rect 51160 6575 51215 6695
rect 51335 6575 51380 6695
rect 51500 6575 51545 6695
rect 51665 6575 51710 6695
rect 51830 6575 51885 6695
rect 52005 6575 52050 6695
rect 52170 6575 52215 6695
rect 52335 6575 52380 6695
rect 52500 6575 52555 6695
rect 52675 6575 52720 6695
rect 52840 6575 52885 6695
rect 53005 6575 53050 6695
rect 53170 6575 53225 6695
rect 53345 6575 53370 6695
rect 30770 6530 53370 6575
rect 30770 6410 30795 6530
rect 30915 6410 30960 6530
rect 31080 6410 31125 6530
rect 31245 6410 31290 6530
rect 31410 6410 31465 6530
rect 31585 6410 31630 6530
rect 31750 6410 31795 6530
rect 31915 6410 31960 6530
rect 32080 6410 32135 6530
rect 32255 6410 32300 6530
rect 32420 6410 32465 6530
rect 32585 6410 32630 6530
rect 32750 6410 32805 6530
rect 32925 6410 32970 6530
rect 33090 6410 33135 6530
rect 33255 6410 33300 6530
rect 33420 6410 33475 6530
rect 33595 6410 33640 6530
rect 33760 6410 33805 6530
rect 33925 6410 33970 6530
rect 34090 6410 34145 6530
rect 34265 6410 34310 6530
rect 34430 6410 34475 6530
rect 34595 6410 34640 6530
rect 34760 6410 34815 6530
rect 34935 6410 34980 6530
rect 35100 6410 35145 6530
rect 35265 6410 35310 6530
rect 35430 6410 35485 6530
rect 35605 6410 35650 6530
rect 35770 6410 35815 6530
rect 35935 6410 35980 6530
rect 36100 6410 36155 6530
rect 36275 6410 36485 6530
rect 36605 6410 36650 6530
rect 36770 6410 36815 6530
rect 36935 6410 36980 6530
rect 37100 6410 37155 6530
rect 37275 6410 37320 6530
rect 37440 6410 37485 6530
rect 37605 6410 37650 6530
rect 37770 6410 37825 6530
rect 37945 6410 37990 6530
rect 38110 6410 38155 6530
rect 38275 6410 38320 6530
rect 38440 6410 38495 6530
rect 38615 6410 38660 6530
rect 38780 6410 38825 6530
rect 38945 6410 38990 6530
rect 39110 6410 39165 6530
rect 39285 6410 39330 6530
rect 39450 6410 39495 6530
rect 39615 6410 39660 6530
rect 39780 6410 39835 6530
rect 39955 6410 40000 6530
rect 40120 6410 40165 6530
rect 40285 6410 40330 6530
rect 40450 6410 40505 6530
rect 40625 6410 40670 6530
rect 40790 6410 40835 6530
rect 40955 6410 41000 6530
rect 41120 6410 41175 6530
rect 41295 6410 41340 6530
rect 41460 6410 41505 6530
rect 41625 6410 41670 6530
rect 41790 6410 41845 6530
rect 41965 6410 42175 6530
rect 42295 6410 42340 6530
rect 42460 6410 42505 6530
rect 42625 6410 42670 6530
rect 42790 6410 42845 6530
rect 42965 6410 43010 6530
rect 43130 6410 43175 6530
rect 43295 6410 43340 6530
rect 43460 6410 43515 6530
rect 43635 6410 43680 6530
rect 43800 6410 43845 6530
rect 43965 6410 44010 6530
rect 44130 6410 44185 6530
rect 44305 6410 44350 6530
rect 44470 6410 44515 6530
rect 44635 6410 44680 6530
rect 44800 6410 44855 6530
rect 44975 6410 45020 6530
rect 45140 6410 45185 6530
rect 45305 6410 45350 6530
rect 45470 6410 45525 6530
rect 45645 6410 45690 6530
rect 45810 6410 45855 6530
rect 45975 6410 46020 6530
rect 46140 6410 46195 6530
rect 46315 6410 46360 6530
rect 46480 6410 46525 6530
rect 46645 6410 46690 6530
rect 46810 6410 46865 6530
rect 46985 6410 47030 6530
rect 47150 6410 47195 6530
rect 47315 6410 47360 6530
rect 47480 6410 47535 6530
rect 47655 6410 47865 6530
rect 47985 6410 48030 6530
rect 48150 6410 48195 6530
rect 48315 6410 48360 6530
rect 48480 6410 48535 6530
rect 48655 6410 48700 6530
rect 48820 6410 48865 6530
rect 48985 6410 49030 6530
rect 49150 6410 49205 6530
rect 49325 6410 49370 6530
rect 49490 6410 49535 6530
rect 49655 6410 49700 6530
rect 49820 6410 49875 6530
rect 49995 6410 50040 6530
rect 50160 6410 50205 6530
rect 50325 6410 50370 6530
rect 50490 6410 50545 6530
rect 50665 6410 50710 6530
rect 50830 6410 50875 6530
rect 50995 6410 51040 6530
rect 51160 6410 51215 6530
rect 51335 6410 51380 6530
rect 51500 6410 51545 6530
rect 51665 6410 51710 6530
rect 51830 6410 51885 6530
rect 52005 6410 52050 6530
rect 52170 6410 52215 6530
rect 52335 6410 52380 6530
rect 52500 6410 52555 6530
rect 52675 6410 52720 6530
rect 52840 6410 52885 6530
rect 53005 6410 53050 6530
rect 53170 6410 53225 6530
rect 53345 6410 53370 6530
rect 30770 6355 53370 6410
rect 30770 6235 30795 6355
rect 30915 6235 30960 6355
rect 31080 6235 31125 6355
rect 31245 6235 31290 6355
rect 31410 6235 31465 6355
rect 31585 6235 31630 6355
rect 31750 6235 31795 6355
rect 31915 6235 31960 6355
rect 32080 6235 32135 6355
rect 32255 6235 32300 6355
rect 32420 6235 32465 6355
rect 32585 6235 32630 6355
rect 32750 6235 32805 6355
rect 32925 6235 32970 6355
rect 33090 6235 33135 6355
rect 33255 6235 33300 6355
rect 33420 6235 33475 6355
rect 33595 6235 33640 6355
rect 33760 6235 33805 6355
rect 33925 6235 33970 6355
rect 34090 6235 34145 6355
rect 34265 6235 34310 6355
rect 34430 6235 34475 6355
rect 34595 6235 34640 6355
rect 34760 6235 34815 6355
rect 34935 6235 34980 6355
rect 35100 6235 35145 6355
rect 35265 6235 35310 6355
rect 35430 6235 35485 6355
rect 35605 6235 35650 6355
rect 35770 6235 35815 6355
rect 35935 6235 35980 6355
rect 36100 6235 36155 6355
rect 36275 6235 36485 6355
rect 36605 6235 36650 6355
rect 36770 6235 36815 6355
rect 36935 6235 36980 6355
rect 37100 6235 37155 6355
rect 37275 6235 37320 6355
rect 37440 6235 37485 6355
rect 37605 6235 37650 6355
rect 37770 6235 37825 6355
rect 37945 6235 37990 6355
rect 38110 6235 38155 6355
rect 38275 6235 38320 6355
rect 38440 6235 38495 6355
rect 38615 6235 38660 6355
rect 38780 6235 38825 6355
rect 38945 6235 38990 6355
rect 39110 6235 39165 6355
rect 39285 6235 39330 6355
rect 39450 6235 39495 6355
rect 39615 6235 39660 6355
rect 39780 6235 39835 6355
rect 39955 6235 40000 6355
rect 40120 6235 40165 6355
rect 40285 6235 40330 6355
rect 40450 6235 40505 6355
rect 40625 6235 40670 6355
rect 40790 6235 40835 6355
rect 40955 6235 41000 6355
rect 41120 6235 41175 6355
rect 41295 6235 41340 6355
rect 41460 6235 41505 6355
rect 41625 6235 41670 6355
rect 41790 6235 41845 6355
rect 41965 6235 42175 6355
rect 42295 6235 42340 6355
rect 42460 6235 42505 6355
rect 42625 6235 42670 6355
rect 42790 6235 42845 6355
rect 42965 6235 43010 6355
rect 43130 6235 43175 6355
rect 43295 6235 43340 6355
rect 43460 6235 43515 6355
rect 43635 6235 43680 6355
rect 43800 6235 43845 6355
rect 43965 6235 44010 6355
rect 44130 6235 44185 6355
rect 44305 6235 44350 6355
rect 44470 6235 44515 6355
rect 44635 6235 44680 6355
rect 44800 6235 44855 6355
rect 44975 6235 45020 6355
rect 45140 6235 45185 6355
rect 45305 6235 45350 6355
rect 45470 6235 45525 6355
rect 45645 6235 45690 6355
rect 45810 6235 45855 6355
rect 45975 6235 46020 6355
rect 46140 6235 46195 6355
rect 46315 6235 46360 6355
rect 46480 6235 46525 6355
rect 46645 6235 46690 6355
rect 46810 6235 46865 6355
rect 46985 6235 47030 6355
rect 47150 6235 47195 6355
rect 47315 6235 47360 6355
rect 47480 6235 47535 6355
rect 47655 6235 47865 6355
rect 47985 6235 48030 6355
rect 48150 6235 48195 6355
rect 48315 6235 48360 6355
rect 48480 6235 48535 6355
rect 48655 6235 48700 6355
rect 48820 6235 48865 6355
rect 48985 6235 49030 6355
rect 49150 6235 49205 6355
rect 49325 6235 49370 6355
rect 49490 6235 49535 6355
rect 49655 6235 49700 6355
rect 49820 6235 49875 6355
rect 49995 6235 50040 6355
rect 50160 6235 50205 6355
rect 50325 6235 50370 6355
rect 50490 6235 50545 6355
rect 50665 6235 50710 6355
rect 50830 6235 50875 6355
rect 50995 6235 51040 6355
rect 51160 6235 51215 6355
rect 51335 6235 51380 6355
rect 51500 6235 51545 6355
rect 51665 6235 51710 6355
rect 51830 6235 51885 6355
rect 52005 6235 52050 6355
rect 52170 6235 52215 6355
rect 52335 6235 52380 6355
rect 52500 6235 52555 6355
rect 52675 6235 52720 6355
rect 52840 6235 52885 6355
rect 53005 6235 53050 6355
rect 53170 6235 53225 6355
rect 53345 6235 53370 6355
rect 30770 6190 53370 6235
rect 30770 6070 30795 6190
rect 30915 6070 30960 6190
rect 31080 6070 31125 6190
rect 31245 6070 31290 6190
rect 31410 6070 31465 6190
rect 31585 6070 31630 6190
rect 31750 6070 31795 6190
rect 31915 6070 31960 6190
rect 32080 6070 32135 6190
rect 32255 6070 32300 6190
rect 32420 6070 32465 6190
rect 32585 6070 32630 6190
rect 32750 6070 32805 6190
rect 32925 6070 32970 6190
rect 33090 6070 33135 6190
rect 33255 6070 33300 6190
rect 33420 6070 33475 6190
rect 33595 6070 33640 6190
rect 33760 6070 33805 6190
rect 33925 6070 33970 6190
rect 34090 6070 34145 6190
rect 34265 6070 34310 6190
rect 34430 6070 34475 6190
rect 34595 6070 34640 6190
rect 34760 6070 34815 6190
rect 34935 6070 34980 6190
rect 35100 6070 35145 6190
rect 35265 6070 35310 6190
rect 35430 6070 35485 6190
rect 35605 6070 35650 6190
rect 35770 6070 35815 6190
rect 35935 6070 35980 6190
rect 36100 6070 36155 6190
rect 36275 6070 36485 6190
rect 36605 6070 36650 6190
rect 36770 6070 36815 6190
rect 36935 6070 36980 6190
rect 37100 6070 37155 6190
rect 37275 6070 37320 6190
rect 37440 6070 37485 6190
rect 37605 6070 37650 6190
rect 37770 6070 37825 6190
rect 37945 6070 37990 6190
rect 38110 6070 38155 6190
rect 38275 6070 38320 6190
rect 38440 6070 38495 6190
rect 38615 6070 38660 6190
rect 38780 6070 38825 6190
rect 38945 6070 38990 6190
rect 39110 6070 39165 6190
rect 39285 6070 39330 6190
rect 39450 6070 39495 6190
rect 39615 6070 39660 6190
rect 39780 6070 39835 6190
rect 39955 6070 40000 6190
rect 40120 6070 40165 6190
rect 40285 6070 40330 6190
rect 40450 6070 40505 6190
rect 40625 6070 40670 6190
rect 40790 6070 40835 6190
rect 40955 6070 41000 6190
rect 41120 6070 41175 6190
rect 41295 6070 41340 6190
rect 41460 6070 41505 6190
rect 41625 6070 41670 6190
rect 41790 6070 41845 6190
rect 41965 6070 42175 6190
rect 42295 6070 42340 6190
rect 42460 6070 42505 6190
rect 42625 6070 42670 6190
rect 42790 6070 42845 6190
rect 42965 6070 43010 6190
rect 43130 6070 43175 6190
rect 43295 6070 43340 6190
rect 43460 6070 43515 6190
rect 43635 6070 43680 6190
rect 43800 6070 43845 6190
rect 43965 6070 44010 6190
rect 44130 6070 44185 6190
rect 44305 6070 44350 6190
rect 44470 6070 44515 6190
rect 44635 6070 44680 6190
rect 44800 6070 44855 6190
rect 44975 6070 45020 6190
rect 45140 6070 45185 6190
rect 45305 6070 45350 6190
rect 45470 6070 45525 6190
rect 45645 6070 45690 6190
rect 45810 6070 45855 6190
rect 45975 6070 46020 6190
rect 46140 6070 46195 6190
rect 46315 6070 46360 6190
rect 46480 6070 46525 6190
rect 46645 6070 46690 6190
rect 46810 6070 46865 6190
rect 46985 6070 47030 6190
rect 47150 6070 47195 6190
rect 47315 6070 47360 6190
rect 47480 6070 47535 6190
rect 47655 6070 47865 6190
rect 47985 6070 48030 6190
rect 48150 6070 48195 6190
rect 48315 6070 48360 6190
rect 48480 6070 48535 6190
rect 48655 6070 48700 6190
rect 48820 6070 48865 6190
rect 48985 6070 49030 6190
rect 49150 6070 49205 6190
rect 49325 6070 49370 6190
rect 49490 6070 49535 6190
rect 49655 6070 49700 6190
rect 49820 6070 49875 6190
rect 49995 6070 50040 6190
rect 50160 6070 50205 6190
rect 50325 6070 50370 6190
rect 50490 6070 50545 6190
rect 50665 6070 50710 6190
rect 50830 6070 50875 6190
rect 50995 6070 51040 6190
rect 51160 6070 51215 6190
rect 51335 6070 51380 6190
rect 51500 6070 51545 6190
rect 51665 6070 51710 6190
rect 51830 6070 51885 6190
rect 52005 6070 52050 6190
rect 52170 6070 52215 6190
rect 52335 6070 52380 6190
rect 52500 6070 52555 6190
rect 52675 6070 52720 6190
rect 52840 6070 52885 6190
rect 53005 6070 53050 6190
rect 53170 6070 53225 6190
rect 53345 6070 53370 6190
rect 30770 6025 53370 6070
rect 30770 5905 30795 6025
rect 30915 5905 30960 6025
rect 31080 5905 31125 6025
rect 31245 5905 31290 6025
rect 31410 5905 31465 6025
rect 31585 5905 31630 6025
rect 31750 5905 31795 6025
rect 31915 5905 31960 6025
rect 32080 5905 32135 6025
rect 32255 5905 32300 6025
rect 32420 5905 32465 6025
rect 32585 5905 32630 6025
rect 32750 5905 32805 6025
rect 32925 5905 32970 6025
rect 33090 5905 33135 6025
rect 33255 5905 33300 6025
rect 33420 5905 33475 6025
rect 33595 5905 33640 6025
rect 33760 5905 33805 6025
rect 33925 5905 33970 6025
rect 34090 5905 34145 6025
rect 34265 5905 34310 6025
rect 34430 5905 34475 6025
rect 34595 5905 34640 6025
rect 34760 5905 34815 6025
rect 34935 5905 34980 6025
rect 35100 5905 35145 6025
rect 35265 5905 35310 6025
rect 35430 5905 35485 6025
rect 35605 5905 35650 6025
rect 35770 5905 35815 6025
rect 35935 5905 35980 6025
rect 36100 5905 36155 6025
rect 36275 5905 36485 6025
rect 36605 5905 36650 6025
rect 36770 5905 36815 6025
rect 36935 5905 36980 6025
rect 37100 5905 37155 6025
rect 37275 5905 37320 6025
rect 37440 5905 37485 6025
rect 37605 5905 37650 6025
rect 37770 5905 37825 6025
rect 37945 5905 37990 6025
rect 38110 5905 38155 6025
rect 38275 5905 38320 6025
rect 38440 5905 38495 6025
rect 38615 5905 38660 6025
rect 38780 5905 38825 6025
rect 38945 5905 38990 6025
rect 39110 5905 39165 6025
rect 39285 5905 39330 6025
rect 39450 5905 39495 6025
rect 39615 5905 39660 6025
rect 39780 5905 39835 6025
rect 39955 5905 40000 6025
rect 40120 5905 40165 6025
rect 40285 5905 40330 6025
rect 40450 5905 40505 6025
rect 40625 5905 40670 6025
rect 40790 5905 40835 6025
rect 40955 5905 41000 6025
rect 41120 5905 41175 6025
rect 41295 5905 41340 6025
rect 41460 5905 41505 6025
rect 41625 5905 41670 6025
rect 41790 5905 41845 6025
rect 41965 5905 42175 6025
rect 42295 5905 42340 6025
rect 42460 5905 42505 6025
rect 42625 5905 42670 6025
rect 42790 5905 42845 6025
rect 42965 5905 43010 6025
rect 43130 5905 43175 6025
rect 43295 5905 43340 6025
rect 43460 5905 43515 6025
rect 43635 5905 43680 6025
rect 43800 5905 43845 6025
rect 43965 5905 44010 6025
rect 44130 5905 44185 6025
rect 44305 5905 44350 6025
rect 44470 5905 44515 6025
rect 44635 5905 44680 6025
rect 44800 5905 44855 6025
rect 44975 5905 45020 6025
rect 45140 5905 45185 6025
rect 45305 5905 45350 6025
rect 45470 5905 45525 6025
rect 45645 5905 45690 6025
rect 45810 5905 45855 6025
rect 45975 5905 46020 6025
rect 46140 5905 46195 6025
rect 46315 5905 46360 6025
rect 46480 5905 46525 6025
rect 46645 5905 46690 6025
rect 46810 5905 46865 6025
rect 46985 5905 47030 6025
rect 47150 5905 47195 6025
rect 47315 5905 47360 6025
rect 47480 5905 47535 6025
rect 47655 5905 47865 6025
rect 47985 5905 48030 6025
rect 48150 5905 48195 6025
rect 48315 5905 48360 6025
rect 48480 5905 48535 6025
rect 48655 5905 48700 6025
rect 48820 5905 48865 6025
rect 48985 5905 49030 6025
rect 49150 5905 49205 6025
rect 49325 5905 49370 6025
rect 49490 5905 49535 6025
rect 49655 5905 49700 6025
rect 49820 5905 49875 6025
rect 49995 5905 50040 6025
rect 50160 5905 50205 6025
rect 50325 5905 50370 6025
rect 50490 5905 50545 6025
rect 50665 5905 50710 6025
rect 50830 5905 50875 6025
rect 50995 5905 51040 6025
rect 51160 5905 51215 6025
rect 51335 5905 51380 6025
rect 51500 5905 51545 6025
rect 51665 5905 51710 6025
rect 51830 5905 51885 6025
rect 52005 5905 52050 6025
rect 52170 5905 52215 6025
rect 52335 5905 52380 6025
rect 52500 5905 52555 6025
rect 52675 5905 52720 6025
rect 52840 5905 52885 6025
rect 53005 5905 53050 6025
rect 53170 5905 53225 6025
rect 53345 5905 53370 6025
rect 30770 5860 53370 5905
rect 30770 5740 30795 5860
rect 30915 5740 30960 5860
rect 31080 5740 31125 5860
rect 31245 5740 31290 5860
rect 31410 5740 31465 5860
rect 31585 5740 31630 5860
rect 31750 5740 31795 5860
rect 31915 5740 31960 5860
rect 32080 5740 32135 5860
rect 32255 5740 32300 5860
rect 32420 5740 32465 5860
rect 32585 5740 32630 5860
rect 32750 5740 32805 5860
rect 32925 5740 32970 5860
rect 33090 5740 33135 5860
rect 33255 5740 33300 5860
rect 33420 5740 33475 5860
rect 33595 5740 33640 5860
rect 33760 5740 33805 5860
rect 33925 5740 33970 5860
rect 34090 5740 34145 5860
rect 34265 5740 34310 5860
rect 34430 5740 34475 5860
rect 34595 5740 34640 5860
rect 34760 5740 34815 5860
rect 34935 5740 34980 5860
rect 35100 5740 35145 5860
rect 35265 5740 35310 5860
rect 35430 5740 35485 5860
rect 35605 5740 35650 5860
rect 35770 5740 35815 5860
rect 35935 5740 35980 5860
rect 36100 5740 36155 5860
rect 36275 5740 36485 5860
rect 36605 5740 36650 5860
rect 36770 5740 36815 5860
rect 36935 5740 36980 5860
rect 37100 5740 37155 5860
rect 37275 5740 37320 5860
rect 37440 5740 37485 5860
rect 37605 5740 37650 5860
rect 37770 5740 37825 5860
rect 37945 5740 37990 5860
rect 38110 5740 38155 5860
rect 38275 5740 38320 5860
rect 38440 5740 38495 5860
rect 38615 5740 38660 5860
rect 38780 5740 38825 5860
rect 38945 5740 38990 5860
rect 39110 5740 39165 5860
rect 39285 5740 39330 5860
rect 39450 5740 39495 5860
rect 39615 5740 39660 5860
rect 39780 5740 39835 5860
rect 39955 5740 40000 5860
rect 40120 5740 40165 5860
rect 40285 5740 40330 5860
rect 40450 5740 40505 5860
rect 40625 5740 40670 5860
rect 40790 5740 40835 5860
rect 40955 5740 41000 5860
rect 41120 5740 41175 5860
rect 41295 5740 41340 5860
rect 41460 5740 41505 5860
rect 41625 5740 41670 5860
rect 41790 5740 41845 5860
rect 41965 5740 42175 5860
rect 42295 5740 42340 5860
rect 42460 5740 42505 5860
rect 42625 5740 42670 5860
rect 42790 5740 42845 5860
rect 42965 5740 43010 5860
rect 43130 5740 43175 5860
rect 43295 5740 43340 5860
rect 43460 5740 43515 5860
rect 43635 5740 43680 5860
rect 43800 5740 43845 5860
rect 43965 5740 44010 5860
rect 44130 5740 44185 5860
rect 44305 5740 44350 5860
rect 44470 5740 44515 5860
rect 44635 5740 44680 5860
rect 44800 5740 44855 5860
rect 44975 5740 45020 5860
rect 45140 5740 45185 5860
rect 45305 5740 45350 5860
rect 45470 5740 45525 5860
rect 45645 5740 45690 5860
rect 45810 5740 45855 5860
rect 45975 5740 46020 5860
rect 46140 5740 46195 5860
rect 46315 5740 46360 5860
rect 46480 5740 46525 5860
rect 46645 5740 46690 5860
rect 46810 5740 46865 5860
rect 46985 5740 47030 5860
rect 47150 5740 47195 5860
rect 47315 5740 47360 5860
rect 47480 5740 47535 5860
rect 47655 5740 47865 5860
rect 47985 5740 48030 5860
rect 48150 5740 48195 5860
rect 48315 5740 48360 5860
rect 48480 5740 48535 5860
rect 48655 5740 48700 5860
rect 48820 5740 48865 5860
rect 48985 5740 49030 5860
rect 49150 5740 49205 5860
rect 49325 5740 49370 5860
rect 49490 5740 49535 5860
rect 49655 5740 49700 5860
rect 49820 5740 49875 5860
rect 49995 5740 50040 5860
rect 50160 5740 50205 5860
rect 50325 5740 50370 5860
rect 50490 5740 50545 5860
rect 50665 5740 50710 5860
rect 50830 5740 50875 5860
rect 50995 5740 51040 5860
rect 51160 5740 51215 5860
rect 51335 5740 51380 5860
rect 51500 5740 51545 5860
rect 51665 5740 51710 5860
rect 51830 5740 51885 5860
rect 52005 5740 52050 5860
rect 52170 5740 52215 5860
rect 52335 5740 52380 5860
rect 52500 5740 52555 5860
rect 52675 5740 52720 5860
rect 52840 5740 52885 5860
rect 53005 5740 53050 5860
rect 53170 5740 53225 5860
rect 53345 5740 53370 5860
rect 30770 5685 53370 5740
rect 30770 5565 30795 5685
rect 30915 5565 30960 5685
rect 31080 5565 31125 5685
rect 31245 5565 31290 5685
rect 31410 5565 31465 5685
rect 31585 5565 31630 5685
rect 31750 5565 31795 5685
rect 31915 5565 31960 5685
rect 32080 5565 32135 5685
rect 32255 5565 32300 5685
rect 32420 5565 32465 5685
rect 32585 5565 32630 5685
rect 32750 5565 32805 5685
rect 32925 5565 32970 5685
rect 33090 5565 33135 5685
rect 33255 5565 33300 5685
rect 33420 5565 33475 5685
rect 33595 5565 33640 5685
rect 33760 5565 33805 5685
rect 33925 5565 33970 5685
rect 34090 5565 34145 5685
rect 34265 5565 34310 5685
rect 34430 5565 34475 5685
rect 34595 5565 34640 5685
rect 34760 5565 34815 5685
rect 34935 5565 34980 5685
rect 35100 5565 35145 5685
rect 35265 5565 35310 5685
rect 35430 5565 35485 5685
rect 35605 5565 35650 5685
rect 35770 5565 35815 5685
rect 35935 5565 35980 5685
rect 36100 5565 36155 5685
rect 36275 5565 36485 5685
rect 36605 5565 36650 5685
rect 36770 5565 36815 5685
rect 36935 5565 36980 5685
rect 37100 5565 37155 5685
rect 37275 5565 37320 5685
rect 37440 5565 37485 5685
rect 37605 5565 37650 5685
rect 37770 5565 37825 5685
rect 37945 5565 37990 5685
rect 38110 5565 38155 5685
rect 38275 5565 38320 5685
rect 38440 5565 38495 5685
rect 38615 5565 38660 5685
rect 38780 5565 38825 5685
rect 38945 5565 38990 5685
rect 39110 5565 39165 5685
rect 39285 5565 39330 5685
rect 39450 5565 39495 5685
rect 39615 5565 39660 5685
rect 39780 5565 39835 5685
rect 39955 5565 40000 5685
rect 40120 5565 40165 5685
rect 40285 5565 40330 5685
rect 40450 5565 40505 5685
rect 40625 5565 40670 5685
rect 40790 5565 40835 5685
rect 40955 5565 41000 5685
rect 41120 5565 41175 5685
rect 41295 5565 41340 5685
rect 41460 5565 41505 5685
rect 41625 5565 41670 5685
rect 41790 5565 41845 5685
rect 41965 5565 42175 5685
rect 42295 5565 42340 5685
rect 42460 5565 42505 5685
rect 42625 5565 42670 5685
rect 42790 5565 42845 5685
rect 42965 5565 43010 5685
rect 43130 5565 43175 5685
rect 43295 5565 43340 5685
rect 43460 5565 43515 5685
rect 43635 5565 43680 5685
rect 43800 5565 43845 5685
rect 43965 5565 44010 5685
rect 44130 5565 44185 5685
rect 44305 5565 44350 5685
rect 44470 5565 44515 5685
rect 44635 5565 44680 5685
rect 44800 5565 44855 5685
rect 44975 5565 45020 5685
rect 45140 5565 45185 5685
rect 45305 5565 45350 5685
rect 45470 5565 45525 5685
rect 45645 5565 45690 5685
rect 45810 5565 45855 5685
rect 45975 5565 46020 5685
rect 46140 5565 46195 5685
rect 46315 5565 46360 5685
rect 46480 5565 46525 5685
rect 46645 5565 46690 5685
rect 46810 5565 46865 5685
rect 46985 5565 47030 5685
rect 47150 5565 47195 5685
rect 47315 5565 47360 5685
rect 47480 5565 47535 5685
rect 47655 5565 47865 5685
rect 47985 5565 48030 5685
rect 48150 5565 48195 5685
rect 48315 5565 48360 5685
rect 48480 5565 48535 5685
rect 48655 5565 48700 5685
rect 48820 5565 48865 5685
rect 48985 5565 49030 5685
rect 49150 5565 49205 5685
rect 49325 5565 49370 5685
rect 49490 5565 49535 5685
rect 49655 5565 49700 5685
rect 49820 5565 49875 5685
rect 49995 5565 50040 5685
rect 50160 5565 50205 5685
rect 50325 5565 50370 5685
rect 50490 5565 50545 5685
rect 50665 5565 50710 5685
rect 50830 5565 50875 5685
rect 50995 5565 51040 5685
rect 51160 5565 51215 5685
rect 51335 5565 51380 5685
rect 51500 5565 51545 5685
rect 51665 5565 51710 5685
rect 51830 5565 51885 5685
rect 52005 5565 52050 5685
rect 52170 5565 52215 5685
rect 52335 5565 52380 5685
rect 52500 5565 52555 5685
rect 52675 5565 52720 5685
rect 52840 5565 52885 5685
rect 53005 5565 53050 5685
rect 53170 5565 53225 5685
rect 53345 5565 53370 5685
rect 30770 5520 53370 5565
rect 30770 5400 30795 5520
rect 30915 5400 30960 5520
rect 31080 5400 31125 5520
rect 31245 5400 31290 5520
rect 31410 5400 31465 5520
rect 31585 5400 31630 5520
rect 31750 5400 31795 5520
rect 31915 5400 31960 5520
rect 32080 5400 32135 5520
rect 32255 5400 32300 5520
rect 32420 5400 32465 5520
rect 32585 5400 32630 5520
rect 32750 5400 32805 5520
rect 32925 5400 32970 5520
rect 33090 5400 33135 5520
rect 33255 5400 33300 5520
rect 33420 5400 33475 5520
rect 33595 5400 33640 5520
rect 33760 5400 33805 5520
rect 33925 5400 33970 5520
rect 34090 5400 34145 5520
rect 34265 5400 34310 5520
rect 34430 5400 34475 5520
rect 34595 5400 34640 5520
rect 34760 5400 34815 5520
rect 34935 5400 34980 5520
rect 35100 5400 35145 5520
rect 35265 5400 35310 5520
rect 35430 5400 35485 5520
rect 35605 5400 35650 5520
rect 35770 5400 35815 5520
rect 35935 5400 35980 5520
rect 36100 5400 36155 5520
rect 36275 5400 36485 5520
rect 36605 5400 36650 5520
rect 36770 5400 36815 5520
rect 36935 5400 36980 5520
rect 37100 5400 37155 5520
rect 37275 5400 37320 5520
rect 37440 5400 37485 5520
rect 37605 5400 37650 5520
rect 37770 5400 37825 5520
rect 37945 5400 37990 5520
rect 38110 5400 38155 5520
rect 38275 5400 38320 5520
rect 38440 5400 38495 5520
rect 38615 5400 38660 5520
rect 38780 5400 38825 5520
rect 38945 5400 38990 5520
rect 39110 5400 39165 5520
rect 39285 5400 39330 5520
rect 39450 5400 39495 5520
rect 39615 5400 39660 5520
rect 39780 5400 39835 5520
rect 39955 5400 40000 5520
rect 40120 5400 40165 5520
rect 40285 5400 40330 5520
rect 40450 5400 40505 5520
rect 40625 5400 40670 5520
rect 40790 5400 40835 5520
rect 40955 5400 41000 5520
rect 41120 5400 41175 5520
rect 41295 5400 41340 5520
rect 41460 5400 41505 5520
rect 41625 5400 41670 5520
rect 41790 5400 41845 5520
rect 41965 5400 42175 5520
rect 42295 5400 42340 5520
rect 42460 5400 42505 5520
rect 42625 5400 42670 5520
rect 42790 5400 42845 5520
rect 42965 5400 43010 5520
rect 43130 5400 43175 5520
rect 43295 5400 43340 5520
rect 43460 5400 43515 5520
rect 43635 5400 43680 5520
rect 43800 5400 43845 5520
rect 43965 5400 44010 5520
rect 44130 5400 44185 5520
rect 44305 5400 44350 5520
rect 44470 5400 44515 5520
rect 44635 5400 44680 5520
rect 44800 5400 44855 5520
rect 44975 5400 45020 5520
rect 45140 5400 45185 5520
rect 45305 5400 45350 5520
rect 45470 5400 45525 5520
rect 45645 5400 45690 5520
rect 45810 5400 45855 5520
rect 45975 5400 46020 5520
rect 46140 5400 46195 5520
rect 46315 5400 46360 5520
rect 46480 5400 46525 5520
rect 46645 5400 46690 5520
rect 46810 5400 46865 5520
rect 46985 5400 47030 5520
rect 47150 5400 47195 5520
rect 47315 5400 47360 5520
rect 47480 5400 47535 5520
rect 47655 5400 47865 5520
rect 47985 5400 48030 5520
rect 48150 5400 48195 5520
rect 48315 5400 48360 5520
rect 48480 5400 48535 5520
rect 48655 5400 48700 5520
rect 48820 5400 48865 5520
rect 48985 5400 49030 5520
rect 49150 5400 49205 5520
rect 49325 5400 49370 5520
rect 49490 5400 49535 5520
rect 49655 5400 49700 5520
rect 49820 5400 49875 5520
rect 49995 5400 50040 5520
rect 50160 5400 50205 5520
rect 50325 5400 50370 5520
rect 50490 5400 50545 5520
rect 50665 5400 50710 5520
rect 50830 5400 50875 5520
rect 50995 5400 51040 5520
rect 51160 5400 51215 5520
rect 51335 5400 51380 5520
rect 51500 5400 51545 5520
rect 51665 5400 51710 5520
rect 51830 5400 51885 5520
rect 52005 5400 52050 5520
rect 52170 5400 52215 5520
rect 52335 5400 52380 5520
rect 52500 5400 52555 5520
rect 52675 5400 52720 5520
rect 52840 5400 52885 5520
rect 53005 5400 53050 5520
rect 53170 5400 53225 5520
rect 53345 5400 53370 5520
rect 30770 5355 53370 5400
rect 30770 5235 30795 5355
rect 30915 5235 30960 5355
rect 31080 5235 31125 5355
rect 31245 5235 31290 5355
rect 31410 5235 31465 5355
rect 31585 5235 31630 5355
rect 31750 5235 31795 5355
rect 31915 5235 31960 5355
rect 32080 5235 32135 5355
rect 32255 5235 32300 5355
rect 32420 5235 32465 5355
rect 32585 5235 32630 5355
rect 32750 5235 32805 5355
rect 32925 5235 32970 5355
rect 33090 5235 33135 5355
rect 33255 5235 33300 5355
rect 33420 5235 33475 5355
rect 33595 5235 33640 5355
rect 33760 5235 33805 5355
rect 33925 5235 33970 5355
rect 34090 5235 34145 5355
rect 34265 5235 34310 5355
rect 34430 5235 34475 5355
rect 34595 5235 34640 5355
rect 34760 5235 34815 5355
rect 34935 5235 34980 5355
rect 35100 5235 35145 5355
rect 35265 5235 35310 5355
rect 35430 5235 35485 5355
rect 35605 5235 35650 5355
rect 35770 5235 35815 5355
rect 35935 5235 35980 5355
rect 36100 5235 36155 5355
rect 36275 5235 36485 5355
rect 36605 5235 36650 5355
rect 36770 5235 36815 5355
rect 36935 5235 36980 5355
rect 37100 5235 37155 5355
rect 37275 5235 37320 5355
rect 37440 5235 37485 5355
rect 37605 5235 37650 5355
rect 37770 5235 37825 5355
rect 37945 5235 37990 5355
rect 38110 5235 38155 5355
rect 38275 5235 38320 5355
rect 38440 5235 38495 5355
rect 38615 5235 38660 5355
rect 38780 5235 38825 5355
rect 38945 5235 38990 5355
rect 39110 5235 39165 5355
rect 39285 5235 39330 5355
rect 39450 5235 39495 5355
rect 39615 5235 39660 5355
rect 39780 5235 39835 5355
rect 39955 5235 40000 5355
rect 40120 5235 40165 5355
rect 40285 5235 40330 5355
rect 40450 5235 40505 5355
rect 40625 5235 40670 5355
rect 40790 5235 40835 5355
rect 40955 5235 41000 5355
rect 41120 5235 41175 5355
rect 41295 5235 41340 5355
rect 41460 5235 41505 5355
rect 41625 5235 41670 5355
rect 41790 5235 41845 5355
rect 41965 5235 42175 5355
rect 42295 5235 42340 5355
rect 42460 5235 42505 5355
rect 42625 5235 42670 5355
rect 42790 5235 42845 5355
rect 42965 5235 43010 5355
rect 43130 5235 43175 5355
rect 43295 5235 43340 5355
rect 43460 5235 43515 5355
rect 43635 5235 43680 5355
rect 43800 5235 43845 5355
rect 43965 5235 44010 5355
rect 44130 5235 44185 5355
rect 44305 5235 44350 5355
rect 44470 5235 44515 5355
rect 44635 5235 44680 5355
rect 44800 5235 44855 5355
rect 44975 5235 45020 5355
rect 45140 5235 45185 5355
rect 45305 5235 45350 5355
rect 45470 5235 45525 5355
rect 45645 5235 45690 5355
rect 45810 5235 45855 5355
rect 45975 5235 46020 5355
rect 46140 5235 46195 5355
rect 46315 5235 46360 5355
rect 46480 5235 46525 5355
rect 46645 5235 46690 5355
rect 46810 5235 46865 5355
rect 46985 5235 47030 5355
rect 47150 5235 47195 5355
rect 47315 5235 47360 5355
rect 47480 5235 47535 5355
rect 47655 5235 47865 5355
rect 47985 5235 48030 5355
rect 48150 5235 48195 5355
rect 48315 5235 48360 5355
rect 48480 5235 48535 5355
rect 48655 5235 48700 5355
rect 48820 5235 48865 5355
rect 48985 5235 49030 5355
rect 49150 5235 49205 5355
rect 49325 5235 49370 5355
rect 49490 5235 49535 5355
rect 49655 5235 49700 5355
rect 49820 5235 49875 5355
rect 49995 5235 50040 5355
rect 50160 5235 50205 5355
rect 50325 5235 50370 5355
rect 50490 5235 50545 5355
rect 50665 5235 50710 5355
rect 50830 5235 50875 5355
rect 50995 5235 51040 5355
rect 51160 5235 51215 5355
rect 51335 5235 51380 5355
rect 51500 5235 51545 5355
rect 51665 5235 51710 5355
rect 51830 5235 51885 5355
rect 52005 5235 52050 5355
rect 52170 5235 52215 5355
rect 52335 5235 52380 5355
rect 52500 5235 52555 5355
rect 52675 5235 52720 5355
rect 52840 5235 52885 5355
rect 53005 5235 53050 5355
rect 53170 5235 53225 5355
rect 53345 5235 53370 5355
rect 30770 5190 53370 5235
rect 30770 5070 30795 5190
rect 30915 5070 30960 5190
rect 31080 5070 31125 5190
rect 31245 5070 31290 5190
rect 31410 5070 31465 5190
rect 31585 5070 31630 5190
rect 31750 5070 31795 5190
rect 31915 5070 31960 5190
rect 32080 5070 32135 5190
rect 32255 5070 32300 5190
rect 32420 5070 32465 5190
rect 32585 5070 32630 5190
rect 32750 5070 32805 5190
rect 32925 5070 32970 5190
rect 33090 5070 33135 5190
rect 33255 5070 33300 5190
rect 33420 5070 33475 5190
rect 33595 5070 33640 5190
rect 33760 5070 33805 5190
rect 33925 5070 33970 5190
rect 34090 5070 34145 5190
rect 34265 5070 34310 5190
rect 34430 5070 34475 5190
rect 34595 5070 34640 5190
rect 34760 5070 34815 5190
rect 34935 5070 34980 5190
rect 35100 5070 35145 5190
rect 35265 5070 35310 5190
rect 35430 5070 35485 5190
rect 35605 5070 35650 5190
rect 35770 5070 35815 5190
rect 35935 5070 35980 5190
rect 36100 5070 36155 5190
rect 36275 5070 36485 5190
rect 36605 5070 36650 5190
rect 36770 5070 36815 5190
rect 36935 5070 36980 5190
rect 37100 5070 37155 5190
rect 37275 5070 37320 5190
rect 37440 5070 37485 5190
rect 37605 5070 37650 5190
rect 37770 5070 37825 5190
rect 37945 5070 37990 5190
rect 38110 5070 38155 5190
rect 38275 5070 38320 5190
rect 38440 5070 38495 5190
rect 38615 5070 38660 5190
rect 38780 5070 38825 5190
rect 38945 5070 38990 5190
rect 39110 5070 39165 5190
rect 39285 5070 39330 5190
rect 39450 5070 39495 5190
rect 39615 5070 39660 5190
rect 39780 5070 39835 5190
rect 39955 5070 40000 5190
rect 40120 5070 40165 5190
rect 40285 5070 40330 5190
rect 40450 5070 40505 5190
rect 40625 5070 40670 5190
rect 40790 5070 40835 5190
rect 40955 5070 41000 5190
rect 41120 5070 41175 5190
rect 41295 5070 41340 5190
rect 41460 5070 41505 5190
rect 41625 5070 41670 5190
rect 41790 5070 41845 5190
rect 41965 5070 42175 5190
rect 42295 5070 42340 5190
rect 42460 5070 42505 5190
rect 42625 5070 42670 5190
rect 42790 5070 42845 5190
rect 42965 5070 43010 5190
rect 43130 5070 43175 5190
rect 43295 5070 43340 5190
rect 43460 5070 43515 5190
rect 43635 5070 43680 5190
rect 43800 5070 43845 5190
rect 43965 5070 44010 5190
rect 44130 5070 44185 5190
rect 44305 5070 44350 5190
rect 44470 5070 44515 5190
rect 44635 5070 44680 5190
rect 44800 5070 44855 5190
rect 44975 5070 45020 5190
rect 45140 5070 45185 5190
rect 45305 5070 45350 5190
rect 45470 5070 45525 5190
rect 45645 5070 45690 5190
rect 45810 5070 45855 5190
rect 45975 5070 46020 5190
rect 46140 5070 46195 5190
rect 46315 5070 46360 5190
rect 46480 5070 46525 5190
rect 46645 5070 46690 5190
rect 46810 5070 46865 5190
rect 46985 5070 47030 5190
rect 47150 5070 47195 5190
rect 47315 5070 47360 5190
rect 47480 5070 47535 5190
rect 47655 5070 47865 5190
rect 47985 5070 48030 5190
rect 48150 5070 48195 5190
rect 48315 5070 48360 5190
rect 48480 5070 48535 5190
rect 48655 5070 48700 5190
rect 48820 5070 48865 5190
rect 48985 5070 49030 5190
rect 49150 5070 49205 5190
rect 49325 5070 49370 5190
rect 49490 5070 49535 5190
rect 49655 5070 49700 5190
rect 49820 5070 49875 5190
rect 49995 5070 50040 5190
rect 50160 5070 50205 5190
rect 50325 5070 50370 5190
rect 50490 5070 50545 5190
rect 50665 5070 50710 5190
rect 50830 5070 50875 5190
rect 50995 5070 51040 5190
rect 51160 5070 51215 5190
rect 51335 5070 51380 5190
rect 51500 5070 51545 5190
rect 51665 5070 51710 5190
rect 51830 5070 51885 5190
rect 52005 5070 52050 5190
rect 52170 5070 52215 5190
rect 52335 5070 52380 5190
rect 52500 5070 52555 5190
rect 52675 5070 52720 5190
rect 52840 5070 52885 5190
rect 53005 5070 53050 5190
rect 53170 5070 53225 5190
rect 53345 5070 53370 5190
rect 30770 5015 53370 5070
rect 30770 4895 30795 5015
rect 30915 4895 30960 5015
rect 31080 4895 31125 5015
rect 31245 4895 31290 5015
rect 31410 4895 31465 5015
rect 31585 4895 31630 5015
rect 31750 4895 31795 5015
rect 31915 4895 31960 5015
rect 32080 4895 32135 5015
rect 32255 4895 32300 5015
rect 32420 4895 32465 5015
rect 32585 4895 32630 5015
rect 32750 4895 32805 5015
rect 32925 4895 32970 5015
rect 33090 4895 33135 5015
rect 33255 4895 33300 5015
rect 33420 4895 33475 5015
rect 33595 4895 33640 5015
rect 33760 4895 33805 5015
rect 33925 4895 33970 5015
rect 34090 4895 34145 5015
rect 34265 4895 34310 5015
rect 34430 4895 34475 5015
rect 34595 4895 34640 5015
rect 34760 4895 34815 5015
rect 34935 4895 34980 5015
rect 35100 4895 35145 5015
rect 35265 4895 35310 5015
rect 35430 4895 35485 5015
rect 35605 4895 35650 5015
rect 35770 4895 35815 5015
rect 35935 4895 35980 5015
rect 36100 4895 36155 5015
rect 36275 4895 36485 5015
rect 36605 4895 36650 5015
rect 36770 4895 36815 5015
rect 36935 4895 36980 5015
rect 37100 4895 37155 5015
rect 37275 4895 37320 5015
rect 37440 4895 37485 5015
rect 37605 4895 37650 5015
rect 37770 4895 37825 5015
rect 37945 4895 37990 5015
rect 38110 4895 38155 5015
rect 38275 4895 38320 5015
rect 38440 4895 38495 5015
rect 38615 4895 38660 5015
rect 38780 4895 38825 5015
rect 38945 4895 38990 5015
rect 39110 4895 39165 5015
rect 39285 4895 39330 5015
rect 39450 4895 39495 5015
rect 39615 4895 39660 5015
rect 39780 4895 39835 5015
rect 39955 4895 40000 5015
rect 40120 4895 40165 5015
rect 40285 4895 40330 5015
rect 40450 4895 40505 5015
rect 40625 4895 40670 5015
rect 40790 4895 40835 5015
rect 40955 4895 41000 5015
rect 41120 4895 41175 5015
rect 41295 4895 41340 5015
rect 41460 4895 41505 5015
rect 41625 4895 41670 5015
rect 41790 4895 41845 5015
rect 41965 4895 42175 5015
rect 42295 4895 42340 5015
rect 42460 4895 42505 5015
rect 42625 4895 42670 5015
rect 42790 4895 42845 5015
rect 42965 4895 43010 5015
rect 43130 4895 43175 5015
rect 43295 4895 43340 5015
rect 43460 4895 43515 5015
rect 43635 4895 43680 5015
rect 43800 4895 43845 5015
rect 43965 4895 44010 5015
rect 44130 4895 44185 5015
rect 44305 4895 44350 5015
rect 44470 4895 44515 5015
rect 44635 4895 44680 5015
rect 44800 4895 44855 5015
rect 44975 4895 45020 5015
rect 45140 4895 45185 5015
rect 45305 4895 45350 5015
rect 45470 4895 45525 5015
rect 45645 4895 45690 5015
rect 45810 4895 45855 5015
rect 45975 4895 46020 5015
rect 46140 4895 46195 5015
rect 46315 4895 46360 5015
rect 46480 4895 46525 5015
rect 46645 4895 46690 5015
rect 46810 4895 46865 5015
rect 46985 4895 47030 5015
rect 47150 4895 47195 5015
rect 47315 4895 47360 5015
rect 47480 4895 47535 5015
rect 47655 4895 47865 5015
rect 47985 4895 48030 5015
rect 48150 4895 48195 5015
rect 48315 4895 48360 5015
rect 48480 4895 48535 5015
rect 48655 4895 48700 5015
rect 48820 4895 48865 5015
rect 48985 4895 49030 5015
rect 49150 4895 49205 5015
rect 49325 4895 49370 5015
rect 49490 4895 49535 5015
rect 49655 4895 49700 5015
rect 49820 4895 49875 5015
rect 49995 4895 50040 5015
rect 50160 4895 50205 5015
rect 50325 4895 50370 5015
rect 50490 4895 50545 5015
rect 50665 4895 50710 5015
rect 50830 4895 50875 5015
rect 50995 4895 51040 5015
rect 51160 4895 51215 5015
rect 51335 4895 51380 5015
rect 51500 4895 51545 5015
rect 51665 4895 51710 5015
rect 51830 4895 51885 5015
rect 52005 4895 52050 5015
rect 52170 4895 52215 5015
rect 52335 4895 52380 5015
rect 52500 4895 52555 5015
rect 52675 4895 52720 5015
rect 52840 4895 52885 5015
rect 53005 4895 53050 5015
rect 53170 4895 53225 5015
rect 53345 4895 53370 5015
rect 30770 4850 53370 4895
rect 30770 4730 30795 4850
rect 30915 4730 30960 4850
rect 31080 4730 31125 4850
rect 31245 4730 31290 4850
rect 31410 4730 31465 4850
rect 31585 4730 31630 4850
rect 31750 4730 31795 4850
rect 31915 4730 31960 4850
rect 32080 4730 32135 4850
rect 32255 4730 32300 4850
rect 32420 4730 32465 4850
rect 32585 4730 32630 4850
rect 32750 4730 32805 4850
rect 32925 4730 32970 4850
rect 33090 4730 33135 4850
rect 33255 4730 33300 4850
rect 33420 4730 33475 4850
rect 33595 4730 33640 4850
rect 33760 4730 33805 4850
rect 33925 4730 33970 4850
rect 34090 4730 34145 4850
rect 34265 4730 34310 4850
rect 34430 4730 34475 4850
rect 34595 4730 34640 4850
rect 34760 4730 34815 4850
rect 34935 4730 34980 4850
rect 35100 4730 35145 4850
rect 35265 4730 35310 4850
rect 35430 4730 35485 4850
rect 35605 4730 35650 4850
rect 35770 4730 35815 4850
rect 35935 4730 35980 4850
rect 36100 4730 36155 4850
rect 36275 4730 36485 4850
rect 36605 4730 36650 4850
rect 36770 4730 36815 4850
rect 36935 4730 36980 4850
rect 37100 4730 37155 4850
rect 37275 4730 37320 4850
rect 37440 4730 37485 4850
rect 37605 4730 37650 4850
rect 37770 4730 37825 4850
rect 37945 4730 37990 4850
rect 38110 4730 38155 4850
rect 38275 4730 38320 4850
rect 38440 4730 38495 4850
rect 38615 4730 38660 4850
rect 38780 4730 38825 4850
rect 38945 4730 38990 4850
rect 39110 4730 39165 4850
rect 39285 4730 39330 4850
rect 39450 4730 39495 4850
rect 39615 4730 39660 4850
rect 39780 4730 39835 4850
rect 39955 4730 40000 4850
rect 40120 4730 40165 4850
rect 40285 4730 40330 4850
rect 40450 4730 40505 4850
rect 40625 4730 40670 4850
rect 40790 4730 40835 4850
rect 40955 4730 41000 4850
rect 41120 4730 41175 4850
rect 41295 4730 41340 4850
rect 41460 4730 41505 4850
rect 41625 4730 41670 4850
rect 41790 4730 41845 4850
rect 41965 4730 42175 4850
rect 42295 4730 42340 4850
rect 42460 4730 42505 4850
rect 42625 4730 42670 4850
rect 42790 4730 42845 4850
rect 42965 4730 43010 4850
rect 43130 4730 43175 4850
rect 43295 4730 43340 4850
rect 43460 4730 43515 4850
rect 43635 4730 43680 4850
rect 43800 4730 43845 4850
rect 43965 4730 44010 4850
rect 44130 4730 44185 4850
rect 44305 4730 44350 4850
rect 44470 4730 44515 4850
rect 44635 4730 44680 4850
rect 44800 4730 44855 4850
rect 44975 4730 45020 4850
rect 45140 4730 45185 4850
rect 45305 4730 45350 4850
rect 45470 4730 45525 4850
rect 45645 4730 45690 4850
rect 45810 4730 45855 4850
rect 45975 4730 46020 4850
rect 46140 4730 46195 4850
rect 46315 4730 46360 4850
rect 46480 4730 46525 4850
rect 46645 4730 46690 4850
rect 46810 4730 46865 4850
rect 46985 4730 47030 4850
rect 47150 4730 47195 4850
rect 47315 4730 47360 4850
rect 47480 4730 47535 4850
rect 47655 4730 47865 4850
rect 47985 4730 48030 4850
rect 48150 4730 48195 4850
rect 48315 4730 48360 4850
rect 48480 4730 48535 4850
rect 48655 4730 48700 4850
rect 48820 4730 48865 4850
rect 48985 4730 49030 4850
rect 49150 4730 49205 4850
rect 49325 4730 49370 4850
rect 49490 4730 49535 4850
rect 49655 4730 49700 4850
rect 49820 4730 49875 4850
rect 49995 4730 50040 4850
rect 50160 4730 50205 4850
rect 50325 4730 50370 4850
rect 50490 4730 50545 4850
rect 50665 4730 50710 4850
rect 50830 4730 50875 4850
rect 50995 4730 51040 4850
rect 51160 4730 51215 4850
rect 51335 4730 51380 4850
rect 51500 4730 51545 4850
rect 51665 4730 51710 4850
rect 51830 4730 51885 4850
rect 52005 4730 52050 4850
rect 52170 4730 52215 4850
rect 52335 4730 52380 4850
rect 52500 4730 52555 4850
rect 52675 4730 52720 4850
rect 52840 4730 52885 4850
rect 53005 4730 53050 4850
rect 53170 4730 53225 4850
rect 53345 4730 53370 4850
rect 30770 4685 53370 4730
rect 30770 4625 30795 4685
rect 30530 4565 30795 4625
rect 30915 4565 30960 4685
rect 31080 4565 31125 4685
rect 31245 4565 31290 4685
rect 31410 4565 31465 4685
rect 31585 4565 31630 4685
rect 31750 4565 31795 4685
rect 31915 4565 31960 4685
rect 32080 4565 32135 4685
rect 32255 4565 32300 4685
rect 32420 4565 32465 4685
rect 32585 4565 32630 4685
rect 32750 4565 32805 4685
rect 32925 4565 32970 4685
rect 33090 4565 33135 4685
rect 33255 4565 33300 4685
rect 33420 4565 33475 4685
rect 33595 4565 33640 4685
rect 33760 4565 33805 4685
rect 33925 4565 33970 4685
rect 34090 4565 34145 4685
rect 34265 4565 34310 4685
rect 34430 4565 34475 4685
rect 34595 4565 34640 4685
rect 34760 4565 34815 4685
rect 34935 4565 34980 4685
rect 35100 4565 35145 4685
rect 35265 4565 35310 4685
rect 35430 4565 35485 4685
rect 35605 4565 35650 4685
rect 35770 4565 35815 4685
rect 35935 4565 35980 4685
rect 36100 4565 36155 4685
rect 36275 4565 36485 4685
rect 36605 4565 36650 4685
rect 36770 4565 36815 4685
rect 36935 4565 36980 4685
rect 37100 4565 37155 4685
rect 37275 4565 37320 4685
rect 37440 4565 37485 4685
rect 37605 4565 37650 4685
rect 37770 4565 37825 4685
rect 37945 4565 37990 4685
rect 38110 4565 38155 4685
rect 38275 4565 38320 4685
rect 38440 4565 38495 4685
rect 38615 4565 38660 4685
rect 38780 4565 38825 4685
rect 38945 4565 38990 4685
rect 39110 4565 39165 4685
rect 39285 4565 39330 4685
rect 39450 4565 39495 4685
rect 39615 4565 39660 4685
rect 39780 4565 39835 4685
rect 39955 4565 40000 4685
rect 40120 4565 40165 4685
rect 40285 4565 40330 4685
rect 40450 4565 40505 4685
rect 40625 4565 40670 4685
rect 40790 4565 40835 4685
rect 40955 4565 41000 4685
rect 41120 4565 41175 4685
rect 41295 4565 41340 4685
rect 41460 4565 41505 4685
rect 41625 4565 41670 4685
rect 41790 4565 41845 4685
rect 41965 4565 42175 4685
rect 42295 4565 42340 4685
rect 42460 4565 42505 4685
rect 42625 4565 42670 4685
rect 42790 4565 42845 4685
rect 42965 4565 43010 4685
rect 43130 4565 43175 4685
rect 43295 4565 43340 4685
rect 43460 4565 43515 4685
rect 43635 4565 43680 4685
rect 43800 4565 43845 4685
rect 43965 4565 44010 4685
rect 44130 4565 44185 4685
rect 44305 4565 44350 4685
rect 44470 4565 44515 4685
rect 44635 4565 44680 4685
rect 44800 4565 44855 4685
rect 44975 4565 45020 4685
rect 45140 4565 45185 4685
rect 45305 4565 45350 4685
rect 45470 4565 45525 4685
rect 45645 4565 45690 4685
rect 45810 4565 45855 4685
rect 45975 4565 46020 4685
rect 46140 4565 46195 4685
rect 46315 4565 46360 4685
rect 46480 4565 46525 4685
rect 46645 4565 46690 4685
rect 46810 4565 46865 4685
rect 46985 4565 47030 4685
rect 47150 4565 47195 4685
rect 47315 4565 47360 4685
rect 47480 4565 47535 4685
rect 47655 4565 47865 4685
rect 47985 4565 48030 4685
rect 48150 4565 48195 4685
rect 48315 4565 48360 4685
rect 48480 4565 48535 4685
rect 48655 4565 48700 4685
rect 48820 4565 48865 4685
rect 48985 4565 49030 4685
rect 49150 4565 49205 4685
rect 49325 4565 49370 4685
rect 49490 4565 49535 4685
rect 49655 4565 49700 4685
rect 49820 4565 49875 4685
rect 49995 4565 50040 4685
rect 50160 4565 50205 4685
rect 50325 4565 50370 4685
rect 50490 4565 50545 4685
rect 50665 4565 50710 4685
rect 50830 4565 50875 4685
rect 50995 4565 51040 4685
rect 51160 4565 51215 4685
rect 51335 4565 51380 4685
rect 51500 4565 51545 4685
rect 51665 4565 51710 4685
rect 51830 4565 51885 4685
rect 52005 4565 52050 4685
rect 52170 4565 52215 4685
rect 52335 4565 52380 4685
rect 52500 4565 52555 4685
rect 52675 4565 52720 4685
rect 52840 4565 52885 4685
rect 53005 4565 53050 4685
rect 53170 4565 53225 4685
rect 53345 4565 53370 4685
rect 30530 4520 53370 4565
rect 30530 4400 30795 4520
rect 30915 4400 30960 4520
rect 31080 4400 31125 4520
rect 31245 4400 31290 4520
rect 31410 4400 31465 4520
rect 31585 4400 31630 4520
rect 31750 4400 31795 4520
rect 31915 4400 31960 4520
rect 32080 4400 32135 4520
rect 32255 4400 32300 4520
rect 32420 4400 32465 4520
rect 32585 4400 32630 4520
rect 32750 4400 32805 4520
rect 32925 4400 32970 4520
rect 33090 4400 33135 4520
rect 33255 4400 33300 4520
rect 33420 4400 33475 4520
rect 33595 4400 33640 4520
rect 33760 4400 33805 4520
rect 33925 4400 33970 4520
rect 34090 4400 34145 4520
rect 34265 4400 34310 4520
rect 34430 4400 34475 4520
rect 34595 4400 34640 4520
rect 34760 4400 34815 4520
rect 34935 4400 34980 4520
rect 35100 4400 35145 4520
rect 35265 4400 35310 4520
rect 35430 4400 35485 4520
rect 35605 4400 35650 4520
rect 35770 4400 35815 4520
rect 35935 4400 35980 4520
rect 36100 4400 36155 4520
rect 36275 4400 36485 4520
rect 36605 4400 36650 4520
rect 36770 4400 36815 4520
rect 36935 4400 36980 4520
rect 37100 4400 37155 4520
rect 37275 4400 37320 4520
rect 37440 4400 37485 4520
rect 37605 4400 37650 4520
rect 37770 4400 37825 4520
rect 37945 4400 37990 4520
rect 38110 4400 38155 4520
rect 38275 4400 38320 4520
rect 38440 4400 38495 4520
rect 38615 4400 38660 4520
rect 38780 4400 38825 4520
rect 38945 4400 38990 4520
rect 39110 4400 39165 4520
rect 39285 4400 39330 4520
rect 39450 4400 39495 4520
rect 39615 4400 39660 4520
rect 39780 4400 39835 4520
rect 39955 4400 40000 4520
rect 40120 4400 40165 4520
rect 40285 4400 40330 4520
rect 40450 4400 40505 4520
rect 40625 4400 40670 4520
rect 40790 4400 40835 4520
rect 40955 4400 41000 4520
rect 41120 4400 41175 4520
rect 41295 4400 41340 4520
rect 41460 4400 41505 4520
rect 41625 4400 41670 4520
rect 41790 4400 41845 4520
rect 41965 4400 42175 4520
rect 42295 4400 42340 4520
rect 42460 4400 42505 4520
rect 42625 4400 42670 4520
rect 42790 4400 42845 4520
rect 42965 4400 43010 4520
rect 43130 4400 43175 4520
rect 43295 4400 43340 4520
rect 43460 4400 43515 4520
rect 43635 4400 43680 4520
rect 43800 4400 43845 4520
rect 43965 4400 44010 4520
rect 44130 4400 44185 4520
rect 44305 4400 44350 4520
rect 44470 4400 44515 4520
rect 44635 4400 44680 4520
rect 44800 4400 44855 4520
rect 44975 4400 45020 4520
rect 45140 4400 45185 4520
rect 45305 4400 45350 4520
rect 45470 4400 45525 4520
rect 45645 4400 45690 4520
rect 45810 4400 45855 4520
rect 45975 4400 46020 4520
rect 46140 4400 46195 4520
rect 46315 4400 46360 4520
rect 46480 4400 46525 4520
rect 46645 4400 46690 4520
rect 46810 4400 46865 4520
rect 46985 4400 47030 4520
rect 47150 4400 47195 4520
rect 47315 4400 47360 4520
rect 47480 4400 47535 4520
rect 47655 4400 47865 4520
rect 47985 4400 48030 4520
rect 48150 4400 48195 4520
rect 48315 4400 48360 4520
rect 48480 4400 48535 4520
rect 48655 4400 48700 4520
rect 48820 4400 48865 4520
rect 48985 4400 49030 4520
rect 49150 4400 49205 4520
rect 49325 4400 49370 4520
rect 49490 4400 49535 4520
rect 49655 4400 49700 4520
rect 49820 4400 49875 4520
rect 49995 4400 50040 4520
rect 50160 4400 50205 4520
rect 50325 4400 50370 4520
rect 50490 4400 50545 4520
rect 50665 4400 50710 4520
rect 50830 4400 50875 4520
rect 50995 4400 51040 4520
rect 51160 4400 51215 4520
rect 51335 4400 51380 4520
rect 51500 4400 51545 4520
rect 51665 4400 51710 4520
rect 51830 4400 51885 4520
rect 52005 4400 52050 4520
rect 52170 4400 52215 4520
rect 52335 4400 52380 4520
rect 52500 4400 52555 4520
rect 52675 4400 52720 4520
rect 52840 4400 52885 4520
rect 53005 4400 53050 4520
rect 53170 4400 53225 4520
rect 53345 4400 53370 4520
rect 30530 4345 53370 4400
rect 30530 4270 30795 4345
rect 30770 4225 30795 4270
rect 30915 4225 30960 4345
rect 31080 4225 31125 4345
rect 31245 4225 31290 4345
rect 31410 4225 31465 4345
rect 31585 4225 31630 4345
rect 31750 4225 31795 4345
rect 31915 4225 31960 4345
rect 32080 4225 32135 4345
rect 32255 4225 32300 4345
rect 32420 4225 32465 4345
rect 32585 4225 32630 4345
rect 32750 4225 32805 4345
rect 32925 4225 32970 4345
rect 33090 4225 33135 4345
rect 33255 4225 33300 4345
rect 33420 4225 33475 4345
rect 33595 4225 33640 4345
rect 33760 4225 33805 4345
rect 33925 4225 33970 4345
rect 34090 4225 34145 4345
rect 34265 4225 34310 4345
rect 34430 4225 34475 4345
rect 34595 4225 34640 4345
rect 34760 4225 34815 4345
rect 34935 4225 34980 4345
rect 35100 4225 35145 4345
rect 35265 4225 35310 4345
rect 35430 4225 35485 4345
rect 35605 4225 35650 4345
rect 35770 4225 35815 4345
rect 35935 4225 35980 4345
rect 36100 4225 36155 4345
rect 36275 4225 36485 4345
rect 36605 4225 36650 4345
rect 36770 4225 36815 4345
rect 36935 4225 36980 4345
rect 37100 4225 37155 4345
rect 37275 4225 37320 4345
rect 37440 4225 37485 4345
rect 37605 4225 37650 4345
rect 37770 4225 37825 4345
rect 37945 4225 37990 4345
rect 38110 4225 38155 4345
rect 38275 4225 38320 4345
rect 38440 4225 38495 4345
rect 38615 4225 38660 4345
rect 38780 4225 38825 4345
rect 38945 4225 38990 4345
rect 39110 4225 39165 4345
rect 39285 4225 39330 4345
rect 39450 4225 39495 4345
rect 39615 4225 39660 4345
rect 39780 4225 39835 4345
rect 39955 4225 40000 4345
rect 40120 4225 40165 4345
rect 40285 4225 40330 4345
rect 40450 4225 40505 4345
rect 40625 4225 40670 4345
rect 40790 4225 40835 4345
rect 40955 4225 41000 4345
rect 41120 4225 41175 4345
rect 41295 4225 41340 4345
rect 41460 4225 41505 4345
rect 41625 4225 41670 4345
rect 41790 4225 41845 4345
rect 41965 4225 42175 4345
rect 42295 4225 42340 4345
rect 42460 4225 42505 4345
rect 42625 4225 42670 4345
rect 42790 4225 42845 4345
rect 42965 4225 43010 4345
rect 43130 4225 43175 4345
rect 43295 4225 43340 4345
rect 43460 4225 43515 4345
rect 43635 4225 43680 4345
rect 43800 4225 43845 4345
rect 43965 4225 44010 4345
rect 44130 4225 44185 4345
rect 44305 4225 44350 4345
rect 44470 4225 44515 4345
rect 44635 4225 44680 4345
rect 44800 4225 44855 4345
rect 44975 4225 45020 4345
rect 45140 4225 45185 4345
rect 45305 4225 45350 4345
rect 45470 4225 45525 4345
rect 45645 4225 45690 4345
rect 45810 4225 45855 4345
rect 45975 4225 46020 4345
rect 46140 4225 46195 4345
rect 46315 4225 46360 4345
rect 46480 4225 46525 4345
rect 46645 4225 46690 4345
rect 46810 4225 46865 4345
rect 46985 4225 47030 4345
rect 47150 4225 47195 4345
rect 47315 4225 47360 4345
rect 47480 4225 47535 4345
rect 47655 4225 47865 4345
rect 47985 4225 48030 4345
rect 48150 4225 48195 4345
rect 48315 4225 48360 4345
rect 48480 4225 48535 4345
rect 48655 4225 48700 4345
rect 48820 4225 48865 4345
rect 48985 4225 49030 4345
rect 49150 4225 49205 4345
rect 49325 4225 49370 4345
rect 49490 4225 49535 4345
rect 49655 4225 49700 4345
rect 49820 4225 49875 4345
rect 49995 4225 50040 4345
rect 50160 4225 50205 4345
rect 50325 4225 50370 4345
rect 50490 4225 50545 4345
rect 50665 4225 50710 4345
rect 50830 4225 50875 4345
rect 50995 4225 51040 4345
rect 51160 4225 51215 4345
rect 51335 4225 51380 4345
rect 51500 4225 51545 4345
rect 51665 4225 51710 4345
rect 51830 4225 51885 4345
rect 52005 4225 52050 4345
rect 52170 4225 52215 4345
rect 52335 4225 52380 4345
rect 52500 4225 52555 4345
rect 52675 4225 52720 4345
rect 52840 4225 52885 4345
rect 53005 4225 53050 4345
rect 53170 4225 53225 4345
rect 53345 4225 53370 4345
rect 30770 4180 53370 4225
rect 30770 4060 30795 4180
rect 30915 4060 30960 4180
rect 31080 4060 31125 4180
rect 31245 4060 31290 4180
rect 31410 4060 31465 4180
rect 31585 4060 31630 4180
rect 31750 4060 31795 4180
rect 31915 4060 31960 4180
rect 32080 4060 32135 4180
rect 32255 4060 32300 4180
rect 32420 4060 32465 4180
rect 32585 4060 32630 4180
rect 32750 4060 32805 4180
rect 32925 4060 32970 4180
rect 33090 4060 33135 4180
rect 33255 4060 33300 4180
rect 33420 4060 33475 4180
rect 33595 4060 33640 4180
rect 33760 4060 33805 4180
rect 33925 4060 33970 4180
rect 34090 4060 34145 4180
rect 34265 4060 34310 4180
rect 34430 4060 34475 4180
rect 34595 4060 34640 4180
rect 34760 4060 34815 4180
rect 34935 4060 34980 4180
rect 35100 4060 35145 4180
rect 35265 4060 35310 4180
rect 35430 4060 35485 4180
rect 35605 4060 35650 4180
rect 35770 4060 35815 4180
rect 35935 4060 35980 4180
rect 36100 4060 36155 4180
rect 36275 4060 36485 4180
rect 36605 4060 36650 4180
rect 36770 4060 36815 4180
rect 36935 4060 36980 4180
rect 37100 4060 37155 4180
rect 37275 4060 37320 4180
rect 37440 4060 37485 4180
rect 37605 4060 37650 4180
rect 37770 4060 37825 4180
rect 37945 4060 37990 4180
rect 38110 4060 38155 4180
rect 38275 4060 38320 4180
rect 38440 4060 38495 4180
rect 38615 4060 38660 4180
rect 38780 4060 38825 4180
rect 38945 4060 38990 4180
rect 39110 4060 39165 4180
rect 39285 4060 39330 4180
rect 39450 4060 39495 4180
rect 39615 4060 39660 4180
rect 39780 4060 39835 4180
rect 39955 4060 40000 4180
rect 40120 4060 40165 4180
rect 40285 4060 40330 4180
rect 40450 4060 40505 4180
rect 40625 4060 40670 4180
rect 40790 4060 40835 4180
rect 40955 4060 41000 4180
rect 41120 4060 41175 4180
rect 41295 4060 41340 4180
rect 41460 4060 41505 4180
rect 41625 4060 41670 4180
rect 41790 4060 41845 4180
rect 41965 4060 42175 4180
rect 42295 4060 42340 4180
rect 42460 4060 42505 4180
rect 42625 4060 42670 4180
rect 42790 4060 42845 4180
rect 42965 4060 43010 4180
rect 43130 4060 43175 4180
rect 43295 4060 43340 4180
rect 43460 4060 43515 4180
rect 43635 4060 43680 4180
rect 43800 4060 43845 4180
rect 43965 4060 44010 4180
rect 44130 4060 44185 4180
rect 44305 4060 44350 4180
rect 44470 4060 44515 4180
rect 44635 4060 44680 4180
rect 44800 4060 44855 4180
rect 44975 4060 45020 4180
rect 45140 4060 45185 4180
rect 45305 4060 45350 4180
rect 45470 4060 45525 4180
rect 45645 4060 45690 4180
rect 45810 4060 45855 4180
rect 45975 4060 46020 4180
rect 46140 4060 46195 4180
rect 46315 4060 46360 4180
rect 46480 4060 46525 4180
rect 46645 4060 46690 4180
rect 46810 4060 46865 4180
rect 46985 4060 47030 4180
rect 47150 4060 47195 4180
rect 47315 4060 47360 4180
rect 47480 4060 47535 4180
rect 47655 4060 47865 4180
rect 47985 4060 48030 4180
rect 48150 4060 48195 4180
rect 48315 4060 48360 4180
rect 48480 4060 48535 4180
rect 48655 4060 48700 4180
rect 48820 4060 48865 4180
rect 48985 4060 49030 4180
rect 49150 4060 49205 4180
rect 49325 4060 49370 4180
rect 49490 4060 49535 4180
rect 49655 4060 49700 4180
rect 49820 4060 49875 4180
rect 49995 4060 50040 4180
rect 50160 4060 50205 4180
rect 50325 4060 50370 4180
rect 50490 4060 50545 4180
rect 50665 4060 50710 4180
rect 50830 4060 50875 4180
rect 50995 4060 51040 4180
rect 51160 4060 51215 4180
rect 51335 4060 51380 4180
rect 51500 4060 51545 4180
rect 51665 4060 51710 4180
rect 51830 4060 51885 4180
rect 52005 4060 52050 4180
rect 52170 4060 52215 4180
rect 52335 4060 52380 4180
rect 52500 4060 52555 4180
rect 52675 4060 52720 4180
rect 52840 4060 52885 4180
rect 53005 4060 53050 4180
rect 53170 4060 53225 4180
rect 53345 4060 53370 4180
rect 30770 4015 53370 4060
rect 30770 3895 30795 4015
rect 30915 3895 30960 4015
rect 31080 3895 31125 4015
rect 31245 3895 31290 4015
rect 31410 3895 31465 4015
rect 31585 3895 31630 4015
rect 31750 3895 31795 4015
rect 31915 3895 31960 4015
rect 32080 3895 32135 4015
rect 32255 3895 32300 4015
rect 32420 3895 32465 4015
rect 32585 3895 32630 4015
rect 32750 3895 32805 4015
rect 32925 3895 32970 4015
rect 33090 3895 33135 4015
rect 33255 3895 33300 4015
rect 33420 3895 33475 4015
rect 33595 3895 33640 4015
rect 33760 3895 33805 4015
rect 33925 3895 33970 4015
rect 34090 3895 34145 4015
rect 34265 3895 34310 4015
rect 34430 3895 34475 4015
rect 34595 3895 34640 4015
rect 34760 3895 34815 4015
rect 34935 3895 34980 4015
rect 35100 3895 35145 4015
rect 35265 3895 35310 4015
rect 35430 3895 35485 4015
rect 35605 3895 35650 4015
rect 35770 3895 35815 4015
rect 35935 3895 35980 4015
rect 36100 3895 36155 4015
rect 36275 3895 36485 4015
rect 36605 3895 36650 4015
rect 36770 3895 36815 4015
rect 36935 3895 36980 4015
rect 37100 3895 37155 4015
rect 37275 3895 37320 4015
rect 37440 3895 37485 4015
rect 37605 3895 37650 4015
rect 37770 3895 37825 4015
rect 37945 3895 37990 4015
rect 38110 3895 38155 4015
rect 38275 3895 38320 4015
rect 38440 3895 38495 4015
rect 38615 3895 38660 4015
rect 38780 3895 38825 4015
rect 38945 3895 38990 4015
rect 39110 3895 39165 4015
rect 39285 3895 39330 4015
rect 39450 3895 39495 4015
rect 39615 3895 39660 4015
rect 39780 3895 39835 4015
rect 39955 3895 40000 4015
rect 40120 3895 40165 4015
rect 40285 3895 40330 4015
rect 40450 3895 40505 4015
rect 40625 3895 40670 4015
rect 40790 3895 40835 4015
rect 40955 3895 41000 4015
rect 41120 3895 41175 4015
rect 41295 3895 41340 4015
rect 41460 3895 41505 4015
rect 41625 3895 41670 4015
rect 41790 3895 41845 4015
rect 41965 3895 42175 4015
rect 42295 3895 42340 4015
rect 42460 3895 42505 4015
rect 42625 3895 42670 4015
rect 42790 3895 42845 4015
rect 42965 3895 43010 4015
rect 43130 3895 43175 4015
rect 43295 3895 43340 4015
rect 43460 3895 43515 4015
rect 43635 3895 43680 4015
rect 43800 3895 43845 4015
rect 43965 3895 44010 4015
rect 44130 3895 44185 4015
rect 44305 3895 44350 4015
rect 44470 3895 44515 4015
rect 44635 3895 44680 4015
rect 44800 3895 44855 4015
rect 44975 3895 45020 4015
rect 45140 3895 45185 4015
rect 45305 3895 45350 4015
rect 45470 3895 45525 4015
rect 45645 3895 45690 4015
rect 45810 3895 45855 4015
rect 45975 3895 46020 4015
rect 46140 3895 46195 4015
rect 46315 3895 46360 4015
rect 46480 3895 46525 4015
rect 46645 3895 46690 4015
rect 46810 3895 46865 4015
rect 46985 3895 47030 4015
rect 47150 3895 47195 4015
rect 47315 3895 47360 4015
rect 47480 3895 47535 4015
rect 47655 3895 47865 4015
rect 47985 3895 48030 4015
rect 48150 3895 48195 4015
rect 48315 3895 48360 4015
rect 48480 3895 48535 4015
rect 48655 3895 48700 4015
rect 48820 3895 48865 4015
rect 48985 3895 49030 4015
rect 49150 3895 49205 4015
rect 49325 3895 49370 4015
rect 49490 3895 49535 4015
rect 49655 3895 49700 4015
rect 49820 3895 49875 4015
rect 49995 3895 50040 4015
rect 50160 3895 50205 4015
rect 50325 3895 50370 4015
rect 50490 3895 50545 4015
rect 50665 3895 50710 4015
rect 50830 3895 50875 4015
rect 50995 3895 51040 4015
rect 51160 3895 51215 4015
rect 51335 3895 51380 4015
rect 51500 3895 51545 4015
rect 51665 3895 51710 4015
rect 51830 3895 51885 4015
rect 52005 3895 52050 4015
rect 52170 3895 52215 4015
rect 52335 3895 52380 4015
rect 52500 3895 52555 4015
rect 52675 3895 52720 4015
rect 52840 3895 52885 4015
rect 53005 3895 53050 4015
rect 53170 3895 53225 4015
rect 53345 3895 53370 4015
rect 30770 3850 53370 3895
rect 30770 3730 30795 3850
rect 30915 3730 30960 3850
rect 31080 3730 31125 3850
rect 31245 3730 31290 3850
rect 31410 3730 31465 3850
rect 31585 3730 31630 3850
rect 31750 3730 31795 3850
rect 31915 3730 31960 3850
rect 32080 3730 32135 3850
rect 32255 3730 32300 3850
rect 32420 3730 32465 3850
rect 32585 3730 32630 3850
rect 32750 3730 32805 3850
rect 32925 3730 32970 3850
rect 33090 3730 33135 3850
rect 33255 3730 33300 3850
rect 33420 3730 33475 3850
rect 33595 3730 33640 3850
rect 33760 3730 33805 3850
rect 33925 3730 33970 3850
rect 34090 3730 34145 3850
rect 34265 3730 34310 3850
rect 34430 3730 34475 3850
rect 34595 3730 34640 3850
rect 34760 3730 34815 3850
rect 34935 3730 34980 3850
rect 35100 3730 35145 3850
rect 35265 3730 35310 3850
rect 35430 3730 35485 3850
rect 35605 3730 35650 3850
rect 35770 3730 35815 3850
rect 35935 3730 35980 3850
rect 36100 3730 36155 3850
rect 36275 3730 36485 3850
rect 36605 3730 36650 3850
rect 36770 3730 36815 3850
rect 36935 3730 36980 3850
rect 37100 3730 37155 3850
rect 37275 3730 37320 3850
rect 37440 3730 37485 3850
rect 37605 3730 37650 3850
rect 37770 3730 37825 3850
rect 37945 3730 37990 3850
rect 38110 3730 38155 3850
rect 38275 3730 38320 3850
rect 38440 3730 38495 3850
rect 38615 3730 38660 3850
rect 38780 3730 38825 3850
rect 38945 3730 38990 3850
rect 39110 3730 39165 3850
rect 39285 3730 39330 3850
rect 39450 3730 39495 3850
rect 39615 3730 39660 3850
rect 39780 3730 39835 3850
rect 39955 3730 40000 3850
rect 40120 3730 40165 3850
rect 40285 3730 40330 3850
rect 40450 3730 40505 3850
rect 40625 3730 40670 3850
rect 40790 3730 40835 3850
rect 40955 3730 41000 3850
rect 41120 3730 41175 3850
rect 41295 3730 41340 3850
rect 41460 3730 41505 3850
rect 41625 3730 41670 3850
rect 41790 3730 41845 3850
rect 41965 3730 42175 3850
rect 42295 3730 42340 3850
rect 42460 3730 42505 3850
rect 42625 3730 42670 3850
rect 42790 3730 42845 3850
rect 42965 3730 43010 3850
rect 43130 3730 43175 3850
rect 43295 3730 43340 3850
rect 43460 3730 43515 3850
rect 43635 3730 43680 3850
rect 43800 3730 43845 3850
rect 43965 3730 44010 3850
rect 44130 3730 44185 3850
rect 44305 3730 44350 3850
rect 44470 3730 44515 3850
rect 44635 3730 44680 3850
rect 44800 3730 44855 3850
rect 44975 3730 45020 3850
rect 45140 3730 45185 3850
rect 45305 3730 45350 3850
rect 45470 3730 45525 3850
rect 45645 3730 45690 3850
rect 45810 3730 45855 3850
rect 45975 3730 46020 3850
rect 46140 3730 46195 3850
rect 46315 3730 46360 3850
rect 46480 3730 46525 3850
rect 46645 3730 46690 3850
rect 46810 3730 46865 3850
rect 46985 3730 47030 3850
rect 47150 3730 47195 3850
rect 47315 3730 47360 3850
rect 47480 3730 47535 3850
rect 47655 3730 47865 3850
rect 47985 3730 48030 3850
rect 48150 3730 48195 3850
rect 48315 3730 48360 3850
rect 48480 3730 48535 3850
rect 48655 3730 48700 3850
rect 48820 3730 48865 3850
rect 48985 3730 49030 3850
rect 49150 3730 49205 3850
rect 49325 3730 49370 3850
rect 49490 3730 49535 3850
rect 49655 3730 49700 3850
rect 49820 3730 49875 3850
rect 49995 3730 50040 3850
rect 50160 3730 50205 3850
rect 50325 3730 50370 3850
rect 50490 3730 50545 3850
rect 50665 3730 50710 3850
rect 50830 3730 50875 3850
rect 50995 3730 51040 3850
rect 51160 3730 51215 3850
rect 51335 3730 51380 3850
rect 51500 3730 51545 3850
rect 51665 3730 51710 3850
rect 51830 3730 51885 3850
rect 52005 3730 52050 3850
rect 52170 3730 52215 3850
rect 52335 3730 52380 3850
rect 52500 3730 52555 3850
rect 52675 3730 52720 3850
rect 52840 3730 52885 3850
rect 53005 3730 53050 3850
rect 53170 3730 53225 3850
rect 53345 3730 53370 3850
rect 30770 3675 53370 3730
rect 30770 3555 30795 3675
rect 30915 3555 30960 3675
rect 31080 3555 31125 3675
rect 31245 3555 31290 3675
rect 31410 3555 31465 3675
rect 31585 3555 31630 3675
rect 31750 3555 31795 3675
rect 31915 3555 31960 3675
rect 32080 3555 32135 3675
rect 32255 3555 32300 3675
rect 32420 3555 32465 3675
rect 32585 3555 32630 3675
rect 32750 3555 32805 3675
rect 32925 3555 32970 3675
rect 33090 3555 33135 3675
rect 33255 3555 33300 3675
rect 33420 3555 33475 3675
rect 33595 3555 33640 3675
rect 33760 3555 33805 3675
rect 33925 3555 33970 3675
rect 34090 3555 34145 3675
rect 34265 3555 34310 3675
rect 34430 3555 34475 3675
rect 34595 3555 34640 3675
rect 34760 3555 34815 3675
rect 34935 3555 34980 3675
rect 35100 3555 35145 3675
rect 35265 3555 35310 3675
rect 35430 3555 35485 3675
rect 35605 3555 35650 3675
rect 35770 3555 35815 3675
rect 35935 3555 35980 3675
rect 36100 3555 36155 3675
rect 36275 3555 36485 3675
rect 36605 3555 36650 3675
rect 36770 3555 36815 3675
rect 36935 3555 36980 3675
rect 37100 3555 37155 3675
rect 37275 3555 37320 3675
rect 37440 3555 37485 3675
rect 37605 3555 37650 3675
rect 37770 3555 37825 3675
rect 37945 3555 37990 3675
rect 38110 3555 38155 3675
rect 38275 3555 38320 3675
rect 38440 3555 38495 3675
rect 38615 3555 38660 3675
rect 38780 3555 38825 3675
rect 38945 3555 38990 3675
rect 39110 3555 39165 3675
rect 39285 3555 39330 3675
rect 39450 3555 39495 3675
rect 39615 3555 39660 3675
rect 39780 3555 39835 3675
rect 39955 3555 40000 3675
rect 40120 3555 40165 3675
rect 40285 3555 40330 3675
rect 40450 3555 40505 3675
rect 40625 3555 40670 3675
rect 40790 3555 40835 3675
rect 40955 3555 41000 3675
rect 41120 3555 41175 3675
rect 41295 3555 41340 3675
rect 41460 3555 41505 3675
rect 41625 3555 41670 3675
rect 41790 3555 41845 3675
rect 41965 3555 42175 3675
rect 42295 3555 42340 3675
rect 42460 3555 42505 3675
rect 42625 3555 42670 3675
rect 42790 3555 42845 3675
rect 42965 3555 43010 3675
rect 43130 3555 43175 3675
rect 43295 3555 43340 3675
rect 43460 3555 43515 3675
rect 43635 3555 43680 3675
rect 43800 3555 43845 3675
rect 43965 3555 44010 3675
rect 44130 3555 44185 3675
rect 44305 3555 44350 3675
rect 44470 3555 44515 3675
rect 44635 3555 44680 3675
rect 44800 3555 44855 3675
rect 44975 3555 45020 3675
rect 45140 3555 45185 3675
rect 45305 3555 45350 3675
rect 45470 3555 45525 3675
rect 45645 3555 45690 3675
rect 45810 3555 45855 3675
rect 45975 3555 46020 3675
rect 46140 3555 46195 3675
rect 46315 3555 46360 3675
rect 46480 3555 46525 3675
rect 46645 3555 46690 3675
rect 46810 3555 46865 3675
rect 46985 3555 47030 3675
rect 47150 3555 47195 3675
rect 47315 3555 47360 3675
rect 47480 3555 47535 3675
rect 47655 3555 47865 3675
rect 47985 3555 48030 3675
rect 48150 3555 48195 3675
rect 48315 3555 48360 3675
rect 48480 3555 48535 3675
rect 48655 3555 48700 3675
rect 48820 3555 48865 3675
rect 48985 3555 49030 3675
rect 49150 3555 49205 3675
rect 49325 3555 49370 3675
rect 49490 3555 49535 3675
rect 49655 3555 49700 3675
rect 49820 3555 49875 3675
rect 49995 3555 50040 3675
rect 50160 3555 50205 3675
rect 50325 3555 50370 3675
rect 50490 3555 50545 3675
rect 50665 3555 50710 3675
rect 50830 3555 50875 3675
rect 50995 3555 51040 3675
rect 51160 3555 51215 3675
rect 51335 3555 51380 3675
rect 51500 3555 51545 3675
rect 51665 3555 51710 3675
rect 51830 3555 51885 3675
rect 52005 3555 52050 3675
rect 52170 3555 52215 3675
rect 52335 3555 52380 3675
rect 52500 3555 52555 3675
rect 52675 3555 52720 3675
rect 52840 3555 52885 3675
rect 53005 3555 53050 3675
rect 53170 3555 53225 3675
rect 53345 3555 53370 3675
rect 30770 3510 53370 3555
rect 30770 3390 30795 3510
rect 30915 3390 30960 3510
rect 31080 3390 31125 3510
rect 31245 3390 31290 3510
rect 31410 3390 31465 3510
rect 31585 3390 31630 3510
rect 31750 3390 31795 3510
rect 31915 3390 31960 3510
rect 32080 3390 32135 3510
rect 32255 3390 32300 3510
rect 32420 3390 32465 3510
rect 32585 3390 32630 3510
rect 32750 3390 32805 3510
rect 32925 3390 32970 3510
rect 33090 3390 33135 3510
rect 33255 3390 33300 3510
rect 33420 3390 33475 3510
rect 33595 3390 33640 3510
rect 33760 3390 33805 3510
rect 33925 3390 33970 3510
rect 34090 3390 34145 3510
rect 34265 3390 34310 3510
rect 34430 3390 34475 3510
rect 34595 3390 34640 3510
rect 34760 3390 34815 3510
rect 34935 3390 34980 3510
rect 35100 3390 35145 3510
rect 35265 3390 35310 3510
rect 35430 3390 35485 3510
rect 35605 3390 35650 3510
rect 35770 3390 35815 3510
rect 35935 3390 35980 3510
rect 36100 3390 36155 3510
rect 36275 3390 36485 3510
rect 36605 3390 36650 3510
rect 36770 3390 36815 3510
rect 36935 3390 36980 3510
rect 37100 3390 37155 3510
rect 37275 3390 37320 3510
rect 37440 3390 37485 3510
rect 37605 3390 37650 3510
rect 37770 3390 37825 3510
rect 37945 3390 37990 3510
rect 38110 3390 38155 3510
rect 38275 3390 38320 3510
rect 38440 3390 38495 3510
rect 38615 3390 38660 3510
rect 38780 3390 38825 3510
rect 38945 3390 38990 3510
rect 39110 3390 39165 3510
rect 39285 3390 39330 3510
rect 39450 3390 39495 3510
rect 39615 3390 39660 3510
rect 39780 3390 39835 3510
rect 39955 3390 40000 3510
rect 40120 3390 40165 3510
rect 40285 3390 40330 3510
rect 40450 3390 40505 3510
rect 40625 3390 40670 3510
rect 40790 3390 40835 3510
rect 40955 3390 41000 3510
rect 41120 3390 41175 3510
rect 41295 3390 41340 3510
rect 41460 3390 41505 3510
rect 41625 3390 41670 3510
rect 41790 3390 41845 3510
rect 41965 3390 42175 3510
rect 42295 3390 42340 3510
rect 42460 3390 42505 3510
rect 42625 3390 42670 3510
rect 42790 3390 42845 3510
rect 42965 3390 43010 3510
rect 43130 3390 43175 3510
rect 43295 3390 43340 3510
rect 43460 3390 43515 3510
rect 43635 3390 43680 3510
rect 43800 3390 43845 3510
rect 43965 3390 44010 3510
rect 44130 3390 44185 3510
rect 44305 3390 44350 3510
rect 44470 3390 44515 3510
rect 44635 3390 44680 3510
rect 44800 3390 44855 3510
rect 44975 3390 45020 3510
rect 45140 3390 45185 3510
rect 45305 3390 45350 3510
rect 45470 3390 45525 3510
rect 45645 3390 45690 3510
rect 45810 3390 45855 3510
rect 45975 3390 46020 3510
rect 46140 3390 46195 3510
rect 46315 3390 46360 3510
rect 46480 3390 46525 3510
rect 46645 3390 46690 3510
rect 46810 3390 46865 3510
rect 46985 3390 47030 3510
rect 47150 3390 47195 3510
rect 47315 3390 47360 3510
rect 47480 3390 47535 3510
rect 47655 3390 47865 3510
rect 47985 3390 48030 3510
rect 48150 3390 48195 3510
rect 48315 3390 48360 3510
rect 48480 3390 48535 3510
rect 48655 3390 48700 3510
rect 48820 3390 48865 3510
rect 48985 3390 49030 3510
rect 49150 3390 49205 3510
rect 49325 3390 49370 3510
rect 49490 3390 49535 3510
rect 49655 3390 49700 3510
rect 49820 3390 49875 3510
rect 49995 3390 50040 3510
rect 50160 3390 50205 3510
rect 50325 3390 50370 3510
rect 50490 3390 50545 3510
rect 50665 3390 50710 3510
rect 50830 3390 50875 3510
rect 50995 3390 51040 3510
rect 51160 3390 51215 3510
rect 51335 3390 51380 3510
rect 51500 3390 51545 3510
rect 51665 3390 51710 3510
rect 51830 3390 51885 3510
rect 52005 3390 52050 3510
rect 52170 3390 52215 3510
rect 52335 3390 52380 3510
rect 52500 3390 52555 3510
rect 52675 3390 52720 3510
rect 52840 3390 52885 3510
rect 53005 3390 53050 3510
rect 53170 3390 53225 3510
rect 53345 3390 53370 3510
rect 30770 3345 53370 3390
rect 30770 3225 30795 3345
rect 30915 3225 30960 3345
rect 31080 3225 31125 3345
rect 31245 3225 31290 3345
rect 31410 3225 31465 3345
rect 31585 3225 31630 3345
rect 31750 3225 31795 3345
rect 31915 3225 31960 3345
rect 32080 3225 32135 3345
rect 32255 3225 32300 3345
rect 32420 3225 32465 3345
rect 32585 3225 32630 3345
rect 32750 3225 32805 3345
rect 32925 3225 32970 3345
rect 33090 3225 33135 3345
rect 33255 3225 33300 3345
rect 33420 3225 33475 3345
rect 33595 3225 33640 3345
rect 33760 3225 33805 3345
rect 33925 3225 33970 3345
rect 34090 3225 34145 3345
rect 34265 3225 34310 3345
rect 34430 3225 34475 3345
rect 34595 3225 34640 3345
rect 34760 3225 34815 3345
rect 34935 3225 34980 3345
rect 35100 3225 35145 3345
rect 35265 3225 35310 3345
rect 35430 3225 35485 3345
rect 35605 3225 35650 3345
rect 35770 3225 35815 3345
rect 35935 3225 35980 3345
rect 36100 3225 36155 3345
rect 36275 3225 36485 3345
rect 36605 3225 36650 3345
rect 36770 3225 36815 3345
rect 36935 3225 36980 3345
rect 37100 3225 37155 3345
rect 37275 3225 37320 3345
rect 37440 3225 37485 3345
rect 37605 3225 37650 3345
rect 37770 3225 37825 3345
rect 37945 3225 37990 3345
rect 38110 3225 38155 3345
rect 38275 3225 38320 3345
rect 38440 3225 38495 3345
rect 38615 3225 38660 3345
rect 38780 3225 38825 3345
rect 38945 3225 38990 3345
rect 39110 3225 39165 3345
rect 39285 3225 39330 3345
rect 39450 3225 39495 3345
rect 39615 3225 39660 3345
rect 39780 3225 39835 3345
rect 39955 3225 40000 3345
rect 40120 3225 40165 3345
rect 40285 3225 40330 3345
rect 40450 3225 40505 3345
rect 40625 3225 40670 3345
rect 40790 3225 40835 3345
rect 40955 3225 41000 3345
rect 41120 3225 41175 3345
rect 41295 3225 41340 3345
rect 41460 3225 41505 3345
rect 41625 3225 41670 3345
rect 41790 3225 41845 3345
rect 41965 3225 42175 3345
rect 42295 3225 42340 3345
rect 42460 3225 42505 3345
rect 42625 3225 42670 3345
rect 42790 3225 42845 3345
rect 42965 3225 43010 3345
rect 43130 3225 43175 3345
rect 43295 3225 43340 3345
rect 43460 3225 43515 3345
rect 43635 3225 43680 3345
rect 43800 3225 43845 3345
rect 43965 3225 44010 3345
rect 44130 3225 44185 3345
rect 44305 3225 44350 3345
rect 44470 3225 44515 3345
rect 44635 3225 44680 3345
rect 44800 3225 44855 3345
rect 44975 3225 45020 3345
rect 45140 3225 45185 3345
rect 45305 3225 45350 3345
rect 45470 3225 45525 3345
rect 45645 3225 45690 3345
rect 45810 3225 45855 3345
rect 45975 3225 46020 3345
rect 46140 3225 46195 3345
rect 46315 3225 46360 3345
rect 46480 3225 46525 3345
rect 46645 3225 46690 3345
rect 46810 3225 46865 3345
rect 46985 3225 47030 3345
rect 47150 3225 47195 3345
rect 47315 3225 47360 3345
rect 47480 3225 47535 3345
rect 47655 3225 47865 3345
rect 47985 3225 48030 3345
rect 48150 3225 48195 3345
rect 48315 3225 48360 3345
rect 48480 3225 48535 3345
rect 48655 3225 48700 3345
rect 48820 3225 48865 3345
rect 48985 3225 49030 3345
rect 49150 3225 49205 3345
rect 49325 3225 49370 3345
rect 49490 3225 49535 3345
rect 49655 3225 49700 3345
rect 49820 3225 49875 3345
rect 49995 3225 50040 3345
rect 50160 3225 50205 3345
rect 50325 3225 50370 3345
rect 50490 3225 50545 3345
rect 50665 3225 50710 3345
rect 50830 3225 50875 3345
rect 50995 3225 51040 3345
rect 51160 3225 51215 3345
rect 51335 3225 51380 3345
rect 51500 3225 51545 3345
rect 51665 3225 51710 3345
rect 51830 3225 51885 3345
rect 52005 3225 52050 3345
rect 52170 3225 52215 3345
rect 52335 3225 52380 3345
rect 52500 3225 52555 3345
rect 52675 3225 52720 3345
rect 52840 3225 52885 3345
rect 53005 3225 53050 3345
rect 53170 3225 53225 3345
rect 53345 3225 53370 3345
rect 30770 3180 53370 3225
rect 30770 3060 30795 3180
rect 30915 3060 30960 3180
rect 31080 3060 31125 3180
rect 31245 3060 31290 3180
rect 31410 3060 31465 3180
rect 31585 3060 31630 3180
rect 31750 3060 31795 3180
rect 31915 3060 31960 3180
rect 32080 3060 32135 3180
rect 32255 3060 32300 3180
rect 32420 3060 32465 3180
rect 32585 3060 32630 3180
rect 32750 3060 32805 3180
rect 32925 3060 32970 3180
rect 33090 3060 33135 3180
rect 33255 3060 33300 3180
rect 33420 3060 33475 3180
rect 33595 3060 33640 3180
rect 33760 3060 33805 3180
rect 33925 3060 33970 3180
rect 34090 3060 34145 3180
rect 34265 3060 34310 3180
rect 34430 3060 34475 3180
rect 34595 3060 34640 3180
rect 34760 3060 34815 3180
rect 34935 3060 34980 3180
rect 35100 3060 35145 3180
rect 35265 3060 35310 3180
rect 35430 3060 35485 3180
rect 35605 3060 35650 3180
rect 35770 3060 35815 3180
rect 35935 3060 35980 3180
rect 36100 3060 36155 3180
rect 36275 3060 36485 3180
rect 36605 3060 36650 3180
rect 36770 3060 36815 3180
rect 36935 3060 36980 3180
rect 37100 3060 37155 3180
rect 37275 3060 37320 3180
rect 37440 3060 37485 3180
rect 37605 3060 37650 3180
rect 37770 3060 37825 3180
rect 37945 3060 37990 3180
rect 38110 3060 38155 3180
rect 38275 3060 38320 3180
rect 38440 3060 38495 3180
rect 38615 3060 38660 3180
rect 38780 3060 38825 3180
rect 38945 3060 38990 3180
rect 39110 3060 39165 3180
rect 39285 3060 39330 3180
rect 39450 3060 39495 3180
rect 39615 3060 39660 3180
rect 39780 3060 39835 3180
rect 39955 3060 40000 3180
rect 40120 3060 40165 3180
rect 40285 3060 40330 3180
rect 40450 3060 40505 3180
rect 40625 3060 40670 3180
rect 40790 3060 40835 3180
rect 40955 3060 41000 3180
rect 41120 3060 41175 3180
rect 41295 3060 41340 3180
rect 41460 3060 41505 3180
rect 41625 3060 41670 3180
rect 41790 3060 41845 3180
rect 41965 3060 42175 3180
rect 42295 3060 42340 3180
rect 42460 3060 42505 3180
rect 42625 3060 42670 3180
rect 42790 3060 42845 3180
rect 42965 3060 43010 3180
rect 43130 3060 43175 3180
rect 43295 3060 43340 3180
rect 43460 3060 43515 3180
rect 43635 3060 43680 3180
rect 43800 3060 43845 3180
rect 43965 3060 44010 3180
rect 44130 3060 44185 3180
rect 44305 3060 44350 3180
rect 44470 3060 44515 3180
rect 44635 3060 44680 3180
rect 44800 3060 44855 3180
rect 44975 3060 45020 3180
rect 45140 3060 45185 3180
rect 45305 3060 45350 3180
rect 45470 3060 45525 3180
rect 45645 3060 45690 3180
rect 45810 3060 45855 3180
rect 45975 3060 46020 3180
rect 46140 3060 46195 3180
rect 46315 3060 46360 3180
rect 46480 3060 46525 3180
rect 46645 3060 46690 3180
rect 46810 3060 46865 3180
rect 46985 3060 47030 3180
rect 47150 3060 47195 3180
rect 47315 3060 47360 3180
rect 47480 3060 47535 3180
rect 47655 3060 47865 3180
rect 47985 3060 48030 3180
rect 48150 3060 48195 3180
rect 48315 3060 48360 3180
rect 48480 3060 48535 3180
rect 48655 3060 48700 3180
rect 48820 3060 48865 3180
rect 48985 3060 49030 3180
rect 49150 3060 49205 3180
rect 49325 3060 49370 3180
rect 49490 3060 49535 3180
rect 49655 3060 49700 3180
rect 49820 3060 49875 3180
rect 49995 3060 50040 3180
rect 50160 3060 50205 3180
rect 50325 3060 50370 3180
rect 50490 3060 50545 3180
rect 50665 3060 50710 3180
rect 50830 3060 50875 3180
rect 50995 3060 51040 3180
rect 51160 3060 51215 3180
rect 51335 3060 51380 3180
rect 51500 3060 51545 3180
rect 51665 3060 51710 3180
rect 51830 3060 51885 3180
rect 52005 3060 52050 3180
rect 52170 3060 52215 3180
rect 52335 3060 52380 3180
rect 52500 3060 52555 3180
rect 52675 3060 52720 3180
rect 52840 3060 52885 3180
rect 53005 3060 53050 3180
rect 53170 3060 53225 3180
rect 53345 3060 53370 3180
rect 30770 3005 53370 3060
rect 30770 2885 30795 3005
rect 30915 2885 30960 3005
rect 31080 2885 31125 3005
rect 31245 2885 31290 3005
rect 31410 2885 31465 3005
rect 31585 2885 31630 3005
rect 31750 2885 31795 3005
rect 31915 2885 31960 3005
rect 32080 2885 32135 3005
rect 32255 2885 32300 3005
rect 32420 2885 32465 3005
rect 32585 2885 32630 3005
rect 32750 2885 32805 3005
rect 32925 2885 32970 3005
rect 33090 2885 33135 3005
rect 33255 2885 33300 3005
rect 33420 2885 33475 3005
rect 33595 2885 33640 3005
rect 33760 2885 33805 3005
rect 33925 2885 33970 3005
rect 34090 2885 34145 3005
rect 34265 2885 34310 3005
rect 34430 2885 34475 3005
rect 34595 2885 34640 3005
rect 34760 2885 34815 3005
rect 34935 2885 34980 3005
rect 35100 2885 35145 3005
rect 35265 2885 35310 3005
rect 35430 2885 35485 3005
rect 35605 2885 35650 3005
rect 35770 2885 35815 3005
rect 35935 2885 35980 3005
rect 36100 2885 36155 3005
rect 36275 2885 36485 3005
rect 36605 2885 36650 3005
rect 36770 2885 36815 3005
rect 36935 2885 36980 3005
rect 37100 2885 37155 3005
rect 37275 2885 37320 3005
rect 37440 2885 37485 3005
rect 37605 2885 37650 3005
rect 37770 2885 37825 3005
rect 37945 2885 37990 3005
rect 38110 2885 38155 3005
rect 38275 2885 38320 3005
rect 38440 2885 38495 3005
rect 38615 2885 38660 3005
rect 38780 2885 38825 3005
rect 38945 2885 38990 3005
rect 39110 2885 39165 3005
rect 39285 2885 39330 3005
rect 39450 2885 39495 3005
rect 39615 2885 39660 3005
rect 39780 2885 39835 3005
rect 39955 2885 40000 3005
rect 40120 2885 40165 3005
rect 40285 2885 40330 3005
rect 40450 2885 40505 3005
rect 40625 2885 40670 3005
rect 40790 2885 40835 3005
rect 40955 2885 41000 3005
rect 41120 2885 41175 3005
rect 41295 2885 41340 3005
rect 41460 2885 41505 3005
rect 41625 2885 41670 3005
rect 41790 2885 41845 3005
rect 41965 2885 42175 3005
rect 42295 2885 42340 3005
rect 42460 2885 42505 3005
rect 42625 2885 42670 3005
rect 42790 2885 42845 3005
rect 42965 2885 43010 3005
rect 43130 2885 43175 3005
rect 43295 2885 43340 3005
rect 43460 2885 43515 3005
rect 43635 2885 43680 3005
rect 43800 2885 43845 3005
rect 43965 2885 44010 3005
rect 44130 2885 44185 3005
rect 44305 2885 44350 3005
rect 44470 2885 44515 3005
rect 44635 2885 44680 3005
rect 44800 2885 44855 3005
rect 44975 2885 45020 3005
rect 45140 2885 45185 3005
rect 45305 2885 45350 3005
rect 45470 2885 45525 3005
rect 45645 2885 45690 3005
rect 45810 2885 45855 3005
rect 45975 2885 46020 3005
rect 46140 2885 46195 3005
rect 46315 2885 46360 3005
rect 46480 2885 46525 3005
rect 46645 2885 46690 3005
rect 46810 2885 46865 3005
rect 46985 2885 47030 3005
rect 47150 2885 47195 3005
rect 47315 2885 47360 3005
rect 47480 2885 47535 3005
rect 47655 2885 47865 3005
rect 47985 2885 48030 3005
rect 48150 2885 48195 3005
rect 48315 2885 48360 3005
rect 48480 2885 48535 3005
rect 48655 2885 48700 3005
rect 48820 2885 48865 3005
rect 48985 2885 49030 3005
rect 49150 2885 49205 3005
rect 49325 2885 49370 3005
rect 49490 2885 49535 3005
rect 49655 2885 49700 3005
rect 49820 2885 49875 3005
rect 49995 2885 50040 3005
rect 50160 2885 50205 3005
rect 50325 2885 50370 3005
rect 50490 2885 50545 3005
rect 50665 2885 50710 3005
rect 50830 2885 50875 3005
rect 50995 2885 51040 3005
rect 51160 2885 51215 3005
rect 51335 2885 51380 3005
rect 51500 2885 51545 3005
rect 51665 2885 51710 3005
rect 51830 2885 51885 3005
rect 52005 2885 52050 3005
rect 52170 2885 52215 3005
rect 52335 2885 52380 3005
rect 52500 2885 52555 3005
rect 52675 2885 52720 3005
rect 52840 2885 52885 3005
rect 53005 2885 53050 3005
rect 53170 2885 53225 3005
rect 53345 2885 53370 3005
rect 30770 2840 53370 2885
rect 30770 2720 30795 2840
rect 30915 2720 30960 2840
rect 31080 2720 31125 2840
rect 31245 2720 31290 2840
rect 31410 2720 31465 2840
rect 31585 2720 31630 2840
rect 31750 2720 31795 2840
rect 31915 2720 31960 2840
rect 32080 2720 32135 2840
rect 32255 2720 32300 2840
rect 32420 2720 32465 2840
rect 32585 2720 32630 2840
rect 32750 2720 32805 2840
rect 32925 2720 32970 2840
rect 33090 2720 33135 2840
rect 33255 2720 33300 2840
rect 33420 2720 33475 2840
rect 33595 2720 33640 2840
rect 33760 2720 33805 2840
rect 33925 2720 33970 2840
rect 34090 2720 34145 2840
rect 34265 2720 34310 2840
rect 34430 2720 34475 2840
rect 34595 2720 34640 2840
rect 34760 2720 34815 2840
rect 34935 2720 34980 2840
rect 35100 2720 35145 2840
rect 35265 2720 35310 2840
rect 35430 2720 35485 2840
rect 35605 2720 35650 2840
rect 35770 2720 35815 2840
rect 35935 2720 35980 2840
rect 36100 2720 36155 2840
rect 36275 2720 36485 2840
rect 36605 2720 36650 2840
rect 36770 2720 36815 2840
rect 36935 2720 36980 2840
rect 37100 2720 37155 2840
rect 37275 2720 37320 2840
rect 37440 2720 37485 2840
rect 37605 2720 37650 2840
rect 37770 2720 37825 2840
rect 37945 2720 37990 2840
rect 38110 2720 38155 2840
rect 38275 2720 38320 2840
rect 38440 2720 38495 2840
rect 38615 2720 38660 2840
rect 38780 2720 38825 2840
rect 38945 2720 38990 2840
rect 39110 2720 39165 2840
rect 39285 2720 39330 2840
rect 39450 2720 39495 2840
rect 39615 2720 39660 2840
rect 39780 2720 39835 2840
rect 39955 2720 40000 2840
rect 40120 2720 40165 2840
rect 40285 2720 40330 2840
rect 40450 2720 40505 2840
rect 40625 2720 40670 2840
rect 40790 2720 40835 2840
rect 40955 2720 41000 2840
rect 41120 2720 41175 2840
rect 41295 2720 41340 2840
rect 41460 2720 41505 2840
rect 41625 2720 41670 2840
rect 41790 2720 41845 2840
rect 41965 2720 42175 2840
rect 42295 2720 42340 2840
rect 42460 2720 42505 2840
rect 42625 2720 42670 2840
rect 42790 2720 42845 2840
rect 42965 2720 43010 2840
rect 43130 2720 43175 2840
rect 43295 2720 43340 2840
rect 43460 2720 43515 2840
rect 43635 2720 43680 2840
rect 43800 2720 43845 2840
rect 43965 2720 44010 2840
rect 44130 2720 44185 2840
rect 44305 2720 44350 2840
rect 44470 2720 44515 2840
rect 44635 2720 44680 2840
rect 44800 2720 44855 2840
rect 44975 2720 45020 2840
rect 45140 2720 45185 2840
rect 45305 2720 45350 2840
rect 45470 2720 45525 2840
rect 45645 2720 45690 2840
rect 45810 2720 45855 2840
rect 45975 2720 46020 2840
rect 46140 2720 46195 2840
rect 46315 2720 46360 2840
rect 46480 2720 46525 2840
rect 46645 2720 46690 2840
rect 46810 2720 46865 2840
rect 46985 2720 47030 2840
rect 47150 2720 47195 2840
rect 47315 2720 47360 2840
rect 47480 2720 47535 2840
rect 47655 2720 47865 2840
rect 47985 2720 48030 2840
rect 48150 2720 48195 2840
rect 48315 2720 48360 2840
rect 48480 2720 48535 2840
rect 48655 2720 48700 2840
rect 48820 2720 48865 2840
rect 48985 2720 49030 2840
rect 49150 2720 49205 2840
rect 49325 2720 49370 2840
rect 49490 2720 49535 2840
rect 49655 2720 49700 2840
rect 49820 2720 49875 2840
rect 49995 2720 50040 2840
rect 50160 2720 50205 2840
rect 50325 2720 50370 2840
rect 50490 2720 50545 2840
rect 50665 2720 50710 2840
rect 50830 2720 50875 2840
rect 50995 2720 51040 2840
rect 51160 2720 51215 2840
rect 51335 2720 51380 2840
rect 51500 2720 51545 2840
rect 51665 2720 51710 2840
rect 51830 2720 51885 2840
rect 52005 2720 52050 2840
rect 52170 2720 52215 2840
rect 52335 2720 52380 2840
rect 52500 2720 52555 2840
rect 52675 2720 52720 2840
rect 52840 2720 52885 2840
rect 53005 2720 53050 2840
rect 53170 2720 53225 2840
rect 53345 2720 53370 2840
rect 30770 2675 53370 2720
rect 30770 2555 30795 2675
rect 30915 2555 30960 2675
rect 31080 2555 31125 2675
rect 31245 2555 31290 2675
rect 31410 2555 31465 2675
rect 31585 2555 31630 2675
rect 31750 2555 31795 2675
rect 31915 2555 31960 2675
rect 32080 2555 32135 2675
rect 32255 2555 32300 2675
rect 32420 2555 32465 2675
rect 32585 2555 32630 2675
rect 32750 2555 32805 2675
rect 32925 2555 32970 2675
rect 33090 2555 33135 2675
rect 33255 2555 33300 2675
rect 33420 2555 33475 2675
rect 33595 2555 33640 2675
rect 33760 2555 33805 2675
rect 33925 2555 33970 2675
rect 34090 2555 34145 2675
rect 34265 2555 34310 2675
rect 34430 2555 34475 2675
rect 34595 2555 34640 2675
rect 34760 2555 34815 2675
rect 34935 2555 34980 2675
rect 35100 2555 35145 2675
rect 35265 2555 35310 2675
rect 35430 2555 35485 2675
rect 35605 2555 35650 2675
rect 35770 2555 35815 2675
rect 35935 2555 35980 2675
rect 36100 2555 36155 2675
rect 36275 2555 36485 2675
rect 36605 2555 36650 2675
rect 36770 2555 36815 2675
rect 36935 2555 36980 2675
rect 37100 2555 37155 2675
rect 37275 2555 37320 2675
rect 37440 2555 37485 2675
rect 37605 2555 37650 2675
rect 37770 2555 37825 2675
rect 37945 2555 37990 2675
rect 38110 2555 38155 2675
rect 38275 2555 38320 2675
rect 38440 2555 38495 2675
rect 38615 2555 38660 2675
rect 38780 2555 38825 2675
rect 38945 2555 38990 2675
rect 39110 2555 39165 2675
rect 39285 2555 39330 2675
rect 39450 2555 39495 2675
rect 39615 2555 39660 2675
rect 39780 2555 39835 2675
rect 39955 2555 40000 2675
rect 40120 2555 40165 2675
rect 40285 2555 40330 2675
rect 40450 2555 40505 2675
rect 40625 2555 40670 2675
rect 40790 2555 40835 2675
rect 40955 2555 41000 2675
rect 41120 2555 41175 2675
rect 41295 2555 41340 2675
rect 41460 2555 41505 2675
rect 41625 2555 41670 2675
rect 41790 2555 41845 2675
rect 41965 2555 42175 2675
rect 42295 2555 42340 2675
rect 42460 2555 42505 2675
rect 42625 2555 42670 2675
rect 42790 2555 42845 2675
rect 42965 2555 43010 2675
rect 43130 2555 43175 2675
rect 43295 2555 43340 2675
rect 43460 2555 43515 2675
rect 43635 2555 43680 2675
rect 43800 2555 43845 2675
rect 43965 2555 44010 2675
rect 44130 2555 44185 2675
rect 44305 2555 44350 2675
rect 44470 2555 44515 2675
rect 44635 2555 44680 2675
rect 44800 2555 44855 2675
rect 44975 2555 45020 2675
rect 45140 2555 45185 2675
rect 45305 2555 45350 2675
rect 45470 2555 45525 2675
rect 45645 2555 45690 2675
rect 45810 2555 45855 2675
rect 45975 2555 46020 2675
rect 46140 2555 46195 2675
rect 46315 2555 46360 2675
rect 46480 2555 46525 2675
rect 46645 2555 46690 2675
rect 46810 2555 46865 2675
rect 46985 2555 47030 2675
rect 47150 2555 47195 2675
rect 47315 2555 47360 2675
rect 47480 2555 47535 2675
rect 47655 2555 47865 2675
rect 47985 2555 48030 2675
rect 48150 2555 48195 2675
rect 48315 2555 48360 2675
rect 48480 2555 48535 2675
rect 48655 2555 48700 2675
rect 48820 2555 48865 2675
rect 48985 2555 49030 2675
rect 49150 2555 49205 2675
rect 49325 2555 49370 2675
rect 49490 2555 49535 2675
rect 49655 2555 49700 2675
rect 49820 2555 49875 2675
rect 49995 2555 50040 2675
rect 50160 2555 50205 2675
rect 50325 2555 50370 2675
rect 50490 2555 50545 2675
rect 50665 2555 50710 2675
rect 50830 2555 50875 2675
rect 50995 2555 51040 2675
rect 51160 2555 51215 2675
rect 51335 2555 51380 2675
rect 51500 2555 51545 2675
rect 51665 2555 51710 2675
rect 51830 2555 51885 2675
rect 52005 2555 52050 2675
rect 52170 2555 52215 2675
rect 52335 2555 52380 2675
rect 52500 2555 52555 2675
rect 52675 2555 52720 2675
rect 52840 2555 52885 2675
rect 53005 2555 53050 2675
rect 53170 2555 53225 2675
rect 53345 2555 53370 2675
rect 30770 2510 53370 2555
rect 30770 2390 30795 2510
rect 30915 2390 30960 2510
rect 31080 2390 31125 2510
rect 31245 2390 31290 2510
rect 31410 2390 31465 2510
rect 31585 2390 31630 2510
rect 31750 2390 31795 2510
rect 31915 2390 31960 2510
rect 32080 2390 32135 2510
rect 32255 2390 32300 2510
rect 32420 2390 32465 2510
rect 32585 2390 32630 2510
rect 32750 2390 32805 2510
rect 32925 2390 32970 2510
rect 33090 2390 33135 2510
rect 33255 2390 33300 2510
rect 33420 2390 33475 2510
rect 33595 2390 33640 2510
rect 33760 2390 33805 2510
rect 33925 2390 33970 2510
rect 34090 2390 34145 2510
rect 34265 2390 34310 2510
rect 34430 2390 34475 2510
rect 34595 2390 34640 2510
rect 34760 2390 34815 2510
rect 34935 2390 34980 2510
rect 35100 2390 35145 2510
rect 35265 2390 35310 2510
rect 35430 2390 35485 2510
rect 35605 2390 35650 2510
rect 35770 2390 35815 2510
rect 35935 2390 35980 2510
rect 36100 2390 36155 2510
rect 36275 2390 36485 2510
rect 36605 2390 36650 2510
rect 36770 2390 36815 2510
rect 36935 2390 36980 2510
rect 37100 2390 37155 2510
rect 37275 2390 37320 2510
rect 37440 2390 37485 2510
rect 37605 2390 37650 2510
rect 37770 2390 37825 2510
rect 37945 2390 37990 2510
rect 38110 2390 38155 2510
rect 38275 2390 38320 2510
rect 38440 2390 38495 2510
rect 38615 2390 38660 2510
rect 38780 2390 38825 2510
rect 38945 2390 38990 2510
rect 39110 2390 39165 2510
rect 39285 2390 39330 2510
rect 39450 2390 39495 2510
rect 39615 2390 39660 2510
rect 39780 2390 39835 2510
rect 39955 2390 40000 2510
rect 40120 2390 40165 2510
rect 40285 2390 40330 2510
rect 40450 2390 40505 2510
rect 40625 2390 40670 2510
rect 40790 2390 40835 2510
rect 40955 2390 41000 2510
rect 41120 2390 41175 2510
rect 41295 2390 41340 2510
rect 41460 2390 41505 2510
rect 41625 2390 41670 2510
rect 41790 2390 41845 2510
rect 41965 2390 42175 2510
rect 42295 2390 42340 2510
rect 42460 2390 42505 2510
rect 42625 2390 42670 2510
rect 42790 2390 42845 2510
rect 42965 2390 43010 2510
rect 43130 2390 43175 2510
rect 43295 2390 43340 2510
rect 43460 2390 43515 2510
rect 43635 2390 43680 2510
rect 43800 2390 43845 2510
rect 43965 2390 44010 2510
rect 44130 2390 44185 2510
rect 44305 2390 44350 2510
rect 44470 2390 44515 2510
rect 44635 2390 44680 2510
rect 44800 2390 44855 2510
rect 44975 2390 45020 2510
rect 45140 2390 45185 2510
rect 45305 2390 45350 2510
rect 45470 2390 45525 2510
rect 45645 2390 45690 2510
rect 45810 2390 45855 2510
rect 45975 2390 46020 2510
rect 46140 2390 46195 2510
rect 46315 2390 46360 2510
rect 46480 2390 46525 2510
rect 46645 2390 46690 2510
rect 46810 2390 46865 2510
rect 46985 2390 47030 2510
rect 47150 2390 47195 2510
rect 47315 2390 47360 2510
rect 47480 2390 47535 2510
rect 47655 2390 47865 2510
rect 47985 2390 48030 2510
rect 48150 2390 48195 2510
rect 48315 2390 48360 2510
rect 48480 2390 48535 2510
rect 48655 2390 48700 2510
rect 48820 2390 48865 2510
rect 48985 2390 49030 2510
rect 49150 2390 49205 2510
rect 49325 2390 49370 2510
rect 49490 2390 49535 2510
rect 49655 2390 49700 2510
rect 49820 2390 49875 2510
rect 49995 2390 50040 2510
rect 50160 2390 50205 2510
rect 50325 2390 50370 2510
rect 50490 2390 50545 2510
rect 50665 2390 50710 2510
rect 50830 2390 50875 2510
rect 50995 2390 51040 2510
rect 51160 2390 51215 2510
rect 51335 2390 51380 2510
rect 51500 2390 51545 2510
rect 51665 2390 51710 2510
rect 51830 2390 51885 2510
rect 52005 2390 52050 2510
rect 52170 2390 52215 2510
rect 52335 2390 52380 2510
rect 52500 2390 52555 2510
rect 52675 2390 52720 2510
rect 52840 2390 52885 2510
rect 53005 2390 53050 2510
rect 53170 2390 53225 2510
rect 53345 2390 53370 2510
rect 30770 2335 53370 2390
rect 30770 2215 30795 2335
rect 30915 2215 30960 2335
rect 31080 2215 31125 2335
rect 31245 2215 31290 2335
rect 31410 2215 31465 2335
rect 31585 2215 31630 2335
rect 31750 2215 31795 2335
rect 31915 2215 31960 2335
rect 32080 2215 32135 2335
rect 32255 2215 32300 2335
rect 32420 2215 32465 2335
rect 32585 2215 32630 2335
rect 32750 2215 32805 2335
rect 32925 2215 32970 2335
rect 33090 2215 33135 2335
rect 33255 2215 33300 2335
rect 33420 2215 33475 2335
rect 33595 2215 33640 2335
rect 33760 2215 33805 2335
rect 33925 2215 33970 2335
rect 34090 2215 34145 2335
rect 34265 2215 34310 2335
rect 34430 2215 34475 2335
rect 34595 2215 34640 2335
rect 34760 2215 34815 2335
rect 34935 2215 34980 2335
rect 35100 2215 35145 2335
rect 35265 2215 35310 2335
rect 35430 2215 35485 2335
rect 35605 2215 35650 2335
rect 35770 2215 35815 2335
rect 35935 2215 35980 2335
rect 36100 2215 36155 2335
rect 36275 2215 36485 2335
rect 36605 2215 36650 2335
rect 36770 2215 36815 2335
rect 36935 2215 36980 2335
rect 37100 2215 37155 2335
rect 37275 2215 37320 2335
rect 37440 2215 37485 2335
rect 37605 2215 37650 2335
rect 37770 2215 37825 2335
rect 37945 2215 37990 2335
rect 38110 2215 38155 2335
rect 38275 2215 38320 2335
rect 38440 2215 38495 2335
rect 38615 2215 38660 2335
rect 38780 2215 38825 2335
rect 38945 2215 38990 2335
rect 39110 2215 39165 2335
rect 39285 2215 39330 2335
rect 39450 2215 39495 2335
rect 39615 2215 39660 2335
rect 39780 2215 39835 2335
rect 39955 2215 40000 2335
rect 40120 2215 40165 2335
rect 40285 2215 40330 2335
rect 40450 2215 40505 2335
rect 40625 2215 40670 2335
rect 40790 2215 40835 2335
rect 40955 2215 41000 2335
rect 41120 2215 41175 2335
rect 41295 2215 41340 2335
rect 41460 2215 41505 2335
rect 41625 2215 41670 2335
rect 41790 2215 41845 2335
rect 41965 2215 42175 2335
rect 42295 2215 42340 2335
rect 42460 2215 42505 2335
rect 42625 2215 42670 2335
rect 42790 2215 42845 2335
rect 42965 2215 43010 2335
rect 43130 2215 43175 2335
rect 43295 2215 43340 2335
rect 43460 2215 43515 2335
rect 43635 2215 43680 2335
rect 43800 2215 43845 2335
rect 43965 2215 44010 2335
rect 44130 2215 44185 2335
rect 44305 2215 44350 2335
rect 44470 2215 44515 2335
rect 44635 2215 44680 2335
rect 44800 2215 44855 2335
rect 44975 2215 45020 2335
rect 45140 2215 45185 2335
rect 45305 2215 45350 2335
rect 45470 2215 45525 2335
rect 45645 2215 45690 2335
rect 45810 2215 45855 2335
rect 45975 2215 46020 2335
rect 46140 2215 46195 2335
rect 46315 2215 46360 2335
rect 46480 2215 46525 2335
rect 46645 2215 46690 2335
rect 46810 2215 46865 2335
rect 46985 2215 47030 2335
rect 47150 2215 47195 2335
rect 47315 2215 47360 2335
rect 47480 2215 47535 2335
rect 47655 2215 47865 2335
rect 47985 2215 48030 2335
rect 48150 2215 48195 2335
rect 48315 2215 48360 2335
rect 48480 2215 48535 2335
rect 48655 2215 48700 2335
rect 48820 2215 48865 2335
rect 48985 2215 49030 2335
rect 49150 2215 49205 2335
rect 49325 2215 49370 2335
rect 49490 2215 49535 2335
rect 49655 2215 49700 2335
rect 49820 2215 49875 2335
rect 49995 2215 50040 2335
rect 50160 2215 50205 2335
rect 50325 2215 50370 2335
rect 50490 2215 50545 2335
rect 50665 2215 50710 2335
rect 50830 2215 50875 2335
rect 50995 2215 51040 2335
rect 51160 2215 51215 2335
rect 51335 2215 51380 2335
rect 51500 2215 51545 2335
rect 51665 2215 51710 2335
rect 51830 2215 51885 2335
rect 52005 2215 52050 2335
rect 52170 2215 52215 2335
rect 52335 2215 52380 2335
rect 52500 2215 52555 2335
rect 52675 2215 52720 2335
rect 52840 2215 52885 2335
rect 53005 2215 53050 2335
rect 53170 2215 53225 2335
rect 53345 2215 53370 2335
rect 30770 2170 53370 2215
rect 30770 2050 30795 2170
rect 30915 2050 30960 2170
rect 31080 2050 31125 2170
rect 31245 2050 31290 2170
rect 31410 2050 31465 2170
rect 31585 2050 31630 2170
rect 31750 2050 31795 2170
rect 31915 2050 31960 2170
rect 32080 2050 32135 2170
rect 32255 2050 32300 2170
rect 32420 2050 32465 2170
rect 32585 2050 32630 2170
rect 32750 2050 32805 2170
rect 32925 2050 32970 2170
rect 33090 2050 33135 2170
rect 33255 2050 33300 2170
rect 33420 2050 33475 2170
rect 33595 2050 33640 2170
rect 33760 2050 33805 2170
rect 33925 2050 33970 2170
rect 34090 2050 34145 2170
rect 34265 2050 34310 2170
rect 34430 2050 34475 2170
rect 34595 2050 34640 2170
rect 34760 2050 34815 2170
rect 34935 2050 34980 2170
rect 35100 2050 35145 2170
rect 35265 2050 35310 2170
rect 35430 2050 35485 2170
rect 35605 2050 35650 2170
rect 35770 2050 35815 2170
rect 35935 2050 35980 2170
rect 36100 2050 36155 2170
rect 36275 2050 36485 2170
rect 36605 2050 36650 2170
rect 36770 2050 36815 2170
rect 36935 2050 36980 2170
rect 37100 2050 37155 2170
rect 37275 2050 37320 2170
rect 37440 2050 37485 2170
rect 37605 2050 37650 2170
rect 37770 2050 37825 2170
rect 37945 2050 37990 2170
rect 38110 2050 38155 2170
rect 38275 2050 38320 2170
rect 38440 2050 38495 2170
rect 38615 2050 38660 2170
rect 38780 2050 38825 2170
rect 38945 2050 38990 2170
rect 39110 2050 39165 2170
rect 39285 2050 39330 2170
rect 39450 2050 39495 2170
rect 39615 2050 39660 2170
rect 39780 2050 39835 2170
rect 39955 2050 40000 2170
rect 40120 2050 40165 2170
rect 40285 2050 40330 2170
rect 40450 2050 40505 2170
rect 40625 2050 40670 2170
rect 40790 2050 40835 2170
rect 40955 2050 41000 2170
rect 41120 2050 41175 2170
rect 41295 2050 41340 2170
rect 41460 2050 41505 2170
rect 41625 2050 41670 2170
rect 41790 2050 41845 2170
rect 41965 2050 42175 2170
rect 42295 2050 42340 2170
rect 42460 2050 42505 2170
rect 42625 2050 42670 2170
rect 42790 2050 42845 2170
rect 42965 2050 43010 2170
rect 43130 2050 43175 2170
rect 43295 2050 43340 2170
rect 43460 2050 43515 2170
rect 43635 2050 43680 2170
rect 43800 2050 43845 2170
rect 43965 2050 44010 2170
rect 44130 2050 44185 2170
rect 44305 2050 44350 2170
rect 44470 2050 44515 2170
rect 44635 2050 44680 2170
rect 44800 2050 44855 2170
rect 44975 2050 45020 2170
rect 45140 2050 45185 2170
rect 45305 2050 45350 2170
rect 45470 2050 45525 2170
rect 45645 2050 45690 2170
rect 45810 2050 45855 2170
rect 45975 2050 46020 2170
rect 46140 2050 46195 2170
rect 46315 2050 46360 2170
rect 46480 2050 46525 2170
rect 46645 2050 46690 2170
rect 46810 2050 46865 2170
rect 46985 2050 47030 2170
rect 47150 2050 47195 2170
rect 47315 2050 47360 2170
rect 47480 2050 47535 2170
rect 47655 2050 47865 2170
rect 47985 2050 48030 2170
rect 48150 2050 48195 2170
rect 48315 2050 48360 2170
rect 48480 2050 48535 2170
rect 48655 2050 48700 2170
rect 48820 2050 48865 2170
rect 48985 2050 49030 2170
rect 49150 2050 49205 2170
rect 49325 2050 49370 2170
rect 49490 2050 49535 2170
rect 49655 2050 49700 2170
rect 49820 2050 49875 2170
rect 49995 2050 50040 2170
rect 50160 2050 50205 2170
rect 50325 2050 50370 2170
rect 50490 2050 50545 2170
rect 50665 2050 50710 2170
rect 50830 2050 50875 2170
rect 50995 2050 51040 2170
rect 51160 2050 51215 2170
rect 51335 2050 51380 2170
rect 51500 2050 51545 2170
rect 51665 2050 51710 2170
rect 51830 2050 51885 2170
rect 52005 2050 52050 2170
rect 52170 2050 52215 2170
rect 52335 2050 52380 2170
rect 52500 2050 52555 2170
rect 52675 2050 52720 2170
rect 52840 2050 52885 2170
rect 53005 2050 53050 2170
rect 53170 2050 53225 2170
rect 53345 2050 53370 2170
rect 30770 2005 53370 2050
rect 30770 1885 30795 2005
rect 30915 1885 30960 2005
rect 31080 1885 31125 2005
rect 31245 1885 31290 2005
rect 31410 1885 31465 2005
rect 31585 1885 31630 2005
rect 31750 1885 31795 2005
rect 31915 1885 31960 2005
rect 32080 1885 32135 2005
rect 32255 1885 32300 2005
rect 32420 1885 32465 2005
rect 32585 1885 32630 2005
rect 32750 1885 32805 2005
rect 32925 1885 32970 2005
rect 33090 1885 33135 2005
rect 33255 1885 33300 2005
rect 33420 1885 33475 2005
rect 33595 1885 33640 2005
rect 33760 1885 33805 2005
rect 33925 1885 33970 2005
rect 34090 1885 34145 2005
rect 34265 1885 34310 2005
rect 34430 1885 34475 2005
rect 34595 1885 34640 2005
rect 34760 1885 34815 2005
rect 34935 1885 34980 2005
rect 35100 1885 35145 2005
rect 35265 1885 35310 2005
rect 35430 1885 35485 2005
rect 35605 1885 35650 2005
rect 35770 1885 35815 2005
rect 35935 1885 35980 2005
rect 36100 1885 36155 2005
rect 36275 1885 36485 2005
rect 36605 1885 36650 2005
rect 36770 1885 36815 2005
rect 36935 1885 36980 2005
rect 37100 1885 37155 2005
rect 37275 1885 37320 2005
rect 37440 1885 37485 2005
rect 37605 1885 37650 2005
rect 37770 1885 37825 2005
rect 37945 1885 37990 2005
rect 38110 1885 38155 2005
rect 38275 1885 38320 2005
rect 38440 1885 38495 2005
rect 38615 1885 38660 2005
rect 38780 1885 38825 2005
rect 38945 1885 38990 2005
rect 39110 1885 39165 2005
rect 39285 1885 39330 2005
rect 39450 1885 39495 2005
rect 39615 1885 39660 2005
rect 39780 1885 39835 2005
rect 39955 1885 40000 2005
rect 40120 1885 40165 2005
rect 40285 1885 40330 2005
rect 40450 1885 40505 2005
rect 40625 1885 40670 2005
rect 40790 1885 40835 2005
rect 40955 1885 41000 2005
rect 41120 1885 41175 2005
rect 41295 1885 41340 2005
rect 41460 1885 41505 2005
rect 41625 1885 41670 2005
rect 41790 1885 41845 2005
rect 41965 1885 42175 2005
rect 42295 1885 42340 2005
rect 42460 1885 42505 2005
rect 42625 1885 42670 2005
rect 42790 1885 42845 2005
rect 42965 1885 43010 2005
rect 43130 1885 43175 2005
rect 43295 1885 43340 2005
rect 43460 1885 43515 2005
rect 43635 1885 43680 2005
rect 43800 1885 43845 2005
rect 43965 1885 44010 2005
rect 44130 1885 44185 2005
rect 44305 1885 44350 2005
rect 44470 1885 44515 2005
rect 44635 1885 44680 2005
rect 44800 1885 44855 2005
rect 44975 1885 45020 2005
rect 45140 1885 45185 2005
rect 45305 1885 45350 2005
rect 45470 1885 45525 2005
rect 45645 1885 45690 2005
rect 45810 1885 45855 2005
rect 45975 1885 46020 2005
rect 46140 1885 46195 2005
rect 46315 1885 46360 2005
rect 46480 1885 46525 2005
rect 46645 1885 46690 2005
rect 46810 1885 46865 2005
rect 46985 1885 47030 2005
rect 47150 1885 47195 2005
rect 47315 1885 47360 2005
rect 47480 1885 47535 2005
rect 47655 1885 47865 2005
rect 47985 1885 48030 2005
rect 48150 1885 48195 2005
rect 48315 1885 48360 2005
rect 48480 1885 48535 2005
rect 48655 1885 48700 2005
rect 48820 1885 48865 2005
rect 48985 1885 49030 2005
rect 49150 1885 49205 2005
rect 49325 1885 49370 2005
rect 49490 1885 49535 2005
rect 49655 1885 49700 2005
rect 49820 1885 49875 2005
rect 49995 1885 50040 2005
rect 50160 1885 50205 2005
rect 50325 1885 50370 2005
rect 50490 1885 50545 2005
rect 50665 1885 50710 2005
rect 50830 1885 50875 2005
rect 50995 1885 51040 2005
rect 51160 1885 51215 2005
rect 51335 1885 51380 2005
rect 51500 1885 51545 2005
rect 51665 1885 51710 2005
rect 51830 1885 51885 2005
rect 52005 1885 52050 2005
rect 52170 1885 52215 2005
rect 52335 1885 52380 2005
rect 52500 1885 52555 2005
rect 52675 1885 52720 2005
rect 52840 1885 52885 2005
rect 53005 1885 53050 2005
rect 53170 1885 53225 2005
rect 53345 1885 53370 2005
rect 30770 1840 53370 1885
rect 30770 1720 30795 1840
rect 30915 1720 30960 1840
rect 31080 1720 31125 1840
rect 31245 1720 31290 1840
rect 31410 1720 31465 1840
rect 31585 1720 31630 1840
rect 31750 1720 31795 1840
rect 31915 1720 31960 1840
rect 32080 1720 32135 1840
rect 32255 1720 32300 1840
rect 32420 1720 32465 1840
rect 32585 1720 32630 1840
rect 32750 1720 32805 1840
rect 32925 1720 32970 1840
rect 33090 1720 33135 1840
rect 33255 1720 33300 1840
rect 33420 1720 33475 1840
rect 33595 1720 33640 1840
rect 33760 1720 33805 1840
rect 33925 1720 33970 1840
rect 34090 1720 34145 1840
rect 34265 1720 34310 1840
rect 34430 1720 34475 1840
rect 34595 1720 34640 1840
rect 34760 1720 34815 1840
rect 34935 1720 34980 1840
rect 35100 1720 35145 1840
rect 35265 1720 35310 1840
rect 35430 1720 35485 1840
rect 35605 1720 35650 1840
rect 35770 1720 35815 1840
rect 35935 1720 35980 1840
rect 36100 1720 36155 1840
rect 36275 1720 36485 1840
rect 36605 1720 36650 1840
rect 36770 1720 36815 1840
rect 36935 1720 36980 1840
rect 37100 1720 37155 1840
rect 37275 1720 37320 1840
rect 37440 1720 37485 1840
rect 37605 1720 37650 1840
rect 37770 1720 37825 1840
rect 37945 1720 37990 1840
rect 38110 1720 38155 1840
rect 38275 1720 38320 1840
rect 38440 1720 38495 1840
rect 38615 1720 38660 1840
rect 38780 1720 38825 1840
rect 38945 1720 38990 1840
rect 39110 1720 39165 1840
rect 39285 1720 39330 1840
rect 39450 1720 39495 1840
rect 39615 1720 39660 1840
rect 39780 1720 39835 1840
rect 39955 1720 40000 1840
rect 40120 1720 40165 1840
rect 40285 1720 40330 1840
rect 40450 1720 40505 1840
rect 40625 1720 40670 1840
rect 40790 1720 40835 1840
rect 40955 1720 41000 1840
rect 41120 1720 41175 1840
rect 41295 1720 41340 1840
rect 41460 1720 41505 1840
rect 41625 1720 41670 1840
rect 41790 1720 41845 1840
rect 41965 1720 42175 1840
rect 42295 1720 42340 1840
rect 42460 1720 42505 1840
rect 42625 1720 42670 1840
rect 42790 1720 42845 1840
rect 42965 1720 43010 1840
rect 43130 1720 43175 1840
rect 43295 1720 43340 1840
rect 43460 1720 43515 1840
rect 43635 1720 43680 1840
rect 43800 1720 43845 1840
rect 43965 1720 44010 1840
rect 44130 1720 44185 1840
rect 44305 1720 44350 1840
rect 44470 1720 44515 1840
rect 44635 1720 44680 1840
rect 44800 1720 44855 1840
rect 44975 1720 45020 1840
rect 45140 1720 45185 1840
rect 45305 1720 45350 1840
rect 45470 1720 45525 1840
rect 45645 1720 45690 1840
rect 45810 1720 45855 1840
rect 45975 1720 46020 1840
rect 46140 1720 46195 1840
rect 46315 1720 46360 1840
rect 46480 1720 46525 1840
rect 46645 1720 46690 1840
rect 46810 1720 46865 1840
rect 46985 1720 47030 1840
rect 47150 1720 47195 1840
rect 47315 1720 47360 1840
rect 47480 1720 47535 1840
rect 47655 1720 47865 1840
rect 47985 1720 48030 1840
rect 48150 1720 48195 1840
rect 48315 1720 48360 1840
rect 48480 1720 48535 1840
rect 48655 1720 48700 1840
rect 48820 1720 48865 1840
rect 48985 1720 49030 1840
rect 49150 1720 49205 1840
rect 49325 1720 49370 1840
rect 49490 1720 49535 1840
rect 49655 1720 49700 1840
rect 49820 1720 49875 1840
rect 49995 1720 50040 1840
rect 50160 1720 50205 1840
rect 50325 1720 50370 1840
rect 50490 1720 50545 1840
rect 50665 1720 50710 1840
rect 50830 1720 50875 1840
rect 50995 1720 51040 1840
rect 51160 1720 51215 1840
rect 51335 1720 51380 1840
rect 51500 1720 51545 1840
rect 51665 1720 51710 1840
rect 51830 1720 51885 1840
rect 52005 1720 52050 1840
rect 52170 1720 52215 1840
rect 52335 1720 52380 1840
rect 52500 1720 52555 1840
rect 52675 1720 52720 1840
rect 52840 1720 52885 1840
rect 53005 1720 53050 1840
rect 53170 1720 53225 1840
rect 53345 1720 53370 1840
rect 30770 1695 53370 1720
rect 36300 1645 36460 1650
rect 41990 1645 42150 1650
rect 47680 1645 47840 1650
rect 30770 1630 53370 1645
rect 30770 1510 30835 1630
rect 30955 1510 31000 1630
rect 31120 1510 31165 1630
rect 31285 1510 31330 1630
rect 31450 1510 31495 1630
rect 31615 1510 31660 1630
rect 31780 1510 31825 1630
rect 31945 1510 31990 1630
rect 32110 1510 32155 1630
rect 32275 1510 32320 1630
rect 32440 1510 32485 1630
rect 32605 1510 32650 1630
rect 32770 1510 32815 1630
rect 32935 1510 32980 1630
rect 33100 1510 33145 1630
rect 33265 1510 33310 1630
rect 33430 1510 33475 1630
rect 33595 1510 33640 1630
rect 33760 1510 33805 1630
rect 33925 1510 33970 1630
rect 34090 1510 34135 1630
rect 34255 1510 34300 1630
rect 34420 1510 34465 1630
rect 34585 1510 34630 1630
rect 34750 1510 34795 1630
rect 34915 1510 34960 1630
rect 35080 1510 35125 1630
rect 35245 1510 35290 1630
rect 35410 1510 35455 1630
rect 35575 1510 35620 1630
rect 35740 1510 35785 1630
rect 35905 1510 35950 1630
rect 36070 1510 36115 1630
rect 36235 1510 36525 1630
rect 36645 1510 36690 1630
rect 36810 1510 36855 1630
rect 36975 1510 37020 1630
rect 37140 1510 37185 1630
rect 37305 1510 37350 1630
rect 37470 1510 37515 1630
rect 37635 1510 37680 1630
rect 37800 1510 37845 1630
rect 37965 1510 38010 1630
rect 38130 1510 38175 1630
rect 38295 1510 38340 1630
rect 38460 1510 38505 1630
rect 38625 1510 38670 1630
rect 38790 1510 38835 1630
rect 38955 1510 39000 1630
rect 39120 1510 39165 1630
rect 39285 1510 39330 1630
rect 39450 1510 39495 1630
rect 39615 1510 39660 1630
rect 39780 1510 39825 1630
rect 39945 1510 39990 1630
rect 40110 1510 40155 1630
rect 40275 1510 40320 1630
rect 40440 1510 40485 1630
rect 40605 1510 40650 1630
rect 40770 1510 40815 1630
rect 40935 1510 40980 1630
rect 41100 1510 41145 1630
rect 41265 1510 41310 1630
rect 41430 1510 41475 1630
rect 41595 1510 41640 1630
rect 41760 1510 41805 1630
rect 41925 1510 42215 1630
rect 42335 1510 42380 1630
rect 42500 1510 42545 1630
rect 42665 1510 42710 1630
rect 42830 1510 42875 1630
rect 42995 1510 43040 1630
rect 43160 1510 43205 1630
rect 43325 1510 43370 1630
rect 43490 1510 43535 1630
rect 43655 1510 43700 1630
rect 43820 1510 43865 1630
rect 43985 1510 44030 1630
rect 44150 1510 44195 1630
rect 44315 1510 44360 1630
rect 44480 1510 44525 1630
rect 44645 1510 44690 1630
rect 44810 1510 44855 1630
rect 44975 1510 45020 1630
rect 45140 1510 45185 1630
rect 45305 1510 45350 1630
rect 45470 1510 45515 1630
rect 45635 1510 45680 1630
rect 45800 1510 45845 1630
rect 45965 1510 46010 1630
rect 46130 1510 46175 1630
rect 46295 1510 46340 1630
rect 46460 1510 46505 1630
rect 46625 1510 46670 1630
rect 46790 1510 46835 1630
rect 46955 1510 47000 1630
rect 47120 1510 47165 1630
rect 47285 1510 47330 1630
rect 47450 1510 47495 1630
rect 47615 1510 47905 1630
rect 48025 1510 48070 1630
rect 48190 1510 48235 1630
rect 48355 1510 48400 1630
rect 48520 1510 48565 1630
rect 48685 1510 48730 1630
rect 48850 1510 48895 1630
rect 49015 1510 49060 1630
rect 49180 1510 49225 1630
rect 49345 1510 49390 1630
rect 49510 1510 49555 1630
rect 49675 1510 49720 1630
rect 49840 1510 49885 1630
rect 50005 1510 50050 1630
rect 50170 1510 50215 1630
rect 50335 1510 50380 1630
rect 50500 1510 50545 1630
rect 50665 1510 50710 1630
rect 50830 1510 50875 1630
rect 50995 1510 51040 1630
rect 51160 1510 51205 1630
rect 51325 1510 51370 1630
rect 51490 1510 51535 1630
rect 51655 1510 51700 1630
rect 51820 1510 51865 1630
rect 51985 1510 52030 1630
rect 52150 1510 52195 1630
rect 52315 1510 52360 1630
rect 52480 1510 52525 1630
rect 52645 1510 52690 1630
rect 52810 1510 52855 1630
rect 52975 1510 53020 1630
rect 53140 1510 53185 1630
rect 53305 1510 53370 1630
rect 30770 1495 53370 1510
rect 36300 1490 36460 1495
rect 41990 1490 42150 1495
rect 47680 1490 47840 1495
rect 30770 1420 53370 1445
rect 30770 1300 30795 1420
rect 30915 1300 30970 1420
rect 31090 1300 31135 1420
rect 31255 1300 31300 1420
rect 31420 1300 31465 1420
rect 31585 1300 31640 1420
rect 31760 1300 31805 1420
rect 31925 1300 31970 1420
rect 32090 1300 32135 1420
rect 32255 1300 32310 1420
rect 32430 1300 32475 1420
rect 32595 1300 32640 1420
rect 32760 1300 32805 1420
rect 32925 1300 32980 1420
rect 33100 1300 33145 1420
rect 33265 1300 33310 1420
rect 33430 1300 33475 1420
rect 33595 1300 33650 1420
rect 33770 1300 33815 1420
rect 33935 1300 33980 1420
rect 34100 1300 34145 1420
rect 34265 1300 34320 1420
rect 34440 1300 34485 1420
rect 34605 1300 34650 1420
rect 34770 1300 34815 1420
rect 34935 1300 34990 1420
rect 35110 1300 35155 1420
rect 35275 1300 35320 1420
rect 35440 1300 35485 1420
rect 35605 1300 35660 1420
rect 35780 1300 35825 1420
rect 35945 1300 35990 1420
rect 36110 1300 36155 1420
rect 36275 1300 36485 1420
rect 36605 1300 36660 1420
rect 36780 1300 36825 1420
rect 36945 1300 36990 1420
rect 37110 1300 37155 1420
rect 37275 1300 37330 1420
rect 37450 1300 37495 1420
rect 37615 1300 37660 1420
rect 37780 1300 37825 1420
rect 37945 1300 38000 1420
rect 38120 1300 38165 1420
rect 38285 1300 38330 1420
rect 38450 1300 38495 1420
rect 38615 1300 38670 1420
rect 38790 1300 38835 1420
rect 38955 1300 39000 1420
rect 39120 1300 39165 1420
rect 39285 1300 39340 1420
rect 39460 1300 39505 1420
rect 39625 1300 39670 1420
rect 39790 1300 39835 1420
rect 39955 1300 40010 1420
rect 40130 1300 40175 1420
rect 40295 1300 40340 1420
rect 40460 1300 40505 1420
rect 40625 1300 40680 1420
rect 40800 1300 40845 1420
rect 40965 1300 41010 1420
rect 41130 1300 41175 1420
rect 41295 1300 41350 1420
rect 41470 1300 41515 1420
rect 41635 1300 41680 1420
rect 41800 1300 41845 1420
rect 41965 1300 42175 1420
rect 42295 1300 42350 1420
rect 42470 1300 42515 1420
rect 42635 1300 42680 1420
rect 42800 1300 42845 1420
rect 42965 1300 43020 1420
rect 43140 1300 43185 1420
rect 43305 1300 43350 1420
rect 43470 1300 43515 1420
rect 43635 1300 43690 1420
rect 43810 1300 43855 1420
rect 43975 1300 44020 1420
rect 44140 1300 44185 1420
rect 44305 1300 44360 1420
rect 44480 1300 44525 1420
rect 44645 1300 44690 1420
rect 44810 1300 44855 1420
rect 44975 1300 45030 1420
rect 45150 1300 45195 1420
rect 45315 1300 45360 1420
rect 45480 1300 45525 1420
rect 45645 1300 45700 1420
rect 45820 1300 45865 1420
rect 45985 1300 46030 1420
rect 46150 1300 46195 1420
rect 46315 1300 46370 1420
rect 46490 1300 46535 1420
rect 46655 1300 46700 1420
rect 46820 1300 46865 1420
rect 46985 1300 47040 1420
rect 47160 1300 47205 1420
rect 47325 1300 47370 1420
rect 47490 1300 47535 1420
rect 47655 1300 47865 1420
rect 47985 1300 48040 1420
rect 48160 1300 48205 1420
rect 48325 1300 48370 1420
rect 48490 1300 48535 1420
rect 48655 1300 48710 1420
rect 48830 1300 48875 1420
rect 48995 1300 49040 1420
rect 49160 1300 49205 1420
rect 49325 1300 49380 1420
rect 49500 1300 49545 1420
rect 49665 1300 49710 1420
rect 49830 1300 49875 1420
rect 49995 1300 50050 1420
rect 50170 1300 50215 1420
rect 50335 1300 50380 1420
rect 50500 1300 50545 1420
rect 50665 1300 50720 1420
rect 50840 1300 50885 1420
rect 51005 1300 51050 1420
rect 51170 1300 51215 1420
rect 51335 1300 51390 1420
rect 51510 1300 51555 1420
rect 51675 1300 51720 1420
rect 51840 1300 51885 1420
rect 52005 1300 52060 1420
rect 52180 1300 52225 1420
rect 52345 1300 52390 1420
rect 52510 1300 52555 1420
rect 52675 1300 52730 1420
rect 52850 1300 52895 1420
rect 53015 1300 53060 1420
rect 53180 1300 53225 1420
rect 53345 1300 53370 1420
rect 30770 1255 53370 1300
rect 30770 1135 30795 1255
rect 30915 1135 30970 1255
rect 31090 1135 31135 1255
rect 31255 1135 31300 1255
rect 31420 1135 31465 1255
rect 31585 1135 31640 1255
rect 31760 1135 31805 1255
rect 31925 1135 31970 1255
rect 32090 1135 32135 1255
rect 32255 1135 32310 1255
rect 32430 1135 32475 1255
rect 32595 1135 32640 1255
rect 32760 1135 32805 1255
rect 32925 1135 32980 1255
rect 33100 1135 33145 1255
rect 33265 1135 33310 1255
rect 33430 1135 33475 1255
rect 33595 1135 33650 1255
rect 33770 1135 33815 1255
rect 33935 1135 33980 1255
rect 34100 1135 34145 1255
rect 34265 1135 34320 1255
rect 34440 1135 34485 1255
rect 34605 1135 34650 1255
rect 34770 1135 34815 1255
rect 34935 1135 34990 1255
rect 35110 1135 35155 1255
rect 35275 1135 35320 1255
rect 35440 1135 35485 1255
rect 35605 1135 35660 1255
rect 35780 1135 35825 1255
rect 35945 1135 35990 1255
rect 36110 1135 36155 1255
rect 36275 1135 36485 1255
rect 36605 1135 36660 1255
rect 36780 1135 36825 1255
rect 36945 1135 36990 1255
rect 37110 1135 37155 1255
rect 37275 1135 37330 1255
rect 37450 1135 37495 1255
rect 37615 1135 37660 1255
rect 37780 1135 37825 1255
rect 37945 1135 38000 1255
rect 38120 1135 38165 1255
rect 38285 1135 38330 1255
rect 38450 1135 38495 1255
rect 38615 1135 38670 1255
rect 38790 1135 38835 1255
rect 38955 1135 39000 1255
rect 39120 1135 39165 1255
rect 39285 1135 39340 1255
rect 39460 1135 39505 1255
rect 39625 1135 39670 1255
rect 39790 1135 39835 1255
rect 39955 1135 40010 1255
rect 40130 1135 40175 1255
rect 40295 1135 40340 1255
rect 40460 1135 40505 1255
rect 40625 1135 40680 1255
rect 40800 1135 40845 1255
rect 40965 1135 41010 1255
rect 41130 1135 41175 1255
rect 41295 1135 41350 1255
rect 41470 1135 41515 1255
rect 41635 1135 41680 1255
rect 41800 1135 41845 1255
rect 41965 1135 42175 1255
rect 42295 1135 42350 1255
rect 42470 1135 42515 1255
rect 42635 1135 42680 1255
rect 42800 1135 42845 1255
rect 42965 1135 43020 1255
rect 43140 1135 43185 1255
rect 43305 1135 43350 1255
rect 43470 1135 43515 1255
rect 43635 1135 43690 1255
rect 43810 1135 43855 1255
rect 43975 1135 44020 1255
rect 44140 1135 44185 1255
rect 44305 1135 44360 1255
rect 44480 1135 44525 1255
rect 44645 1135 44690 1255
rect 44810 1135 44855 1255
rect 44975 1135 45030 1255
rect 45150 1135 45195 1255
rect 45315 1135 45360 1255
rect 45480 1135 45525 1255
rect 45645 1135 45700 1255
rect 45820 1135 45865 1255
rect 45985 1135 46030 1255
rect 46150 1135 46195 1255
rect 46315 1135 46370 1255
rect 46490 1135 46535 1255
rect 46655 1135 46700 1255
rect 46820 1135 46865 1255
rect 46985 1135 47040 1255
rect 47160 1135 47205 1255
rect 47325 1135 47370 1255
rect 47490 1135 47535 1255
rect 47655 1135 47865 1255
rect 47985 1135 48040 1255
rect 48160 1135 48205 1255
rect 48325 1135 48370 1255
rect 48490 1135 48535 1255
rect 48655 1135 48710 1255
rect 48830 1135 48875 1255
rect 48995 1135 49040 1255
rect 49160 1135 49205 1255
rect 49325 1135 49380 1255
rect 49500 1135 49545 1255
rect 49665 1135 49710 1255
rect 49830 1135 49875 1255
rect 49995 1135 50050 1255
rect 50170 1135 50215 1255
rect 50335 1135 50380 1255
rect 50500 1135 50545 1255
rect 50665 1135 50720 1255
rect 50840 1135 50885 1255
rect 51005 1135 51050 1255
rect 51170 1135 51215 1255
rect 51335 1135 51390 1255
rect 51510 1135 51555 1255
rect 51675 1135 51720 1255
rect 51840 1135 51885 1255
rect 52005 1135 52060 1255
rect 52180 1135 52225 1255
rect 52345 1135 52390 1255
rect 52510 1135 52555 1255
rect 52675 1135 52730 1255
rect 52850 1135 52895 1255
rect 53015 1135 53060 1255
rect 53180 1135 53225 1255
rect 53345 1135 53370 1255
rect 30770 1090 53370 1135
rect 30770 970 30795 1090
rect 30915 970 30970 1090
rect 31090 970 31135 1090
rect 31255 970 31300 1090
rect 31420 970 31465 1090
rect 31585 970 31640 1090
rect 31760 970 31805 1090
rect 31925 970 31970 1090
rect 32090 970 32135 1090
rect 32255 970 32310 1090
rect 32430 970 32475 1090
rect 32595 970 32640 1090
rect 32760 970 32805 1090
rect 32925 970 32980 1090
rect 33100 970 33145 1090
rect 33265 970 33310 1090
rect 33430 970 33475 1090
rect 33595 970 33650 1090
rect 33770 970 33815 1090
rect 33935 970 33980 1090
rect 34100 970 34145 1090
rect 34265 970 34320 1090
rect 34440 970 34485 1090
rect 34605 970 34650 1090
rect 34770 970 34815 1090
rect 34935 970 34990 1090
rect 35110 970 35155 1090
rect 35275 970 35320 1090
rect 35440 970 35485 1090
rect 35605 970 35660 1090
rect 35780 970 35825 1090
rect 35945 970 35990 1090
rect 36110 970 36155 1090
rect 36275 970 36485 1090
rect 36605 970 36660 1090
rect 36780 970 36825 1090
rect 36945 970 36990 1090
rect 37110 970 37155 1090
rect 37275 970 37330 1090
rect 37450 970 37495 1090
rect 37615 970 37660 1090
rect 37780 970 37825 1090
rect 37945 970 38000 1090
rect 38120 970 38165 1090
rect 38285 970 38330 1090
rect 38450 970 38495 1090
rect 38615 970 38670 1090
rect 38790 970 38835 1090
rect 38955 970 39000 1090
rect 39120 970 39165 1090
rect 39285 970 39340 1090
rect 39460 970 39505 1090
rect 39625 970 39670 1090
rect 39790 970 39835 1090
rect 39955 970 40010 1090
rect 40130 970 40175 1090
rect 40295 970 40340 1090
rect 40460 970 40505 1090
rect 40625 970 40680 1090
rect 40800 970 40845 1090
rect 40965 970 41010 1090
rect 41130 970 41175 1090
rect 41295 970 41350 1090
rect 41470 970 41515 1090
rect 41635 970 41680 1090
rect 41800 970 41845 1090
rect 41965 970 42175 1090
rect 42295 970 42350 1090
rect 42470 970 42515 1090
rect 42635 970 42680 1090
rect 42800 970 42845 1090
rect 42965 970 43020 1090
rect 43140 970 43185 1090
rect 43305 970 43350 1090
rect 43470 970 43515 1090
rect 43635 970 43690 1090
rect 43810 970 43855 1090
rect 43975 970 44020 1090
rect 44140 970 44185 1090
rect 44305 970 44360 1090
rect 44480 970 44525 1090
rect 44645 970 44690 1090
rect 44810 970 44855 1090
rect 44975 970 45030 1090
rect 45150 970 45195 1090
rect 45315 970 45360 1090
rect 45480 970 45525 1090
rect 45645 970 45700 1090
rect 45820 970 45865 1090
rect 45985 970 46030 1090
rect 46150 970 46195 1090
rect 46315 970 46370 1090
rect 46490 970 46535 1090
rect 46655 970 46700 1090
rect 46820 970 46865 1090
rect 46985 970 47040 1090
rect 47160 970 47205 1090
rect 47325 970 47370 1090
rect 47490 970 47535 1090
rect 47655 970 47865 1090
rect 47985 970 48040 1090
rect 48160 970 48205 1090
rect 48325 970 48370 1090
rect 48490 970 48535 1090
rect 48655 970 48710 1090
rect 48830 970 48875 1090
rect 48995 970 49040 1090
rect 49160 970 49205 1090
rect 49325 970 49380 1090
rect 49500 970 49545 1090
rect 49665 970 49710 1090
rect 49830 970 49875 1090
rect 49995 970 50050 1090
rect 50170 970 50215 1090
rect 50335 970 50380 1090
rect 50500 970 50545 1090
rect 50665 970 50720 1090
rect 50840 970 50885 1090
rect 51005 970 51050 1090
rect 51170 970 51215 1090
rect 51335 970 51390 1090
rect 51510 970 51555 1090
rect 51675 970 51720 1090
rect 51840 970 51885 1090
rect 52005 970 52060 1090
rect 52180 970 52225 1090
rect 52345 970 52390 1090
rect 52510 970 52555 1090
rect 52675 970 52730 1090
rect 52850 970 52895 1090
rect 53015 970 53060 1090
rect 53180 970 53225 1090
rect 53345 970 53370 1090
rect 30770 925 53370 970
rect 30770 805 30795 925
rect 30915 805 30970 925
rect 31090 805 31135 925
rect 31255 805 31300 925
rect 31420 805 31465 925
rect 31585 805 31640 925
rect 31760 805 31805 925
rect 31925 805 31970 925
rect 32090 805 32135 925
rect 32255 805 32310 925
rect 32430 805 32475 925
rect 32595 805 32640 925
rect 32760 805 32805 925
rect 32925 805 32980 925
rect 33100 805 33145 925
rect 33265 805 33310 925
rect 33430 805 33475 925
rect 33595 805 33650 925
rect 33770 805 33815 925
rect 33935 805 33980 925
rect 34100 805 34145 925
rect 34265 805 34320 925
rect 34440 805 34485 925
rect 34605 805 34650 925
rect 34770 805 34815 925
rect 34935 805 34990 925
rect 35110 805 35155 925
rect 35275 805 35320 925
rect 35440 805 35485 925
rect 35605 805 35660 925
rect 35780 805 35825 925
rect 35945 805 35990 925
rect 36110 805 36155 925
rect 36275 805 36485 925
rect 36605 805 36660 925
rect 36780 805 36825 925
rect 36945 805 36990 925
rect 37110 805 37155 925
rect 37275 805 37330 925
rect 37450 805 37495 925
rect 37615 805 37660 925
rect 37780 805 37825 925
rect 37945 805 38000 925
rect 38120 805 38165 925
rect 38285 805 38330 925
rect 38450 805 38495 925
rect 38615 805 38670 925
rect 38790 805 38835 925
rect 38955 805 39000 925
rect 39120 805 39165 925
rect 39285 805 39340 925
rect 39460 805 39505 925
rect 39625 805 39670 925
rect 39790 805 39835 925
rect 39955 805 40010 925
rect 40130 805 40175 925
rect 40295 805 40340 925
rect 40460 805 40505 925
rect 40625 805 40680 925
rect 40800 805 40845 925
rect 40965 805 41010 925
rect 41130 805 41175 925
rect 41295 805 41350 925
rect 41470 805 41515 925
rect 41635 805 41680 925
rect 41800 805 41845 925
rect 41965 805 42175 925
rect 42295 805 42350 925
rect 42470 805 42515 925
rect 42635 805 42680 925
rect 42800 805 42845 925
rect 42965 805 43020 925
rect 43140 805 43185 925
rect 43305 805 43350 925
rect 43470 805 43515 925
rect 43635 805 43690 925
rect 43810 805 43855 925
rect 43975 805 44020 925
rect 44140 805 44185 925
rect 44305 805 44360 925
rect 44480 805 44525 925
rect 44645 805 44690 925
rect 44810 805 44855 925
rect 44975 805 45030 925
rect 45150 805 45195 925
rect 45315 805 45360 925
rect 45480 805 45525 925
rect 45645 805 45700 925
rect 45820 805 45865 925
rect 45985 805 46030 925
rect 46150 805 46195 925
rect 46315 805 46370 925
rect 46490 805 46535 925
rect 46655 805 46700 925
rect 46820 805 46865 925
rect 46985 805 47040 925
rect 47160 805 47205 925
rect 47325 805 47370 925
rect 47490 805 47535 925
rect 47655 805 47865 925
rect 47985 805 48040 925
rect 48160 805 48205 925
rect 48325 805 48370 925
rect 48490 805 48535 925
rect 48655 805 48710 925
rect 48830 805 48875 925
rect 48995 805 49040 925
rect 49160 805 49205 925
rect 49325 805 49380 925
rect 49500 805 49545 925
rect 49665 805 49710 925
rect 49830 805 49875 925
rect 49995 805 50050 925
rect 50170 805 50215 925
rect 50335 805 50380 925
rect 50500 805 50545 925
rect 50665 805 50720 925
rect 50840 805 50885 925
rect 51005 805 51050 925
rect 51170 805 51215 925
rect 51335 805 51390 925
rect 51510 805 51555 925
rect 51675 805 51720 925
rect 51840 805 51885 925
rect 52005 805 52060 925
rect 52180 805 52225 925
rect 52345 805 52390 925
rect 52510 805 52555 925
rect 52675 805 52730 925
rect 52850 805 52895 925
rect 53015 805 53060 925
rect 53180 805 53225 925
rect 53345 805 53370 925
rect 30770 750 53370 805
rect 30770 630 30795 750
rect 30915 630 30970 750
rect 31090 630 31135 750
rect 31255 630 31300 750
rect 31420 630 31465 750
rect 31585 630 31640 750
rect 31760 630 31805 750
rect 31925 630 31970 750
rect 32090 630 32135 750
rect 32255 630 32310 750
rect 32430 630 32475 750
rect 32595 630 32640 750
rect 32760 630 32805 750
rect 32925 630 32980 750
rect 33100 630 33145 750
rect 33265 630 33310 750
rect 33430 630 33475 750
rect 33595 630 33650 750
rect 33770 630 33815 750
rect 33935 630 33980 750
rect 34100 630 34145 750
rect 34265 630 34320 750
rect 34440 630 34485 750
rect 34605 630 34650 750
rect 34770 630 34815 750
rect 34935 630 34990 750
rect 35110 630 35155 750
rect 35275 630 35320 750
rect 35440 630 35485 750
rect 35605 630 35660 750
rect 35780 630 35825 750
rect 35945 630 35990 750
rect 36110 630 36155 750
rect 36275 630 36485 750
rect 36605 630 36660 750
rect 36780 630 36825 750
rect 36945 630 36990 750
rect 37110 630 37155 750
rect 37275 630 37330 750
rect 37450 630 37495 750
rect 37615 630 37660 750
rect 37780 630 37825 750
rect 37945 630 38000 750
rect 38120 630 38165 750
rect 38285 630 38330 750
rect 38450 630 38495 750
rect 38615 630 38670 750
rect 38790 630 38835 750
rect 38955 630 39000 750
rect 39120 630 39165 750
rect 39285 630 39340 750
rect 39460 630 39505 750
rect 39625 630 39670 750
rect 39790 630 39835 750
rect 39955 630 40010 750
rect 40130 630 40175 750
rect 40295 630 40340 750
rect 40460 630 40505 750
rect 40625 630 40680 750
rect 40800 630 40845 750
rect 40965 630 41010 750
rect 41130 630 41175 750
rect 41295 630 41350 750
rect 41470 630 41515 750
rect 41635 630 41680 750
rect 41800 630 41845 750
rect 41965 630 42175 750
rect 42295 630 42350 750
rect 42470 630 42515 750
rect 42635 630 42680 750
rect 42800 630 42845 750
rect 42965 630 43020 750
rect 43140 630 43185 750
rect 43305 630 43350 750
rect 43470 630 43515 750
rect 43635 630 43690 750
rect 43810 630 43855 750
rect 43975 630 44020 750
rect 44140 630 44185 750
rect 44305 630 44360 750
rect 44480 630 44525 750
rect 44645 630 44690 750
rect 44810 630 44855 750
rect 44975 630 45030 750
rect 45150 630 45195 750
rect 45315 630 45360 750
rect 45480 630 45525 750
rect 45645 630 45700 750
rect 45820 630 45865 750
rect 45985 630 46030 750
rect 46150 630 46195 750
rect 46315 630 46370 750
rect 46490 630 46535 750
rect 46655 630 46700 750
rect 46820 630 46865 750
rect 46985 630 47040 750
rect 47160 630 47205 750
rect 47325 630 47370 750
rect 47490 630 47535 750
rect 47655 630 47865 750
rect 47985 630 48040 750
rect 48160 630 48205 750
rect 48325 630 48370 750
rect 48490 630 48535 750
rect 48655 630 48710 750
rect 48830 630 48875 750
rect 48995 630 49040 750
rect 49160 630 49205 750
rect 49325 630 49380 750
rect 49500 630 49545 750
rect 49665 630 49710 750
rect 49830 630 49875 750
rect 49995 630 50050 750
rect 50170 630 50215 750
rect 50335 630 50380 750
rect 50500 630 50545 750
rect 50665 630 50720 750
rect 50840 630 50885 750
rect 51005 630 51050 750
rect 51170 630 51215 750
rect 51335 630 51390 750
rect 51510 630 51555 750
rect 51675 630 51720 750
rect 51840 630 51885 750
rect 52005 630 52060 750
rect 52180 630 52225 750
rect 52345 630 52390 750
rect 52510 630 52555 750
rect 52675 630 52730 750
rect 52850 630 52895 750
rect 53015 630 53060 750
rect 53180 630 53225 750
rect 53345 630 53370 750
rect 30770 585 53370 630
rect 30770 465 30795 585
rect 30915 465 30970 585
rect 31090 465 31135 585
rect 31255 465 31300 585
rect 31420 465 31465 585
rect 31585 465 31640 585
rect 31760 465 31805 585
rect 31925 465 31970 585
rect 32090 465 32135 585
rect 32255 465 32310 585
rect 32430 465 32475 585
rect 32595 465 32640 585
rect 32760 465 32805 585
rect 32925 465 32980 585
rect 33100 465 33145 585
rect 33265 465 33310 585
rect 33430 465 33475 585
rect 33595 465 33650 585
rect 33770 465 33815 585
rect 33935 465 33980 585
rect 34100 465 34145 585
rect 34265 465 34320 585
rect 34440 465 34485 585
rect 34605 465 34650 585
rect 34770 465 34815 585
rect 34935 465 34990 585
rect 35110 465 35155 585
rect 35275 465 35320 585
rect 35440 465 35485 585
rect 35605 465 35660 585
rect 35780 465 35825 585
rect 35945 465 35990 585
rect 36110 465 36155 585
rect 36275 465 36485 585
rect 36605 465 36660 585
rect 36780 465 36825 585
rect 36945 465 36990 585
rect 37110 465 37155 585
rect 37275 465 37330 585
rect 37450 465 37495 585
rect 37615 465 37660 585
rect 37780 465 37825 585
rect 37945 465 38000 585
rect 38120 465 38165 585
rect 38285 465 38330 585
rect 38450 465 38495 585
rect 38615 465 38670 585
rect 38790 465 38835 585
rect 38955 465 39000 585
rect 39120 465 39165 585
rect 39285 465 39340 585
rect 39460 465 39505 585
rect 39625 465 39670 585
rect 39790 465 39835 585
rect 39955 465 40010 585
rect 40130 465 40175 585
rect 40295 465 40340 585
rect 40460 465 40505 585
rect 40625 465 40680 585
rect 40800 465 40845 585
rect 40965 465 41010 585
rect 41130 465 41175 585
rect 41295 465 41350 585
rect 41470 465 41515 585
rect 41635 465 41680 585
rect 41800 465 41845 585
rect 41965 465 42175 585
rect 42295 465 42350 585
rect 42470 465 42515 585
rect 42635 465 42680 585
rect 42800 465 42845 585
rect 42965 465 43020 585
rect 43140 465 43185 585
rect 43305 465 43350 585
rect 43470 465 43515 585
rect 43635 465 43690 585
rect 43810 465 43855 585
rect 43975 465 44020 585
rect 44140 465 44185 585
rect 44305 465 44360 585
rect 44480 465 44525 585
rect 44645 465 44690 585
rect 44810 465 44855 585
rect 44975 465 45030 585
rect 45150 465 45195 585
rect 45315 465 45360 585
rect 45480 465 45525 585
rect 45645 465 45700 585
rect 45820 465 45865 585
rect 45985 465 46030 585
rect 46150 465 46195 585
rect 46315 465 46370 585
rect 46490 465 46535 585
rect 46655 465 46700 585
rect 46820 465 46865 585
rect 46985 465 47040 585
rect 47160 465 47205 585
rect 47325 465 47370 585
rect 47490 465 47535 585
rect 47655 465 47865 585
rect 47985 465 48040 585
rect 48160 465 48205 585
rect 48325 465 48370 585
rect 48490 465 48535 585
rect 48655 465 48710 585
rect 48830 465 48875 585
rect 48995 465 49040 585
rect 49160 465 49205 585
rect 49325 465 49380 585
rect 49500 465 49545 585
rect 49665 465 49710 585
rect 49830 465 49875 585
rect 49995 465 50050 585
rect 50170 465 50215 585
rect 50335 465 50380 585
rect 50500 465 50545 585
rect 50665 465 50720 585
rect 50840 465 50885 585
rect 51005 465 51050 585
rect 51170 465 51215 585
rect 51335 465 51390 585
rect 51510 465 51555 585
rect 51675 465 51720 585
rect 51840 465 51885 585
rect 52005 465 52060 585
rect 52180 465 52225 585
rect 52345 465 52390 585
rect 52510 465 52555 585
rect 52675 465 52730 585
rect 52850 465 52895 585
rect 53015 465 53060 585
rect 53180 465 53225 585
rect 53345 465 53370 585
rect 30770 420 53370 465
rect 30770 300 30795 420
rect 30915 300 30970 420
rect 31090 300 31135 420
rect 31255 300 31300 420
rect 31420 300 31465 420
rect 31585 300 31640 420
rect 31760 300 31805 420
rect 31925 300 31970 420
rect 32090 300 32135 420
rect 32255 300 32310 420
rect 32430 300 32475 420
rect 32595 300 32640 420
rect 32760 300 32805 420
rect 32925 300 32980 420
rect 33100 300 33145 420
rect 33265 300 33310 420
rect 33430 300 33475 420
rect 33595 300 33650 420
rect 33770 300 33815 420
rect 33935 300 33980 420
rect 34100 300 34145 420
rect 34265 300 34320 420
rect 34440 300 34485 420
rect 34605 300 34650 420
rect 34770 300 34815 420
rect 34935 300 34990 420
rect 35110 300 35155 420
rect 35275 300 35320 420
rect 35440 300 35485 420
rect 35605 300 35660 420
rect 35780 300 35825 420
rect 35945 300 35990 420
rect 36110 300 36155 420
rect 36275 300 36485 420
rect 36605 300 36660 420
rect 36780 300 36825 420
rect 36945 300 36990 420
rect 37110 300 37155 420
rect 37275 300 37330 420
rect 37450 300 37495 420
rect 37615 300 37660 420
rect 37780 300 37825 420
rect 37945 300 38000 420
rect 38120 300 38165 420
rect 38285 300 38330 420
rect 38450 300 38495 420
rect 38615 300 38670 420
rect 38790 300 38835 420
rect 38955 300 39000 420
rect 39120 300 39165 420
rect 39285 300 39340 420
rect 39460 300 39505 420
rect 39625 300 39670 420
rect 39790 300 39835 420
rect 39955 300 40010 420
rect 40130 300 40175 420
rect 40295 300 40340 420
rect 40460 300 40505 420
rect 40625 300 40680 420
rect 40800 300 40845 420
rect 40965 300 41010 420
rect 41130 300 41175 420
rect 41295 300 41350 420
rect 41470 300 41515 420
rect 41635 300 41680 420
rect 41800 300 41845 420
rect 41965 300 42175 420
rect 42295 300 42350 420
rect 42470 300 42515 420
rect 42635 300 42680 420
rect 42800 300 42845 420
rect 42965 300 43020 420
rect 43140 300 43185 420
rect 43305 300 43350 420
rect 43470 300 43515 420
rect 43635 300 43690 420
rect 43810 300 43855 420
rect 43975 300 44020 420
rect 44140 300 44185 420
rect 44305 300 44360 420
rect 44480 300 44525 420
rect 44645 300 44690 420
rect 44810 300 44855 420
rect 44975 300 45030 420
rect 45150 300 45195 420
rect 45315 300 45360 420
rect 45480 300 45525 420
rect 45645 300 45700 420
rect 45820 300 45865 420
rect 45985 300 46030 420
rect 46150 300 46195 420
rect 46315 300 46370 420
rect 46490 300 46535 420
rect 46655 300 46700 420
rect 46820 300 46865 420
rect 46985 300 47040 420
rect 47160 300 47205 420
rect 47325 300 47370 420
rect 47490 300 47535 420
rect 47655 300 47865 420
rect 47985 300 48040 420
rect 48160 300 48205 420
rect 48325 300 48370 420
rect 48490 300 48535 420
rect 48655 300 48710 420
rect 48830 300 48875 420
rect 48995 300 49040 420
rect 49160 300 49205 420
rect 49325 300 49380 420
rect 49500 300 49545 420
rect 49665 300 49710 420
rect 49830 300 49875 420
rect 49995 300 50050 420
rect 50170 300 50215 420
rect 50335 300 50380 420
rect 50500 300 50545 420
rect 50665 300 50720 420
rect 50840 300 50885 420
rect 51005 300 51050 420
rect 51170 300 51215 420
rect 51335 300 51390 420
rect 51510 300 51555 420
rect 51675 300 51720 420
rect 51840 300 51885 420
rect 52005 300 52060 420
rect 52180 300 52225 420
rect 52345 300 52390 420
rect 52510 300 52555 420
rect 52675 300 52730 420
rect 52850 300 52895 420
rect 53015 300 53060 420
rect 53180 300 53225 420
rect 53345 300 53370 420
rect 30770 255 53370 300
rect 30770 135 30795 255
rect 30915 135 30970 255
rect 31090 135 31135 255
rect 31255 135 31300 255
rect 31420 135 31465 255
rect 31585 135 31640 255
rect 31760 135 31805 255
rect 31925 135 31970 255
rect 32090 135 32135 255
rect 32255 135 32310 255
rect 32430 135 32475 255
rect 32595 135 32640 255
rect 32760 135 32805 255
rect 32925 135 32980 255
rect 33100 135 33145 255
rect 33265 135 33310 255
rect 33430 135 33475 255
rect 33595 135 33650 255
rect 33770 135 33815 255
rect 33935 135 33980 255
rect 34100 135 34145 255
rect 34265 135 34320 255
rect 34440 135 34485 255
rect 34605 135 34650 255
rect 34770 135 34815 255
rect 34935 135 34990 255
rect 35110 135 35155 255
rect 35275 135 35320 255
rect 35440 135 35485 255
rect 35605 135 35660 255
rect 35780 135 35825 255
rect 35945 135 35990 255
rect 36110 135 36155 255
rect 36275 135 36485 255
rect 36605 135 36660 255
rect 36780 135 36825 255
rect 36945 135 36990 255
rect 37110 135 37155 255
rect 37275 135 37330 255
rect 37450 135 37495 255
rect 37615 135 37660 255
rect 37780 135 37825 255
rect 37945 135 38000 255
rect 38120 135 38165 255
rect 38285 135 38330 255
rect 38450 135 38495 255
rect 38615 135 38670 255
rect 38790 135 38835 255
rect 38955 135 39000 255
rect 39120 135 39165 255
rect 39285 135 39340 255
rect 39460 135 39505 255
rect 39625 135 39670 255
rect 39790 135 39835 255
rect 39955 135 40010 255
rect 40130 135 40175 255
rect 40295 135 40340 255
rect 40460 135 40505 255
rect 40625 135 40680 255
rect 40800 135 40845 255
rect 40965 135 41010 255
rect 41130 135 41175 255
rect 41295 135 41350 255
rect 41470 135 41515 255
rect 41635 135 41680 255
rect 41800 135 41845 255
rect 41965 135 42175 255
rect 42295 135 42350 255
rect 42470 135 42515 255
rect 42635 135 42680 255
rect 42800 135 42845 255
rect 42965 135 43020 255
rect 43140 135 43185 255
rect 43305 135 43350 255
rect 43470 135 43515 255
rect 43635 135 43690 255
rect 43810 135 43855 255
rect 43975 135 44020 255
rect 44140 135 44185 255
rect 44305 135 44360 255
rect 44480 135 44525 255
rect 44645 135 44690 255
rect 44810 135 44855 255
rect 44975 135 45030 255
rect 45150 135 45195 255
rect 45315 135 45360 255
rect 45480 135 45525 255
rect 45645 135 45700 255
rect 45820 135 45865 255
rect 45985 135 46030 255
rect 46150 135 46195 255
rect 46315 135 46370 255
rect 46490 135 46535 255
rect 46655 135 46700 255
rect 46820 135 46865 255
rect 46985 135 47040 255
rect 47160 135 47205 255
rect 47325 135 47370 255
rect 47490 135 47535 255
rect 47655 135 47865 255
rect 47985 135 48040 255
rect 48160 135 48205 255
rect 48325 135 48370 255
rect 48490 135 48535 255
rect 48655 135 48710 255
rect 48830 135 48875 255
rect 48995 135 49040 255
rect 49160 135 49205 255
rect 49325 135 49380 255
rect 49500 135 49545 255
rect 49665 135 49710 255
rect 49830 135 49875 255
rect 49995 135 50050 255
rect 50170 135 50215 255
rect 50335 135 50380 255
rect 50500 135 50545 255
rect 50665 135 50720 255
rect 50840 135 50885 255
rect 51005 135 51050 255
rect 51170 135 51215 255
rect 51335 135 51390 255
rect 51510 135 51555 255
rect 51675 135 51720 255
rect 51840 135 51885 255
rect 52005 135 52060 255
rect 52180 135 52225 255
rect 52345 135 52390 255
rect 52510 135 52555 255
rect 52675 135 52730 255
rect 52850 135 52895 255
rect 53015 135 53060 255
rect 53180 135 53225 255
rect 53345 135 53370 255
rect 30770 80 53370 135
rect 30770 -40 30795 80
rect 30915 -40 30970 80
rect 31090 -40 31135 80
rect 31255 -40 31300 80
rect 31420 -40 31465 80
rect 31585 -40 31640 80
rect 31760 -40 31805 80
rect 31925 -40 31970 80
rect 32090 -40 32135 80
rect 32255 -40 32310 80
rect 32430 -40 32475 80
rect 32595 -40 32640 80
rect 32760 -40 32805 80
rect 32925 -40 32980 80
rect 33100 -40 33145 80
rect 33265 -40 33310 80
rect 33430 -40 33475 80
rect 33595 -40 33650 80
rect 33770 -40 33815 80
rect 33935 -40 33980 80
rect 34100 -40 34145 80
rect 34265 -40 34320 80
rect 34440 -40 34485 80
rect 34605 -40 34650 80
rect 34770 -40 34815 80
rect 34935 -40 34990 80
rect 35110 -40 35155 80
rect 35275 -40 35320 80
rect 35440 -40 35485 80
rect 35605 -40 35660 80
rect 35780 -40 35825 80
rect 35945 -40 35990 80
rect 36110 -40 36155 80
rect 36275 -40 36485 80
rect 36605 -40 36660 80
rect 36780 -40 36825 80
rect 36945 -40 36990 80
rect 37110 -40 37155 80
rect 37275 -40 37330 80
rect 37450 -40 37495 80
rect 37615 -40 37660 80
rect 37780 -40 37825 80
rect 37945 -40 38000 80
rect 38120 -40 38165 80
rect 38285 -40 38330 80
rect 38450 -40 38495 80
rect 38615 -40 38670 80
rect 38790 -40 38835 80
rect 38955 -40 39000 80
rect 39120 -40 39165 80
rect 39285 -40 39340 80
rect 39460 -40 39505 80
rect 39625 -40 39670 80
rect 39790 -40 39835 80
rect 39955 -40 40010 80
rect 40130 -40 40175 80
rect 40295 -40 40340 80
rect 40460 -40 40505 80
rect 40625 -40 40680 80
rect 40800 -40 40845 80
rect 40965 -40 41010 80
rect 41130 -40 41175 80
rect 41295 -40 41350 80
rect 41470 -40 41515 80
rect 41635 -40 41680 80
rect 41800 -40 41845 80
rect 41965 -40 42175 80
rect 42295 -40 42350 80
rect 42470 -40 42515 80
rect 42635 -40 42680 80
rect 42800 -40 42845 80
rect 42965 -40 43020 80
rect 43140 -40 43185 80
rect 43305 -40 43350 80
rect 43470 -40 43515 80
rect 43635 -40 43690 80
rect 43810 -40 43855 80
rect 43975 -40 44020 80
rect 44140 -40 44185 80
rect 44305 -40 44360 80
rect 44480 -40 44525 80
rect 44645 -40 44690 80
rect 44810 -40 44855 80
rect 44975 -40 45030 80
rect 45150 -40 45195 80
rect 45315 -40 45360 80
rect 45480 -40 45525 80
rect 45645 -40 45700 80
rect 45820 -40 45865 80
rect 45985 -40 46030 80
rect 46150 -40 46195 80
rect 46315 -40 46370 80
rect 46490 -40 46535 80
rect 46655 -40 46700 80
rect 46820 -40 46865 80
rect 46985 -40 47040 80
rect 47160 -40 47205 80
rect 47325 -40 47370 80
rect 47490 -40 47535 80
rect 47655 -40 47865 80
rect 47985 -40 48040 80
rect 48160 -40 48205 80
rect 48325 -40 48370 80
rect 48490 -40 48535 80
rect 48655 -40 48710 80
rect 48830 -40 48875 80
rect 48995 -40 49040 80
rect 49160 -40 49205 80
rect 49325 -40 49380 80
rect 49500 -40 49545 80
rect 49665 -40 49710 80
rect 49830 -40 49875 80
rect 49995 -40 50050 80
rect 50170 -40 50215 80
rect 50335 -40 50380 80
rect 50500 -40 50545 80
rect 50665 -40 50720 80
rect 50840 -40 50885 80
rect 51005 -40 51050 80
rect 51170 -40 51215 80
rect 51335 -40 51390 80
rect 51510 -40 51555 80
rect 51675 -40 51720 80
rect 51840 -40 51885 80
rect 52005 -40 52060 80
rect 52180 -40 52225 80
rect 52345 -40 52390 80
rect 52510 -40 52555 80
rect 52675 -40 52730 80
rect 52850 -40 52895 80
rect 53015 -40 53060 80
rect 53180 -40 53225 80
rect 53345 -40 53370 80
rect 30770 -85 53370 -40
rect 30770 -205 30795 -85
rect 30915 -205 30970 -85
rect 31090 -205 31135 -85
rect 31255 -205 31300 -85
rect 31420 -205 31465 -85
rect 31585 -205 31640 -85
rect 31760 -205 31805 -85
rect 31925 -205 31970 -85
rect 32090 -205 32135 -85
rect 32255 -205 32310 -85
rect 32430 -205 32475 -85
rect 32595 -205 32640 -85
rect 32760 -205 32805 -85
rect 32925 -205 32980 -85
rect 33100 -205 33145 -85
rect 33265 -205 33310 -85
rect 33430 -205 33475 -85
rect 33595 -205 33650 -85
rect 33770 -205 33815 -85
rect 33935 -205 33980 -85
rect 34100 -205 34145 -85
rect 34265 -205 34320 -85
rect 34440 -205 34485 -85
rect 34605 -205 34650 -85
rect 34770 -205 34815 -85
rect 34935 -205 34990 -85
rect 35110 -205 35155 -85
rect 35275 -205 35320 -85
rect 35440 -205 35485 -85
rect 35605 -205 35660 -85
rect 35780 -205 35825 -85
rect 35945 -205 35990 -85
rect 36110 -205 36155 -85
rect 36275 -205 36485 -85
rect 36605 -205 36660 -85
rect 36780 -205 36825 -85
rect 36945 -205 36990 -85
rect 37110 -205 37155 -85
rect 37275 -205 37330 -85
rect 37450 -205 37495 -85
rect 37615 -205 37660 -85
rect 37780 -205 37825 -85
rect 37945 -205 38000 -85
rect 38120 -205 38165 -85
rect 38285 -205 38330 -85
rect 38450 -205 38495 -85
rect 38615 -205 38670 -85
rect 38790 -205 38835 -85
rect 38955 -205 39000 -85
rect 39120 -205 39165 -85
rect 39285 -205 39340 -85
rect 39460 -205 39505 -85
rect 39625 -205 39670 -85
rect 39790 -205 39835 -85
rect 39955 -205 40010 -85
rect 40130 -205 40175 -85
rect 40295 -205 40340 -85
rect 40460 -205 40505 -85
rect 40625 -205 40680 -85
rect 40800 -205 40845 -85
rect 40965 -205 41010 -85
rect 41130 -205 41175 -85
rect 41295 -205 41350 -85
rect 41470 -205 41515 -85
rect 41635 -205 41680 -85
rect 41800 -205 41845 -85
rect 41965 -205 42175 -85
rect 42295 -205 42350 -85
rect 42470 -205 42515 -85
rect 42635 -205 42680 -85
rect 42800 -205 42845 -85
rect 42965 -205 43020 -85
rect 43140 -205 43185 -85
rect 43305 -205 43350 -85
rect 43470 -205 43515 -85
rect 43635 -205 43690 -85
rect 43810 -205 43855 -85
rect 43975 -205 44020 -85
rect 44140 -205 44185 -85
rect 44305 -205 44360 -85
rect 44480 -205 44525 -85
rect 44645 -205 44690 -85
rect 44810 -205 44855 -85
rect 44975 -205 45030 -85
rect 45150 -205 45195 -85
rect 45315 -205 45360 -85
rect 45480 -205 45525 -85
rect 45645 -205 45700 -85
rect 45820 -205 45865 -85
rect 45985 -205 46030 -85
rect 46150 -205 46195 -85
rect 46315 -205 46370 -85
rect 46490 -205 46535 -85
rect 46655 -205 46700 -85
rect 46820 -205 46865 -85
rect 46985 -205 47040 -85
rect 47160 -205 47205 -85
rect 47325 -205 47370 -85
rect 47490 -205 47535 -85
rect 47655 -205 47865 -85
rect 47985 -205 48040 -85
rect 48160 -205 48205 -85
rect 48325 -205 48370 -85
rect 48490 -205 48535 -85
rect 48655 -205 48710 -85
rect 48830 -205 48875 -85
rect 48995 -205 49040 -85
rect 49160 -205 49205 -85
rect 49325 -205 49380 -85
rect 49500 -205 49545 -85
rect 49665 -205 49710 -85
rect 49830 -205 49875 -85
rect 49995 -205 50050 -85
rect 50170 -205 50215 -85
rect 50335 -205 50380 -85
rect 50500 -205 50545 -85
rect 50665 -205 50720 -85
rect 50840 -205 50885 -85
rect 51005 -205 51050 -85
rect 51170 -205 51215 -85
rect 51335 -205 51390 -85
rect 51510 -205 51555 -85
rect 51675 -205 51720 -85
rect 51840 -205 51885 -85
rect 52005 -205 52060 -85
rect 52180 -205 52225 -85
rect 52345 -205 52390 -85
rect 52510 -205 52555 -85
rect 52675 -205 52730 -85
rect 52850 -205 52895 -85
rect 53015 -205 53060 -85
rect 53180 -205 53225 -85
rect 53345 -205 53370 -85
rect 30770 -250 53370 -205
rect 30770 -370 30795 -250
rect 30915 -370 30970 -250
rect 31090 -370 31135 -250
rect 31255 -370 31300 -250
rect 31420 -370 31465 -250
rect 31585 -370 31640 -250
rect 31760 -370 31805 -250
rect 31925 -370 31970 -250
rect 32090 -370 32135 -250
rect 32255 -370 32310 -250
rect 32430 -370 32475 -250
rect 32595 -370 32640 -250
rect 32760 -370 32805 -250
rect 32925 -370 32980 -250
rect 33100 -370 33145 -250
rect 33265 -370 33310 -250
rect 33430 -370 33475 -250
rect 33595 -370 33650 -250
rect 33770 -370 33815 -250
rect 33935 -370 33980 -250
rect 34100 -370 34145 -250
rect 34265 -370 34320 -250
rect 34440 -370 34485 -250
rect 34605 -370 34650 -250
rect 34770 -370 34815 -250
rect 34935 -370 34990 -250
rect 35110 -370 35155 -250
rect 35275 -370 35320 -250
rect 35440 -370 35485 -250
rect 35605 -370 35660 -250
rect 35780 -370 35825 -250
rect 35945 -370 35990 -250
rect 36110 -370 36155 -250
rect 36275 -370 36485 -250
rect 36605 -370 36660 -250
rect 36780 -370 36825 -250
rect 36945 -370 36990 -250
rect 37110 -370 37155 -250
rect 37275 -370 37330 -250
rect 37450 -370 37495 -250
rect 37615 -370 37660 -250
rect 37780 -370 37825 -250
rect 37945 -370 38000 -250
rect 38120 -370 38165 -250
rect 38285 -370 38330 -250
rect 38450 -370 38495 -250
rect 38615 -370 38670 -250
rect 38790 -370 38835 -250
rect 38955 -370 39000 -250
rect 39120 -370 39165 -250
rect 39285 -370 39340 -250
rect 39460 -370 39505 -250
rect 39625 -370 39670 -250
rect 39790 -370 39835 -250
rect 39955 -370 40010 -250
rect 40130 -370 40175 -250
rect 40295 -370 40340 -250
rect 40460 -370 40505 -250
rect 40625 -370 40680 -250
rect 40800 -370 40845 -250
rect 40965 -370 41010 -250
rect 41130 -370 41175 -250
rect 41295 -370 41350 -250
rect 41470 -370 41515 -250
rect 41635 -370 41680 -250
rect 41800 -370 41845 -250
rect 41965 -370 42175 -250
rect 42295 -370 42350 -250
rect 42470 -370 42515 -250
rect 42635 -370 42680 -250
rect 42800 -370 42845 -250
rect 42965 -370 43020 -250
rect 43140 -370 43185 -250
rect 43305 -370 43350 -250
rect 43470 -370 43515 -250
rect 43635 -370 43690 -250
rect 43810 -370 43855 -250
rect 43975 -370 44020 -250
rect 44140 -370 44185 -250
rect 44305 -370 44360 -250
rect 44480 -370 44525 -250
rect 44645 -370 44690 -250
rect 44810 -370 44855 -250
rect 44975 -370 45030 -250
rect 45150 -370 45195 -250
rect 45315 -370 45360 -250
rect 45480 -370 45525 -250
rect 45645 -370 45700 -250
rect 45820 -370 45865 -250
rect 45985 -370 46030 -250
rect 46150 -370 46195 -250
rect 46315 -370 46370 -250
rect 46490 -370 46535 -250
rect 46655 -370 46700 -250
rect 46820 -370 46865 -250
rect 46985 -370 47040 -250
rect 47160 -370 47205 -250
rect 47325 -370 47370 -250
rect 47490 -370 47535 -250
rect 47655 -370 47865 -250
rect 47985 -370 48040 -250
rect 48160 -370 48205 -250
rect 48325 -370 48370 -250
rect 48490 -370 48535 -250
rect 48655 -370 48710 -250
rect 48830 -370 48875 -250
rect 48995 -370 49040 -250
rect 49160 -370 49205 -250
rect 49325 -370 49380 -250
rect 49500 -370 49545 -250
rect 49665 -370 49710 -250
rect 49830 -370 49875 -250
rect 49995 -370 50050 -250
rect 50170 -370 50215 -250
rect 50335 -370 50380 -250
rect 50500 -370 50545 -250
rect 50665 -370 50720 -250
rect 50840 -370 50885 -250
rect 51005 -370 51050 -250
rect 51170 -370 51215 -250
rect 51335 -370 51390 -250
rect 51510 -370 51555 -250
rect 51675 -370 51720 -250
rect 51840 -370 51885 -250
rect 52005 -370 52060 -250
rect 52180 -370 52225 -250
rect 52345 -370 52390 -250
rect 52510 -370 52555 -250
rect 52675 -370 52730 -250
rect 52850 -370 52895 -250
rect 53015 -370 53060 -250
rect 53180 -370 53225 -250
rect 53345 -370 53370 -250
rect 30770 -415 53370 -370
rect 30770 -535 30795 -415
rect 30915 -535 30970 -415
rect 31090 -535 31135 -415
rect 31255 -535 31300 -415
rect 31420 -535 31465 -415
rect 31585 -535 31640 -415
rect 31760 -535 31805 -415
rect 31925 -535 31970 -415
rect 32090 -535 32135 -415
rect 32255 -535 32310 -415
rect 32430 -535 32475 -415
rect 32595 -535 32640 -415
rect 32760 -535 32805 -415
rect 32925 -535 32980 -415
rect 33100 -535 33145 -415
rect 33265 -535 33310 -415
rect 33430 -535 33475 -415
rect 33595 -535 33650 -415
rect 33770 -535 33815 -415
rect 33935 -535 33980 -415
rect 34100 -535 34145 -415
rect 34265 -535 34320 -415
rect 34440 -535 34485 -415
rect 34605 -535 34650 -415
rect 34770 -535 34815 -415
rect 34935 -535 34990 -415
rect 35110 -535 35155 -415
rect 35275 -535 35320 -415
rect 35440 -535 35485 -415
rect 35605 -535 35660 -415
rect 35780 -535 35825 -415
rect 35945 -535 35990 -415
rect 36110 -535 36155 -415
rect 36275 -535 36485 -415
rect 36605 -535 36660 -415
rect 36780 -535 36825 -415
rect 36945 -535 36990 -415
rect 37110 -535 37155 -415
rect 37275 -535 37330 -415
rect 37450 -535 37495 -415
rect 37615 -535 37660 -415
rect 37780 -535 37825 -415
rect 37945 -535 38000 -415
rect 38120 -535 38165 -415
rect 38285 -535 38330 -415
rect 38450 -535 38495 -415
rect 38615 -535 38670 -415
rect 38790 -535 38835 -415
rect 38955 -535 39000 -415
rect 39120 -535 39165 -415
rect 39285 -535 39340 -415
rect 39460 -535 39505 -415
rect 39625 -535 39670 -415
rect 39790 -535 39835 -415
rect 39955 -535 40010 -415
rect 40130 -535 40175 -415
rect 40295 -535 40340 -415
rect 40460 -535 40505 -415
rect 40625 -535 40680 -415
rect 40800 -535 40845 -415
rect 40965 -535 41010 -415
rect 41130 -535 41175 -415
rect 41295 -535 41350 -415
rect 41470 -535 41515 -415
rect 41635 -535 41680 -415
rect 41800 -535 41845 -415
rect 41965 -535 42175 -415
rect 42295 -535 42350 -415
rect 42470 -535 42515 -415
rect 42635 -535 42680 -415
rect 42800 -535 42845 -415
rect 42965 -535 43020 -415
rect 43140 -535 43185 -415
rect 43305 -535 43350 -415
rect 43470 -535 43515 -415
rect 43635 -535 43690 -415
rect 43810 -535 43855 -415
rect 43975 -535 44020 -415
rect 44140 -535 44185 -415
rect 44305 -535 44360 -415
rect 44480 -535 44525 -415
rect 44645 -535 44690 -415
rect 44810 -535 44855 -415
rect 44975 -535 45030 -415
rect 45150 -535 45195 -415
rect 45315 -535 45360 -415
rect 45480 -535 45525 -415
rect 45645 -535 45700 -415
rect 45820 -535 45865 -415
rect 45985 -535 46030 -415
rect 46150 -535 46195 -415
rect 46315 -535 46370 -415
rect 46490 -535 46535 -415
rect 46655 -535 46700 -415
rect 46820 -535 46865 -415
rect 46985 -535 47040 -415
rect 47160 -535 47205 -415
rect 47325 -535 47370 -415
rect 47490 -535 47535 -415
rect 47655 -535 47865 -415
rect 47985 -535 48040 -415
rect 48160 -535 48205 -415
rect 48325 -535 48370 -415
rect 48490 -535 48535 -415
rect 48655 -535 48710 -415
rect 48830 -535 48875 -415
rect 48995 -535 49040 -415
rect 49160 -535 49205 -415
rect 49325 -535 49380 -415
rect 49500 -535 49545 -415
rect 49665 -535 49710 -415
rect 49830 -535 49875 -415
rect 49995 -535 50050 -415
rect 50170 -535 50215 -415
rect 50335 -535 50380 -415
rect 50500 -535 50545 -415
rect 50665 -535 50720 -415
rect 50840 -535 50885 -415
rect 51005 -535 51050 -415
rect 51170 -535 51215 -415
rect 51335 -535 51390 -415
rect 51510 -535 51555 -415
rect 51675 -535 51720 -415
rect 51840 -535 51885 -415
rect 52005 -535 52060 -415
rect 52180 -535 52225 -415
rect 52345 -535 52390 -415
rect 52510 -535 52555 -415
rect 52675 -535 52730 -415
rect 52850 -535 52895 -415
rect 53015 -535 53060 -415
rect 53180 -535 53225 -415
rect 53345 -535 53370 -415
rect 30770 -590 53370 -535
rect 30770 -710 30795 -590
rect 30915 -710 30970 -590
rect 31090 -710 31135 -590
rect 31255 -710 31300 -590
rect 31420 -710 31465 -590
rect 31585 -710 31640 -590
rect 31760 -710 31805 -590
rect 31925 -710 31970 -590
rect 32090 -710 32135 -590
rect 32255 -710 32310 -590
rect 32430 -710 32475 -590
rect 32595 -710 32640 -590
rect 32760 -710 32805 -590
rect 32925 -710 32980 -590
rect 33100 -710 33145 -590
rect 33265 -710 33310 -590
rect 33430 -710 33475 -590
rect 33595 -710 33650 -590
rect 33770 -710 33815 -590
rect 33935 -710 33980 -590
rect 34100 -710 34145 -590
rect 34265 -710 34320 -590
rect 34440 -710 34485 -590
rect 34605 -710 34650 -590
rect 34770 -710 34815 -590
rect 34935 -710 34990 -590
rect 35110 -710 35155 -590
rect 35275 -710 35320 -590
rect 35440 -710 35485 -590
rect 35605 -710 35660 -590
rect 35780 -710 35825 -590
rect 35945 -710 35990 -590
rect 36110 -710 36155 -590
rect 36275 -710 36485 -590
rect 36605 -710 36660 -590
rect 36780 -710 36825 -590
rect 36945 -710 36990 -590
rect 37110 -710 37155 -590
rect 37275 -710 37330 -590
rect 37450 -710 37495 -590
rect 37615 -710 37660 -590
rect 37780 -710 37825 -590
rect 37945 -710 38000 -590
rect 38120 -710 38165 -590
rect 38285 -710 38330 -590
rect 38450 -710 38495 -590
rect 38615 -710 38670 -590
rect 38790 -710 38835 -590
rect 38955 -710 39000 -590
rect 39120 -710 39165 -590
rect 39285 -710 39340 -590
rect 39460 -710 39505 -590
rect 39625 -710 39670 -590
rect 39790 -710 39835 -590
rect 39955 -710 40010 -590
rect 40130 -710 40175 -590
rect 40295 -710 40340 -590
rect 40460 -710 40505 -590
rect 40625 -710 40680 -590
rect 40800 -710 40845 -590
rect 40965 -710 41010 -590
rect 41130 -710 41175 -590
rect 41295 -710 41350 -590
rect 41470 -710 41515 -590
rect 41635 -710 41680 -590
rect 41800 -710 41845 -590
rect 41965 -710 42175 -590
rect 42295 -710 42350 -590
rect 42470 -710 42515 -590
rect 42635 -710 42680 -590
rect 42800 -710 42845 -590
rect 42965 -710 43020 -590
rect 43140 -710 43185 -590
rect 43305 -710 43350 -590
rect 43470 -710 43515 -590
rect 43635 -710 43690 -590
rect 43810 -710 43855 -590
rect 43975 -710 44020 -590
rect 44140 -710 44185 -590
rect 44305 -710 44360 -590
rect 44480 -710 44525 -590
rect 44645 -710 44690 -590
rect 44810 -710 44855 -590
rect 44975 -710 45030 -590
rect 45150 -710 45195 -590
rect 45315 -710 45360 -590
rect 45480 -710 45525 -590
rect 45645 -710 45700 -590
rect 45820 -710 45865 -590
rect 45985 -710 46030 -590
rect 46150 -710 46195 -590
rect 46315 -710 46370 -590
rect 46490 -710 46535 -590
rect 46655 -710 46700 -590
rect 46820 -710 46865 -590
rect 46985 -710 47040 -590
rect 47160 -710 47205 -590
rect 47325 -710 47370 -590
rect 47490 -710 47535 -590
rect 47655 -710 47865 -590
rect 47985 -710 48040 -590
rect 48160 -710 48205 -590
rect 48325 -710 48370 -590
rect 48490 -710 48535 -590
rect 48655 -710 48710 -590
rect 48830 -710 48875 -590
rect 48995 -710 49040 -590
rect 49160 -710 49205 -590
rect 49325 -710 49380 -590
rect 49500 -710 49545 -590
rect 49665 -710 49710 -590
rect 49830 -710 49875 -590
rect 49995 -710 50050 -590
rect 50170 -710 50215 -590
rect 50335 -710 50380 -590
rect 50500 -710 50545 -590
rect 50665 -710 50720 -590
rect 50840 -710 50885 -590
rect 51005 -710 51050 -590
rect 51170 -710 51215 -590
rect 51335 -710 51390 -590
rect 51510 -710 51555 -590
rect 51675 -710 51720 -590
rect 51840 -710 51885 -590
rect 52005 -710 52060 -590
rect 52180 -710 52225 -590
rect 52345 -710 52390 -590
rect 52510 -710 52555 -590
rect 52675 -710 52730 -590
rect 52850 -710 52895 -590
rect 53015 -710 53060 -590
rect 53180 -710 53225 -590
rect 53345 -710 53370 -590
rect 30770 -755 53370 -710
rect 30770 -875 30795 -755
rect 30915 -875 30970 -755
rect 31090 -875 31135 -755
rect 31255 -875 31300 -755
rect 31420 -875 31465 -755
rect 31585 -875 31640 -755
rect 31760 -875 31805 -755
rect 31925 -875 31970 -755
rect 32090 -875 32135 -755
rect 32255 -875 32310 -755
rect 32430 -875 32475 -755
rect 32595 -875 32640 -755
rect 32760 -875 32805 -755
rect 32925 -875 32980 -755
rect 33100 -875 33145 -755
rect 33265 -875 33310 -755
rect 33430 -875 33475 -755
rect 33595 -875 33650 -755
rect 33770 -875 33815 -755
rect 33935 -875 33980 -755
rect 34100 -875 34145 -755
rect 34265 -875 34320 -755
rect 34440 -875 34485 -755
rect 34605 -875 34650 -755
rect 34770 -875 34815 -755
rect 34935 -875 34990 -755
rect 35110 -875 35155 -755
rect 35275 -875 35320 -755
rect 35440 -875 35485 -755
rect 35605 -875 35660 -755
rect 35780 -875 35825 -755
rect 35945 -875 35990 -755
rect 36110 -875 36155 -755
rect 36275 -875 36485 -755
rect 36605 -875 36660 -755
rect 36780 -875 36825 -755
rect 36945 -875 36990 -755
rect 37110 -875 37155 -755
rect 37275 -875 37330 -755
rect 37450 -875 37495 -755
rect 37615 -875 37660 -755
rect 37780 -875 37825 -755
rect 37945 -875 38000 -755
rect 38120 -875 38165 -755
rect 38285 -875 38330 -755
rect 38450 -875 38495 -755
rect 38615 -875 38670 -755
rect 38790 -875 38835 -755
rect 38955 -875 39000 -755
rect 39120 -875 39165 -755
rect 39285 -875 39340 -755
rect 39460 -875 39505 -755
rect 39625 -875 39670 -755
rect 39790 -875 39835 -755
rect 39955 -875 40010 -755
rect 40130 -875 40175 -755
rect 40295 -875 40340 -755
rect 40460 -875 40505 -755
rect 40625 -875 40680 -755
rect 40800 -875 40845 -755
rect 40965 -875 41010 -755
rect 41130 -875 41175 -755
rect 41295 -875 41350 -755
rect 41470 -875 41515 -755
rect 41635 -875 41680 -755
rect 41800 -875 41845 -755
rect 41965 -875 42175 -755
rect 42295 -875 42350 -755
rect 42470 -875 42515 -755
rect 42635 -875 42680 -755
rect 42800 -875 42845 -755
rect 42965 -875 43020 -755
rect 43140 -875 43185 -755
rect 43305 -875 43350 -755
rect 43470 -875 43515 -755
rect 43635 -875 43690 -755
rect 43810 -875 43855 -755
rect 43975 -875 44020 -755
rect 44140 -875 44185 -755
rect 44305 -875 44360 -755
rect 44480 -875 44525 -755
rect 44645 -875 44690 -755
rect 44810 -875 44855 -755
rect 44975 -875 45030 -755
rect 45150 -875 45195 -755
rect 45315 -875 45360 -755
rect 45480 -875 45525 -755
rect 45645 -875 45700 -755
rect 45820 -875 45865 -755
rect 45985 -875 46030 -755
rect 46150 -875 46195 -755
rect 46315 -875 46370 -755
rect 46490 -875 46535 -755
rect 46655 -875 46700 -755
rect 46820 -875 46865 -755
rect 46985 -875 47040 -755
rect 47160 -875 47205 -755
rect 47325 -875 47370 -755
rect 47490 -875 47535 -755
rect 47655 -875 47865 -755
rect 47985 -875 48040 -755
rect 48160 -875 48205 -755
rect 48325 -875 48370 -755
rect 48490 -875 48535 -755
rect 48655 -875 48710 -755
rect 48830 -875 48875 -755
rect 48995 -875 49040 -755
rect 49160 -875 49205 -755
rect 49325 -875 49380 -755
rect 49500 -875 49545 -755
rect 49665 -875 49710 -755
rect 49830 -875 49875 -755
rect 49995 -875 50050 -755
rect 50170 -875 50215 -755
rect 50335 -875 50380 -755
rect 50500 -875 50545 -755
rect 50665 -875 50720 -755
rect 50840 -875 50885 -755
rect 51005 -875 51050 -755
rect 51170 -875 51215 -755
rect 51335 -875 51390 -755
rect 51510 -875 51555 -755
rect 51675 -875 51720 -755
rect 51840 -875 51885 -755
rect 52005 -875 52060 -755
rect 52180 -875 52225 -755
rect 52345 -875 52390 -755
rect 52510 -875 52555 -755
rect 52675 -875 52730 -755
rect 52850 -875 52895 -755
rect 53015 -875 53060 -755
rect 53180 -875 53225 -755
rect 53345 -875 53370 -755
rect 30770 -920 53370 -875
rect 30770 -1040 30795 -920
rect 30915 -1040 30970 -920
rect 31090 -1040 31135 -920
rect 31255 -1040 31300 -920
rect 31420 -1040 31465 -920
rect 31585 -1040 31640 -920
rect 31760 -1040 31805 -920
rect 31925 -1040 31970 -920
rect 32090 -1040 32135 -920
rect 32255 -1040 32310 -920
rect 32430 -1040 32475 -920
rect 32595 -1040 32640 -920
rect 32760 -1040 32805 -920
rect 32925 -1040 32980 -920
rect 33100 -1040 33145 -920
rect 33265 -1040 33310 -920
rect 33430 -1040 33475 -920
rect 33595 -1040 33650 -920
rect 33770 -1040 33815 -920
rect 33935 -1040 33980 -920
rect 34100 -1040 34145 -920
rect 34265 -1040 34320 -920
rect 34440 -1040 34485 -920
rect 34605 -1040 34650 -920
rect 34770 -1040 34815 -920
rect 34935 -1040 34990 -920
rect 35110 -1040 35155 -920
rect 35275 -1040 35320 -920
rect 35440 -1040 35485 -920
rect 35605 -1040 35660 -920
rect 35780 -1040 35825 -920
rect 35945 -1040 35990 -920
rect 36110 -1040 36155 -920
rect 36275 -1040 36485 -920
rect 36605 -1040 36660 -920
rect 36780 -1040 36825 -920
rect 36945 -1040 36990 -920
rect 37110 -1040 37155 -920
rect 37275 -1040 37330 -920
rect 37450 -1040 37495 -920
rect 37615 -1040 37660 -920
rect 37780 -1040 37825 -920
rect 37945 -1040 38000 -920
rect 38120 -1040 38165 -920
rect 38285 -1040 38330 -920
rect 38450 -1040 38495 -920
rect 38615 -1040 38670 -920
rect 38790 -1040 38835 -920
rect 38955 -1040 39000 -920
rect 39120 -1040 39165 -920
rect 39285 -1040 39340 -920
rect 39460 -1040 39505 -920
rect 39625 -1040 39670 -920
rect 39790 -1040 39835 -920
rect 39955 -1040 40010 -920
rect 40130 -1040 40175 -920
rect 40295 -1040 40340 -920
rect 40460 -1040 40505 -920
rect 40625 -1040 40680 -920
rect 40800 -1040 40845 -920
rect 40965 -1040 41010 -920
rect 41130 -1040 41175 -920
rect 41295 -1040 41350 -920
rect 41470 -1040 41515 -920
rect 41635 -1040 41680 -920
rect 41800 -1040 41845 -920
rect 41965 -1040 42175 -920
rect 42295 -1040 42350 -920
rect 42470 -1040 42515 -920
rect 42635 -1040 42680 -920
rect 42800 -1040 42845 -920
rect 42965 -1040 43020 -920
rect 43140 -1040 43185 -920
rect 43305 -1040 43350 -920
rect 43470 -1040 43515 -920
rect 43635 -1040 43690 -920
rect 43810 -1040 43855 -920
rect 43975 -1040 44020 -920
rect 44140 -1040 44185 -920
rect 44305 -1040 44360 -920
rect 44480 -1040 44525 -920
rect 44645 -1040 44690 -920
rect 44810 -1040 44855 -920
rect 44975 -1040 45030 -920
rect 45150 -1040 45195 -920
rect 45315 -1040 45360 -920
rect 45480 -1040 45525 -920
rect 45645 -1040 45700 -920
rect 45820 -1040 45865 -920
rect 45985 -1040 46030 -920
rect 46150 -1040 46195 -920
rect 46315 -1040 46370 -920
rect 46490 -1040 46535 -920
rect 46655 -1040 46700 -920
rect 46820 -1040 46865 -920
rect 46985 -1040 47040 -920
rect 47160 -1040 47205 -920
rect 47325 -1040 47370 -920
rect 47490 -1040 47535 -920
rect 47655 -1040 47865 -920
rect 47985 -1040 48040 -920
rect 48160 -1040 48205 -920
rect 48325 -1040 48370 -920
rect 48490 -1040 48535 -920
rect 48655 -1040 48710 -920
rect 48830 -1040 48875 -920
rect 48995 -1040 49040 -920
rect 49160 -1040 49205 -920
rect 49325 -1040 49380 -920
rect 49500 -1040 49545 -920
rect 49665 -1040 49710 -920
rect 49830 -1040 49875 -920
rect 49995 -1040 50050 -920
rect 50170 -1040 50215 -920
rect 50335 -1040 50380 -920
rect 50500 -1040 50545 -920
rect 50665 -1040 50720 -920
rect 50840 -1040 50885 -920
rect 51005 -1040 51050 -920
rect 51170 -1040 51215 -920
rect 51335 -1040 51390 -920
rect 51510 -1040 51555 -920
rect 51675 -1040 51720 -920
rect 51840 -1040 51885 -920
rect 52005 -1040 52060 -920
rect 52180 -1040 52225 -920
rect 52345 -1040 52390 -920
rect 52510 -1040 52555 -920
rect 52675 -1040 52730 -920
rect 52850 -1040 52895 -920
rect 53015 -1040 53060 -920
rect 53180 -1040 53225 -920
rect 53345 -1040 53370 -920
rect 30770 -1085 53370 -1040
rect 30770 -1205 30795 -1085
rect 30915 -1205 30970 -1085
rect 31090 -1205 31135 -1085
rect 31255 -1205 31300 -1085
rect 31420 -1205 31465 -1085
rect 31585 -1205 31640 -1085
rect 31760 -1205 31805 -1085
rect 31925 -1205 31970 -1085
rect 32090 -1205 32135 -1085
rect 32255 -1205 32310 -1085
rect 32430 -1205 32475 -1085
rect 32595 -1205 32640 -1085
rect 32760 -1205 32805 -1085
rect 32925 -1205 32980 -1085
rect 33100 -1205 33145 -1085
rect 33265 -1205 33310 -1085
rect 33430 -1205 33475 -1085
rect 33595 -1205 33650 -1085
rect 33770 -1205 33815 -1085
rect 33935 -1205 33980 -1085
rect 34100 -1205 34145 -1085
rect 34265 -1205 34320 -1085
rect 34440 -1205 34485 -1085
rect 34605 -1205 34650 -1085
rect 34770 -1205 34815 -1085
rect 34935 -1205 34990 -1085
rect 35110 -1205 35155 -1085
rect 35275 -1205 35320 -1085
rect 35440 -1205 35485 -1085
rect 35605 -1205 35660 -1085
rect 35780 -1205 35825 -1085
rect 35945 -1205 35990 -1085
rect 36110 -1205 36155 -1085
rect 36275 -1205 36485 -1085
rect 36605 -1205 36660 -1085
rect 36780 -1205 36825 -1085
rect 36945 -1205 36990 -1085
rect 37110 -1205 37155 -1085
rect 37275 -1205 37330 -1085
rect 37450 -1205 37495 -1085
rect 37615 -1205 37660 -1085
rect 37780 -1205 37825 -1085
rect 37945 -1205 38000 -1085
rect 38120 -1205 38165 -1085
rect 38285 -1205 38330 -1085
rect 38450 -1205 38495 -1085
rect 38615 -1205 38670 -1085
rect 38790 -1205 38835 -1085
rect 38955 -1205 39000 -1085
rect 39120 -1205 39165 -1085
rect 39285 -1205 39340 -1085
rect 39460 -1205 39505 -1085
rect 39625 -1205 39670 -1085
rect 39790 -1205 39835 -1085
rect 39955 -1205 40010 -1085
rect 40130 -1205 40175 -1085
rect 40295 -1205 40340 -1085
rect 40460 -1205 40505 -1085
rect 40625 -1205 40680 -1085
rect 40800 -1205 40845 -1085
rect 40965 -1205 41010 -1085
rect 41130 -1205 41175 -1085
rect 41295 -1205 41350 -1085
rect 41470 -1205 41515 -1085
rect 41635 -1205 41680 -1085
rect 41800 -1205 41845 -1085
rect 41965 -1205 42175 -1085
rect 42295 -1205 42350 -1085
rect 42470 -1205 42515 -1085
rect 42635 -1205 42680 -1085
rect 42800 -1205 42845 -1085
rect 42965 -1205 43020 -1085
rect 43140 -1205 43185 -1085
rect 43305 -1205 43350 -1085
rect 43470 -1205 43515 -1085
rect 43635 -1205 43690 -1085
rect 43810 -1205 43855 -1085
rect 43975 -1205 44020 -1085
rect 44140 -1205 44185 -1085
rect 44305 -1205 44360 -1085
rect 44480 -1205 44525 -1085
rect 44645 -1205 44690 -1085
rect 44810 -1205 44855 -1085
rect 44975 -1205 45030 -1085
rect 45150 -1205 45195 -1085
rect 45315 -1205 45360 -1085
rect 45480 -1205 45525 -1085
rect 45645 -1205 45700 -1085
rect 45820 -1205 45865 -1085
rect 45985 -1205 46030 -1085
rect 46150 -1205 46195 -1085
rect 46315 -1205 46370 -1085
rect 46490 -1205 46535 -1085
rect 46655 -1205 46700 -1085
rect 46820 -1205 46865 -1085
rect 46985 -1205 47040 -1085
rect 47160 -1205 47205 -1085
rect 47325 -1205 47370 -1085
rect 47490 -1205 47535 -1085
rect 47655 -1205 47865 -1085
rect 47985 -1205 48040 -1085
rect 48160 -1205 48205 -1085
rect 48325 -1205 48370 -1085
rect 48490 -1205 48535 -1085
rect 48655 -1205 48710 -1085
rect 48830 -1205 48875 -1085
rect 48995 -1205 49040 -1085
rect 49160 -1205 49205 -1085
rect 49325 -1205 49380 -1085
rect 49500 -1205 49545 -1085
rect 49665 -1205 49710 -1085
rect 49830 -1205 49875 -1085
rect 49995 -1205 50050 -1085
rect 50170 -1205 50215 -1085
rect 50335 -1205 50380 -1085
rect 50500 -1205 50545 -1085
rect 50665 -1205 50720 -1085
rect 50840 -1205 50885 -1085
rect 51005 -1205 51050 -1085
rect 51170 -1205 51215 -1085
rect 51335 -1205 51390 -1085
rect 51510 -1205 51555 -1085
rect 51675 -1205 51720 -1085
rect 51840 -1205 51885 -1085
rect 52005 -1205 52060 -1085
rect 52180 -1205 52225 -1085
rect 52345 -1205 52390 -1085
rect 52510 -1205 52555 -1085
rect 52675 -1205 52730 -1085
rect 52850 -1205 52895 -1085
rect 53015 -1205 53060 -1085
rect 53180 -1205 53225 -1085
rect 53345 -1205 53370 -1085
rect 30770 -1260 53370 -1205
rect 30770 -1380 30795 -1260
rect 30915 -1380 30970 -1260
rect 31090 -1380 31135 -1260
rect 31255 -1380 31300 -1260
rect 31420 -1380 31465 -1260
rect 31585 -1380 31640 -1260
rect 31760 -1380 31805 -1260
rect 31925 -1380 31970 -1260
rect 32090 -1380 32135 -1260
rect 32255 -1380 32310 -1260
rect 32430 -1380 32475 -1260
rect 32595 -1380 32640 -1260
rect 32760 -1380 32805 -1260
rect 32925 -1380 32980 -1260
rect 33100 -1380 33145 -1260
rect 33265 -1380 33310 -1260
rect 33430 -1380 33475 -1260
rect 33595 -1380 33650 -1260
rect 33770 -1380 33815 -1260
rect 33935 -1380 33980 -1260
rect 34100 -1380 34145 -1260
rect 34265 -1380 34320 -1260
rect 34440 -1380 34485 -1260
rect 34605 -1380 34650 -1260
rect 34770 -1380 34815 -1260
rect 34935 -1380 34990 -1260
rect 35110 -1380 35155 -1260
rect 35275 -1380 35320 -1260
rect 35440 -1380 35485 -1260
rect 35605 -1380 35660 -1260
rect 35780 -1380 35825 -1260
rect 35945 -1380 35990 -1260
rect 36110 -1380 36155 -1260
rect 36275 -1380 36485 -1260
rect 36605 -1380 36660 -1260
rect 36780 -1380 36825 -1260
rect 36945 -1380 36990 -1260
rect 37110 -1380 37155 -1260
rect 37275 -1380 37330 -1260
rect 37450 -1380 37495 -1260
rect 37615 -1380 37660 -1260
rect 37780 -1380 37825 -1260
rect 37945 -1380 38000 -1260
rect 38120 -1380 38165 -1260
rect 38285 -1380 38330 -1260
rect 38450 -1380 38495 -1260
rect 38615 -1380 38670 -1260
rect 38790 -1380 38835 -1260
rect 38955 -1380 39000 -1260
rect 39120 -1380 39165 -1260
rect 39285 -1380 39340 -1260
rect 39460 -1380 39505 -1260
rect 39625 -1380 39670 -1260
rect 39790 -1380 39835 -1260
rect 39955 -1380 40010 -1260
rect 40130 -1380 40175 -1260
rect 40295 -1380 40340 -1260
rect 40460 -1380 40505 -1260
rect 40625 -1380 40680 -1260
rect 40800 -1380 40845 -1260
rect 40965 -1380 41010 -1260
rect 41130 -1380 41175 -1260
rect 41295 -1380 41350 -1260
rect 41470 -1380 41515 -1260
rect 41635 -1380 41680 -1260
rect 41800 -1380 41845 -1260
rect 41965 -1380 42175 -1260
rect 42295 -1380 42350 -1260
rect 42470 -1380 42515 -1260
rect 42635 -1380 42680 -1260
rect 42800 -1380 42845 -1260
rect 42965 -1380 43020 -1260
rect 43140 -1380 43185 -1260
rect 43305 -1380 43350 -1260
rect 43470 -1380 43515 -1260
rect 43635 -1380 43690 -1260
rect 43810 -1380 43855 -1260
rect 43975 -1380 44020 -1260
rect 44140 -1380 44185 -1260
rect 44305 -1380 44360 -1260
rect 44480 -1380 44525 -1260
rect 44645 -1380 44690 -1260
rect 44810 -1380 44855 -1260
rect 44975 -1380 45030 -1260
rect 45150 -1380 45195 -1260
rect 45315 -1380 45360 -1260
rect 45480 -1380 45525 -1260
rect 45645 -1380 45700 -1260
rect 45820 -1380 45865 -1260
rect 45985 -1380 46030 -1260
rect 46150 -1380 46195 -1260
rect 46315 -1380 46370 -1260
rect 46490 -1380 46535 -1260
rect 46655 -1380 46700 -1260
rect 46820 -1380 46865 -1260
rect 46985 -1380 47040 -1260
rect 47160 -1380 47205 -1260
rect 47325 -1380 47370 -1260
rect 47490 -1380 47535 -1260
rect 47655 -1380 47865 -1260
rect 47985 -1380 48040 -1260
rect 48160 -1380 48205 -1260
rect 48325 -1380 48370 -1260
rect 48490 -1380 48535 -1260
rect 48655 -1380 48710 -1260
rect 48830 -1380 48875 -1260
rect 48995 -1380 49040 -1260
rect 49160 -1380 49205 -1260
rect 49325 -1380 49380 -1260
rect 49500 -1380 49545 -1260
rect 49665 -1380 49710 -1260
rect 49830 -1380 49875 -1260
rect 49995 -1380 50050 -1260
rect 50170 -1380 50215 -1260
rect 50335 -1380 50380 -1260
rect 50500 -1380 50545 -1260
rect 50665 -1380 50720 -1260
rect 50840 -1380 50885 -1260
rect 51005 -1380 51050 -1260
rect 51170 -1380 51215 -1260
rect 51335 -1380 51390 -1260
rect 51510 -1380 51555 -1260
rect 51675 -1380 51720 -1260
rect 51840 -1380 51885 -1260
rect 52005 -1380 52060 -1260
rect 52180 -1380 52225 -1260
rect 52345 -1380 52390 -1260
rect 52510 -1380 52555 -1260
rect 52675 -1380 52730 -1260
rect 52850 -1380 52895 -1260
rect 53015 -1380 53060 -1260
rect 53180 -1380 53225 -1260
rect 53345 -1380 53370 -1260
rect 30770 -1425 53370 -1380
rect 30770 -1545 30795 -1425
rect 30915 -1545 30970 -1425
rect 31090 -1545 31135 -1425
rect 31255 -1545 31300 -1425
rect 31420 -1545 31465 -1425
rect 31585 -1545 31640 -1425
rect 31760 -1545 31805 -1425
rect 31925 -1545 31970 -1425
rect 32090 -1545 32135 -1425
rect 32255 -1545 32310 -1425
rect 32430 -1545 32475 -1425
rect 32595 -1545 32640 -1425
rect 32760 -1545 32805 -1425
rect 32925 -1545 32980 -1425
rect 33100 -1545 33145 -1425
rect 33265 -1545 33310 -1425
rect 33430 -1545 33475 -1425
rect 33595 -1545 33650 -1425
rect 33770 -1545 33815 -1425
rect 33935 -1545 33980 -1425
rect 34100 -1545 34145 -1425
rect 34265 -1545 34320 -1425
rect 34440 -1545 34485 -1425
rect 34605 -1545 34650 -1425
rect 34770 -1545 34815 -1425
rect 34935 -1545 34990 -1425
rect 35110 -1545 35155 -1425
rect 35275 -1545 35320 -1425
rect 35440 -1545 35485 -1425
rect 35605 -1545 35660 -1425
rect 35780 -1545 35825 -1425
rect 35945 -1545 35990 -1425
rect 36110 -1545 36155 -1425
rect 36275 -1545 36485 -1425
rect 36605 -1545 36660 -1425
rect 36780 -1545 36825 -1425
rect 36945 -1545 36990 -1425
rect 37110 -1545 37155 -1425
rect 37275 -1545 37330 -1425
rect 37450 -1545 37495 -1425
rect 37615 -1545 37660 -1425
rect 37780 -1545 37825 -1425
rect 37945 -1545 38000 -1425
rect 38120 -1545 38165 -1425
rect 38285 -1545 38330 -1425
rect 38450 -1545 38495 -1425
rect 38615 -1545 38670 -1425
rect 38790 -1545 38835 -1425
rect 38955 -1545 39000 -1425
rect 39120 -1545 39165 -1425
rect 39285 -1545 39340 -1425
rect 39460 -1545 39505 -1425
rect 39625 -1545 39670 -1425
rect 39790 -1545 39835 -1425
rect 39955 -1545 40010 -1425
rect 40130 -1545 40175 -1425
rect 40295 -1545 40340 -1425
rect 40460 -1545 40505 -1425
rect 40625 -1545 40680 -1425
rect 40800 -1545 40845 -1425
rect 40965 -1545 41010 -1425
rect 41130 -1545 41175 -1425
rect 41295 -1545 41350 -1425
rect 41470 -1545 41515 -1425
rect 41635 -1545 41680 -1425
rect 41800 -1545 41845 -1425
rect 41965 -1545 42175 -1425
rect 42295 -1545 42350 -1425
rect 42470 -1545 42515 -1425
rect 42635 -1545 42680 -1425
rect 42800 -1545 42845 -1425
rect 42965 -1545 43020 -1425
rect 43140 -1545 43185 -1425
rect 43305 -1545 43350 -1425
rect 43470 -1545 43515 -1425
rect 43635 -1545 43690 -1425
rect 43810 -1545 43855 -1425
rect 43975 -1545 44020 -1425
rect 44140 -1545 44185 -1425
rect 44305 -1545 44360 -1425
rect 44480 -1545 44525 -1425
rect 44645 -1545 44690 -1425
rect 44810 -1545 44855 -1425
rect 44975 -1545 45030 -1425
rect 45150 -1545 45195 -1425
rect 45315 -1545 45360 -1425
rect 45480 -1545 45525 -1425
rect 45645 -1545 45700 -1425
rect 45820 -1545 45865 -1425
rect 45985 -1545 46030 -1425
rect 46150 -1545 46195 -1425
rect 46315 -1545 46370 -1425
rect 46490 -1545 46535 -1425
rect 46655 -1545 46700 -1425
rect 46820 -1545 46865 -1425
rect 46985 -1545 47040 -1425
rect 47160 -1545 47205 -1425
rect 47325 -1545 47370 -1425
rect 47490 -1545 47535 -1425
rect 47655 -1545 47865 -1425
rect 47985 -1545 48040 -1425
rect 48160 -1545 48205 -1425
rect 48325 -1545 48370 -1425
rect 48490 -1545 48535 -1425
rect 48655 -1545 48710 -1425
rect 48830 -1545 48875 -1425
rect 48995 -1545 49040 -1425
rect 49160 -1545 49205 -1425
rect 49325 -1545 49380 -1425
rect 49500 -1545 49545 -1425
rect 49665 -1545 49710 -1425
rect 49830 -1545 49875 -1425
rect 49995 -1545 50050 -1425
rect 50170 -1545 50215 -1425
rect 50335 -1545 50380 -1425
rect 50500 -1545 50545 -1425
rect 50665 -1545 50720 -1425
rect 50840 -1545 50885 -1425
rect 51005 -1545 51050 -1425
rect 51170 -1545 51215 -1425
rect 51335 -1545 51390 -1425
rect 51510 -1545 51555 -1425
rect 51675 -1545 51720 -1425
rect 51840 -1545 51885 -1425
rect 52005 -1545 52060 -1425
rect 52180 -1545 52225 -1425
rect 52345 -1545 52390 -1425
rect 52510 -1545 52555 -1425
rect 52675 -1545 52730 -1425
rect 52850 -1545 52895 -1425
rect 53015 -1545 53060 -1425
rect 53180 -1545 53225 -1425
rect 53345 -1545 53370 -1425
rect 30770 -1590 53370 -1545
rect 30770 -1710 30795 -1590
rect 30915 -1710 30970 -1590
rect 31090 -1710 31135 -1590
rect 31255 -1710 31300 -1590
rect 31420 -1710 31465 -1590
rect 31585 -1710 31640 -1590
rect 31760 -1710 31805 -1590
rect 31925 -1710 31970 -1590
rect 32090 -1710 32135 -1590
rect 32255 -1710 32310 -1590
rect 32430 -1710 32475 -1590
rect 32595 -1710 32640 -1590
rect 32760 -1710 32805 -1590
rect 32925 -1710 32980 -1590
rect 33100 -1710 33145 -1590
rect 33265 -1710 33310 -1590
rect 33430 -1710 33475 -1590
rect 33595 -1710 33650 -1590
rect 33770 -1710 33815 -1590
rect 33935 -1710 33980 -1590
rect 34100 -1710 34145 -1590
rect 34265 -1710 34320 -1590
rect 34440 -1710 34485 -1590
rect 34605 -1710 34650 -1590
rect 34770 -1710 34815 -1590
rect 34935 -1710 34990 -1590
rect 35110 -1710 35155 -1590
rect 35275 -1710 35320 -1590
rect 35440 -1710 35485 -1590
rect 35605 -1710 35660 -1590
rect 35780 -1710 35825 -1590
rect 35945 -1710 35990 -1590
rect 36110 -1710 36155 -1590
rect 36275 -1710 36485 -1590
rect 36605 -1710 36660 -1590
rect 36780 -1710 36825 -1590
rect 36945 -1710 36990 -1590
rect 37110 -1710 37155 -1590
rect 37275 -1710 37330 -1590
rect 37450 -1710 37495 -1590
rect 37615 -1710 37660 -1590
rect 37780 -1710 37825 -1590
rect 37945 -1710 38000 -1590
rect 38120 -1710 38165 -1590
rect 38285 -1710 38330 -1590
rect 38450 -1710 38495 -1590
rect 38615 -1710 38670 -1590
rect 38790 -1710 38835 -1590
rect 38955 -1710 39000 -1590
rect 39120 -1710 39165 -1590
rect 39285 -1710 39340 -1590
rect 39460 -1710 39505 -1590
rect 39625 -1710 39670 -1590
rect 39790 -1710 39835 -1590
rect 39955 -1710 40010 -1590
rect 40130 -1710 40175 -1590
rect 40295 -1710 40340 -1590
rect 40460 -1710 40505 -1590
rect 40625 -1710 40680 -1590
rect 40800 -1710 40845 -1590
rect 40965 -1710 41010 -1590
rect 41130 -1710 41175 -1590
rect 41295 -1710 41350 -1590
rect 41470 -1710 41515 -1590
rect 41635 -1710 41680 -1590
rect 41800 -1710 41845 -1590
rect 41965 -1710 42175 -1590
rect 42295 -1710 42350 -1590
rect 42470 -1710 42515 -1590
rect 42635 -1710 42680 -1590
rect 42800 -1710 42845 -1590
rect 42965 -1710 43020 -1590
rect 43140 -1710 43185 -1590
rect 43305 -1710 43350 -1590
rect 43470 -1710 43515 -1590
rect 43635 -1710 43690 -1590
rect 43810 -1710 43855 -1590
rect 43975 -1710 44020 -1590
rect 44140 -1710 44185 -1590
rect 44305 -1710 44360 -1590
rect 44480 -1710 44525 -1590
rect 44645 -1710 44690 -1590
rect 44810 -1710 44855 -1590
rect 44975 -1710 45030 -1590
rect 45150 -1710 45195 -1590
rect 45315 -1710 45360 -1590
rect 45480 -1710 45525 -1590
rect 45645 -1710 45700 -1590
rect 45820 -1710 45865 -1590
rect 45985 -1710 46030 -1590
rect 46150 -1710 46195 -1590
rect 46315 -1710 46370 -1590
rect 46490 -1710 46535 -1590
rect 46655 -1710 46700 -1590
rect 46820 -1710 46865 -1590
rect 46985 -1710 47040 -1590
rect 47160 -1710 47205 -1590
rect 47325 -1710 47370 -1590
rect 47490 -1710 47535 -1590
rect 47655 -1710 47865 -1590
rect 47985 -1710 48040 -1590
rect 48160 -1710 48205 -1590
rect 48325 -1710 48370 -1590
rect 48490 -1710 48535 -1590
rect 48655 -1710 48710 -1590
rect 48830 -1710 48875 -1590
rect 48995 -1710 49040 -1590
rect 49160 -1710 49205 -1590
rect 49325 -1710 49380 -1590
rect 49500 -1710 49545 -1590
rect 49665 -1710 49710 -1590
rect 49830 -1710 49875 -1590
rect 49995 -1710 50050 -1590
rect 50170 -1710 50215 -1590
rect 50335 -1710 50380 -1590
rect 50500 -1710 50545 -1590
rect 50665 -1710 50720 -1590
rect 50840 -1710 50885 -1590
rect 51005 -1710 51050 -1590
rect 51170 -1710 51215 -1590
rect 51335 -1710 51390 -1590
rect 51510 -1710 51555 -1590
rect 51675 -1710 51720 -1590
rect 51840 -1710 51885 -1590
rect 52005 -1710 52060 -1590
rect 52180 -1710 52225 -1590
rect 52345 -1710 52390 -1590
rect 52510 -1710 52555 -1590
rect 52675 -1710 52730 -1590
rect 52850 -1710 52895 -1590
rect 53015 -1710 53060 -1590
rect 53180 -1710 53225 -1590
rect 53345 -1710 53370 -1590
rect 30770 -1755 53370 -1710
rect 30770 -1875 30795 -1755
rect 30915 -1875 30970 -1755
rect 31090 -1875 31135 -1755
rect 31255 -1875 31300 -1755
rect 31420 -1875 31465 -1755
rect 31585 -1875 31640 -1755
rect 31760 -1875 31805 -1755
rect 31925 -1875 31970 -1755
rect 32090 -1875 32135 -1755
rect 32255 -1875 32310 -1755
rect 32430 -1875 32475 -1755
rect 32595 -1875 32640 -1755
rect 32760 -1875 32805 -1755
rect 32925 -1875 32980 -1755
rect 33100 -1875 33145 -1755
rect 33265 -1875 33310 -1755
rect 33430 -1875 33475 -1755
rect 33595 -1875 33650 -1755
rect 33770 -1875 33815 -1755
rect 33935 -1875 33980 -1755
rect 34100 -1875 34145 -1755
rect 34265 -1875 34320 -1755
rect 34440 -1875 34485 -1755
rect 34605 -1875 34650 -1755
rect 34770 -1875 34815 -1755
rect 34935 -1875 34990 -1755
rect 35110 -1875 35155 -1755
rect 35275 -1875 35320 -1755
rect 35440 -1875 35485 -1755
rect 35605 -1875 35660 -1755
rect 35780 -1875 35825 -1755
rect 35945 -1875 35990 -1755
rect 36110 -1875 36155 -1755
rect 36275 -1875 36485 -1755
rect 36605 -1875 36660 -1755
rect 36780 -1875 36825 -1755
rect 36945 -1875 36990 -1755
rect 37110 -1875 37155 -1755
rect 37275 -1875 37330 -1755
rect 37450 -1875 37495 -1755
rect 37615 -1875 37660 -1755
rect 37780 -1875 37825 -1755
rect 37945 -1875 38000 -1755
rect 38120 -1875 38165 -1755
rect 38285 -1875 38330 -1755
rect 38450 -1875 38495 -1755
rect 38615 -1875 38670 -1755
rect 38790 -1875 38835 -1755
rect 38955 -1875 39000 -1755
rect 39120 -1875 39165 -1755
rect 39285 -1875 39340 -1755
rect 39460 -1875 39505 -1755
rect 39625 -1875 39670 -1755
rect 39790 -1875 39835 -1755
rect 39955 -1875 40010 -1755
rect 40130 -1875 40175 -1755
rect 40295 -1875 40340 -1755
rect 40460 -1875 40505 -1755
rect 40625 -1875 40680 -1755
rect 40800 -1875 40845 -1755
rect 40965 -1875 41010 -1755
rect 41130 -1875 41175 -1755
rect 41295 -1875 41350 -1755
rect 41470 -1875 41515 -1755
rect 41635 -1875 41680 -1755
rect 41800 -1875 41845 -1755
rect 41965 -1875 42175 -1755
rect 42295 -1875 42350 -1755
rect 42470 -1875 42515 -1755
rect 42635 -1875 42680 -1755
rect 42800 -1875 42845 -1755
rect 42965 -1875 43020 -1755
rect 43140 -1875 43185 -1755
rect 43305 -1875 43350 -1755
rect 43470 -1875 43515 -1755
rect 43635 -1875 43690 -1755
rect 43810 -1875 43855 -1755
rect 43975 -1875 44020 -1755
rect 44140 -1875 44185 -1755
rect 44305 -1875 44360 -1755
rect 44480 -1875 44525 -1755
rect 44645 -1875 44690 -1755
rect 44810 -1875 44855 -1755
rect 44975 -1875 45030 -1755
rect 45150 -1875 45195 -1755
rect 45315 -1875 45360 -1755
rect 45480 -1875 45525 -1755
rect 45645 -1875 45700 -1755
rect 45820 -1875 45865 -1755
rect 45985 -1875 46030 -1755
rect 46150 -1875 46195 -1755
rect 46315 -1875 46370 -1755
rect 46490 -1875 46535 -1755
rect 46655 -1875 46700 -1755
rect 46820 -1875 46865 -1755
rect 46985 -1875 47040 -1755
rect 47160 -1875 47205 -1755
rect 47325 -1875 47370 -1755
rect 47490 -1875 47535 -1755
rect 47655 -1875 47865 -1755
rect 47985 -1875 48040 -1755
rect 48160 -1875 48205 -1755
rect 48325 -1875 48370 -1755
rect 48490 -1875 48535 -1755
rect 48655 -1875 48710 -1755
rect 48830 -1875 48875 -1755
rect 48995 -1875 49040 -1755
rect 49160 -1875 49205 -1755
rect 49325 -1875 49380 -1755
rect 49500 -1875 49545 -1755
rect 49665 -1875 49710 -1755
rect 49830 -1875 49875 -1755
rect 49995 -1875 50050 -1755
rect 50170 -1875 50215 -1755
rect 50335 -1875 50380 -1755
rect 50500 -1875 50545 -1755
rect 50665 -1875 50720 -1755
rect 50840 -1875 50885 -1755
rect 51005 -1875 51050 -1755
rect 51170 -1875 51215 -1755
rect 51335 -1875 51390 -1755
rect 51510 -1875 51555 -1755
rect 51675 -1875 51720 -1755
rect 51840 -1875 51885 -1755
rect 52005 -1875 52060 -1755
rect 52180 -1875 52225 -1755
rect 52345 -1875 52390 -1755
rect 52510 -1875 52555 -1755
rect 52675 -1875 52730 -1755
rect 52850 -1875 52895 -1755
rect 53015 -1875 53060 -1755
rect 53180 -1875 53225 -1755
rect 53345 -1875 53370 -1755
rect 30770 -1930 53370 -1875
rect 30770 -2005 30795 -1930
rect 30665 -2050 30795 -2005
rect 30915 -2050 30970 -1930
rect 31090 -2050 31135 -1930
rect 31255 -2050 31300 -1930
rect 31420 -2050 31465 -1930
rect 31585 -2050 31640 -1930
rect 31760 -2050 31805 -1930
rect 31925 -2050 31970 -1930
rect 32090 -2050 32135 -1930
rect 32255 -2050 32310 -1930
rect 32430 -2050 32475 -1930
rect 32595 -2050 32640 -1930
rect 32760 -2050 32805 -1930
rect 32925 -2050 32980 -1930
rect 33100 -2050 33145 -1930
rect 33265 -2050 33310 -1930
rect 33430 -2050 33475 -1930
rect 33595 -2050 33650 -1930
rect 33770 -2050 33815 -1930
rect 33935 -2050 33980 -1930
rect 34100 -2050 34145 -1930
rect 34265 -2050 34320 -1930
rect 34440 -2050 34485 -1930
rect 34605 -2050 34650 -1930
rect 34770 -2050 34815 -1930
rect 34935 -2050 34990 -1930
rect 35110 -2050 35155 -1930
rect 35275 -2050 35320 -1930
rect 35440 -2050 35485 -1930
rect 35605 -2050 35660 -1930
rect 35780 -2050 35825 -1930
rect 35945 -2050 35990 -1930
rect 36110 -2050 36155 -1930
rect 36275 -2050 36485 -1930
rect 36605 -2050 36660 -1930
rect 36780 -2050 36825 -1930
rect 36945 -2050 36990 -1930
rect 37110 -2050 37155 -1930
rect 37275 -2050 37330 -1930
rect 37450 -2050 37495 -1930
rect 37615 -2050 37660 -1930
rect 37780 -2050 37825 -1930
rect 37945 -2050 38000 -1930
rect 38120 -2050 38165 -1930
rect 38285 -2050 38330 -1930
rect 38450 -2050 38495 -1930
rect 38615 -2050 38670 -1930
rect 38790 -2050 38835 -1930
rect 38955 -2050 39000 -1930
rect 39120 -2050 39165 -1930
rect 39285 -2050 39340 -1930
rect 39460 -2050 39505 -1930
rect 39625 -2050 39670 -1930
rect 39790 -2050 39835 -1930
rect 39955 -2050 40010 -1930
rect 40130 -2050 40175 -1930
rect 40295 -2050 40340 -1930
rect 40460 -2050 40505 -1930
rect 40625 -2050 40680 -1930
rect 40800 -2050 40845 -1930
rect 40965 -2050 41010 -1930
rect 41130 -2050 41175 -1930
rect 41295 -2050 41350 -1930
rect 41470 -2050 41515 -1930
rect 41635 -2050 41680 -1930
rect 41800 -2050 41845 -1930
rect 41965 -2050 42175 -1930
rect 42295 -2050 42350 -1930
rect 42470 -2050 42515 -1930
rect 42635 -2050 42680 -1930
rect 42800 -2050 42845 -1930
rect 42965 -2050 43020 -1930
rect 43140 -2050 43185 -1930
rect 43305 -2050 43350 -1930
rect 43470 -2050 43515 -1930
rect 43635 -2050 43690 -1930
rect 43810 -2050 43855 -1930
rect 43975 -2050 44020 -1930
rect 44140 -2050 44185 -1930
rect 44305 -2050 44360 -1930
rect 44480 -2050 44525 -1930
rect 44645 -2050 44690 -1930
rect 44810 -2050 44855 -1930
rect 44975 -2050 45030 -1930
rect 45150 -2050 45195 -1930
rect 45315 -2050 45360 -1930
rect 45480 -2050 45525 -1930
rect 45645 -2050 45700 -1930
rect 45820 -2050 45865 -1930
rect 45985 -2050 46030 -1930
rect 46150 -2050 46195 -1930
rect 46315 -2050 46370 -1930
rect 46490 -2050 46535 -1930
rect 46655 -2050 46700 -1930
rect 46820 -2050 46865 -1930
rect 46985 -2050 47040 -1930
rect 47160 -2050 47205 -1930
rect 47325 -2050 47370 -1930
rect 47490 -2050 47535 -1930
rect 47655 -2050 47865 -1930
rect 47985 -2050 48040 -1930
rect 48160 -2050 48205 -1930
rect 48325 -2050 48370 -1930
rect 48490 -2050 48535 -1930
rect 48655 -2050 48710 -1930
rect 48830 -2050 48875 -1930
rect 48995 -2050 49040 -1930
rect 49160 -2050 49205 -1930
rect 49325 -2050 49380 -1930
rect 49500 -2050 49545 -1930
rect 49665 -2050 49710 -1930
rect 49830 -2050 49875 -1930
rect 49995 -2050 50050 -1930
rect 50170 -2050 50215 -1930
rect 50335 -2050 50380 -1930
rect 50500 -2050 50545 -1930
rect 50665 -2050 50720 -1930
rect 50840 -2050 50885 -1930
rect 51005 -2050 51050 -1930
rect 51170 -2050 51215 -1930
rect 51335 -2050 51390 -1930
rect 51510 -2050 51555 -1930
rect 51675 -2050 51720 -1930
rect 51840 -2050 51885 -1930
rect 52005 -2050 52060 -1930
rect 52180 -2050 52225 -1930
rect 52345 -2050 52390 -1930
rect 52510 -2050 52555 -1930
rect 52675 -2050 52730 -1930
rect 52850 -2050 52895 -1930
rect 53015 -2050 53060 -1930
rect 53180 -2050 53225 -1930
rect 53345 -2050 53370 -1930
rect 30665 -2095 53370 -2050
rect 30665 -2215 30795 -2095
rect 30915 -2215 30970 -2095
rect 31090 -2215 31135 -2095
rect 31255 -2215 31300 -2095
rect 31420 -2215 31465 -2095
rect 31585 -2215 31640 -2095
rect 31760 -2215 31805 -2095
rect 31925 -2215 31970 -2095
rect 32090 -2215 32135 -2095
rect 32255 -2215 32310 -2095
rect 32430 -2215 32475 -2095
rect 32595 -2215 32640 -2095
rect 32760 -2215 32805 -2095
rect 32925 -2215 32980 -2095
rect 33100 -2215 33145 -2095
rect 33265 -2215 33310 -2095
rect 33430 -2215 33475 -2095
rect 33595 -2215 33650 -2095
rect 33770 -2215 33815 -2095
rect 33935 -2215 33980 -2095
rect 34100 -2215 34145 -2095
rect 34265 -2215 34320 -2095
rect 34440 -2215 34485 -2095
rect 34605 -2215 34650 -2095
rect 34770 -2215 34815 -2095
rect 34935 -2215 34990 -2095
rect 35110 -2215 35155 -2095
rect 35275 -2215 35320 -2095
rect 35440 -2215 35485 -2095
rect 35605 -2215 35660 -2095
rect 35780 -2215 35825 -2095
rect 35945 -2215 35990 -2095
rect 36110 -2215 36155 -2095
rect 36275 -2215 36485 -2095
rect 36605 -2215 36660 -2095
rect 36780 -2215 36825 -2095
rect 36945 -2215 36990 -2095
rect 37110 -2215 37155 -2095
rect 37275 -2215 37330 -2095
rect 37450 -2215 37495 -2095
rect 37615 -2215 37660 -2095
rect 37780 -2215 37825 -2095
rect 37945 -2215 38000 -2095
rect 38120 -2215 38165 -2095
rect 38285 -2215 38330 -2095
rect 38450 -2215 38495 -2095
rect 38615 -2215 38670 -2095
rect 38790 -2215 38835 -2095
rect 38955 -2215 39000 -2095
rect 39120 -2215 39165 -2095
rect 39285 -2215 39340 -2095
rect 39460 -2215 39505 -2095
rect 39625 -2215 39670 -2095
rect 39790 -2215 39835 -2095
rect 39955 -2215 40010 -2095
rect 40130 -2215 40175 -2095
rect 40295 -2215 40340 -2095
rect 40460 -2215 40505 -2095
rect 40625 -2215 40680 -2095
rect 40800 -2215 40845 -2095
rect 40965 -2215 41010 -2095
rect 41130 -2215 41175 -2095
rect 41295 -2215 41350 -2095
rect 41470 -2215 41515 -2095
rect 41635 -2215 41680 -2095
rect 41800 -2215 41845 -2095
rect 41965 -2215 42175 -2095
rect 42295 -2215 42350 -2095
rect 42470 -2215 42515 -2095
rect 42635 -2215 42680 -2095
rect 42800 -2215 42845 -2095
rect 42965 -2215 43020 -2095
rect 43140 -2215 43185 -2095
rect 43305 -2215 43350 -2095
rect 43470 -2215 43515 -2095
rect 43635 -2215 43690 -2095
rect 43810 -2215 43855 -2095
rect 43975 -2215 44020 -2095
rect 44140 -2215 44185 -2095
rect 44305 -2215 44360 -2095
rect 44480 -2215 44525 -2095
rect 44645 -2215 44690 -2095
rect 44810 -2215 44855 -2095
rect 44975 -2215 45030 -2095
rect 45150 -2215 45195 -2095
rect 45315 -2215 45360 -2095
rect 45480 -2215 45525 -2095
rect 45645 -2215 45700 -2095
rect 45820 -2215 45865 -2095
rect 45985 -2215 46030 -2095
rect 46150 -2215 46195 -2095
rect 46315 -2215 46370 -2095
rect 46490 -2215 46535 -2095
rect 46655 -2215 46700 -2095
rect 46820 -2215 46865 -2095
rect 46985 -2215 47040 -2095
rect 47160 -2215 47205 -2095
rect 47325 -2215 47370 -2095
rect 47490 -2215 47535 -2095
rect 47655 -2215 47865 -2095
rect 47985 -2215 48040 -2095
rect 48160 -2215 48205 -2095
rect 48325 -2215 48370 -2095
rect 48490 -2215 48535 -2095
rect 48655 -2215 48710 -2095
rect 48830 -2215 48875 -2095
rect 48995 -2215 49040 -2095
rect 49160 -2215 49205 -2095
rect 49325 -2215 49380 -2095
rect 49500 -2215 49545 -2095
rect 49665 -2215 49710 -2095
rect 49830 -2215 49875 -2095
rect 49995 -2215 50050 -2095
rect 50170 -2215 50215 -2095
rect 50335 -2215 50380 -2095
rect 50500 -2215 50545 -2095
rect 50665 -2215 50720 -2095
rect 50840 -2215 50885 -2095
rect 51005 -2215 51050 -2095
rect 51170 -2215 51215 -2095
rect 51335 -2215 51390 -2095
rect 51510 -2215 51555 -2095
rect 51675 -2215 51720 -2095
rect 51840 -2215 51885 -2095
rect 52005 -2215 52060 -2095
rect 52180 -2215 52225 -2095
rect 52345 -2215 52390 -2095
rect 52510 -2215 52555 -2095
rect 52675 -2215 52730 -2095
rect 52850 -2215 52895 -2095
rect 53015 -2215 53060 -2095
rect 53180 -2215 53225 -2095
rect 53345 -2215 53370 -2095
rect 30665 -2255 53370 -2215
rect 30770 -2260 53370 -2255
rect 30770 -2380 30795 -2260
rect 30915 -2380 30970 -2260
rect 31090 -2380 31135 -2260
rect 31255 -2380 31300 -2260
rect 31420 -2380 31465 -2260
rect 31585 -2380 31640 -2260
rect 31760 -2380 31805 -2260
rect 31925 -2380 31970 -2260
rect 32090 -2380 32135 -2260
rect 32255 -2380 32310 -2260
rect 32430 -2380 32475 -2260
rect 32595 -2380 32640 -2260
rect 32760 -2380 32805 -2260
rect 32925 -2380 32980 -2260
rect 33100 -2380 33145 -2260
rect 33265 -2380 33310 -2260
rect 33430 -2380 33475 -2260
rect 33595 -2380 33650 -2260
rect 33770 -2380 33815 -2260
rect 33935 -2380 33980 -2260
rect 34100 -2380 34145 -2260
rect 34265 -2380 34320 -2260
rect 34440 -2380 34485 -2260
rect 34605 -2380 34650 -2260
rect 34770 -2380 34815 -2260
rect 34935 -2380 34990 -2260
rect 35110 -2380 35155 -2260
rect 35275 -2380 35320 -2260
rect 35440 -2380 35485 -2260
rect 35605 -2380 35660 -2260
rect 35780 -2380 35825 -2260
rect 35945 -2380 35990 -2260
rect 36110 -2380 36155 -2260
rect 36275 -2380 36485 -2260
rect 36605 -2380 36660 -2260
rect 36780 -2380 36825 -2260
rect 36945 -2380 36990 -2260
rect 37110 -2380 37155 -2260
rect 37275 -2380 37330 -2260
rect 37450 -2380 37495 -2260
rect 37615 -2380 37660 -2260
rect 37780 -2380 37825 -2260
rect 37945 -2380 38000 -2260
rect 38120 -2380 38165 -2260
rect 38285 -2380 38330 -2260
rect 38450 -2380 38495 -2260
rect 38615 -2380 38670 -2260
rect 38790 -2380 38835 -2260
rect 38955 -2380 39000 -2260
rect 39120 -2380 39165 -2260
rect 39285 -2380 39340 -2260
rect 39460 -2380 39505 -2260
rect 39625 -2380 39670 -2260
rect 39790 -2380 39835 -2260
rect 39955 -2380 40010 -2260
rect 40130 -2380 40175 -2260
rect 40295 -2380 40340 -2260
rect 40460 -2380 40505 -2260
rect 40625 -2380 40680 -2260
rect 40800 -2380 40845 -2260
rect 40965 -2380 41010 -2260
rect 41130 -2380 41175 -2260
rect 41295 -2380 41350 -2260
rect 41470 -2380 41515 -2260
rect 41635 -2380 41680 -2260
rect 41800 -2380 41845 -2260
rect 41965 -2380 42175 -2260
rect 42295 -2380 42350 -2260
rect 42470 -2380 42515 -2260
rect 42635 -2380 42680 -2260
rect 42800 -2380 42845 -2260
rect 42965 -2380 43020 -2260
rect 43140 -2380 43185 -2260
rect 43305 -2380 43350 -2260
rect 43470 -2380 43515 -2260
rect 43635 -2380 43690 -2260
rect 43810 -2380 43855 -2260
rect 43975 -2380 44020 -2260
rect 44140 -2380 44185 -2260
rect 44305 -2380 44360 -2260
rect 44480 -2380 44525 -2260
rect 44645 -2380 44690 -2260
rect 44810 -2380 44855 -2260
rect 44975 -2380 45030 -2260
rect 45150 -2380 45195 -2260
rect 45315 -2380 45360 -2260
rect 45480 -2380 45525 -2260
rect 45645 -2380 45700 -2260
rect 45820 -2380 45865 -2260
rect 45985 -2380 46030 -2260
rect 46150 -2380 46195 -2260
rect 46315 -2380 46370 -2260
rect 46490 -2380 46535 -2260
rect 46655 -2380 46700 -2260
rect 46820 -2380 46865 -2260
rect 46985 -2380 47040 -2260
rect 47160 -2380 47205 -2260
rect 47325 -2380 47370 -2260
rect 47490 -2380 47535 -2260
rect 47655 -2380 47865 -2260
rect 47985 -2380 48040 -2260
rect 48160 -2380 48205 -2260
rect 48325 -2380 48370 -2260
rect 48490 -2380 48535 -2260
rect 48655 -2380 48710 -2260
rect 48830 -2380 48875 -2260
rect 48995 -2380 49040 -2260
rect 49160 -2380 49205 -2260
rect 49325 -2380 49380 -2260
rect 49500 -2380 49545 -2260
rect 49665 -2380 49710 -2260
rect 49830 -2380 49875 -2260
rect 49995 -2380 50050 -2260
rect 50170 -2380 50215 -2260
rect 50335 -2380 50380 -2260
rect 50500 -2380 50545 -2260
rect 50665 -2380 50720 -2260
rect 50840 -2380 50885 -2260
rect 51005 -2380 51050 -2260
rect 51170 -2380 51215 -2260
rect 51335 -2380 51390 -2260
rect 51510 -2380 51555 -2260
rect 51675 -2380 51720 -2260
rect 51840 -2380 51885 -2260
rect 52005 -2380 52060 -2260
rect 52180 -2380 52225 -2260
rect 52345 -2380 52390 -2260
rect 52510 -2380 52555 -2260
rect 52675 -2380 52730 -2260
rect 52850 -2380 52895 -2260
rect 53015 -2380 53060 -2260
rect 53180 -2380 53225 -2260
rect 53345 -2380 53370 -2260
rect 30770 -2425 53370 -2380
rect 30770 -2545 30795 -2425
rect 30915 -2545 30970 -2425
rect 31090 -2545 31135 -2425
rect 31255 -2545 31300 -2425
rect 31420 -2545 31465 -2425
rect 31585 -2545 31640 -2425
rect 31760 -2545 31805 -2425
rect 31925 -2545 31970 -2425
rect 32090 -2545 32135 -2425
rect 32255 -2545 32310 -2425
rect 32430 -2545 32475 -2425
rect 32595 -2545 32640 -2425
rect 32760 -2545 32805 -2425
rect 32925 -2545 32980 -2425
rect 33100 -2545 33145 -2425
rect 33265 -2545 33310 -2425
rect 33430 -2545 33475 -2425
rect 33595 -2545 33650 -2425
rect 33770 -2545 33815 -2425
rect 33935 -2545 33980 -2425
rect 34100 -2545 34145 -2425
rect 34265 -2545 34320 -2425
rect 34440 -2545 34485 -2425
rect 34605 -2545 34650 -2425
rect 34770 -2545 34815 -2425
rect 34935 -2545 34990 -2425
rect 35110 -2545 35155 -2425
rect 35275 -2545 35320 -2425
rect 35440 -2545 35485 -2425
rect 35605 -2545 35660 -2425
rect 35780 -2545 35825 -2425
rect 35945 -2545 35990 -2425
rect 36110 -2545 36155 -2425
rect 36275 -2545 36485 -2425
rect 36605 -2545 36660 -2425
rect 36780 -2545 36825 -2425
rect 36945 -2545 36990 -2425
rect 37110 -2545 37155 -2425
rect 37275 -2545 37330 -2425
rect 37450 -2545 37495 -2425
rect 37615 -2545 37660 -2425
rect 37780 -2545 37825 -2425
rect 37945 -2545 38000 -2425
rect 38120 -2545 38165 -2425
rect 38285 -2545 38330 -2425
rect 38450 -2545 38495 -2425
rect 38615 -2545 38670 -2425
rect 38790 -2545 38835 -2425
rect 38955 -2545 39000 -2425
rect 39120 -2545 39165 -2425
rect 39285 -2545 39340 -2425
rect 39460 -2545 39505 -2425
rect 39625 -2545 39670 -2425
rect 39790 -2545 39835 -2425
rect 39955 -2545 40010 -2425
rect 40130 -2545 40175 -2425
rect 40295 -2545 40340 -2425
rect 40460 -2545 40505 -2425
rect 40625 -2545 40680 -2425
rect 40800 -2545 40845 -2425
rect 40965 -2545 41010 -2425
rect 41130 -2545 41175 -2425
rect 41295 -2545 41350 -2425
rect 41470 -2545 41515 -2425
rect 41635 -2545 41680 -2425
rect 41800 -2545 41845 -2425
rect 41965 -2545 42175 -2425
rect 42295 -2545 42350 -2425
rect 42470 -2545 42515 -2425
rect 42635 -2545 42680 -2425
rect 42800 -2545 42845 -2425
rect 42965 -2545 43020 -2425
rect 43140 -2545 43185 -2425
rect 43305 -2545 43350 -2425
rect 43470 -2545 43515 -2425
rect 43635 -2545 43690 -2425
rect 43810 -2545 43855 -2425
rect 43975 -2545 44020 -2425
rect 44140 -2545 44185 -2425
rect 44305 -2545 44360 -2425
rect 44480 -2545 44525 -2425
rect 44645 -2545 44690 -2425
rect 44810 -2545 44855 -2425
rect 44975 -2545 45030 -2425
rect 45150 -2545 45195 -2425
rect 45315 -2545 45360 -2425
rect 45480 -2545 45525 -2425
rect 45645 -2545 45700 -2425
rect 45820 -2545 45865 -2425
rect 45985 -2545 46030 -2425
rect 46150 -2545 46195 -2425
rect 46315 -2545 46370 -2425
rect 46490 -2545 46535 -2425
rect 46655 -2545 46700 -2425
rect 46820 -2545 46865 -2425
rect 46985 -2545 47040 -2425
rect 47160 -2545 47205 -2425
rect 47325 -2545 47370 -2425
rect 47490 -2545 47535 -2425
rect 47655 -2545 47865 -2425
rect 47985 -2545 48040 -2425
rect 48160 -2545 48205 -2425
rect 48325 -2545 48370 -2425
rect 48490 -2545 48535 -2425
rect 48655 -2545 48710 -2425
rect 48830 -2545 48875 -2425
rect 48995 -2545 49040 -2425
rect 49160 -2545 49205 -2425
rect 49325 -2545 49380 -2425
rect 49500 -2545 49545 -2425
rect 49665 -2545 49710 -2425
rect 49830 -2545 49875 -2425
rect 49995 -2545 50050 -2425
rect 50170 -2545 50215 -2425
rect 50335 -2545 50380 -2425
rect 50500 -2545 50545 -2425
rect 50665 -2545 50720 -2425
rect 50840 -2545 50885 -2425
rect 51005 -2545 51050 -2425
rect 51170 -2545 51215 -2425
rect 51335 -2545 51390 -2425
rect 51510 -2545 51555 -2425
rect 51675 -2545 51720 -2425
rect 51840 -2545 51885 -2425
rect 52005 -2545 52060 -2425
rect 52180 -2545 52225 -2425
rect 52345 -2545 52390 -2425
rect 52510 -2545 52555 -2425
rect 52675 -2545 52730 -2425
rect 52850 -2545 52895 -2425
rect 53015 -2545 53060 -2425
rect 53180 -2545 53225 -2425
rect 53345 -2545 53370 -2425
rect 30770 -2600 53370 -2545
rect 30770 -2720 30795 -2600
rect 30915 -2720 30970 -2600
rect 31090 -2720 31135 -2600
rect 31255 -2720 31300 -2600
rect 31420 -2720 31465 -2600
rect 31585 -2720 31640 -2600
rect 31760 -2720 31805 -2600
rect 31925 -2720 31970 -2600
rect 32090 -2720 32135 -2600
rect 32255 -2720 32310 -2600
rect 32430 -2720 32475 -2600
rect 32595 -2720 32640 -2600
rect 32760 -2720 32805 -2600
rect 32925 -2720 32980 -2600
rect 33100 -2720 33145 -2600
rect 33265 -2720 33310 -2600
rect 33430 -2720 33475 -2600
rect 33595 -2720 33650 -2600
rect 33770 -2720 33815 -2600
rect 33935 -2720 33980 -2600
rect 34100 -2720 34145 -2600
rect 34265 -2720 34320 -2600
rect 34440 -2720 34485 -2600
rect 34605 -2720 34650 -2600
rect 34770 -2720 34815 -2600
rect 34935 -2720 34990 -2600
rect 35110 -2720 35155 -2600
rect 35275 -2720 35320 -2600
rect 35440 -2720 35485 -2600
rect 35605 -2720 35660 -2600
rect 35780 -2720 35825 -2600
rect 35945 -2720 35990 -2600
rect 36110 -2720 36155 -2600
rect 36275 -2720 36485 -2600
rect 36605 -2720 36660 -2600
rect 36780 -2720 36825 -2600
rect 36945 -2720 36990 -2600
rect 37110 -2720 37155 -2600
rect 37275 -2720 37330 -2600
rect 37450 -2720 37495 -2600
rect 37615 -2720 37660 -2600
rect 37780 -2720 37825 -2600
rect 37945 -2720 38000 -2600
rect 38120 -2720 38165 -2600
rect 38285 -2720 38330 -2600
rect 38450 -2720 38495 -2600
rect 38615 -2720 38670 -2600
rect 38790 -2720 38835 -2600
rect 38955 -2720 39000 -2600
rect 39120 -2720 39165 -2600
rect 39285 -2720 39340 -2600
rect 39460 -2720 39505 -2600
rect 39625 -2720 39670 -2600
rect 39790 -2720 39835 -2600
rect 39955 -2720 40010 -2600
rect 40130 -2720 40175 -2600
rect 40295 -2720 40340 -2600
rect 40460 -2720 40505 -2600
rect 40625 -2720 40680 -2600
rect 40800 -2720 40845 -2600
rect 40965 -2720 41010 -2600
rect 41130 -2720 41175 -2600
rect 41295 -2720 41350 -2600
rect 41470 -2720 41515 -2600
rect 41635 -2720 41680 -2600
rect 41800 -2720 41845 -2600
rect 41965 -2720 42175 -2600
rect 42295 -2720 42350 -2600
rect 42470 -2720 42515 -2600
rect 42635 -2720 42680 -2600
rect 42800 -2720 42845 -2600
rect 42965 -2720 43020 -2600
rect 43140 -2720 43185 -2600
rect 43305 -2720 43350 -2600
rect 43470 -2720 43515 -2600
rect 43635 -2720 43690 -2600
rect 43810 -2720 43855 -2600
rect 43975 -2720 44020 -2600
rect 44140 -2720 44185 -2600
rect 44305 -2720 44360 -2600
rect 44480 -2720 44525 -2600
rect 44645 -2720 44690 -2600
rect 44810 -2720 44855 -2600
rect 44975 -2720 45030 -2600
rect 45150 -2720 45195 -2600
rect 45315 -2720 45360 -2600
rect 45480 -2720 45525 -2600
rect 45645 -2720 45700 -2600
rect 45820 -2720 45865 -2600
rect 45985 -2720 46030 -2600
rect 46150 -2720 46195 -2600
rect 46315 -2720 46370 -2600
rect 46490 -2720 46535 -2600
rect 46655 -2720 46700 -2600
rect 46820 -2720 46865 -2600
rect 46985 -2720 47040 -2600
rect 47160 -2720 47205 -2600
rect 47325 -2720 47370 -2600
rect 47490 -2720 47535 -2600
rect 47655 -2720 47865 -2600
rect 47985 -2720 48040 -2600
rect 48160 -2720 48205 -2600
rect 48325 -2720 48370 -2600
rect 48490 -2720 48535 -2600
rect 48655 -2720 48710 -2600
rect 48830 -2720 48875 -2600
rect 48995 -2720 49040 -2600
rect 49160 -2720 49205 -2600
rect 49325 -2720 49380 -2600
rect 49500 -2720 49545 -2600
rect 49665 -2720 49710 -2600
rect 49830 -2720 49875 -2600
rect 49995 -2720 50050 -2600
rect 50170 -2720 50215 -2600
rect 50335 -2720 50380 -2600
rect 50500 -2720 50545 -2600
rect 50665 -2720 50720 -2600
rect 50840 -2720 50885 -2600
rect 51005 -2720 51050 -2600
rect 51170 -2720 51215 -2600
rect 51335 -2720 51390 -2600
rect 51510 -2720 51555 -2600
rect 51675 -2720 51720 -2600
rect 51840 -2720 51885 -2600
rect 52005 -2720 52060 -2600
rect 52180 -2720 52225 -2600
rect 52345 -2720 52390 -2600
rect 52510 -2720 52555 -2600
rect 52675 -2720 52730 -2600
rect 52850 -2720 52895 -2600
rect 53015 -2720 53060 -2600
rect 53180 -2720 53225 -2600
rect 53345 -2720 53370 -2600
rect 30770 -2765 53370 -2720
rect 30770 -2885 30795 -2765
rect 30915 -2885 30970 -2765
rect 31090 -2885 31135 -2765
rect 31255 -2885 31300 -2765
rect 31420 -2885 31465 -2765
rect 31585 -2885 31640 -2765
rect 31760 -2885 31805 -2765
rect 31925 -2885 31970 -2765
rect 32090 -2885 32135 -2765
rect 32255 -2885 32310 -2765
rect 32430 -2885 32475 -2765
rect 32595 -2885 32640 -2765
rect 32760 -2885 32805 -2765
rect 32925 -2885 32980 -2765
rect 33100 -2885 33145 -2765
rect 33265 -2885 33310 -2765
rect 33430 -2885 33475 -2765
rect 33595 -2885 33650 -2765
rect 33770 -2885 33815 -2765
rect 33935 -2885 33980 -2765
rect 34100 -2885 34145 -2765
rect 34265 -2885 34320 -2765
rect 34440 -2885 34485 -2765
rect 34605 -2885 34650 -2765
rect 34770 -2885 34815 -2765
rect 34935 -2885 34990 -2765
rect 35110 -2885 35155 -2765
rect 35275 -2885 35320 -2765
rect 35440 -2885 35485 -2765
rect 35605 -2885 35660 -2765
rect 35780 -2885 35825 -2765
rect 35945 -2885 35990 -2765
rect 36110 -2885 36155 -2765
rect 36275 -2885 36485 -2765
rect 36605 -2885 36660 -2765
rect 36780 -2885 36825 -2765
rect 36945 -2885 36990 -2765
rect 37110 -2885 37155 -2765
rect 37275 -2885 37330 -2765
rect 37450 -2885 37495 -2765
rect 37615 -2885 37660 -2765
rect 37780 -2885 37825 -2765
rect 37945 -2885 38000 -2765
rect 38120 -2885 38165 -2765
rect 38285 -2885 38330 -2765
rect 38450 -2885 38495 -2765
rect 38615 -2885 38670 -2765
rect 38790 -2885 38835 -2765
rect 38955 -2885 39000 -2765
rect 39120 -2885 39165 -2765
rect 39285 -2885 39340 -2765
rect 39460 -2885 39505 -2765
rect 39625 -2885 39670 -2765
rect 39790 -2885 39835 -2765
rect 39955 -2885 40010 -2765
rect 40130 -2885 40175 -2765
rect 40295 -2885 40340 -2765
rect 40460 -2885 40505 -2765
rect 40625 -2885 40680 -2765
rect 40800 -2885 40845 -2765
rect 40965 -2885 41010 -2765
rect 41130 -2885 41175 -2765
rect 41295 -2885 41350 -2765
rect 41470 -2885 41515 -2765
rect 41635 -2885 41680 -2765
rect 41800 -2885 41845 -2765
rect 41965 -2885 42175 -2765
rect 42295 -2885 42350 -2765
rect 42470 -2885 42515 -2765
rect 42635 -2885 42680 -2765
rect 42800 -2885 42845 -2765
rect 42965 -2885 43020 -2765
rect 43140 -2885 43185 -2765
rect 43305 -2885 43350 -2765
rect 43470 -2885 43515 -2765
rect 43635 -2885 43690 -2765
rect 43810 -2885 43855 -2765
rect 43975 -2885 44020 -2765
rect 44140 -2885 44185 -2765
rect 44305 -2885 44360 -2765
rect 44480 -2885 44525 -2765
rect 44645 -2885 44690 -2765
rect 44810 -2885 44855 -2765
rect 44975 -2885 45030 -2765
rect 45150 -2885 45195 -2765
rect 45315 -2885 45360 -2765
rect 45480 -2885 45525 -2765
rect 45645 -2885 45700 -2765
rect 45820 -2885 45865 -2765
rect 45985 -2885 46030 -2765
rect 46150 -2885 46195 -2765
rect 46315 -2885 46370 -2765
rect 46490 -2885 46535 -2765
rect 46655 -2885 46700 -2765
rect 46820 -2885 46865 -2765
rect 46985 -2885 47040 -2765
rect 47160 -2885 47205 -2765
rect 47325 -2885 47370 -2765
rect 47490 -2885 47535 -2765
rect 47655 -2885 47865 -2765
rect 47985 -2885 48040 -2765
rect 48160 -2885 48205 -2765
rect 48325 -2885 48370 -2765
rect 48490 -2885 48535 -2765
rect 48655 -2885 48710 -2765
rect 48830 -2885 48875 -2765
rect 48995 -2885 49040 -2765
rect 49160 -2885 49205 -2765
rect 49325 -2885 49380 -2765
rect 49500 -2885 49545 -2765
rect 49665 -2885 49710 -2765
rect 49830 -2885 49875 -2765
rect 49995 -2885 50050 -2765
rect 50170 -2885 50215 -2765
rect 50335 -2885 50380 -2765
rect 50500 -2885 50545 -2765
rect 50665 -2885 50720 -2765
rect 50840 -2885 50885 -2765
rect 51005 -2885 51050 -2765
rect 51170 -2885 51215 -2765
rect 51335 -2885 51390 -2765
rect 51510 -2885 51555 -2765
rect 51675 -2885 51720 -2765
rect 51840 -2885 51885 -2765
rect 52005 -2885 52060 -2765
rect 52180 -2885 52225 -2765
rect 52345 -2885 52390 -2765
rect 52510 -2885 52555 -2765
rect 52675 -2885 52730 -2765
rect 52850 -2885 52895 -2765
rect 53015 -2885 53060 -2765
rect 53180 -2885 53225 -2765
rect 53345 -2885 53370 -2765
rect 30770 -2930 53370 -2885
rect 30770 -3050 30795 -2930
rect 30915 -3050 30970 -2930
rect 31090 -3050 31135 -2930
rect 31255 -3050 31300 -2930
rect 31420 -3050 31465 -2930
rect 31585 -3050 31640 -2930
rect 31760 -3050 31805 -2930
rect 31925 -3050 31970 -2930
rect 32090 -3050 32135 -2930
rect 32255 -3050 32310 -2930
rect 32430 -3050 32475 -2930
rect 32595 -3050 32640 -2930
rect 32760 -3050 32805 -2930
rect 32925 -3050 32980 -2930
rect 33100 -3050 33145 -2930
rect 33265 -3050 33310 -2930
rect 33430 -3050 33475 -2930
rect 33595 -3050 33650 -2930
rect 33770 -3050 33815 -2930
rect 33935 -3050 33980 -2930
rect 34100 -3050 34145 -2930
rect 34265 -3050 34320 -2930
rect 34440 -3050 34485 -2930
rect 34605 -3050 34650 -2930
rect 34770 -3050 34815 -2930
rect 34935 -3050 34990 -2930
rect 35110 -3050 35155 -2930
rect 35275 -3050 35320 -2930
rect 35440 -3050 35485 -2930
rect 35605 -3050 35660 -2930
rect 35780 -3050 35825 -2930
rect 35945 -3050 35990 -2930
rect 36110 -3050 36155 -2930
rect 36275 -3050 36485 -2930
rect 36605 -3050 36660 -2930
rect 36780 -3050 36825 -2930
rect 36945 -3050 36990 -2930
rect 37110 -3050 37155 -2930
rect 37275 -3050 37330 -2930
rect 37450 -3050 37495 -2930
rect 37615 -3050 37660 -2930
rect 37780 -3050 37825 -2930
rect 37945 -3050 38000 -2930
rect 38120 -3050 38165 -2930
rect 38285 -3050 38330 -2930
rect 38450 -3050 38495 -2930
rect 38615 -3050 38670 -2930
rect 38790 -3050 38835 -2930
rect 38955 -3050 39000 -2930
rect 39120 -3050 39165 -2930
rect 39285 -3050 39340 -2930
rect 39460 -3050 39505 -2930
rect 39625 -3050 39670 -2930
rect 39790 -3050 39835 -2930
rect 39955 -3050 40010 -2930
rect 40130 -3050 40175 -2930
rect 40295 -3050 40340 -2930
rect 40460 -3050 40505 -2930
rect 40625 -3050 40680 -2930
rect 40800 -3050 40845 -2930
rect 40965 -3050 41010 -2930
rect 41130 -3050 41175 -2930
rect 41295 -3050 41350 -2930
rect 41470 -3050 41515 -2930
rect 41635 -3050 41680 -2930
rect 41800 -3050 41845 -2930
rect 41965 -3050 42175 -2930
rect 42295 -3050 42350 -2930
rect 42470 -3050 42515 -2930
rect 42635 -3050 42680 -2930
rect 42800 -3050 42845 -2930
rect 42965 -3050 43020 -2930
rect 43140 -3050 43185 -2930
rect 43305 -3050 43350 -2930
rect 43470 -3050 43515 -2930
rect 43635 -3050 43690 -2930
rect 43810 -3050 43855 -2930
rect 43975 -3050 44020 -2930
rect 44140 -3050 44185 -2930
rect 44305 -3050 44360 -2930
rect 44480 -3050 44525 -2930
rect 44645 -3050 44690 -2930
rect 44810 -3050 44855 -2930
rect 44975 -3050 45030 -2930
rect 45150 -3050 45195 -2930
rect 45315 -3050 45360 -2930
rect 45480 -3050 45525 -2930
rect 45645 -3050 45700 -2930
rect 45820 -3050 45865 -2930
rect 45985 -3050 46030 -2930
rect 46150 -3050 46195 -2930
rect 46315 -3050 46370 -2930
rect 46490 -3050 46535 -2930
rect 46655 -3050 46700 -2930
rect 46820 -3050 46865 -2930
rect 46985 -3050 47040 -2930
rect 47160 -3050 47205 -2930
rect 47325 -3050 47370 -2930
rect 47490 -3050 47535 -2930
rect 47655 -3050 47865 -2930
rect 47985 -3050 48040 -2930
rect 48160 -3050 48205 -2930
rect 48325 -3050 48370 -2930
rect 48490 -3050 48535 -2930
rect 48655 -3050 48710 -2930
rect 48830 -3050 48875 -2930
rect 48995 -3050 49040 -2930
rect 49160 -3050 49205 -2930
rect 49325 -3050 49380 -2930
rect 49500 -3050 49545 -2930
rect 49665 -3050 49710 -2930
rect 49830 -3050 49875 -2930
rect 49995 -3050 50050 -2930
rect 50170 -3050 50215 -2930
rect 50335 -3050 50380 -2930
rect 50500 -3050 50545 -2930
rect 50665 -3050 50720 -2930
rect 50840 -3050 50885 -2930
rect 51005 -3050 51050 -2930
rect 51170 -3050 51215 -2930
rect 51335 -3050 51390 -2930
rect 51510 -3050 51555 -2930
rect 51675 -3050 51720 -2930
rect 51840 -3050 51885 -2930
rect 52005 -3050 52060 -2930
rect 52180 -3050 52225 -2930
rect 52345 -3050 52390 -2930
rect 52510 -3050 52555 -2930
rect 52675 -3050 52730 -2930
rect 52850 -3050 52895 -2930
rect 53015 -3050 53060 -2930
rect 53180 -3050 53225 -2930
rect 53345 -3050 53370 -2930
rect 30770 -3095 53370 -3050
rect 30770 -3215 30795 -3095
rect 30915 -3215 30970 -3095
rect 31090 -3215 31135 -3095
rect 31255 -3215 31300 -3095
rect 31420 -3215 31465 -3095
rect 31585 -3215 31640 -3095
rect 31760 -3215 31805 -3095
rect 31925 -3215 31970 -3095
rect 32090 -3215 32135 -3095
rect 32255 -3215 32310 -3095
rect 32430 -3215 32475 -3095
rect 32595 -3215 32640 -3095
rect 32760 -3215 32805 -3095
rect 32925 -3215 32980 -3095
rect 33100 -3215 33145 -3095
rect 33265 -3215 33310 -3095
rect 33430 -3215 33475 -3095
rect 33595 -3215 33650 -3095
rect 33770 -3215 33815 -3095
rect 33935 -3215 33980 -3095
rect 34100 -3215 34145 -3095
rect 34265 -3215 34320 -3095
rect 34440 -3215 34485 -3095
rect 34605 -3215 34650 -3095
rect 34770 -3215 34815 -3095
rect 34935 -3215 34990 -3095
rect 35110 -3215 35155 -3095
rect 35275 -3215 35320 -3095
rect 35440 -3215 35485 -3095
rect 35605 -3215 35660 -3095
rect 35780 -3215 35825 -3095
rect 35945 -3215 35990 -3095
rect 36110 -3215 36155 -3095
rect 36275 -3215 36485 -3095
rect 36605 -3215 36660 -3095
rect 36780 -3215 36825 -3095
rect 36945 -3215 36990 -3095
rect 37110 -3215 37155 -3095
rect 37275 -3215 37330 -3095
rect 37450 -3215 37495 -3095
rect 37615 -3215 37660 -3095
rect 37780 -3215 37825 -3095
rect 37945 -3215 38000 -3095
rect 38120 -3215 38165 -3095
rect 38285 -3215 38330 -3095
rect 38450 -3215 38495 -3095
rect 38615 -3215 38670 -3095
rect 38790 -3215 38835 -3095
rect 38955 -3215 39000 -3095
rect 39120 -3215 39165 -3095
rect 39285 -3215 39340 -3095
rect 39460 -3215 39505 -3095
rect 39625 -3215 39670 -3095
rect 39790 -3215 39835 -3095
rect 39955 -3215 40010 -3095
rect 40130 -3215 40175 -3095
rect 40295 -3215 40340 -3095
rect 40460 -3215 40505 -3095
rect 40625 -3215 40680 -3095
rect 40800 -3215 40845 -3095
rect 40965 -3215 41010 -3095
rect 41130 -3215 41175 -3095
rect 41295 -3215 41350 -3095
rect 41470 -3215 41515 -3095
rect 41635 -3215 41680 -3095
rect 41800 -3215 41845 -3095
rect 41965 -3215 42175 -3095
rect 42295 -3215 42350 -3095
rect 42470 -3215 42515 -3095
rect 42635 -3215 42680 -3095
rect 42800 -3215 42845 -3095
rect 42965 -3215 43020 -3095
rect 43140 -3215 43185 -3095
rect 43305 -3215 43350 -3095
rect 43470 -3215 43515 -3095
rect 43635 -3215 43690 -3095
rect 43810 -3215 43855 -3095
rect 43975 -3215 44020 -3095
rect 44140 -3215 44185 -3095
rect 44305 -3215 44360 -3095
rect 44480 -3215 44525 -3095
rect 44645 -3215 44690 -3095
rect 44810 -3215 44855 -3095
rect 44975 -3215 45030 -3095
rect 45150 -3215 45195 -3095
rect 45315 -3215 45360 -3095
rect 45480 -3215 45525 -3095
rect 45645 -3215 45700 -3095
rect 45820 -3215 45865 -3095
rect 45985 -3215 46030 -3095
rect 46150 -3215 46195 -3095
rect 46315 -3215 46370 -3095
rect 46490 -3215 46535 -3095
rect 46655 -3215 46700 -3095
rect 46820 -3215 46865 -3095
rect 46985 -3215 47040 -3095
rect 47160 -3215 47205 -3095
rect 47325 -3215 47370 -3095
rect 47490 -3215 47535 -3095
rect 47655 -3215 47865 -3095
rect 47985 -3215 48040 -3095
rect 48160 -3215 48205 -3095
rect 48325 -3215 48370 -3095
rect 48490 -3215 48535 -3095
rect 48655 -3215 48710 -3095
rect 48830 -3215 48875 -3095
rect 48995 -3215 49040 -3095
rect 49160 -3215 49205 -3095
rect 49325 -3215 49380 -3095
rect 49500 -3215 49545 -3095
rect 49665 -3215 49710 -3095
rect 49830 -3215 49875 -3095
rect 49995 -3215 50050 -3095
rect 50170 -3215 50215 -3095
rect 50335 -3215 50380 -3095
rect 50500 -3215 50545 -3095
rect 50665 -3215 50720 -3095
rect 50840 -3215 50885 -3095
rect 51005 -3215 51050 -3095
rect 51170 -3215 51215 -3095
rect 51335 -3215 51390 -3095
rect 51510 -3215 51555 -3095
rect 51675 -3215 51720 -3095
rect 51840 -3215 51885 -3095
rect 52005 -3215 52060 -3095
rect 52180 -3215 52225 -3095
rect 52345 -3215 52390 -3095
rect 52510 -3215 52555 -3095
rect 52675 -3215 52730 -3095
rect 52850 -3215 52895 -3095
rect 53015 -3215 53060 -3095
rect 53180 -3215 53225 -3095
rect 53345 -3215 53370 -3095
rect 30770 -3270 53370 -3215
rect 30770 -3390 30795 -3270
rect 30915 -3390 30970 -3270
rect 31090 -3390 31135 -3270
rect 31255 -3390 31300 -3270
rect 31420 -3390 31465 -3270
rect 31585 -3390 31640 -3270
rect 31760 -3390 31805 -3270
rect 31925 -3390 31970 -3270
rect 32090 -3390 32135 -3270
rect 32255 -3390 32310 -3270
rect 32430 -3390 32475 -3270
rect 32595 -3390 32640 -3270
rect 32760 -3390 32805 -3270
rect 32925 -3390 32980 -3270
rect 33100 -3390 33145 -3270
rect 33265 -3390 33310 -3270
rect 33430 -3390 33475 -3270
rect 33595 -3390 33650 -3270
rect 33770 -3390 33815 -3270
rect 33935 -3390 33980 -3270
rect 34100 -3390 34145 -3270
rect 34265 -3390 34320 -3270
rect 34440 -3390 34485 -3270
rect 34605 -3390 34650 -3270
rect 34770 -3390 34815 -3270
rect 34935 -3390 34990 -3270
rect 35110 -3390 35155 -3270
rect 35275 -3390 35320 -3270
rect 35440 -3390 35485 -3270
rect 35605 -3390 35660 -3270
rect 35780 -3390 35825 -3270
rect 35945 -3390 35990 -3270
rect 36110 -3390 36155 -3270
rect 36275 -3390 36485 -3270
rect 36605 -3390 36660 -3270
rect 36780 -3390 36825 -3270
rect 36945 -3390 36990 -3270
rect 37110 -3390 37155 -3270
rect 37275 -3390 37330 -3270
rect 37450 -3390 37495 -3270
rect 37615 -3390 37660 -3270
rect 37780 -3390 37825 -3270
rect 37945 -3390 38000 -3270
rect 38120 -3390 38165 -3270
rect 38285 -3390 38330 -3270
rect 38450 -3390 38495 -3270
rect 38615 -3390 38670 -3270
rect 38790 -3390 38835 -3270
rect 38955 -3390 39000 -3270
rect 39120 -3390 39165 -3270
rect 39285 -3390 39340 -3270
rect 39460 -3390 39505 -3270
rect 39625 -3390 39670 -3270
rect 39790 -3390 39835 -3270
rect 39955 -3390 40010 -3270
rect 40130 -3390 40175 -3270
rect 40295 -3390 40340 -3270
rect 40460 -3390 40505 -3270
rect 40625 -3390 40680 -3270
rect 40800 -3390 40845 -3270
rect 40965 -3390 41010 -3270
rect 41130 -3390 41175 -3270
rect 41295 -3390 41350 -3270
rect 41470 -3390 41515 -3270
rect 41635 -3390 41680 -3270
rect 41800 -3390 41845 -3270
rect 41965 -3390 42175 -3270
rect 42295 -3390 42350 -3270
rect 42470 -3390 42515 -3270
rect 42635 -3390 42680 -3270
rect 42800 -3390 42845 -3270
rect 42965 -3390 43020 -3270
rect 43140 -3390 43185 -3270
rect 43305 -3390 43350 -3270
rect 43470 -3390 43515 -3270
rect 43635 -3390 43690 -3270
rect 43810 -3390 43855 -3270
rect 43975 -3390 44020 -3270
rect 44140 -3390 44185 -3270
rect 44305 -3390 44360 -3270
rect 44480 -3390 44525 -3270
rect 44645 -3390 44690 -3270
rect 44810 -3390 44855 -3270
rect 44975 -3390 45030 -3270
rect 45150 -3390 45195 -3270
rect 45315 -3390 45360 -3270
rect 45480 -3390 45525 -3270
rect 45645 -3390 45700 -3270
rect 45820 -3390 45865 -3270
rect 45985 -3390 46030 -3270
rect 46150 -3390 46195 -3270
rect 46315 -3390 46370 -3270
rect 46490 -3390 46535 -3270
rect 46655 -3390 46700 -3270
rect 46820 -3390 46865 -3270
rect 46985 -3390 47040 -3270
rect 47160 -3390 47205 -3270
rect 47325 -3390 47370 -3270
rect 47490 -3390 47535 -3270
rect 47655 -3390 47865 -3270
rect 47985 -3390 48040 -3270
rect 48160 -3390 48205 -3270
rect 48325 -3390 48370 -3270
rect 48490 -3390 48535 -3270
rect 48655 -3390 48710 -3270
rect 48830 -3390 48875 -3270
rect 48995 -3390 49040 -3270
rect 49160 -3390 49205 -3270
rect 49325 -3390 49380 -3270
rect 49500 -3390 49545 -3270
rect 49665 -3390 49710 -3270
rect 49830 -3390 49875 -3270
rect 49995 -3390 50050 -3270
rect 50170 -3390 50215 -3270
rect 50335 -3390 50380 -3270
rect 50500 -3390 50545 -3270
rect 50665 -3390 50720 -3270
rect 50840 -3390 50885 -3270
rect 51005 -3390 51050 -3270
rect 51170 -3390 51215 -3270
rect 51335 -3390 51390 -3270
rect 51510 -3390 51555 -3270
rect 51675 -3390 51720 -3270
rect 51840 -3390 51885 -3270
rect 52005 -3390 52060 -3270
rect 52180 -3390 52225 -3270
rect 52345 -3390 52390 -3270
rect 52510 -3390 52555 -3270
rect 52675 -3390 52730 -3270
rect 52850 -3390 52895 -3270
rect 53015 -3390 53060 -3270
rect 53180 -3390 53225 -3270
rect 53345 -3390 53370 -3270
rect 30770 -3435 53370 -3390
rect 30770 -3555 30795 -3435
rect 30915 -3555 30970 -3435
rect 31090 -3555 31135 -3435
rect 31255 -3555 31300 -3435
rect 31420 -3555 31465 -3435
rect 31585 -3555 31640 -3435
rect 31760 -3555 31805 -3435
rect 31925 -3555 31970 -3435
rect 32090 -3555 32135 -3435
rect 32255 -3555 32310 -3435
rect 32430 -3555 32475 -3435
rect 32595 -3555 32640 -3435
rect 32760 -3555 32805 -3435
rect 32925 -3555 32980 -3435
rect 33100 -3555 33145 -3435
rect 33265 -3555 33310 -3435
rect 33430 -3555 33475 -3435
rect 33595 -3555 33650 -3435
rect 33770 -3555 33815 -3435
rect 33935 -3555 33980 -3435
rect 34100 -3555 34145 -3435
rect 34265 -3555 34320 -3435
rect 34440 -3555 34485 -3435
rect 34605 -3555 34650 -3435
rect 34770 -3555 34815 -3435
rect 34935 -3555 34990 -3435
rect 35110 -3555 35155 -3435
rect 35275 -3555 35320 -3435
rect 35440 -3555 35485 -3435
rect 35605 -3555 35660 -3435
rect 35780 -3555 35825 -3435
rect 35945 -3555 35990 -3435
rect 36110 -3555 36155 -3435
rect 36275 -3555 36485 -3435
rect 36605 -3555 36660 -3435
rect 36780 -3555 36825 -3435
rect 36945 -3555 36990 -3435
rect 37110 -3555 37155 -3435
rect 37275 -3555 37330 -3435
rect 37450 -3555 37495 -3435
rect 37615 -3555 37660 -3435
rect 37780 -3555 37825 -3435
rect 37945 -3555 38000 -3435
rect 38120 -3555 38165 -3435
rect 38285 -3555 38330 -3435
rect 38450 -3555 38495 -3435
rect 38615 -3555 38670 -3435
rect 38790 -3555 38835 -3435
rect 38955 -3555 39000 -3435
rect 39120 -3555 39165 -3435
rect 39285 -3555 39340 -3435
rect 39460 -3555 39505 -3435
rect 39625 -3555 39670 -3435
rect 39790 -3555 39835 -3435
rect 39955 -3555 40010 -3435
rect 40130 -3555 40175 -3435
rect 40295 -3555 40340 -3435
rect 40460 -3555 40505 -3435
rect 40625 -3555 40680 -3435
rect 40800 -3555 40845 -3435
rect 40965 -3555 41010 -3435
rect 41130 -3555 41175 -3435
rect 41295 -3555 41350 -3435
rect 41470 -3555 41515 -3435
rect 41635 -3555 41680 -3435
rect 41800 -3555 41845 -3435
rect 41965 -3555 42175 -3435
rect 42295 -3555 42350 -3435
rect 42470 -3555 42515 -3435
rect 42635 -3555 42680 -3435
rect 42800 -3555 42845 -3435
rect 42965 -3555 43020 -3435
rect 43140 -3555 43185 -3435
rect 43305 -3555 43350 -3435
rect 43470 -3555 43515 -3435
rect 43635 -3555 43690 -3435
rect 43810 -3555 43855 -3435
rect 43975 -3555 44020 -3435
rect 44140 -3555 44185 -3435
rect 44305 -3555 44360 -3435
rect 44480 -3555 44525 -3435
rect 44645 -3555 44690 -3435
rect 44810 -3555 44855 -3435
rect 44975 -3555 45030 -3435
rect 45150 -3555 45195 -3435
rect 45315 -3555 45360 -3435
rect 45480 -3555 45525 -3435
rect 45645 -3555 45700 -3435
rect 45820 -3555 45865 -3435
rect 45985 -3555 46030 -3435
rect 46150 -3555 46195 -3435
rect 46315 -3555 46370 -3435
rect 46490 -3555 46535 -3435
rect 46655 -3555 46700 -3435
rect 46820 -3555 46865 -3435
rect 46985 -3555 47040 -3435
rect 47160 -3555 47205 -3435
rect 47325 -3555 47370 -3435
rect 47490 -3555 47535 -3435
rect 47655 -3555 47865 -3435
rect 47985 -3555 48040 -3435
rect 48160 -3555 48205 -3435
rect 48325 -3555 48370 -3435
rect 48490 -3555 48535 -3435
rect 48655 -3555 48710 -3435
rect 48830 -3555 48875 -3435
rect 48995 -3555 49040 -3435
rect 49160 -3555 49205 -3435
rect 49325 -3555 49380 -3435
rect 49500 -3555 49545 -3435
rect 49665 -3555 49710 -3435
rect 49830 -3555 49875 -3435
rect 49995 -3555 50050 -3435
rect 50170 -3555 50215 -3435
rect 50335 -3555 50380 -3435
rect 50500 -3555 50545 -3435
rect 50665 -3555 50720 -3435
rect 50840 -3555 50885 -3435
rect 51005 -3555 51050 -3435
rect 51170 -3555 51215 -3435
rect 51335 -3555 51390 -3435
rect 51510 -3555 51555 -3435
rect 51675 -3555 51720 -3435
rect 51840 -3555 51885 -3435
rect 52005 -3555 52060 -3435
rect 52180 -3555 52225 -3435
rect 52345 -3555 52390 -3435
rect 52510 -3555 52555 -3435
rect 52675 -3555 52730 -3435
rect 52850 -3555 52895 -3435
rect 53015 -3555 53060 -3435
rect 53180 -3555 53225 -3435
rect 53345 -3555 53370 -3435
rect 30770 -3600 53370 -3555
rect 30770 -3720 30795 -3600
rect 30915 -3720 30970 -3600
rect 31090 -3720 31135 -3600
rect 31255 -3720 31300 -3600
rect 31420 -3720 31465 -3600
rect 31585 -3720 31640 -3600
rect 31760 -3720 31805 -3600
rect 31925 -3720 31970 -3600
rect 32090 -3720 32135 -3600
rect 32255 -3720 32310 -3600
rect 32430 -3720 32475 -3600
rect 32595 -3720 32640 -3600
rect 32760 -3720 32805 -3600
rect 32925 -3720 32980 -3600
rect 33100 -3720 33145 -3600
rect 33265 -3720 33310 -3600
rect 33430 -3720 33475 -3600
rect 33595 -3720 33650 -3600
rect 33770 -3720 33815 -3600
rect 33935 -3720 33980 -3600
rect 34100 -3720 34145 -3600
rect 34265 -3720 34320 -3600
rect 34440 -3720 34485 -3600
rect 34605 -3720 34650 -3600
rect 34770 -3720 34815 -3600
rect 34935 -3720 34990 -3600
rect 35110 -3720 35155 -3600
rect 35275 -3720 35320 -3600
rect 35440 -3720 35485 -3600
rect 35605 -3720 35660 -3600
rect 35780 -3720 35825 -3600
rect 35945 -3720 35990 -3600
rect 36110 -3720 36155 -3600
rect 36275 -3720 36485 -3600
rect 36605 -3720 36660 -3600
rect 36780 -3720 36825 -3600
rect 36945 -3720 36990 -3600
rect 37110 -3720 37155 -3600
rect 37275 -3720 37330 -3600
rect 37450 -3720 37495 -3600
rect 37615 -3720 37660 -3600
rect 37780 -3720 37825 -3600
rect 37945 -3720 38000 -3600
rect 38120 -3720 38165 -3600
rect 38285 -3720 38330 -3600
rect 38450 -3720 38495 -3600
rect 38615 -3720 38670 -3600
rect 38790 -3720 38835 -3600
rect 38955 -3720 39000 -3600
rect 39120 -3720 39165 -3600
rect 39285 -3720 39340 -3600
rect 39460 -3720 39505 -3600
rect 39625 -3720 39670 -3600
rect 39790 -3720 39835 -3600
rect 39955 -3720 40010 -3600
rect 40130 -3720 40175 -3600
rect 40295 -3720 40340 -3600
rect 40460 -3720 40505 -3600
rect 40625 -3720 40680 -3600
rect 40800 -3720 40845 -3600
rect 40965 -3720 41010 -3600
rect 41130 -3720 41175 -3600
rect 41295 -3720 41350 -3600
rect 41470 -3720 41515 -3600
rect 41635 -3720 41680 -3600
rect 41800 -3720 41845 -3600
rect 41965 -3720 42175 -3600
rect 42295 -3720 42350 -3600
rect 42470 -3720 42515 -3600
rect 42635 -3720 42680 -3600
rect 42800 -3720 42845 -3600
rect 42965 -3720 43020 -3600
rect 43140 -3720 43185 -3600
rect 43305 -3720 43350 -3600
rect 43470 -3720 43515 -3600
rect 43635 -3720 43690 -3600
rect 43810 -3720 43855 -3600
rect 43975 -3720 44020 -3600
rect 44140 -3720 44185 -3600
rect 44305 -3720 44360 -3600
rect 44480 -3720 44525 -3600
rect 44645 -3720 44690 -3600
rect 44810 -3720 44855 -3600
rect 44975 -3720 45030 -3600
rect 45150 -3720 45195 -3600
rect 45315 -3720 45360 -3600
rect 45480 -3720 45525 -3600
rect 45645 -3720 45700 -3600
rect 45820 -3720 45865 -3600
rect 45985 -3720 46030 -3600
rect 46150 -3720 46195 -3600
rect 46315 -3720 46370 -3600
rect 46490 -3720 46535 -3600
rect 46655 -3720 46700 -3600
rect 46820 -3720 46865 -3600
rect 46985 -3720 47040 -3600
rect 47160 -3720 47205 -3600
rect 47325 -3720 47370 -3600
rect 47490 -3720 47535 -3600
rect 47655 -3720 47865 -3600
rect 47985 -3720 48040 -3600
rect 48160 -3720 48205 -3600
rect 48325 -3720 48370 -3600
rect 48490 -3720 48535 -3600
rect 48655 -3720 48710 -3600
rect 48830 -3720 48875 -3600
rect 48995 -3720 49040 -3600
rect 49160 -3720 49205 -3600
rect 49325 -3720 49380 -3600
rect 49500 -3720 49545 -3600
rect 49665 -3720 49710 -3600
rect 49830 -3720 49875 -3600
rect 49995 -3720 50050 -3600
rect 50170 -3720 50215 -3600
rect 50335 -3720 50380 -3600
rect 50500 -3720 50545 -3600
rect 50665 -3720 50720 -3600
rect 50840 -3720 50885 -3600
rect 51005 -3720 51050 -3600
rect 51170 -3720 51215 -3600
rect 51335 -3720 51390 -3600
rect 51510 -3720 51555 -3600
rect 51675 -3720 51720 -3600
rect 51840 -3720 51885 -3600
rect 52005 -3720 52060 -3600
rect 52180 -3720 52225 -3600
rect 52345 -3720 52390 -3600
rect 52510 -3720 52555 -3600
rect 52675 -3720 52730 -3600
rect 52850 -3720 52895 -3600
rect 53015 -3720 53060 -3600
rect 53180 -3720 53225 -3600
rect 53345 -3720 53370 -3600
rect 30770 -3765 53370 -3720
rect 30770 -3885 30795 -3765
rect 30915 -3885 30970 -3765
rect 31090 -3885 31135 -3765
rect 31255 -3885 31300 -3765
rect 31420 -3885 31465 -3765
rect 31585 -3885 31640 -3765
rect 31760 -3885 31805 -3765
rect 31925 -3885 31970 -3765
rect 32090 -3885 32135 -3765
rect 32255 -3885 32310 -3765
rect 32430 -3885 32475 -3765
rect 32595 -3885 32640 -3765
rect 32760 -3885 32805 -3765
rect 32925 -3885 32980 -3765
rect 33100 -3885 33145 -3765
rect 33265 -3885 33310 -3765
rect 33430 -3885 33475 -3765
rect 33595 -3885 33650 -3765
rect 33770 -3885 33815 -3765
rect 33935 -3885 33980 -3765
rect 34100 -3885 34145 -3765
rect 34265 -3885 34320 -3765
rect 34440 -3885 34485 -3765
rect 34605 -3885 34650 -3765
rect 34770 -3885 34815 -3765
rect 34935 -3885 34990 -3765
rect 35110 -3885 35155 -3765
rect 35275 -3885 35320 -3765
rect 35440 -3885 35485 -3765
rect 35605 -3885 35660 -3765
rect 35780 -3885 35825 -3765
rect 35945 -3885 35990 -3765
rect 36110 -3885 36155 -3765
rect 36275 -3885 36485 -3765
rect 36605 -3885 36660 -3765
rect 36780 -3885 36825 -3765
rect 36945 -3885 36990 -3765
rect 37110 -3885 37155 -3765
rect 37275 -3885 37330 -3765
rect 37450 -3885 37495 -3765
rect 37615 -3885 37660 -3765
rect 37780 -3885 37825 -3765
rect 37945 -3885 38000 -3765
rect 38120 -3885 38165 -3765
rect 38285 -3885 38330 -3765
rect 38450 -3885 38495 -3765
rect 38615 -3885 38670 -3765
rect 38790 -3885 38835 -3765
rect 38955 -3885 39000 -3765
rect 39120 -3885 39165 -3765
rect 39285 -3885 39340 -3765
rect 39460 -3885 39505 -3765
rect 39625 -3885 39670 -3765
rect 39790 -3885 39835 -3765
rect 39955 -3885 40010 -3765
rect 40130 -3885 40175 -3765
rect 40295 -3885 40340 -3765
rect 40460 -3885 40505 -3765
rect 40625 -3885 40680 -3765
rect 40800 -3885 40845 -3765
rect 40965 -3885 41010 -3765
rect 41130 -3885 41175 -3765
rect 41295 -3885 41350 -3765
rect 41470 -3885 41515 -3765
rect 41635 -3885 41680 -3765
rect 41800 -3885 41845 -3765
rect 41965 -3885 42175 -3765
rect 42295 -3885 42350 -3765
rect 42470 -3885 42515 -3765
rect 42635 -3885 42680 -3765
rect 42800 -3885 42845 -3765
rect 42965 -3885 43020 -3765
rect 43140 -3885 43185 -3765
rect 43305 -3885 43350 -3765
rect 43470 -3885 43515 -3765
rect 43635 -3885 43690 -3765
rect 43810 -3885 43855 -3765
rect 43975 -3885 44020 -3765
rect 44140 -3885 44185 -3765
rect 44305 -3885 44360 -3765
rect 44480 -3885 44525 -3765
rect 44645 -3885 44690 -3765
rect 44810 -3885 44855 -3765
rect 44975 -3885 45030 -3765
rect 45150 -3885 45195 -3765
rect 45315 -3885 45360 -3765
rect 45480 -3885 45525 -3765
rect 45645 -3885 45700 -3765
rect 45820 -3885 45865 -3765
rect 45985 -3885 46030 -3765
rect 46150 -3885 46195 -3765
rect 46315 -3885 46370 -3765
rect 46490 -3885 46535 -3765
rect 46655 -3885 46700 -3765
rect 46820 -3885 46865 -3765
rect 46985 -3885 47040 -3765
rect 47160 -3885 47205 -3765
rect 47325 -3885 47370 -3765
rect 47490 -3885 47535 -3765
rect 47655 -3885 47865 -3765
rect 47985 -3885 48040 -3765
rect 48160 -3885 48205 -3765
rect 48325 -3885 48370 -3765
rect 48490 -3885 48535 -3765
rect 48655 -3885 48710 -3765
rect 48830 -3885 48875 -3765
rect 48995 -3885 49040 -3765
rect 49160 -3885 49205 -3765
rect 49325 -3885 49380 -3765
rect 49500 -3885 49545 -3765
rect 49665 -3885 49710 -3765
rect 49830 -3885 49875 -3765
rect 49995 -3885 50050 -3765
rect 50170 -3885 50215 -3765
rect 50335 -3885 50380 -3765
rect 50500 -3885 50545 -3765
rect 50665 -3885 50720 -3765
rect 50840 -3885 50885 -3765
rect 51005 -3885 51050 -3765
rect 51170 -3885 51215 -3765
rect 51335 -3885 51390 -3765
rect 51510 -3885 51555 -3765
rect 51675 -3885 51720 -3765
rect 51840 -3885 51885 -3765
rect 52005 -3885 52060 -3765
rect 52180 -3885 52225 -3765
rect 52345 -3885 52390 -3765
rect 52510 -3885 52555 -3765
rect 52675 -3885 52730 -3765
rect 52850 -3885 52895 -3765
rect 53015 -3885 53060 -3765
rect 53180 -3885 53225 -3765
rect 53345 -3885 53370 -3765
rect 30770 -3940 53370 -3885
rect 30770 -4060 30795 -3940
rect 30915 -4060 30970 -3940
rect 31090 -4060 31135 -3940
rect 31255 -4060 31300 -3940
rect 31420 -4060 31465 -3940
rect 31585 -4060 31640 -3940
rect 31760 -4060 31805 -3940
rect 31925 -4060 31970 -3940
rect 32090 -4060 32135 -3940
rect 32255 -4060 32310 -3940
rect 32430 -4060 32475 -3940
rect 32595 -4060 32640 -3940
rect 32760 -4060 32805 -3940
rect 32925 -4060 32980 -3940
rect 33100 -4060 33145 -3940
rect 33265 -4060 33310 -3940
rect 33430 -4060 33475 -3940
rect 33595 -4060 33650 -3940
rect 33770 -4060 33815 -3940
rect 33935 -4060 33980 -3940
rect 34100 -4060 34145 -3940
rect 34265 -4060 34320 -3940
rect 34440 -4060 34485 -3940
rect 34605 -4060 34650 -3940
rect 34770 -4060 34815 -3940
rect 34935 -4060 34990 -3940
rect 35110 -4060 35155 -3940
rect 35275 -4060 35320 -3940
rect 35440 -4060 35485 -3940
rect 35605 -4060 35660 -3940
rect 35780 -4060 35825 -3940
rect 35945 -4060 35990 -3940
rect 36110 -4060 36155 -3940
rect 36275 -4060 36485 -3940
rect 36605 -4060 36660 -3940
rect 36780 -4060 36825 -3940
rect 36945 -4060 36990 -3940
rect 37110 -4060 37155 -3940
rect 37275 -4060 37330 -3940
rect 37450 -4060 37495 -3940
rect 37615 -4060 37660 -3940
rect 37780 -4060 37825 -3940
rect 37945 -4060 38000 -3940
rect 38120 -4060 38165 -3940
rect 38285 -4060 38330 -3940
rect 38450 -4060 38495 -3940
rect 38615 -4060 38670 -3940
rect 38790 -4060 38835 -3940
rect 38955 -4060 39000 -3940
rect 39120 -4060 39165 -3940
rect 39285 -4060 39340 -3940
rect 39460 -4060 39505 -3940
rect 39625 -4060 39670 -3940
rect 39790 -4060 39835 -3940
rect 39955 -4060 40010 -3940
rect 40130 -4060 40175 -3940
rect 40295 -4060 40340 -3940
rect 40460 -4060 40505 -3940
rect 40625 -4060 40680 -3940
rect 40800 -4060 40845 -3940
rect 40965 -4060 41010 -3940
rect 41130 -4060 41175 -3940
rect 41295 -4060 41350 -3940
rect 41470 -4060 41515 -3940
rect 41635 -4060 41680 -3940
rect 41800 -4060 41845 -3940
rect 41965 -4060 42175 -3940
rect 42295 -4060 42350 -3940
rect 42470 -4060 42515 -3940
rect 42635 -4060 42680 -3940
rect 42800 -4060 42845 -3940
rect 42965 -4060 43020 -3940
rect 43140 -4060 43185 -3940
rect 43305 -4060 43350 -3940
rect 43470 -4060 43515 -3940
rect 43635 -4060 43690 -3940
rect 43810 -4060 43855 -3940
rect 43975 -4060 44020 -3940
rect 44140 -4060 44185 -3940
rect 44305 -4060 44360 -3940
rect 44480 -4060 44525 -3940
rect 44645 -4060 44690 -3940
rect 44810 -4060 44855 -3940
rect 44975 -4060 45030 -3940
rect 45150 -4060 45195 -3940
rect 45315 -4060 45360 -3940
rect 45480 -4060 45525 -3940
rect 45645 -4060 45700 -3940
rect 45820 -4060 45865 -3940
rect 45985 -4060 46030 -3940
rect 46150 -4060 46195 -3940
rect 46315 -4060 46370 -3940
rect 46490 -4060 46535 -3940
rect 46655 -4060 46700 -3940
rect 46820 -4060 46865 -3940
rect 46985 -4060 47040 -3940
rect 47160 -4060 47205 -3940
rect 47325 -4060 47370 -3940
rect 47490 -4060 47535 -3940
rect 47655 -4060 47865 -3940
rect 47985 -4060 48040 -3940
rect 48160 -4060 48205 -3940
rect 48325 -4060 48370 -3940
rect 48490 -4060 48535 -3940
rect 48655 -4060 48710 -3940
rect 48830 -4060 48875 -3940
rect 48995 -4060 49040 -3940
rect 49160 -4060 49205 -3940
rect 49325 -4060 49380 -3940
rect 49500 -4060 49545 -3940
rect 49665 -4060 49710 -3940
rect 49830 -4060 49875 -3940
rect 49995 -4060 50050 -3940
rect 50170 -4060 50215 -3940
rect 50335 -4060 50380 -3940
rect 50500 -4060 50545 -3940
rect 50665 -4060 50720 -3940
rect 50840 -4060 50885 -3940
rect 51005 -4060 51050 -3940
rect 51170 -4060 51215 -3940
rect 51335 -4060 51390 -3940
rect 51510 -4060 51555 -3940
rect 51675 -4060 51720 -3940
rect 51840 -4060 51885 -3940
rect 52005 -4060 52060 -3940
rect 52180 -4060 52225 -3940
rect 52345 -4060 52390 -3940
rect 52510 -4060 52555 -3940
rect 52675 -4060 52730 -3940
rect 52850 -4060 52895 -3940
rect 53015 -4060 53060 -3940
rect 53180 -4060 53225 -3940
rect 53345 -4060 53370 -3940
rect 30770 -4270 53370 -4060
rect 30770 -4390 30795 -4270
rect 30915 -4390 30960 -4270
rect 31080 -4390 31125 -4270
rect 31245 -4390 31290 -4270
rect 31410 -4390 31465 -4270
rect 31585 -4390 31630 -4270
rect 31750 -4390 31795 -4270
rect 31915 -4390 31960 -4270
rect 32080 -4390 32135 -4270
rect 32255 -4390 32300 -4270
rect 32420 -4390 32465 -4270
rect 32585 -4390 32630 -4270
rect 32750 -4390 32805 -4270
rect 32925 -4390 32970 -4270
rect 33090 -4390 33135 -4270
rect 33255 -4390 33300 -4270
rect 33420 -4390 33475 -4270
rect 33595 -4390 33640 -4270
rect 33760 -4390 33805 -4270
rect 33925 -4390 33970 -4270
rect 34090 -4390 34145 -4270
rect 34265 -4390 34310 -4270
rect 34430 -4390 34475 -4270
rect 34595 -4390 34640 -4270
rect 34760 -4390 34815 -4270
rect 34935 -4390 34980 -4270
rect 35100 -4390 35145 -4270
rect 35265 -4390 35310 -4270
rect 35430 -4390 35485 -4270
rect 35605 -4390 35650 -4270
rect 35770 -4390 35815 -4270
rect 35935 -4390 35980 -4270
rect 36100 -4390 36155 -4270
rect 36275 -4390 36485 -4270
rect 36605 -4390 36650 -4270
rect 36770 -4390 36815 -4270
rect 36935 -4390 36980 -4270
rect 37100 -4390 37155 -4270
rect 37275 -4390 37320 -4270
rect 37440 -4390 37485 -4270
rect 37605 -4390 37650 -4270
rect 37770 -4390 37825 -4270
rect 37945 -4390 37990 -4270
rect 38110 -4390 38155 -4270
rect 38275 -4390 38320 -4270
rect 38440 -4390 38495 -4270
rect 38615 -4390 38660 -4270
rect 38780 -4390 38825 -4270
rect 38945 -4390 38990 -4270
rect 39110 -4390 39165 -4270
rect 39285 -4390 39330 -4270
rect 39450 -4390 39495 -4270
rect 39615 -4390 39660 -4270
rect 39780 -4390 39835 -4270
rect 39955 -4390 40000 -4270
rect 40120 -4390 40165 -4270
rect 40285 -4390 40330 -4270
rect 40450 -4390 40505 -4270
rect 40625 -4390 40670 -4270
rect 40790 -4390 40835 -4270
rect 40955 -4390 41000 -4270
rect 41120 -4390 41175 -4270
rect 41295 -4390 41340 -4270
rect 41460 -4390 41505 -4270
rect 41625 -4390 41670 -4270
rect 41790 -4390 41845 -4270
rect 41965 -4390 42175 -4270
rect 42295 -4390 42340 -4270
rect 42460 -4390 42505 -4270
rect 42625 -4390 42670 -4270
rect 42790 -4390 42845 -4270
rect 42965 -4390 43010 -4270
rect 43130 -4390 43175 -4270
rect 43295 -4390 43340 -4270
rect 43460 -4390 43515 -4270
rect 43635 -4390 43680 -4270
rect 43800 -4390 43845 -4270
rect 43965 -4390 44010 -4270
rect 44130 -4390 44185 -4270
rect 44305 -4390 44350 -4270
rect 44470 -4390 44515 -4270
rect 44635 -4390 44680 -4270
rect 44800 -4390 44855 -4270
rect 44975 -4390 45020 -4270
rect 45140 -4390 45185 -4270
rect 45305 -4390 45350 -4270
rect 45470 -4390 45525 -4270
rect 45645 -4390 45690 -4270
rect 45810 -4390 45855 -4270
rect 45975 -4390 46020 -4270
rect 46140 -4390 46195 -4270
rect 46315 -4390 46360 -4270
rect 46480 -4390 46525 -4270
rect 46645 -4390 46690 -4270
rect 46810 -4390 46865 -4270
rect 46985 -4390 47030 -4270
rect 47150 -4390 47195 -4270
rect 47315 -4390 47360 -4270
rect 47480 -4390 47535 -4270
rect 47655 -4390 47865 -4270
rect 47985 -4390 48030 -4270
rect 48150 -4390 48195 -4270
rect 48315 -4390 48360 -4270
rect 48480 -4390 48535 -4270
rect 48655 -4390 48700 -4270
rect 48820 -4390 48865 -4270
rect 48985 -4390 49030 -4270
rect 49150 -4390 49205 -4270
rect 49325 -4390 49370 -4270
rect 49490 -4390 49535 -4270
rect 49655 -4390 49700 -4270
rect 49820 -4390 49875 -4270
rect 49995 -4390 50040 -4270
rect 50160 -4390 50205 -4270
rect 50325 -4390 50370 -4270
rect 50490 -4390 50545 -4270
rect 50665 -4390 50710 -4270
rect 50830 -4390 50875 -4270
rect 50995 -4390 51040 -4270
rect 51160 -4390 51215 -4270
rect 51335 -4390 51380 -4270
rect 51500 -4390 51545 -4270
rect 51665 -4390 51710 -4270
rect 51830 -4390 51885 -4270
rect 52005 -4390 52050 -4270
rect 52170 -4390 52215 -4270
rect 52335 -4390 52380 -4270
rect 52500 -4390 52555 -4270
rect 52675 -4390 52720 -4270
rect 52840 -4390 52885 -4270
rect 53005 -4390 53050 -4270
rect 53170 -4390 53225 -4270
rect 53345 -4390 53370 -4270
rect 30770 -4445 53370 -4390
rect 30770 -4565 30795 -4445
rect 30915 -4565 30960 -4445
rect 31080 -4565 31125 -4445
rect 31245 -4565 31290 -4445
rect 31410 -4565 31465 -4445
rect 31585 -4565 31630 -4445
rect 31750 -4565 31795 -4445
rect 31915 -4565 31960 -4445
rect 32080 -4565 32135 -4445
rect 32255 -4565 32300 -4445
rect 32420 -4565 32465 -4445
rect 32585 -4565 32630 -4445
rect 32750 -4565 32805 -4445
rect 32925 -4565 32970 -4445
rect 33090 -4565 33135 -4445
rect 33255 -4565 33300 -4445
rect 33420 -4565 33475 -4445
rect 33595 -4565 33640 -4445
rect 33760 -4565 33805 -4445
rect 33925 -4565 33970 -4445
rect 34090 -4565 34145 -4445
rect 34265 -4565 34310 -4445
rect 34430 -4565 34475 -4445
rect 34595 -4565 34640 -4445
rect 34760 -4565 34815 -4445
rect 34935 -4565 34980 -4445
rect 35100 -4565 35145 -4445
rect 35265 -4565 35310 -4445
rect 35430 -4565 35485 -4445
rect 35605 -4565 35650 -4445
rect 35770 -4565 35815 -4445
rect 35935 -4565 35980 -4445
rect 36100 -4565 36155 -4445
rect 36275 -4565 36485 -4445
rect 36605 -4565 36650 -4445
rect 36770 -4565 36815 -4445
rect 36935 -4565 36980 -4445
rect 37100 -4565 37155 -4445
rect 37275 -4565 37320 -4445
rect 37440 -4565 37485 -4445
rect 37605 -4565 37650 -4445
rect 37770 -4565 37825 -4445
rect 37945 -4565 37990 -4445
rect 38110 -4565 38155 -4445
rect 38275 -4565 38320 -4445
rect 38440 -4565 38495 -4445
rect 38615 -4565 38660 -4445
rect 38780 -4565 38825 -4445
rect 38945 -4565 38990 -4445
rect 39110 -4565 39165 -4445
rect 39285 -4565 39330 -4445
rect 39450 -4565 39495 -4445
rect 39615 -4565 39660 -4445
rect 39780 -4565 39835 -4445
rect 39955 -4565 40000 -4445
rect 40120 -4565 40165 -4445
rect 40285 -4565 40330 -4445
rect 40450 -4565 40505 -4445
rect 40625 -4565 40670 -4445
rect 40790 -4565 40835 -4445
rect 40955 -4565 41000 -4445
rect 41120 -4565 41175 -4445
rect 41295 -4565 41340 -4445
rect 41460 -4565 41505 -4445
rect 41625 -4565 41670 -4445
rect 41790 -4565 41845 -4445
rect 41965 -4565 42175 -4445
rect 42295 -4565 42340 -4445
rect 42460 -4565 42505 -4445
rect 42625 -4565 42670 -4445
rect 42790 -4565 42845 -4445
rect 42965 -4565 43010 -4445
rect 43130 -4565 43175 -4445
rect 43295 -4565 43340 -4445
rect 43460 -4565 43515 -4445
rect 43635 -4565 43680 -4445
rect 43800 -4565 43845 -4445
rect 43965 -4565 44010 -4445
rect 44130 -4565 44185 -4445
rect 44305 -4565 44350 -4445
rect 44470 -4565 44515 -4445
rect 44635 -4565 44680 -4445
rect 44800 -4565 44855 -4445
rect 44975 -4565 45020 -4445
rect 45140 -4565 45185 -4445
rect 45305 -4565 45350 -4445
rect 45470 -4565 45525 -4445
rect 45645 -4565 45690 -4445
rect 45810 -4565 45855 -4445
rect 45975 -4565 46020 -4445
rect 46140 -4565 46195 -4445
rect 46315 -4565 46360 -4445
rect 46480 -4565 46525 -4445
rect 46645 -4565 46690 -4445
rect 46810 -4565 46865 -4445
rect 46985 -4565 47030 -4445
rect 47150 -4565 47195 -4445
rect 47315 -4565 47360 -4445
rect 47480 -4565 47535 -4445
rect 47655 -4565 47865 -4445
rect 47985 -4565 48030 -4445
rect 48150 -4565 48195 -4445
rect 48315 -4565 48360 -4445
rect 48480 -4565 48535 -4445
rect 48655 -4565 48700 -4445
rect 48820 -4565 48865 -4445
rect 48985 -4565 49030 -4445
rect 49150 -4565 49205 -4445
rect 49325 -4565 49370 -4445
rect 49490 -4565 49535 -4445
rect 49655 -4565 49700 -4445
rect 49820 -4565 49875 -4445
rect 49995 -4565 50040 -4445
rect 50160 -4565 50205 -4445
rect 50325 -4565 50370 -4445
rect 50490 -4565 50545 -4445
rect 50665 -4565 50710 -4445
rect 50830 -4565 50875 -4445
rect 50995 -4565 51040 -4445
rect 51160 -4565 51215 -4445
rect 51335 -4565 51380 -4445
rect 51500 -4565 51545 -4445
rect 51665 -4565 51710 -4445
rect 51830 -4565 51885 -4445
rect 52005 -4565 52050 -4445
rect 52170 -4565 52215 -4445
rect 52335 -4565 52380 -4445
rect 52500 -4565 52555 -4445
rect 52675 -4565 52720 -4445
rect 52840 -4565 52885 -4445
rect 53005 -4565 53050 -4445
rect 53170 -4565 53225 -4445
rect 53345 -4565 53370 -4445
rect 30770 -4610 53370 -4565
rect 30770 -4730 30795 -4610
rect 30915 -4730 30960 -4610
rect 31080 -4730 31125 -4610
rect 31245 -4730 31290 -4610
rect 31410 -4730 31465 -4610
rect 31585 -4730 31630 -4610
rect 31750 -4730 31795 -4610
rect 31915 -4730 31960 -4610
rect 32080 -4730 32135 -4610
rect 32255 -4730 32300 -4610
rect 32420 -4730 32465 -4610
rect 32585 -4730 32630 -4610
rect 32750 -4730 32805 -4610
rect 32925 -4730 32970 -4610
rect 33090 -4730 33135 -4610
rect 33255 -4730 33300 -4610
rect 33420 -4730 33475 -4610
rect 33595 -4730 33640 -4610
rect 33760 -4730 33805 -4610
rect 33925 -4730 33970 -4610
rect 34090 -4730 34145 -4610
rect 34265 -4730 34310 -4610
rect 34430 -4730 34475 -4610
rect 34595 -4730 34640 -4610
rect 34760 -4730 34815 -4610
rect 34935 -4730 34980 -4610
rect 35100 -4730 35145 -4610
rect 35265 -4730 35310 -4610
rect 35430 -4730 35485 -4610
rect 35605 -4730 35650 -4610
rect 35770 -4730 35815 -4610
rect 35935 -4730 35980 -4610
rect 36100 -4730 36155 -4610
rect 36275 -4730 36485 -4610
rect 36605 -4730 36650 -4610
rect 36770 -4730 36815 -4610
rect 36935 -4730 36980 -4610
rect 37100 -4730 37155 -4610
rect 37275 -4730 37320 -4610
rect 37440 -4730 37485 -4610
rect 37605 -4730 37650 -4610
rect 37770 -4730 37825 -4610
rect 37945 -4730 37990 -4610
rect 38110 -4730 38155 -4610
rect 38275 -4730 38320 -4610
rect 38440 -4730 38495 -4610
rect 38615 -4730 38660 -4610
rect 38780 -4730 38825 -4610
rect 38945 -4730 38990 -4610
rect 39110 -4730 39165 -4610
rect 39285 -4730 39330 -4610
rect 39450 -4730 39495 -4610
rect 39615 -4730 39660 -4610
rect 39780 -4730 39835 -4610
rect 39955 -4730 40000 -4610
rect 40120 -4730 40165 -4610
rect 40285 -4730 40330 -4610
rect 40450 -4730 40505 -4610
rect 40625 -4730 40670 -4610
rect 40790 -4730 40835 -4610
rect 40955 -4730 41000 -4610
rect 41120 -4730 41175 -4610
rect 41295 -4730 41340 -4610
rect 41460 -4730 41505 -4610
rect 41625 -4730 41670 -4610
rect 41790 -4730 41845 -4610
rect 41965 -4730 42175 -4610
rect 42295 -4730 42340 -4610
rect 42460 -4730 42505 -4610
rect 42625 -4730 42670 -4610
rect 42790 -4730 42845 -4610
rect 42965 -4730 43010 -4610
rect 43130 -4730 43175 -4610
rect 43295 -4730 43340 -4610
rect 43460 -4730 43515 -4610
rect 43635 -4730 43680 -4610
rect 43800 -4730 43845 -4610
rect 43965 -4730 44010 -4610
rect 44130 -4730 44185 -4610
rect 44305 -4730 44350 -4610
rect 44470 -4730 44515 -4610
rect 44635 -4730 44680 -4610
rect 44800 -4730 44855 -4610
rect 44975 -4730 45020 -4610
rect 45140 -4730 45185 -4610
rect 45305 -4730 45350 -4610
rect 45470 -4730 45525 -4610
rect 45645 -4730 45690 -4610
rect 45810 -4730 45855 -4610
rect 45975 -4730 46020 -4610
rect 46140 -4730 46195 -4610
rect 46315 -4730 46360 -4610
rect 46480 -4730 46525 -4610
rect 46645 -4730 46690 -4610
rect 46810 -4730 46865 -4610
rect 46985 -4730 47030 -4610
rect 47150 -4730 47195 -4610
rect 47315 -4730 47360 -4610
rect 47480 -4730 47535 -4610
rect 47655 -4730 47865 -4610
rect 47985 -4730 48030 -4610
rect 48150 -4730 48195 -4610
rect 48315 -4730 48360 -4610
rect 48480 -4730 48535 -4610
rect 48655 -4730 48700 -4610
rect 48820 -4730 48865 -4610
rect 48985 -4730 49030 -4610
rect 49150 -4730 49205 -4610
rect 49325 -4730 49370 -4610
rect 49490 -4730 49535 -4610
rect 49655 -4730 49700 -4610
rect 49820 -4730 49875 -4610
rect 49995 -4730 50040 -4610
rect 50160 -4730 50205 -4610
rect 50325 -4730 50370 -4610
rect 50490 -4730 50545 -4610
rect 50665 -4730 50710 -4610
rect 50830 -4730 50875 -4610
rect 50995 -4730 51040 -4610
rect 51160 -4730 51215 -4610
rect 51335 -4730 51380 -4610
rect 51500 -4730 51545 -4610
rect 51665 -4730 51710 -4610
rect 51830 -4730 51885 -4610
rect 52005 -4730 52050 -4610
rect 52170 -4730 52215 -4610
rect 52335 -4730 52380 -4610
rect 52500 -4730 52555 -4610
rect 52675 -4730 52720 -4610
rect 52840 -4730 52885 -4610
rect 53005 -4730 53050 -4610
rect 53170 -4730 53225 -4610
rect 53345 -4730 53370 -4610
rect 30770 -4775 53370 -4730
rect 30770 -4895 30795 -4775
rect 30915 -4895 30960 -4775
rect 31080 -4895 31125 -4775
rect 31245 -4895 31290 -4775
rect 31410 -4895 31465 -4775
rect 31585 -4895 31630 -4775
rect 31750 -4895 31795 -4775
rect 31915 -4895 31960 -4775
rect 32080 -4895 32135 -4775
rect 32255 -4895 32300 -4775
rect 32420 -4895 32465 -4775
rect 32585 -4895 32630 -4775
rect 32750 -4895 32805 -4775
rect 32925 -4895 32970 -4775
rect 33090 -4895 33135 -4775
rect 33255 -4895 33300 -4775
rect 33420 -4895 33475 -4775
rect 33595 -4895 33640 -4775
rect 33760 -4895 33805 -4775
rect 33925 -4895 33970 -4775
rect 34090 -4895 34145 -4775
rect 34265 -4895 34310 -4775
rect 34430 -4895 34475 -4775
rect 34595 -4895 34640 -4775
rect 34760 -4895 34815 -4775
rect 34935 -4895 34980 -4775
rect 35100 -4895 35145 -4775
rect 35265 -4895 35310 -4775
rect 35430 -4895 35485 -4775
rect 35605 -4895 35650 -4775
rect 35770 -4895 35815 -4775
rect 35935 -4895 35980 -4775
rect 36100 -4895 36155 -4775
rect 36275 -4895 36485 -4775
rect 36605 -4895 36650 -4775
rect 36770 -4895 36815 -4775
rect 36935 -4895 36980 -4775
rect 37100 -4895 37155 -4775
rect 37275 -4895 37320 -4775
rect 37440 -4895 37485 -4775
rect 37605 -4895 37650 -4775
rect 37770 -4895 37825 -4775
rect 37945 -4895 37990 -4775
rect 38110 -4895 38155 -4775
rect 38275 -4895 38320 -4775
rect 38440 -4895 38495 -4775
rect 38615 -4895 38660 -4775
rect 38780 -4895 38825 -4775
rect 38945 -4895 38990 -4775
rect 39110 -4895 39165 -4775
rect 39285 -4895 39330 -4775
rect 39450 -4895 39495 -4775
rect 39615 -4895 39660 -4775
rect 39780 -4895 39835 -4775
rect 39955 -4895 40000 -4775
rect 40120 -4895 40165 -4775
rect 40285 -4895 40330 -4775
rect 40450 -4895 40505 -4775
rect 40625 -4895 40670 -4775
rect 40790 -4895 40835 -4775
rect 40955 -4895 41000 -4775
rect 41120 -4895 41175 -4775
rect 41295 -4895 41340 -4775
rect 41460 -4895 41505 -4775
rect 41625 -4895 41670 -4775
rect 41790 -4895 41845 -4775
rect 41965 -4895 42175 -4775
rect 42295 -4895 42340 -4775
rect 42460 -4895 42505 -4775
rect 42625 -4895 42670 -4775
rect 42790 -4895 42845 -4775
rect 42965 -4895 43010 -4775
rect 43130 -4895 43175 -4775
rect 43295 -4895 43340 -4775
rect 43460 -4895 43515 -4775
rect 43635 -4895 43680 -4775
rect 43800 -4895 43845 -4775
rect 43965 -4895 44010 -4775
rect 44130 -4895 44185 -4775
rect 44305 -4895 44350 -4775
rect 44470 -4895 44515 -4775
rect 44635 -4895 44680 -4775
rect 44800 -4895 44855 -4775
rect 44975 -4895 45020 -4775
rect 45140 -4895 45185 -4775
rect 45305 -4895 45350 -4775
rect 45470 -4895 45525 -4775
rect 45645 -4895 45690 -4775
rect 45810 -4895 45855 -4775
rect 45975 -4895 46020 -4775
rect 46140 -4895 46195 -4775
rect 46315 -4895 46360 -4775
rect 46480 -4895 46525 -4775
rect 46645 -4895 46690 -4775
rect 46810 -4895 46865 -4775
rect 46985 -4895 47030 -4775
rect 47150 -4895 47195 -4775
rect 47315 -4895 47360 -4775
rect 47480 -4895 47535 -4775
rect 47655 -4895 47865 -4775
rect 47985 -4895 48030 -4775
rect 48150 -4895 48195 -4775
rect 48315 -4895 48360 -4775
rect 48480 -4895 48535 -4775
rect 48655 -4895 48700 -4775
rect 48820 -4895 48865 -4775
rect 48985 -4895 49030 -4775
rect 49150 -4895 49205 -4775
rect 49325 -4895 49370 -4775
rect 49490 -4895 49535 -4775
rect 49655 -4895 49700 -4775
rect 49820 -4895 49875 -4775
rect 49995 -4895 50040 -4775
rect 50160 -4895 50205 -4775
rect 50325 -4895 50370 -4775
rect 50490 -4895 50545 -4775
rect 50665 -4895 50710 -4775
rect 50830 -4895 50875 -4775
rect 50995 -4895 51040 -4775
rect 51160 -4895 51215 -4775
rect 51335 -4895 51380 -4775
rect 51500 -4895 51545 -4775
rect 51665 -4895 51710 -4775
rect 51830 -4895 51885 -4775
rect 52005 -4895 52050 -4775
rect 52170 -4895 52215 -4775
rect 52335 -4895 52380 -4775
rect 52500 -4895 52555 -4775
rect 52675 -4895 52720 -4775
rect 52840 -4895 52885 -4775
rect 53005 -4895 53050 -4775
rect 53170 -4895 53225 -4775
rect 53345 -4895 53370 -4775
rect 30770 -4940 53370 -4895
rect 30770 -5060 30795 -4940
rect 30915 -5060 30960 -4940
rect 31080 -5060 31125 -4940
rect 31245 -5060 31290 -4940
rect 31410 -5060 31465 -4940
rect 31585 -5060 31630 -4940
rect 31750 -5060 31795 -4940
rect 31915 -5060 31960 -4940
rect 32080 -5060 32135 -4940
rect 32255 -5060 32300 -4940
rect 32420 -5060 32465 -4940
rect 32585 -5060 32630 -4940
rect 32750 -5060 32805 -4940
rect 32925 -5060 32970 -4940
rect 33090 -5060 33135 -4940
rect 33255 -5060 33300 -4940
rect 33420 -5060 33475 -4940
rect 33595 -5060 33640 -4940
rect 33760 -5060 33805 -4940
rect 33925 -5060 33970 -4940
rect 34090 -5060 34145 -4940
rect 34265 -5060 34310 -4940
rect 34430 -5060 34475 -4940
rect 34595 -5060 34640 -4940
rect 34760 -5060 34815 -4940
rect 34935 -5060 34980 -4940
rect 35100 -5060 35145 -4940
rect 35265 -5060 35310 -4940
rect 35430 -5060 35485 -4940
rect 35605 -5060 35650 -4940
rect 35770 -5060 35815 -4940
rect 35935 -5060 35980 -4940
rect 36100 -5060 36155 -4940
rect 36275 -5060 36485 -4940
rect 36605 -5060 36650 -4940
rect 36770 -5060 36815 -4940
rect 36935 -5060 36980 -4940
rect 37100 -5060 37155 -4940
rect 37275 -5060 37320 -4940
rect 37440 -5060 37485 -4940
rect 37605 -5060 37650 -4940
rect 37770 -5060 37825 -4940
rect 37945 -5060 37990 -4940
rect 38110 -5060 38155 -4940
rect 38275 -5060 38320 -4940
rect 38440 -5060 38495 -4940
rect 38615 -5060 38660 -4940
rect 38780 -5060 38825 -4940
rect 38945 -5060 38990 -4940
rect 39110 -5060 39165 -4940
rect 39285 -5060 39330 -4940
rect 39450 -5060 39495 -4940
rect 39615 -5060 39660 -4940
rect 39780 -5060 39835 -4940
rect 39955 -5060 40000 -4940
rect 40120 -5060 40165 -4940
rect 40285 -5060 40330 -4940
rect 40450 -5060 40505 -4940
rect 40625 -5060 40670 -4940
rect 40790 -5060 40835 -4940
rect 40955 -5060 41000 -4940
rect 41120 -5060 41175 -4940
rect 41295 -5060 41340 -4940
rect 41460 -5060 41505 -4940
rect 41625 -5060 41670 -4940
rect 41790 -5060 41845 -4940
rect 41965 -5060 42175 -4940
rect 42295 -5060 42340 -4940
rect 42460 -5060 42505 -4940
rect 42625 -5060 42670 -4940
rect 42790 -5060 42845 -4940
rect 42965 -5060 43010 -4940
rect 43130 -5060 43175 -4940
rect 43295 -5060 43340 -4940
rect 43460 -5060 43515 -4940
rect 43635 -5060 43680 -4940
rect 43800 -5060 43845 -4940
rect 43965 -5060 44010 -4940
rect 44130 -5060 44185 -4940
rect 44305 -5060 44350 -4940
rect 44470 -5060 44515 -4940
rect 44635 -5060 44680 -4940
rect 44800 -5060 44855 -4940
rect 44975 -5060 45020 -4940
rect 45140 -5060 45185 -4940
rect 45305 -5060 45350 -4940
rect 45470 -5060 45525 -4940
rect 45645 -5060 45690 -4940
rect 45810 -5060 45855 -4940
rect 45975 -5060 46020 -4940
rect 46140 -5060 46195 -4940
rect 46315 -5060 46360 -4940
rect 46480 -5060 46525 -4940
rect 46645 -5060 46690 -4940
rect 46810 -5060 46865 -4940
rect 46985 -5060 47030 -4940
rect 47150 -5060 47195 -4940
rect 47315 -5060 47360 -4940
rect 47480 -5060 47535 -4940
rect 47655 -5060 47865 -4940
rect 47985 -5060 48030 -4940
rect 48150 -5060 48195 -4940
rect 48315 -5060 48360 -4940
rect 48480 -5060 48535 -4940
rect 48655 -5060 48700 -4940
rect 48820 -5060 48865 -4940
rect 48985 -5060 49030 -4940
rect 49150 -5060 49205 -4940
rect 49325 -5060 49370 -4940
rect 49490 -5060 49535 -4940
rect 49655 -5060 49700 -4940
rect 49820 -5060 49875 -4940
rect 49995 -5060 50040 -4940
rect 50160 -5060 50205 -4940
rect 50325 -5060 50370 -4940
rect 50490 -5060 50545 -4940
rect 50665 -5060 50710 -4940
rect 50830 -5060 50875 -4940
rect 50995 -5060 51040 -4940
rect 51160 -5060 51215 -4940
rect 51335 -5060 51380 -4940
rect 51500 -5060 51545 -4940
rect 51665 -5060 51710 -4940
rect 51830 -5060 51885 -4940
rect 52005 -5060 52050 -4940
rect 52170 -5060 52215 -4940
rect 52335 -5060 52380 -4940
rect 52500 -5060 52555 -4940
rect 52675 -5060 52720 -4940
rect 52840 -5060 52885 -4940
rect 53005 -5060 53050 -4940
rect 53170 -5060 53225 -4940
rect 53345 -5060 53370 -4940
rect 30770 -5115 53370 -5060
rect 30770 -5235 30795 -5115
rect 30915 -5235 30960 -5115
rect 31080 -5235 31125 -5115
rect 31245 -5235 31290 -5115
rect 31410 -5235 31465 -5115
rect 31585 -5235 31630 -5115
rect 31750 -5235 31795 -5115
rect 31915 -5235 31960 -5115
rect 32080 -5235 32135 -5115
rect 32255 -5235 32300 -5115
rect 32420 -5235 32465 -5115
rect 32585 -5235 32630 -5115
rect 32750 -5235 32805 -5115
rect 32925 -5235 32970 -5115
rect 33090 -5235 33135 -5115
rect 33255 -5235 33300 -5115
rect 33420 -5235 33475 -5115
rect 33595 -5235 33640 -5115
rect 33760 -5235 33805 -5115
rect 33925 -5235 33970 -5115
rect 34090 -5235 34145 -5115
rect 34265 -5235 34310 -5115
rect 34430 -5235 34475 -5115
rect 34595 -5235 34640 -5115
rect 34760 -5235 34815 -5115
rect 34935 -5235 34980 -5115
rect 35100 -5235 35145 -5115
rect 35265 -5235 35310 -5115
rect 35430 -5235 35485 -5115
rect 35605 -5235 35650 -5115
rect 35770 -5235 35815 -5115
rect 35935 -5235 35980 -5115
rect 36100 -5235 36155 -5115
rect 36275 -5235 36485 -5115
rect 36605 -5235 36650 -5115
rect 36770 -5235 36815 -5115
rect 36935 -5235 36980 -5115
rect 37100 -5235 37155 -5115
rect 37275 -5235 37320 -5115
rect 37440 -5235 37485 -5115
rect 37605 -5235 37650 -5115
rect 37770 -5235 37825 -5115
rect 37945 -5235 37990 -5115
rect 38110 -5235 38155 -5115
rect 38275 -5235 38320 -5115
rect 38440 -5235 38495 -5115
rect 38615 -5235 38660 -5115
rect 38780 -5235 38825 -5115
rect 38945 -5235 38990 -5115
rect 39110 -5235 39165 -5115
rect 39285 -5235 39330 -5115
rect 39450 -5235 39495 -5115
rect 39615 -5235 39660 -5115
rect 39780 -5235 39835 -5115
rect 39955 -5235 40000 -5115
rect 40120 -5235 40165 -5115
rect 40285 -5235 40330 -5115
rect 40450 -5235 40505 -5115
rect 40625 -5235 40670 -5115
rect 40790 -5235 40835 -5115
rect 40955 -5235 41000 -5115
rect 41120 -5235 41175 -5115
rect 41295 -5235 41340 -5115
rect 41460 -5235 41505 -5115
rect 41625 -5235 41670 -5115
rect 41790 -5235 41845 -5115
rect 41965 -5235 42175 -5115
rect 42295 -5235 42340 -5115
rect 42460 -5235 42505 -5115
rect 42625 -5235 42670 -5115
rect 42790 -5235 42845 -5115
rect 42965 -5235 43010 -5115
rect 43130 -5235 43175 -5115
rect 43295 -5235 43340 -5115
rect 43460 -5235 43515 -5115
rect 43635 -5235 43680 -5115
rect 43800 -5235 43845 -5115
rect 43965 -5235 44010 -5115
rect 44130 -5235 44185 -5115
rect 44305 -5235 44350 -5115
rect 44470 -5235 44515 -5115
rect 44635 -5235 44680 -5115
rect 44800 -5235 44855 -5115
rect 44975 -5235 45020 -5115
rect 45140 -5235 45185 -5115
rect 45305 -5235 45350 -5115
rect 45470 -5235 45525 -5115
rect 45645 -5235 45690 -5115
rect 45810 -5235 45855 -5115
rect 45975 -5235 46020 -5115
rect 46140 -5235 46195 -5115
rect 46315 -5235 46360 -5115
rect 46480 -5235 46525 -5115
rect 46645 -5235 46690 -5115
rect 46810 -5235 46865 -5115
rect 46985 -5235 47030 -5115
rect 47150 -5235 47195 -5115
rect 47315 -5235 47360 -5115
rect 47480 -5235 47535 -5115
rect 47655 -5235 47865 -5115
rect 47985 -5235 48030 -5115
rect 48150 -5235 48195 -5115
rect 48315 -5235 48360 -5115
rect 48480 -5235 48535 -5115
rect 48655 -5235 48700 -5115
rect 48820 -5235 48865 -5115
rect 48985 -5235 49030 -5115
rect 49150 -5235 49205 -5115
rect 49325 -5235 49370 -5115
rect 49490 -5235 49535 -5115
rect 49655 -5235 49700 -5115
rect 49820 -5235 49875 -5115
rect 49995 -5235 50040 -5115
rect 50160 -5235 50205 -5115
rect 50325 -5235 50370 -5115
rect 50490 -5235 50545 -5115
rect 50665 -5235 50710 -5115
rect 50830 -5235 50875 -5115
rect 50995 -5235 51040 -5115
rect 51160 -5235 51215 -5115
rect 51335 -5235 51380 -5115
rect 51500 -5235 51545 -5115
rect 51665 -5235 51710 -5115
rect 51830 -5235 51885 -5115
rect 52005 -5235 52050 -5115
rect 52170 -5235 52215 -5115
rect 52335 -5235 52380 -5115
rect 52500 -5235 52555 -5115
rect 52675 -5235 52720 -5115
rect 52840 -5235 52885 -5115
rect 53005 -5235 53050 -5115
rect 53170 -5235 53225 -5115
rect 53345 -5235 53370 -5115
rect 30770 -5280 53370 -5235
rect 30770 -5400 30795 -5280
rect 30915 -5400 30960 -5280
rect 31080 -5400 31125 -5280
rect 31245 -5400 31290 -5280
rect 31410 -5400 31465 -5280
rect 31585 -5400 31630 -5280
rect 31750 -5400 31795 -5280
rect 31915 -5400 31960 -5280
rect 32080 -5400 32135 -5280
rect 32255 -5400 32300 -5280
rect 32420 -5400 32465 -5280
rect 32585 -5400 32630 -5280
rect 32750 -5400 32805 -5280
rect 32925 -5400 32970 -5280
rect 33090 -5400 33135 -5280
rect 33255 -5400 33300 -5280
rect 33420 -5400 33475 -5280
rect 33595 -5400 33640 -5280
rect 33760 -5400 33805 -5280
rect 33925 -5400 33970 -5280
rect 34090 -5400 34145 -5280
rect 34265 -5400 34310 -5280
rect 34430 -5400 34475 -5280
rect 34595 -5400 34640 -5280
rect 34760 -5400 34815 -5280
rect 34935 -5400 34980 -5280
rect 35100 -5400 35145 -5280
rect 35265 -5400 35310 -5280
rect 35430 -5400 35485 -5280
rect 35605 -5400 35650 -5280
rect 35770 -5400 35815 -5280
rect 35935 -5400 35980 -5280
rect 36100 -5400 36155 -5280
rect 36275 -5400 36485 -5280
rect 36605 -5400 36650 -5280
rect 36770 -5400 36815 -5280
rect 36935 -5400 36980 -5280
rect 37100 -5400 37155 -5280
rect 37275 -5400 37320 -5280
rect 37440 -5400 37485 -5280
rect 37605 -5400 37650 -5280
rect 37770 -5400 37825 -5280
rect 37945 -5400 37990 -5280
rect 38110 -5400 38155 -5280
rect 38275 -5400 38320 -5280
rect 38440 -5400 38495 -5280
rect 38615 -5400 38660 -5280
rect 38780 -5400 38825 -5280
rect 38945 -5400 38990 -5280
rect 39110 -5400 39165 -5280
rect 39285 -5400 39330 -5280
rect 39450 -5400 39495 -5280
rect 39615 -5400 39660 -5280
rect 39780 -5400 39835 -5280
rect 39955 -5400 40000 -5280
rect 40120 -5400 40165 -5280
rect 40285 -5400 40330 -5280
rect 40450 -5400 40505 -5280
rect 40625 -5400 40670 -5280
rect 40790 -5400 40835 -5280
rect 40955 -5400 41000 -5280
rect 41120 -5400 41175 -5280
rect 41295 -5400 41340 -5280
rect 41460 -5400 41505 -5280
rect 41625 -5400 41670 -5280
rect 41790 -5400 41845 -5280
rect 41965 -5400 42175 -5280
rect 42295 -5400 42340 -5280
rect 42460 -5400 42505 -5280
rect 42625 -5400 42670 -5280
rect 42790 -5400 42845 -5280
rect 42965 -5400 43010 -5280
rect 43130 -5400 43175 -5280
rect 43295 -5400 43340 -5280
rect 43460 -5400 43515 -5280
rect 43635 -5400 43680 -5280
rect 43800 -5400 43845 -5280
rect 43965 -5400 44010 -5280
rect 44130 -5400 44185 -5280
rect 44305 -5400 44350 -5280
rect 44470 -5400 44515 -5280
rect 44635 -5400 44680 -5280
rect 44800 -5400 44855 -5280
rect 44975 -5400 45020 -5280
rect 45140 -5400 45185 -5280
rect 45305 -5400 45350 -5280
rect 45470 -5400 45525 -5280
rect 45645 -5400 45690 -5280
rect 45810 -5400 45855 -5280
rect 45975 -5400 46020 -5280
rect 46140 -5400 46195 -5280
rect 46315 -5400 46360 -5280
rect 46480 -5400 46525 -5280
rect 46645 -5400 46690 -5280
rect 46810 -5400 46865 -5280
rect 46985 -5400 47030 -5280
rect 47150 -5400 47195 -5280
rect 47315 -5400 47360 -5280
rect 47480 -5400 47535 -5280
rect 47655 -5400 47865 -5280
rect 47985 -5400 48030 -5280
rect 48150 -5400 48195 -5280
rect 48315 -5400 48360 -5280
rect 48480 -5400 48535 -5280
rect 48655 -5400 48700 -5280
rect 48820 -5400 48865 -5280
rect 48985 -5400 49030 -5280
rect 49150 -5400 49205 -5280
rect 49325 -5400 49370 -5280
rect 49490 -5400 49535 -5280
rect 49655 -5400 49700 -5280
rect 49820 -5400 49875 -5280
rect 49995 -5400 50040 -5280
rect 50160 -5400 50205 -5280
rect 50325 -5400 50370 -5280
rect 50490 -5400 50545 -5280
rect 50665 -5400 50710 -5280
rect 50830 -5400 50875 -5280
rect 50995 -5400 51040 -5280
rect 51160 -5400 51215 -5280
rect 51335 -5400 51380 -5280
rect 51500 -5400 51545 -5280
rect 51665 -5400 51710 -5280
rect 51830 -5400 51885 -5280
rect 52005 -5400 52050 -5280
rect 52170 -5400 52215 -5280
rect 52335 -5400 52380 -5280
rect 52500 -5400 52555 -5280
rect 52675 -5400 52720 -5280
rect 52840 -5400 52885 -5280
rect 53005 -5400 53050 -5280
rect 53170 -5400 53225 -5280
rect 53345 -5400 53370 -5280
rect 30770 -5445 53370 -5400
rect 30770 -5565 30795 -5445
rect 30915 -5565 30960 -5445
rect 31080 -5565 31125 -5445
rect 31245 -5565 31290 -5445
rect 31410 -5565 31465 -5445
rect 31585 -5565 31630 -5445
rect 31750 -5565 31795 -5445
rect 31915 -5565 31960 -5445
rect 32080 -5565 32135 -5445
rect 32255 -5565 32300 -5445
rect 32420 -5565 32465 -5445
rect 32585 -5565 32630 -5445
rect 32750 -5565 32805 -5445
rect 32925 -5565 32970 -5445
rect 33090 -5565 33135 -5445
rect 33255 -5565 33300 -5445
rect 33420 -5565 33475 -5445
rect 33595 -5565 33640 -5445
rect 33760 -5565 33805 -5445
rect 33925 -5565 33970 -5445
rect 34090 -5565 34145 -5445
rect 34265 -5565 34310 -5445
rect 34430 -5565 34475 -5445
rect 34595 -5565 34640 -5445
rect 34760 -5565 34815 -5445
rect 34935 -5565 34980 -5445
rect 35100 -5565 35145 -5445
rect 35265 -5565 35310 -5445
rect 35430 -5565 35485 -5445
rect 35605 -5565 35650 -5445
rect 35770 -5565 35815 -5445
rect 35935 -5565 35980 -5445
rect 36100 -5565 36155 -5445
rect 36275 -5565 36485 -5445
rect 36605 -5565 36650 -5445
rect 36770 -5565 36815 -5445
rect 36935 -5565 36980 -5445
rect 37100 -5565 37155 -5445
rect 37275 -5565 37320 -5445
rect 37440 -5565 37485 -5445
rect 37605 -5565 37650 -5445
rect 37770 -5565 37825 -5445
rect 37945 -5565 37990 -5445
rect 38110 -5565 38155 -5445
rect 38275 -5565 38320 -5445
rect 38440 -5565 38495 -5445
rect 38615 -5565 38660 -5445
rect 38780 -5565 38825 -5445
rect 38945 -5565 38990 -5445
rect 39110 -5565 39165 -5445
rect 39285 -5565 39330 -5445
rect 39450 -5565 39495 -5445
rect 39615 -5565 39660 -5445
rect 39780 -5565 39835 -5445
rect 39955 -5565 40000 -5445
rect 40120 -5565 40165 -5445
rect 40285 -5565 40330 -5445
rect 40450 -5565 40505 -5445
rect 40625 -5565 40670 -5445
rect 40790 -5565 40835 -5445
rect 40955 -5565 41000 -5445
rect 41120 -5565 41175 -5445
rect 41295 -5565 41340 -5445
rect 41460 -5565 41505 -5445
rect 41625 -5565 41670 -5445
rect 41790 -5565 41845 -5445
rect 41965 -5565 42175 -5445
rect 42295 -5565 42340 -5445
rect 42460 -5565 42505 -5445
rect 42625 -5565 42670 -5445
rect 42790 -5565 42845 -5445
rect 42965 -5565 43010 -5445
rect 43130 -5565 43175 -5445
rect 43295 -5565 43340 -5445
rect 43460 -5565 43515 -5445
rect 43635 -5565 43680 -5445
rect 43800 -5565 43845 -5445
rect 43965 -5565 44010 -5445
rect 44130 -5565 44185 -5445
rect 44305 -5565 44350 -5445
rect 44470 -5565 44515 -5445
rect 44635 -5565 44680 -5445
rect 44800 -5565 44855 -5445
rect 44975 -5565 45020 -5445
rect 45140 -5565 45185 -5445
rect 45305 -5565 45350 -5445
rect 45470 -5565 45525 -5445
rect 45645 -5565 45690 -5445
rect 45810 -5565 45855 -5445
rect 45975 -5565 46020 -5445
rect 46140 -5565 46195 -5445
rect 46315 -5565 46360 -5445
rect 46480 -5565 46525 -5445
rect 46645 -5565 46690 -5445
rect 46810 -5565 46865 -5445
rect 46985 -5565 47030 -5445
rect 47150 -5565 47195 -5445
rect 47315 -5565 47360 -5445
rect 47480 -5565 47535 -5445
rect 47655 -5565 47865 -5445
rect 47985 -5565 48030 -5445
rect 48150 -5565 48195 -5445
rect 48315 -5565 48360 -5445
rect 48480 -5565 48535 -5445
rect 48655 -5565 48700 -5445
rect 48820 -5565 48865 -5445
rect 48985 -5565 49030 -5445
rect 49150 -5565 49205 -5445
rect 49325 -5565 49370 -5445
rect 49490 -5565 49535 -5445
rect 49655 -5565 49700 -5445
rect 49820 -5565 49875 -5445
rect 49995 -5565 50040 -5445
rect 50160 -5565 50205 -5445
rect 50325 -5565 50370 -5445
rect 50490 -5565 50545 -5445
rect 50665 -5565 50710 -5445
rect 50830 -5565 50875 -5445
rect 50995 -5565 51040 -5445
rect 51160 -5565 51215 -5445
rect 51335 -5565 51380 -5445
rect 51500 -5565 51545 -5445
rect 51665 -5565 51710 -5445
rect 51830 -5565 51885 -5445
rect 52005 -5565 52050 -5445
rect 52170 -5565 52215 -5445
rect 52335 -5565 52380 -5445
rect 52500 -5565 52555 -5445
rect 52675 -5565 52720 -5445
rect 52840 -5565 52885 -5445
rect 53005 -5565 53050 -5445
rect 53170 -5565 53225 -5445
rect 53345 -5565 53370 -5445
rect 30770 -5610 53370 -5565
rect 30770 -5730 30795 -5610
rect 30915 -5730 30960 -5610
rect 31080 -5730 31125 -5610
rect 31245 -5730 31290 -5610
rect 31410 -5730 31465 -5610
rect 31585 -5730 31630 -5610
rect 31750 -5730 31795 -5610
rect 31915 -5730 31960 -5610
rect 32080 -5730 32135 -5610
rect 32255 -5730 32300 -5610
rect 32420 -5730 32465 -5610
rect 32585 -5730 32630 -5610
rect 32750 -5730 32805 -5610
rect 32925 -5730 32970 -5610
rect 33090 -5730 33135 -5610
rect 33255 -5730 33300 -5610
rect 33420 -5730 33475 -5610
rect 33595 -5730 33640 -5610
rect 33760 -5730 33805 -5610
rect 33925 -5730 33970 -5610
rect 34090 -5730 34145 -5610
rect 34265 -5730 34310 -5610
rect 34430 -5730 34475 -5610
rect 34595 -5730 34640 -5610
rect 34760 -5730 34815 -5610
rect 34935 -5730 34980 -5610
rect 35100 -5730 35145 -5610
rect 35265 -5730 35310 -5610
rect 35430 -5730 35485 -5610
rect 35605 -5730 35650 -5610
rect 35770 -5730 35815 -5610
rect 35935 -5730 35980 -5610
rect 36100 -5730 36155 -5610
rect 36275 -5730 36485 -5610
rect 36605 -5730 36650 -5610
rect 36770 -5730 36815 -5610
rect 36935 -5730 36980 -5610
rect 37100 -5730 37155 -5610
rect 37275 -5730 37320 -5610
rect 37440 -5730 37485 -5610
rect 37605 -5730 37650 -5610
rect 37770 -5730 37825 -5610
rect 37945 -5730 37990 -5610
rect 38110 -5730 38155 -5610
rect 38275 -5730 38320 -5610
rect 38440 -5730 38495 -5610
rect 38615 -5730 38660 -5610
rect 38780 -5730 38825 -5610
rect 38945 -5730 38990 -5610
rect 39110 -5730 39165 -5610
rect 39285 -5730 39330 -5610
rect 39450 -5730 39495 -5610
rect 39615 -5730 39660 -5610
rect 39780 -5730 39835 -5610
rect 39955 -5730 40000 -5610
rect 40120 -5730 40165 -5610
rect 40285 -5730 40330 -5610
rect 40450 -5730 40505 -5610
rect 40625 -5730 40670 -5610
rect 40790 -5730 40835 -5610
rect 40955 -5730 41000 -5610
rect 41120 -5730 41175 -5610
rect 41295 -5730 41340 -5610
rect 41460 -5730 41505 -5610
rect 41625 -5730 41670 -5610
rect 41790 -5730 41845 -5610
rect 41965 -5730 42175 -5610
rect 42295 -5730 42340 -5610
rect 42460 -5730 42505 -5610
rect 42625 -5730 42670 -5610
rect 42790 -5730 42845 -5610
rect 42965 -5730 43010 -5610
rect 43130 -5730 43175 -5610
rect 43295 -5730 43340 -5610
rect 43460 -5730 43515 -5610
rect 43635 -5730 43680 -5610
rect 43800 -5730 43845 -5610
rect 43965 -5730 44010 -5610
rect 44130 -5730 44185 -5610
rect 44305 -5730 44350 -5610
rect 44470 -5730 44515 -5610
rect 44635 -5730 44680 -5610
rect 44800 -5730 44855 -5610
rect 44975 -5730 45020 -5610
rect 45140 -5730 45185 -5610
rect 45305 -5730 45350 -5610
rect 45470 -5730 45525 -5610
rect 45645 -5730 45690 -5610
rect 45810 -5730 45855 -5610
rect 45975 -5730 46020 -5610
rect 46140 -5730 46195 -5610
rect 46315 -5730 46360 -5610
rect 46480 -5730 46525 -5610
rect 46645 -5730 46690 -5610
rect 46810 -5730 46865 -5610
rect 46985 -5730 47030 -5610
rect 47150 -5730 47195 -5610
rect 47315 -5730 47360 -5610
rect 47480 -5730 47535 -5610
rect 47655 -5730 47865 -5610
rect 47985 -5730 48030 -5610
rect 48150 -5730 48195 -5610
rect 48315 -5730 48360 -5610
rect 48480 -5730 48535 -5610
rect 48655 -5730 48700 -5610
rect 48820 -5730 48865 -5610
rect 48985 -5730 49030 -5610
rect 49150 -5730 49205 -5610
rect 49325 -5730 49370 -5610
rect 49490 -5730 49535 -5610
rect 49655 -5730 49700 -5610
rect 49820 -5730 49875 -5610
rect 49995 -5730 50040 -5610
rect 50160 -5730 50205 -5610
rect 50325 -5730 50370 -5610
rect 50490 -5730 50545 -5610
rect 50665 -5730 50710 -5610
rect 50830 -5730 50875 -5610
rect 50995 -5730 51040 -5610
rect 51160 -5730 51215 -5610
rect 51335 -5730 51380 -5610
rect 51500 -5730 51545 -5610
rect 51665 -5730 51710 -5610
rect 51830 -5730 51885 -5610
rect 52005 -5730 52050 -5610
rect 52170 -5730 52215 -5610
rect 52335 -5730 52380 -5610
rect 52500 -5730 52555 -5610
rect 52675 -5730 52720 -5610
rect 52840 -5730 52885 -5610
rect 53005 -5730 53050 -5610
rect 53170 -5730 53225 -5610
rect 53345 -5730 53370 -5610
rect 30770 -5785 53370 -5730
rect 30770 -5905 30795 -5785
rect 30915 -5905 30960 -5785
rect 31080 -5905 31125 -5785
rect 31245 -5905 31290 -5785
rect 31410 -5905 31465 -5785
rect 31585 -5905 31630 -5785
rect 31750 -5905 31795 -5785
rect 31915 -5905 31960 -5785
rect 32080 -5905 32135 -5785
rect 32255 -5905 32300 -5785
rect 32420 -5905 32465 -5785
rect 32585 -5905 32630 -5785
rect 32750 -5905 32805 -5785
rect 32925 -5905 32970 -5785
rect 33090 -5905 33135 -5785
rect 33255 -5905 33300 -5785
rect 33420 -5905 33475 -5785
rect 33595 -5905 33640 -5785
rect 33760 -5905 33805 -5785
rect 33925 -5905 33970 -5785
rect 34090 -5905 34145 -5785
rect 34265 -5905 34310 -5785
rect 34430 -5905 34475 -5785
rect 34595 -5905 34640 -5785
rect 34760 -5905 34815 -5785
rect 34935 -5905 34980 -5785
rect 35100 -5905 35145 -5785
rect 35265 -5905 35310 -5785
rect 35430 -5905 35485 -5785
rect 35605 -5905 35650 -5785
rect 35770 -5905 35815 -5785
rect 35935 -5905 35980 -5785
rect 36100 -5905 36155 -5785
rect 36275 -5905 36485 -5785
rect 36605 -5905 36650 -5785
rect 36770 -5905 36815 -5785
rect 36935 -5905 36980 -5785
rect 37100 -5905 37155 -5785
rect 37275 -5905 37320 -5785
rect 37440 -5905 37485 -5785
rect 37605 -5905 37650 -5785
rect 37770 -5905 37825 -5785
rect 37945 -5905 37990 -5785
rect 38110 -5905 38155 -5785
rect 38275 -5905 38320 -5785
rect 38440 -5905 38495 -5785
rect 38615 -5905 38660 -5785
rect 38780 -5905 38825 -5785
rect 38945 -5905 38990 -5785
rect 39110 -5905 39165 -5785
rect 39285 -5905 39330 -5785
rect 39450 -5905 39495 -5785
rect 39615 -5905 39660 -5785
rect 39780 -5905 39835 -5785
rect 39955 -5905 40000 -5785
rect 40120 -5905 40165 -5785
rect 40285 -5905 40330 -5785
rect 40450 -5905 40505 -5785
rect 40625 -5905 40670 -5785
rect 40790 -5905 40835 -5785
rect 40955 -5905 41000 -5785
rect 41120 -5905 41175 -5785
rect 41295 -5905 41340 -5785
rect 41460 -5905 41505 -5785
rect 41625 -5905 41670 -5785
rect 41790 -5905 41845 -5785
rect 41965 -5905 42175 -5785
rect 42295 -5905 42340 -5785
rect 42460 -5905 42505 -5785
rect 42625 -5905 42670 -5785
rect 42790 -5905 42845 -5785
rect 42965 -5905 43010 -5785
rect 43130 -5905 43175 -5785
rect 43295 -5905 43340 -5785
rect 43460 -5905 43515 -5785
rect 43635 -5905 43680 -5785
rect 43800 -5905 43845 -5785
rect 43965 -5905 44010 -5785
rect 44130 -5905 44185 -5785
rect 44305 -5905 44350 -5785
rect 44470 -5905 44515 -5785
rect 44635 -5905 44680 -5785
rect 44800 -5905 44855 -5785
rect 44975 -5905 45020 -5785
rect 45140 -5905 45185 -5785
rect 45305 -5905 45350 -5785
rect 45470 -5905 45525 -5785
rect 45645 -5905 45690 -5785
rect 45810 -5905 45855 -5785
rect 45975 -5905 46020 -5785
rect 46140 -5905 46195 -5785
rect 46315 -5905 46360 -5785
rect 46480 -5905 46525 -5785
rect 46645 -5905 46690 -5785
rect 46810 -5905 46865 -5785
rect 46985 -5905 47030 -5785
rect 47150 -5905 47195 -5785
rect 47315 -5905 47360 -5785
rect 47480 -5905 47535 -5785
rect 47655 -5905 47865 -5785
rect 47985 -5905 48030 -5785
rect 48150 -5905 48195 -5785
rect 48315 -5905 48360 -5785
rect 48480 -5905 48535 -5785
rect 48655 -5905 48700 -5785
rect 48820 -5905 48865 -5785
rect 48985 -5905 49030 -5785
rect 49150 -5905 49205 -5785
rect 49325 -5905 49370 -5785
rect 49490 -5905 49535 -5785
rect 49655 -5905 49700 -5785
rect 49820 -5905 49875 -5785
rect 49995 -5905 50040 -5785
rect 50160 -5905 50205 -5785
rect 50325 -5905 50370 -5785
rect 50490 -5905 50545 -5785
rect 50665 -5905 50710 -5785
rect 50830 -5905 50875 -5785
rect 50995 -5905 51040 -5785
rect 51160 -5905 51215 -5785
rect 51335 -5905 51380 -5785
rect 51500 -5905 51545 -5785
rect 51665 -5905 51710 -5785
rect 51830 -5905 51885 -5785
rect 52005 -5905 52050 -5785
rect 52170 -5905 52215 -5785
rect 52335 -5905 52380 -5785
rect 52500 -5905 52555 -5785
rect 52675 -5905 52720 -5785
rect 52840 -5905 52885 -5785
rect 53005 -5905 53050 -5785
rect 53170 -5905 53225 -5785
rect 53345 -5905 53370 -5785
rect 30770 -5950 53370 -5905
rect 30770 -6070 30795 -5950
rect 30915 -6070 30960 -5950
rect 31080 -6070 31125 -5950
rect 31245 -6070 31290 -5950
rect 31410 -6070 31465 -5950
rect 31585 -6070 31630 -5950
rect 31750 -6070 31795 -5950
rect 31915 -6070 31960 -5950
rect 32080 -6070 32135 -5950
rect 32255 -6070 32300 -5950
rect 32420 -6070 32465 -5950
rect 32585 -6070 32630 -5950
rect 32750 -6070 32805 -5950
rect 32925 -6070 32970 -5950
rect 33090 -6070 33135 -5950
rect 33255 -6070 33300 -5950
rect 33420 -6070 33475 -5950
rect 33595 -6070 33640 -5950
rect 33760 -6070 33805 -5950
rect 33925 -6070 33970 -5950
rect 34090 -6070 34145 -5950
rect 34265 -6070 34310 -5950
rect 34430 -6070 34475 -5950
rect 34595 -6070 34640 -5950
rect 34760 -6070 34815 -5950
rect 34935 -6070 34980 -5950
rect 35100 -6070 35145 -5950
rect 35265 -6070 35310 -5950
rect 35430 -6070 35485 -5950
rect 35605 -6070 35650 -5950
rect 35770 -6070 35815 -5950
rect 35935 -6070 35980 -5950
rect 36100 -6070 36155 -5950
rect 36275 -6070 36485 -5950
rect 36605 -6070 36650 -5950
rect 36770 -6070 36815 -5950
rect 36935 -6070 36980 -5950
rect 37100 -6070 37155 -5950
rect 37275 -6070 37320 -5950
rect 37440 -6070 37485 -5950
rect 37605 -6070 37650 -5950
rect 37770 -6070 37825 -5950
rect 37945 -6070 37990 -5950
rect 38110 -6070 38155 -5950
rect 38275 -6070 38320 -5950
rect 38440 -6070 38495 -5950
rect 38615 -6070 38660 -5950
rect 38780 -6070 38825 -5950
rect 38945 -6070 38990 -5950
rect 39110 -6070 39165 -5950
rect 39285 -6070 39330 -5950
rect 39450 -6070 39495 -5950
rect 39615 -6070 39660 -5950
rect 39780 -6070 39835 -5950
rect 39955 -6070 40000 -5950
rect 40120 -6070 40165 -5950
rect 40285 -6070 40330 -5950
rect 40450 -6070 40505 -5950
rect 40625 -6070 40670 -5950
rect 40790 -6070 40835 -5950
rect 40955 -6070 41000 -5950
rect 41120 -6070 41175 -5950
rect 41295 -6070 41340 -5950
rect 41460 -6070 41505 -5950
rect 41625 -6070 41670 -5950
rect 41790 -6070 41845 -5950
rect 41965 -6070 42175 -5950
rect 42295 -6070 42340 -5950
rect 42460 -6070 42505 -5950
rect 42625 -6070 42670 -5950
rect 42790 -6070 42845 -5950
rect 42965 -6070 43010 -5950
rect 43130 -6070 43175 -5950
rect 43295 -6070 43340 -5950
rect 43460 -6070 43515 -5950
rect 43635 -6070 43680 -5950
rect 43800 -6070 43845 -5950
rect 43965 -6070 44010 -5950
rect 44130 -6070 44185 -5950
rect 44305 -6070 44350 -5950
rect 44470 -6070 44515 -5950
rect 44635 -6070 44680 -5950
rect 44800 -6070 44855 -5950
rect 44975 -6070 45020 -5950
rect 45140 -6070 45185 -5950
rect 45305 -6070 45350 -5950
rect 45470 -6070 45525 -5950
rect 45645 -6070 45690 -5950
rect 45810 -6070 45855 -5950
rect 45975 -6070 46020 -5950
rect 46140 -6070 46195 -5950
rect 46315 -6070 46360 -5950
rect 46480 -6070 46525 -5950
rect 46645 -6070 46690 -5950
rect 46810 -6070 46865 -5950
rect 46985 -6070 47030 -5950
rect 47150 -6070 47195 -5950
rect 47315 -6070 47360 -5950
rect 47480 -6070 47535 -5950
rect 47655 -6070 47865 -5950
rect 47985 -6070 48030 -5950
rect 48150 -6070 48195 -5950
rect 48315 -6070 48360 -5950
rect 48480 -6070 48535 -5950
rect 48655 -6070 48700 -5950
rect 48820 -6070 48865 -5950
rect 48985 -6070 49030 -5950
rect 49150 -6070 49205 -5950
rect 49325 -6070 49370 -5950
rect 49490 -6070 49535 -5950
rect 49655 -6070 49700 -5950
rect 49820 -6070 49875 -5950
rect 49995 -6070 50040 -5950
rect 50160 -6070 50205 -5950
rect 50325 -6070 50370 -5950
rect 50490 -6070 50545 -5950
rect 50665 -6070 50710 -5950
rect 50830 -6070 50875 -5950
rect 50995 -6070 51040 -5950
rect 51160 -6070 51215 -5950
rect 51335 -6070 51380 -5950
rect 51500 -6070 51545 -5950
rect 51665 -6070 51710 -5950
rect 51830 -6070 51885 -5950
rect 52005 -6070 52050 -5950
rect 52170 -6070 52215 -5950
rect 52335 -6070 52380 -5950
rect 52500 -6070 52555 -5950
rect 52675 -6070 52720 -5950
rect 52840 -6070 52885 -5950
rect 53005 -6070 53050 -5950
rect 53170 -6070 53225 -5950
rect 53345 -6070 53370 -5950
rect 30770 -6115 53370 -6070
rect 30770 -6235 30795 -6115
rect 30915 -6235 30960 -6115
rect 31080 -6235 31125 -6115
rect 31245 -6235 31290 -6115
rect 31410 -6235 31465 -6115
rect 31585 -6235 31630 -6115
rect 31750 -6235 31795 -6115
rect 31915 -6235 31960 -6115
rect 32080 -6235 32135 -6115
rect 32255 -6235 32300 -6115
rect 32420 -6235 32465 -6115
rect 32585 -6235 32630 -6115
rect 32750 -6235 32805 -6115
rect 32925 -6235 32970 -6115
rect 33090 -6235 33135 -6115
rect 33255 -6235 33300 -6115
rect 33420 -6235 33475 -6115
rect 33595 -6235 33640 -6115
rect 33760 -6235 33805 -6115
rect 33925 -6235 33970 -6115
rect 34090 -6235 34145 -6115
rect 34265 -6235 34310 -6115
rect 34430 -6235 34475 -6115
rect 34595 -6235 34640 -6115
rect 34760 -6235 34815 -6115
rect 34935 -6235 34980 -6115
rect 35100 -6235 35145 -6115
rect 35265 -6235 35310 -6115
rect 35430 -6235 35485 -6115
rect 35605 -6235 35650 -6115
rect 35770 -6235 35815 -6115
rect 35935 -6235 35980 -6115
rect 36100 -6235 36155 -6115
rect 36275 -6235 36485 -6115
rect 36605 -6235 36650 -6115
rect 36770 -6235 36815 -6115
rect 36935 -6235 36980 -6115
rect 37100 -6235 37155 -6115
rect 37275 -6235 37320 -6115
rect 37440 -6235 37485 -6115
rect 37605 -6235 37650 -6115
rect 37770 -6235 37825 -6115
rect 37945 -6235 37990 -6115
rect 38110 -6235 38155 -6115
rect 38275 -6235 38320 -6115
rect 38440 -6235 38495 -6115
rect 38615 -6235 38660 -6115
rect 38780 -6235 38825 -6115
rect 38945 -6235 38990 -6115
rect 39110 -6235 39165 -6115
rect 39285 -6235 39330 -6115
rect 39450 -6235 39495 -6115
rect 39615 -6235 39660 -6115
rect 39780 -6235 39835 -6115
rect 39955 -6235 40000 -6115
rect 40120 -6235 40165 -6115
rect 40285 -6235 40330 -6115
rect 40450 -6235 40505 -6115
rect 40625 -6235 40670 -6115
rect 40790 -6235 40835 -6115
rect 40955 -6235 41000 -6115
rect 41120 -6235 41175 -6115
rect 41295 -6235 41340 -6115
rect 41460 -6235 41505 -6115
rect 41625 -6235 41670 -6115
rect 41790 -6235 41845 -6115
rect 41965 -6235 42175 -6115
rect 42295 -6235 42340 -6115
rect 42460 -6235 42505 -6115
rect 42625 -6235 42670 -6115
rect 42790 -6235 42845 -6115
rect 42965 -6235 43010 -6115
rect 43130 -6235 43175 -6115
rect 43295 -6235 43340 -6115
rect 43460 -6235 43515 -6115
rect 43635 -6235 43680 -6115
rect 43800 -6235 43845 -6115
rect 43965 -6235 44010 -6115
rect 44130 -6235 44185 -6115
rect 44305 -6235 44350 -6115
rect 44470 -6235 44515 -6115
rect 44635 -6235 44680 -6115
rect 44800 -6235 44855 -6115
rect 44975 -6235 45020 -6115
rect 45140 -6235 45185 -6115
rect 45305 -6235 45350 -6115
rect 45470 -6235 45525 -6115
rect 45645 -6235 45690 -6115
rect 45810 -6235 45855 -6115
rect 45975 -6235 46020 -6115
rect 46140 -6235 46195 -6115
rect 46315 -6235 46360 -6115
rect 46480 -6235 46525 -6115
rect 46645 -6235 46690 -6115
rect 46810 -6235 46865 -6115
rect 46985 -6235 47030 -6115
rect 47150 -6235 47195 -6115
rect 47315 -6235 47360 -6115
rect 47480 -6235 47535 -6115
rect 47655 -6235 47865 -6115
rect 47985 -6235 48030 -6115
rect 48150 -6235 48195 -6115
rect 48315 -6235 48360 -6115
rect 48480 -6235 48535 -6115
rect 48655 -6235 48700 -6115
rect 48820 -6235 48865 -6115
rect 48985 -6235 49030 -6115
rect 49150 -6235 49205 -6115
rect 49325 -6235 49370 -6115
rect 49490 -6235 49535 -6115
rect 49655 -6235 49700 -6115
rect 49820 -6235 49875 -6115
rect 49995 -6235 50040 -6115
rect 50160 -6235 50205 -6115
rect 50325 -6235 50370 -6115
rect 50490 -6235 50545 -6115
rect 50665 -6235 50710 -6115
rect 50830 -6235 50875 -6115
rect 50995 -6235 51040 -6115
rect 51160 -6235 51215 -6115
rect 51335 -6235 51380 -6115
rect 51500 -6235 51545 -6115
rect 51665 -6235 51710 -6115
rect 51830 -6235 51885 -6115
rect 52005 -6235 52050 -6115
rect 52170 -6235 52215 -6115
rect 52335 -6235 52380 -6115
rect 52500 -6235 52555 -6115
rect 52675 -6235 52720 -6115
rect 52840 -6235 52885 -6115
rect 53005 -6235 53050 -6115
rect 53170 -6235 53225 -6115
rect 53345 -6235 53370 -6115
rect 30770 -6280 53370 -6235
rect 30770 -6400 30795 -6280
rect 30915 -6400 30960 -6280
rect 31080 -6400 31125 -6280
rect 31245 -6400 31290 -6280
rect 31410 -6400 31465 -6280
rect 31585 -6400 31630 -6280
rect 31750 -6400 31795 -6280
rect 31915 -6400 31960 -6280
rect 32080 -6400 32135 -6280
rect 32255 -6400 32300 -6280
rect 32420 -6400 32465 -6280
rect 32585 -6400 32630 -6280
rect 32750 -6400 32805 -6280
rect 32925 -6400 32970 -6280
rect 33090 -6400 33135 -6280
rect 33255 -6400 33300 -6280
rect 33420 -6400 33475 -6280
rect 33595 -6400 33640 -6280
rect 33760 -6400 33805 -6280
rect 33925 -6400 33970 -6280
rect 34090 -6400 34145 -6280
rect 34265 -6400 34310 -6280
rect 34430 -6400 34475 -6280
rect 34595 -6400 34640 -6280
rect 34760 -6400 34815 -6280
rect 34935 -6400 34980 -6280
rect 35100 -6400 35145 -6280
rect 35265 -6400 35310 -6280
rect 35430 -6400 35485 -6280
rect 35605 -6400 35650 -6280
rect 35770 -6400 35815 -6280
rect 35935 -6400 35980 -6280
rect 36100 -6400 36155 -6280
rect 36275 -6400 36485 -6280
rect 36605 -6400 36650 -6280
rect 36770 -6400 36815 -6280
rect 36935 -6400 36980 -6280
rect 37100 -6400 37155 -6280
rect 37275 -6400 37320 -6280
rect 37440 -6400 37485 -6280
rect 37605 -6400 37650 -6280
rect 37770 -6400 37825 -6280
rect 37945 -6400 37990 -6280
rect 38110 -6400 38155 -6280
rect 38275 -6400 38320 -6280
rect 38440 -6400 38495 -6280
rect 38615 -6400 38660 -6280
rect 38780 -6400 38825 -6280
rect 38945 -6400 38990 -6280
rect 39110 -6400 39165 -6280
rect 39285 -6400 39330 -6280
rect 39450 -6400 39495 -6280
rect 39615 -6400 39660 -6280
rect 39780 -6400 39835 -6280
rect 39955 -6400 40000 -6280
rect 40120 -6400 40165 -6280
rect 40285 -6400 40330 -6280
rect 40450 -6400 40505 -6280
rect 40625 -6400 40670 -6280
rect 40790 -6400 40835 -6280
rect 40955 -6400 41000 -6280
rect 41120 -6400 41175 -6280
rect 41295 -6400 41340 -6280
rect 41460 -6400 41505 -6280
rect 41625 -6400 41670 -6280
rect 41790 -6400 41845 -6280
rect 41965 -6400 42175 -6280
rect 42295 -6400 42340 -6280
rect 42460 -6400 42505 -6280
rect 42625 -6400 42670 -6280
rect 42790 -6400 42845 -6280
rect 42965 -6400 43010 -6280
rect 43130 -6400 43175 -6280
rect 43295 -6400 43340 -6280
rect 43460 -6400 43515 -6280
rect 43635 -6400 43680 -6280
rect 43800 -6400 43845 -6280
rect 43965 -6400 44010 -6280
rect 44130 -6400 44185 -6280
rect 44305 -6400 44350 -6280
rect 44470 -6400 44515 -6280
rect 44635 -6400 44680 -6280
rect 44800 -6400 44855 -6280
rect 44975 -6400 45020 -6280
rect 45140 -6400 45185 -6280
rect 45305 -6400 45350 -6280
rect 45470 -6400 45525 -6280
rect 45645 -6400 45690 -6280
rect 45810 -6400 45855 -6280
rect 45975 -6400 46020 -6280
rect 46140 -6400 46195 -6280
rect 46315 -6400 46360 -6280
rect 46480 -6400 46525 -6280
rect 46645 -6400 46690 -6280
rect 46810 -6400 46865 -6280
rect 46985 -6400 47030 -6280
rect 47150 -6400 47195 -6280
rect 47315 -6400 47360 -6280
rect 47480 -6400 47535 -6280
rect 47655 -6400 47865 -6280
rect 47985 -6400 48030 -6280
rect 48150 -6400 48195 -6280
rect 48315 -6400 48360 -6280
rect 48480 -6400 48535 -6280
rect 48655 -6400 48700 -6280
rect 48820 -6400 48865 -6280
rect 48985 -6400 49030 -6280
rect 49150 -6400 49205 -6280
rect 49325 -6400 49370 -6280
rect 49490 -6400 49535 -6280
rect 49655 -6400 49700 -6280
rect 49820 -6400 49875 -6280
rect 49995 -6400 50040 -6280
rect 50160 -6400 50205 -6280
rect 50325 -6400 50370 -6280
rect 50490 -6400 50545 -6280
rect 50665 -6400 50710 -6280
rect 50830 -6400 50875 -6280
rect 50995 -6400 51040 -6280
rect 51160 -6400 51215 -6280
rect 51335 -6400 51380 -6280
rect 51500 -6400 51545 -6280
rect 51665 -6400 51710 -6280
rect 51830 -6400 51885 -6280
rect 52005 -6400 52050 -6280
rect 52170 -6400 52215 -6280
rect 52335 -6400 52380 -6280
rect 52500 -6400 52555 -6280
rect 52675 -6400 52720 -6280
rect 52840 -6400 52885 -6280
rect 53005 -6400 53050 -6280
rect 53170 -6400 53225 -6280
rect 53345 -6400 53370 -6280
rect 30770 -6455 53370 -6400
rect 30770 -6575 30795 -6455
rect 30915 -6575 30960 -6455
rect 31080 -6575 31125 -6455
rect 31245 -6575 31290 -6455
rect 31410 -6575 31465 -6455
rect 31585 -6575 31630 -6455
rect 31750 -6575 31795 -6455
rect 31915 -6575 31960 -6455
rect 32080 -6575 32135 -6455
rect 32255 -6575 32300 -6455
rect 32420 -6575 32465 -6455
rect 32585 -6575 32630 -6455
rect 32750 -6575 32805 -6455
rect 32925 -6575 32970 -6455
rect 33090 -6575 33135 -6455
rect 33255 -6575 33300 -6455
rect 33420 -6575 33475 -6455
rect 33595 -6575 33640 -6455
rect 33760 -6575 33805 -6455
rect 33925 -6575 33970 -6455
rect 34090 -6575 34145 -6455
rect 34265 -6575 34310 -6455
rect 34430 -6575 34475 -6455
rect 34595 -6575 34640 -6455
rect 34760 -6575 34815 -6455
rect 34935 -6575 34980 -6455
rect 35100 -6575 35145 -6455
rect 35265 -6575 35310 -6455
rect 35430 -6575 35485 -6455
rect 35605 -6575 35650 -6455
rect 35770 -6575 35815 -6455
rect 35935 -6575 35980 -6455
rect 36100 -6575 36155 -6455
rect 36275 -6575 36485 -6455
rect 36605 -6575 36650 -6455
rect 36770 -6575 36815 -6455
rect 36935 -6575 36980 -6455
rect 37100 -6575 37155 -6455
rect 37275 -6575 37320 -6455
rect 37440 -6575 37485 -6455
rect 37605 -6575 37650 -6455
rect 37770 -6575 37825 -6455
rect 37945 -6575 37990 -6455
rect 38110 -6575 38155 -6455
rect 38275 -6575 38320 -6455
rect 38440 -6575 38495 -6455
rect 38615 -6575 38660 -6455
rect 38780 -6575 38825 -6455
rect 38945 -6575 38990 -6455
rect 39110 -6575 39165 -6455
rect 39285 -6575 39330 -6455
rect 39450 -6575 39495 -6455
rect 39615 -6575 39660 -6455
rect 39780 -6575 39835 -6455
rect 39955 -6575 40000 -6455
rect 40120 -6575 40165 -6455
rect 40285 -6575 40330 -6455
rect 40450 -6575 40505 -6455
rect 40625 -6575 40670 -6455
rect 40790 -6575 40835 -6455
rect 40955 -6575 41000 -6455
rect 41120 -6575 41175 -6455
rect 41295 -6575 41340 -6455
rect 41460 -6575 41505 -6455
rect 41625 -6575 41670 -6455
rect 41790 -6575 41845 -6455
rect 41965 -6575 42175 -6455
rect 42295 -6575 42340 -6455
rect 42460 -6575 42505 -6455
rect 42625 -6575 42670 -6455
rect 42790 -6575 42845 -6455
rect 42965 -6575 43010 -6455
rect 43130 -6575 43175 -6455
rect 43295 -6575 43340 -6455
rect 43460 -6575 43515 -6455
rect 43635 -6575 43680 -6455
rect 43800 -6575 43845 -6455
rect 43965 -6575 44010 -6455
rect 44130 -6575 44185 -6455
rect 44305 -6575 44350 -6455
rect 44470 -6575 44515 -6455
rect 44635 -6575 44680 -6455
rect 44800 -6575 44855 -6455
rect 44975 -6575 45020 -6455
rect 45140 -6575 45185 -6455
rect 45305 -6575 45350 -6455
rect 45470 -6575 45525 -6455
rect 45645 -6575 45690 -6455
rect 45810 -6575 45855 -6455
rect 45975 -6575 46020 -6455
rect 46140 -6575 46195 -6455
rect 46315 -6575 46360 -6455
rect 46480 -6575 46525 -6455
rect 46645 -6575 46690 -6455
rect 46810 -6575 46865 -6455
rect 46985 -6575 47030 -6455
rect 47150 -6575 47195 -6455
rect 47315 -6575 47360 -6455
rect 47480 -6575 47535 -6455
rect 47655 -6575 47865 -6455
rect 47985 -6575 48030 -6455
rect 48150 -6575 48195 -6455
rect 48315 -6575 48360 -6455
rect 48480 -6575 48535 -6455
rect 48655 -6575 48700 -6455
rect 48820 -6575 48865 -6455
rect 48985 -6575 49030 -6455
rect 49150 -6575 49205 -6455
rect 49325 -6575 49370 -6455
rect 49490 -6575 49535 -6455
rect 49655 -6575 49700 -6455
rect 49820 -6575 49875 -6455
rect 49995 -6575 50040 -6455
rect 50160 -6575 50205 -6455
rect 50325 -6575 50370 -6455
rect 50490 -6575 50545 -6455
rect 50665 -6575 50710 -6455
rect 50830 -6575 50875 -6455
rect 50995 -6575 51040 -6455
rect 51160 -6575 51215 -6455
rect 51335 -6575 51380 -6455
rect 51500 -6575 51545 -6455
rect 51665 -6575 51710 -6455
rect 51830 -6575 51885 -6455
rect 52005 -6575 52050 -6455
rect 52170 -6575 52215 -6455
rect 52335 -6575 52380 -6455
rect 52500 -6575 52555 -6455
rect 52675 -6575 52720 -6455
rect 52840 -6575 52885 -6455
rect 53005 -6575 53050 -6455
rect 53170 -6575 53225 -6455
rect 53345 -6575 53370 -6455
rect 30770 -6620 53370 -6575
rect 30770 -6740 30795 -6620
rect 30915 -6740 30960 -6620
rect 31080 -6740 31125 -6620
rect 31245 -6740 31290 -6620
rect 31410 -6740 31465 -6620
rect 31585 -6740 31630 -6620
rect 31750 -6740 31795 -6620
rect 31915 -6740 31960 -6620
rect 32080 -6740 32135 -6620
rect 32255 -6740 32300 -6620
rect 32420 -6740 32465 -6620
rect 32585 -6740 32630 -6620
rect 32750 -6740 32805 -6620
rect 32925 -6740 32970 -6620
rect 33090 -6740 33135 -6620
rect 33255 -6740 33300 -6620
rect 33420 -6740 33475 -6620
rect 33595 -6740 33640 -6620
rect 33760 -6740 33805 -6620
rect 33925 -6740 33970 -6620
rect 34090 -6740 34145 -6620
rect 34265 -6740 34310 -6620
rect 34430 -6740 34475 -6620
rect 34595 -6740 34640 -6620
rect 34760 -6740 34815 -6620
rect 34935 -6740 34980 -6620
rect 35100 -6740 35145 -6620
rect 35265 -6740 35310 -6620
rect 35430 -6740 35485 -6620
rect 35605 -6740 35650 -6620
rect 35770 -6740 35815 -6620
rect 35935 -6740 35980 -6620
rect 36100 -6740 36155 -6620
rect 36275 -6740 36485 -6620
rect 36605 -6740 36650 -6620
rect 36770 -6740 36815 -6620
rect 36935 -6740 36980 -6620
rect 37100 -6740 37155 -6620
rect 37275 -6740 37320 -6620
rect 37440 -6740 37485 -6620
rect 37605 -6740 37650 -6620
rect 37770 -6740 37825 -6620
rect 37945 -6740 37990 -6620
rect 38110 -6740 38155 -6620
rect 38275 -6740 38320 -6620
rect 38440 -6740 38495 -6620
rect 38615 -6740 38660 -6620
rect 38780 -6740 38825 -6620
rect 38945 -6740 38990 -6620
rect 39110 -6740 39165 -6620
rect 39285 -6740 39330 -6620
rect 39450 -6740 39495 -6620
rect 39615 -6740 39660 -6620
rect 39780 -6740 39835 -6620
rect 39955 -6740 40000 -6620
rect 40120 -6740 40165 -6620
rect 40285 -6740 40330 -6620
rect 40450 -6740 40505 -6620
rect 40625 -6740 40670 -6620
rect 40790 -6740 40835 -6620
rect 40955 -6740 41000 -6620
rect 41120 -6740 41175 -6620
rect 41295 -6740 41340 -6620
rect 41460 -6740 41505 -6620
rect 41625 -6740 41670 -6620
rect 41790 -6740 41845 -6620
rect 41965 -6740 42175 -6620
rect 42295 -6740 42340 -6620
rect 42460 -6740 42505 -6620
rect 42625 -6740 42670 -6620
rect 42790 -6740 42845 -6620
rect 42965 -6740 43010 -6620
rect 43130 -6740 43175 -6620
rect 43295 -6740 43340 -6620
rect 43460 -6740 43515 -6620
rect 43635 -6740 43680 -6620
rect 43800 -6740 43845 -6620
rect 43965 -6740 44010 -6620
rect 44130 -6740 44185 -6620
rect 44305 -6740 44350 -6620
rect 44470 -6740 44515 -6620
rect 44635 -6740 44680 -6620
rect 44800 -6740 44855 -6620
rect 44975 -6740 45020 -6620
rect 45140 -6740 45185 -6620
rect 45305 -6740 45350 -6620
rect 45470 -6740 45525 -6620
rect 45645 -6740 45690 -6620
rect 45810 -6740 45855 -6620
rect 45975 -6740 46020 -6620
rect 46140 -6740 46195 -6620
rect 46315 -6740 46360 -6620
rect 46480 -6740 46525 -6620
rect 46645 -6740 46690 -6620
rect 46810 -6740 46865 -6620
rect 46985 -6740 47030 -6620
rect 47150 -6740 47195 -6620
rect 47315 -6740 47360 -6620
rect 47480 -6740 47535 -6620
rect 47655 -6740 47865 -6620
rect 47985 -6740 48030 -6620
rect 48150 -6740 48195 -6620
rect 48315 -6740 48360 -6620
rect 48480 -6740 48535 -6620
rect 48655 -6740 48700 -6620
rect 48820 -6740 48865 -6620
rect 48985 -6740 49030 -6620
rect 49150 -6740 49205 -6620
rect 49325 -6740 49370 -6620
rect 49490 -6740 49535 -6620
rect 49655 -6740 49700 -6620
rect 49820 -6740 49875 -6620
rect 49995 -6740 50040 -6620
rect 50160 -6740 50205 -6620
rect 50325 -6740 50370 -6620
rect 50490 -6740 50545 -6620
rect 50665 -6740 50710 -6620
rect 50830 -6740 50875 -6620
rect 50995 -6740 51040 -6620
rect 51160 -6740 51215 -6620
rect 51335 -6740 51380 -6620
rect 51500 -6740 51545 -6620
rect 51665 -6740 51710 -6620
rect 51830 -6740 51885 -6620
rect 52005 -6740 52050 -6620
rect 52170 -6740 52215 -6620
rect 52335 -6740 52380 -6620
rect 52500 -6740 52555 -6620
rect 52675 -6740 52720 -6620
rect 52840 -6740 52885 -6620
rect 53005 -6740 53050 -6620
rect 53170 -6740 53225 -6620
rect 53345 -6740 53370 -6620
rect 30770 -6785 53370 -6740
rect 30770 -6905 30795 -6785
rect 30915 -6905 30960 -6785
rect 31080 -6905 31125 -6785
rect 31245 -6905 31290 -6785
rect 31410 -6905 31465 -6785
rect 31585 -6905 31630 -6785
rect 31750 -6905 31795 -6785
rect 31915 -6905 31960 -6785
rect 32080 -6905 32135 -6785
rect 32255 -6905 32300 -6785
rect 32420 -6905 32465 -6785
rect 32585 -6905 32630 -6785
rect 32750 -6905 32805 -6785
rect 32925 -6905 32970 -6785
rect 33090 -6905 33135 -6785
rect 33255 -6905 33300 -6785
rect 33420 -6905 33475 -6785
rect 33595 -6905 33640 -6785
rect 33760 -6905 33805 -6785
rect 33925 -6905 33970 -6785
rect 34090 -6905 34145 -6785
rect 34265 -6905 34310 -6785
rect 34430 -6905 34475 -6785
rect 34595 -6905 34640 -6785
rect 34760 -6905 34815 -6785
rect 34935 -6905 34980 -6785
rect 35100 -6905 35145 -6785
rect 35265 -6905 35310 -6785
rect 35430 -6905 35485 -6785
rect 35605 -6905 35650 -6785
rect 35770 -6905 35815 -6785
rect 35935 -6905 35980 -6785
rect 36100 -6905 36155 -6785
rect 36275 -6905 36485 -6785
rect 36605 -6905 36650 -6785
rect 36770 -6905 36815 -6785
rect 36935 -6905 36980 -6785
rect 37100 -6905 37155 -6785
rect 37275 -6905 37320 -6785
rect 37440 -6905 37485 -6785
rect 37605 -6905 37650 -6785
rect 37770 -6905 37825 -6785
rect 37945 -6905 37990 -6785
rect 38110 -6905 38155 -6785
rect 38275 -6905 38320 -6785
rect 38440 -6905 38495 -6785
rect 38615 -6905 38660 -6785
rect 38780 -6905 38825 -6785
rect 38945 -6905 38990 -6785
rect 39110 -6905 39165 -6785
rect 39285 -6905 39330 -6785
rect 39450 -6905 39495 -6785
rect 39615 -6905 39660 -6785
rect 39780 -6905 39835 -6785
rect 39955 -6905 40000 -6785
rect 40120 -6905 40165 -6785
rect 40285 -6905 40330 -6785
rect 40450 -6905 40505 -6785
rect 40625 -6905 40670 -6785
rect 40790 -6905 40835 -6785
rect 40955 -6905 41000 -6785
rect 41120 -6905 41175 -6785
rect 41295 -6905 41340 -6785
rect 41460 -6905 41505 -6785
rect 41625 -6905 41670 -6785
rect 41790 -6905 41845 -6785
rect 41965 -6905 42175 -6785
rect 42295 -6905 42340 -6785
rect 42460 -6905 42505 -6785
rect 42625 -6905 42670 -6785
rect 42790 -6905 42845 -6785
rect 42965 -6905 43010 -6785
rect 43130 -6905 43175 -6785
rect 43295 -6905 43340 -6785
rect 43460 -6905 43515 -6785
rect 43635 -6905 43680 -6785
rect 43800 -6905 43845 -6785
rect 43965 -6905 44010 -6785
rect 44130 -6905 44185 -6785
rect 44305 -6905 44350 -6785
rect 44470 -6905 44515 -6785
rect 44635 -6905 44680 -6785
rect 44800 -6905 44855 -6785
rect 44975 -6905 45020 -6785
rect 45140 -6905 45185 -6785
rect 45305 -6905 45350 -6785
rect 45470 -6905 45525 -6785
rect 45645 -6905 45690 -6785
rect 45810 -6905 45855 -6785
rect 45975 -6905 46020 -6785
rect 46140 -6905 46195 -6785
rect 46315 -6905 46360 -6785
rect 46480 -6905 46525 -6785
rect 46645 -6905 46690 -6785
rect 46810 -6905 46865 -6785
rect 46985 -6905 47030 -6785
rect 47150 -6905 47195 -6785
rect 47315 -6905 47360 -6785
rect 47480 -6905 47535 -6785
rect 47655 -6905 47865 -6785
rect 47985 -6905 48030 -6785
rect 48150 -6905 48195 -6785
rect 48315 -6905 48360 -6785
rect 48480 -6905 48535 -6785
rect 48655 -6905 48700 -6785
rect 48820 -6905 48865 -6785
rect 48985 -6905 49030 -6785
rect 49150 -6905 49205 -6785
rect 49325 -6905 49370 -6785
rect 49490 -6905 49535 -6785
rect 49655 -6905 49700 -6785
rect 49820 -6905 49875 -6785
rect 49995 -6905 50040 -6785
rect 50160 -6905 50205 -6785
rect 50325 -6905 50370 -6785
rect 50490 -6905 50545 -6785
rect 50665 -6905 50710 -6785
rect 50830 -6905 50875 -6785
rect 50995 -6905 51040 -6785
rect 51160 -6905 51215 -6785
rect 51335 -6905 51380 -6785
rect 51500 -6905 51545 -6785
rect 51665 -6905 51710 -6785
rect 51830 -6905 51885 -6785
rect 52005 -6905 52050 -6785
rect 52170 -6905 52215 -6785
rect 52335 -6905 52380 -6785
rect 52500 -6905 52555 -6785
rect 52675 -6905 52720 -6785
rect 52840 -6905 52885 -6785
rect 53005 -6905 53050 -6785
rect 53170 -6905 53225 -6785
rect 53345 -6905 53370 -6785
rect 30770 -6950 53370 -6905
rect 30770 -7070 30795 -6950
rect 30915 -7070 30960 -6950
rect 31080 -7070 31125 -6950
rect 31245 -7070 31290 -6950
rect 31410 -7070 31465 -6950
rect 31585 -7070 31630 -6950
rect 31750 -7070 31795 -6950
rect 31915 -7070 31960 -6950
rect 32080 -7070 32135 -6950
rect 32255 -7070 32300 -6950
rect 32420 -7070 32465 -6950
rect 32585 -7070 32630 -6950
rect 32750 -7070 32805 -6950
rect 32925 -7070 32970 -6950
rect 33090 -7070 33135 -6950
rect 33255 -7070 33300 -6950
rect 33420 -7070 33475 -6950
rect 33595 -7070 33640 -6950
rect 33760 -7070 33805 -6950
rect 33925 -7070 33970 -6950
rect 34090 -7070 34145 -6950
rect 34265 -7070 34310 -6950
rect 34430 -7070 34475 -6950
rect 34595 -7070 34640 -6950
rect 34760 -7070 34815 -6950
rect 34935 -7070 34980 -6950
rect 35100 -7070 35145 -6950
rect 35265 -7070 35310 -6950
rect 35430 -7070 35485 -6950
rect 35605 -7070 35650 -6950
rect 35770 -7070 35815 -6950
rect 35935 -7070 35980 -6950
rect 36100 -7070 36155 -6950
rect 36275 -7070 36485 -6950
rect 36605 -7070 36650 -6950
rect 36770 -7070 36815 -6950
rect 36935 -7070 36980 -6950
rect 37100 -7070 37155 -6950
rect 37275 -7070 37320 -6950
rect 37440 -7070 37485 -6950
rect 37605 -7070 37650 -6950
rect 37770 -7070 37825 -6950
rect 37945 -7070 37990 -6950
rect 38110 -7070 38155 -6950
rect 38275 -7070 38320 -6950
rect 38440 -7070 38495 -6950
rect 38615 -7070 38660 -6950
rect 38780 -7070 38825 -6950
rect 38945 -7070 38990 -6950
rect 39110 -7070 39165 -6950
rect 39285 -7070 39330 -6950
rect 39450 -7070 39495 -6950
rect 39615 -7070 39660 -6950
rect 39780 -7070 39835 -6950
rect 39955 -7070 40000 -6950
rect 40120 -7070 40165 -6950
rect 40285 -7070 40330 -6950
rect 40450 -7070 40505 -6950
rect 40625 -7070 40670 -6950
rect 40790 -7070 40835 -6950
rect 40955 -7070 41000 -6950
rect 41120 -7070 41175 -6950
rect 41295 -7070 41340 -6950
rect 41460 -7070 41505 -6950
rect 41625 -7070 41670 -6950
rect 41790 -7070 41845 -6950
rect 41965 -7070 42175 -6950
rect 42295 -7070 42340 -6950
rect 42460 -7070 42505 -6950
rect 42625 -7070 42670 -6950
rect 42790 -7070 42845 -6950
rect 42965 -7070 43010 -6950
rect 43130 -7070 43175 -6950
rect 43295 -7070 43340 -6950
rect 43460 -7070 43515 -6950
rect 43635 -7070 43680 -6950
rect 43800 -7070 43845 -6950
rect 43965 -7070 44010 -6950
rect 44130 -7070 44185 -6950
rect 44305 -7070 44350 -6950
rect 44470 -7070 44515 -6950
rect 44635 -7070 44680 -6950
rect 44800 -7070 44855 -6950
rect 44975 -7070 45020 -6950
rect 45140 -7070 45185 -6950
rect 45305 -7070 45350 -6950
rect 45470 -7070 45525 -6950
rect 45645 -7070 45690 -6950
rect 45810 -7070 45855 -6950
rect 45975 -7070 46020 -6950
rect 46140 -7070 46195 -6950
rect 46315 -7070 46360 -6950
rect 46480 -7070 46525 -6950
rect 46645 -7070 46690 -6950
rect 46810 -7070 46865 -6950
rect 46985 -7070 47030 -6950
rect 47150 -7070 47195 -6950
rect 47315 -7070 47360 -6950
rect 47480 -7070 47535 -6950
rect 47655 -7070 47865 -6950
rect 47985 -7070 48030 -6950
rect 48150 -7070 48195 -6950
rect 48315 -7070 48360 -6950
rect 48480 -7070 48535 -6950
rect 48655 -7070 48700 -6950
rect 48820 -7070 48865 -6950
rect 48985 -7070 49030 -6950
rect 49150 -7070 49205 -6950
rect 49325 -7070 49370 -6950
rect 49490 -7070 49535 -6950
rect 49655 -7070 49700 -6950
rect 49820 -7070 49875 -6950
rect 49995 -7070 50040 -6950
rect 50160 -7070 50205 -6950
rect 50325 -7070 50370 -6950
rect 50490 -7070 50545 -6950
rect 50665 -7070 50710 -6950
rect 50830 -7070 50875 -6950
rect 50995 -7070 51040 -6950
rect 51160 -7070 51215 -6950
rect 51335 -7070 51380 -6950
rect 51500 -7070 51545 -6950
rect 51665 -7070 51710 -6950
rect 51830 -7070 51885 -6950
rect 52005 -7070 52050 -6950
rect 52170 -7070 52215 -6950
rect 52335 -7070 52380 -6950
rect 52500 -7070 52555 -6950
rect 52675 -7070 52720 -6950
rect 52840 -7070 52885 -6950
rect 53005 -7070 53050 -6950
rect 53170 -7070 53225 -6950
rect 53345 -7070 53370 -6950
rect 30770 -7125 53370 -7070
rect 30770 -7245 30795 -7125
rect 30915 -7245 30960 -7125
rect 31080 -7245 31125 -7125
rect 31245 -7245 31290 -7125
rect 31410 -7245 31465 -7125
rect 31585 -7245 31630 -7125
rect 31750 -7245 31795 -7125
rect 31915 -7245 31960 -7125
rect 32080 -7245 32135 -7125
rect 32255 -7245 32300 -7125
rect 32420 -7245 32465 -7125
rect 32585 -7245 32630 -7125
rect 32750 -7245 32805 -7125
rect 32925 -7245 32970 -7125
rect 33090 -7245 33135 -7125
rect 33255 -7245 33300 -7125
rect 33420 -7245 33475 -7125
rect 33595 -7245 33640 -7125
rect 33760 -7245 33805 -7125
rect 33925 -7245 33970 -7125
rect 34090 -7245 34145 -7125
rect 34265 -7245 34310 -7125
rect 34430 -7245 34475 -7125
rect 34595 -7245 34640 -7125
rect 34760 -7245 34815 -7125
rect 34935 -7245 34980 -7125
rect 35100 -7245 35145 -7125
rect 35265 -7245 35310 -7125
rect 35430 -7245 35485 -7125
rect 35605 -7245 35650 -7125
rect 35770 -7245 35815 -7125
rect 35935 -7245 35980 -7125
rect 36100 -7245 36155 -7125
rect 36275 -7245 36485 -7125
rect 36605 -7245 36650 -7125
rect 36770 -7245 36815 -7125
rect 36935 -7245 36980 -7125
rect 37100 -7245 37155 -7125
rect 37275 -7245 37320 -7125
rect 37440 -7245 37485 -7125
rect 37605 -7245 37650 -7125
rect 37770 -7245 37825 -7125
rect 37945 -7245 37990 -7125
rect 38110 -7245 38155 -7125
rect 38275 -7245 38320 -7125
rect 38440 -7245 38495 -7125
rect 38615 -7245 38660 -7125
rect 38780 -7245 38825 -7125
rect 38945 -7245 38990 -7125
rect 39110 -7245 39165 -7125
rect 39285 -7245 39330 -7125
rect 39450 -7245 39495 -7125
rect 39615 -7245 39660 -7125
rect 39780 -7245 39835 -7125
rect 39955 -7245 40000 -7125
rect 40120 -7245 40165 -7125
rect 40285 -7245 40330 -7125
rect 40450 -7245 40505 -7125
rect 40625 -7245 40670 -7125
rect 40790 -7245 40835 -7125
rect 40955 -7245 41000 -7125
rect 41120 -7245 41175 -7125
rect 41295 -7245 41340 -7125
rect 41460 -7245 41505 -7125
rect 41625 -7245 41670 -7125
rect 41790 -7245 41845 -7125
rect 41965 -7245 42175 -7125
rect 42295 -7245 42340 -7125
rect 42460 -7245 42505 -7125
rect 42625 -7245 42670 -7125
rect 42790 -7245 42845 -7125
rect 42965 -7245 43010 -7125
rect 43130 -7245 43175 -7125
rect 43295 -7245 43340 -7125
rect 43460 -7245 43515 -7125
rect 43635 -7245 43680 -7125
rect 43800 -7245 43845 -7125
rect 43965 -7245 44010 -7125
rect 44130 -7245 44185 -7125
rect 44305 -7245 44350 -7125
rect 44470 -7245 44515 -7125
rect 44635 -7245 44680 -7125
rect 44800 -7245 44855 -7125
rect 44975 -7245 45020 -7125
rect 45140 -7245 45185 -7125
rect 45305 -7245 45350 -7125
rect 45470 -7245 45525 -7125
rect 45645 -7245 45690 -7125
rect 45810 -7245 45855 -7125
rect 45975 -7245 46020 -7125
rect 46140 -7245 46195 -7125
rect 46315 -7245 46360 -7125
rect 46480 -7245 46525 -7125
rect 46645 -7245 46690 -7125
rect 46810 -7245 46865 -7125
rect 46985 -7245 47030 -7125
rect 47150 -7245 47195 -7125
rect 47315 -7245 47360 -7125
rect 47480 -7245 47535 -7125
rect 47655 -7245 47865 -7125
rect 47985 -7245 48030 -7125
rect 48150 -7245 48195 -7125
rect 48315 -7245 48360 -7125
rect 48480 -7245 48535 -7125
rect 48655 -7245 48700 -7125
rect 48820 -7245 48865 -7125
rect 48985 -7245 49030 -7125
rect 49150 -7245 49205 -7125
rect 49325 -7245 49370 -7125
rect 49490 -7245 49535 -7125
rect 49655 -7245 49700 -7125
rect 49820 -7245 49875 -7125
rect 49995 -7245 50040 -7125
rect 50160 -7245 50205 -7125
rect 50325 -7245 50370 -7125
rect 50490 -7245 50545 -7125
rect 50665 -7245 50710 -7125
rect 50830 -7245 50875 -7125
rect 50995 -7245 51040 -7125
rect 51160 -7245 51215 -7125
rect 51335 -7245 51380 -7125
rect 51500 -7245 51545 -7125
rect 51665 -7245 51710 -7125
rect 51830 -7245 51885 -7125
rect 52005 -7245 52050 -7125
rect 52170 -7245 52215 -7125
rect 52335 -7245 52380 -7125
rect 52500 -7245 52555 -7125
rect 52675 -7245 52720 -7125
rect 52840 -7245 52885 -7125
rect 53005 -7245 53050 -7125
rect 53170 -7245 53225 -7125
rect 53345 -7245 53370 -7125
rect 30770 -7290 53370 -7245
rect 30770 -7410 30795 -7290
rect 30915 -7410 30960 -7290
rect 31080 -7410 31125 -7290
rect 31245 -7410 31290 -7290
rect 31410 -7410 31465 -7290
rect 31585 -7410 31630 -7290
rect 31750 -7410 31795 -7290
rect 31915 -7410 31960 -7290
rect 32080 -7410 32135 -7290
rect 32255 -7410 32300 -7290
rect 32420 -7410 32465 -7290
rect 32585 -7410 32630 -7290
rect 32750 -7410 32805 -7290
rect 32925 -7410 32970 -7290
rect 33090 -7410 33135 -7290
rect 33255 -7410 33300 -7290
rect 33420 -7410 33475 -7290
rect 33595 -7410 33640 -7290
rect 33760 -7410 33805 -7290
rect 33925 -7410 33970 -7290
rect 34090 -7410 34145 -7290
rect 34265 -7410 34310 -7290
rect 34430 -7410 34475 -7290
rect 34595 -7410 34640 -7290
rect 34760 -7410 34815 -7290
rect 34935 -7410 34980 -7290
rect 35100 -7410 35145 -7290
rect 35265 -7410 35310 -7290
rect 35430 -7410 35485 -7290
rect 35605 -7410 35650 -7290
rect 35770 -7410 35815 -7290
rect 35935 -7410 35980 -7290
rect 36100 -7410 36155 -7290
rect 36275 -7410 36485 -7290
rect 36605 -7410 36650 -7290
rect 36770 -7410 36815 -7290
rect 36935 -7410 36980 -7290
rect 37100 -7410 37155 -7290
rect 37275 -7410 37320 -7290
rect 37440 -7410 37485 -7290
rect 37605 -7410 37650 -7290
rect 37770 -7410 37825 -7290
rect 37945 -7410 37990 -7290
rect 38110 -7410 38155 -7290
rect 38275 -7410 38320 -7290
rect 38440 -7410 38495 -7290
rect 38615 -7410 38660 -7290
rect 38780 -7410 38825 -7290
rect 38945 -7410 38990 -7290
rect 39110 -7410 39165 -7290
rect 39285 -7410 39330 -7290
rect 39450 -7410 39495 -7290
rect 39615 -7410 39660 -7290
rect 39780 -7410 39835 -7290
rect 39955 -7410 40000 -7290
rect 40120 -7410 40165 -7290
rect 40285 -7410 40330 -7290
rect 40450 -7410 40505 -7290
rect 40625 -7410 40670 -7290
rect 40790 -7410 40835 -7290
rect 40955 -7410 41000 -7290
rect 41120 -7410 41175 -7290
rect 41295 -7410 41340 -7290
rect 41460 -7410 41505 -7290
rect 41625 -7410 41670 -7290
rect 41790 -7410 41845 -7290
rect 41965 -7410 42175 -7290
rect 42295 -7410 42340 -7290
rect 42460 -7410 42505 -7290
rect 42625 -7410 42670 -7290
rect 42790 -7410 42845 -7290
rect 42965 -7410 43010 -7290
rect 43130 -7410 43175 -7290
rect 43295 -7410 43340 -7290
rect 43460 -7410 43515 -7290
rect 43635 -7410 43680 -7290
rect 43800 -7410 43845 -7290
rect 43965 -7410 44010 -7290
rect 44130 -7410 44185 -7290
rect 44305 -7410 44350 -7290
rect 44470 -7410 44515 -7290
rect 44635 -7410 44680 -7290
rect 44800 -7410 44855 -7290
rect 44975 -7410 45020 -7290
rect 45140 -7410 45185 -7290
rect 45305 -7410 45350 -7290
rect 45470 -7410 45525 -7290
rect 45645 -7410 45690 -7290
rect 45810 -7410 45855 -7290
rect 45975 -7410 46020 -7290
rect 46140 -7410 46195 -7290
rect 46315 -7410 46360 -7290
rect 46480 -7410 46525 -7290
rect 46645 -7410 46690 -7290
rect 46810 -7410 46865 -7290
rect 46985 -7410 47030 -7290
rect 47150 -7410 47195 -7290
rect 47315 -7410 47360 -7290
rect 47480 -7410 47535 -7290
rect 47655 -7410 47865 -7290
rect 47985 -7410 48030 -7290
rect 48150 -7410 48195 -7290
rect 48315 -7410 48360 -7290
rect 48480 -7410 48535 -7290
rect 48655 -7410 48700 -7290
rect 48820 -7410 48865 -7290
rect 48985 -7410 49030 -7290
rect 49150 -7410 49205 -7290
rect 49325 -7410 49370 -7290
rect 49490 -7410 49535 -7290
rect 49655 -7410 49700 -7290
rect 49820 -7410 49875 -7290
rect 49995 -7410 50040 -7290
rect 50160 -7410 50205 -7290
rect 50325 -7410 50370 -7290
rect 50490 -7410 50545 -7290
rect 50665 -7410 50710 -7290
rect 50830 -7410 50875 -7290
rect 50995 -7410 51040 -7290
rect 51160 -7410 51215 -7290
rect 51335 -7410 51380 -7290
rect 51500 -7410 51545 -7290
rect 51665 -7410 51710 -7290
rect 51830 -7410 51885 -7290
rect 52005 -7410 52050 -7290
rect 52170 -7410 52215 -7290
rect 52335 -7410 52380 -7290
rect 52500 -7410 52555 -7290
rect 52675 -7410 52720 -7290
rect 52840 -7410 52885 -7290
rect 53005 -7410 53050 -7290
rect 53170 -7410 53225 -7290
rect 53345 -7410 53370 -7290
rect 30770 -7455 53370 -7410
rect 30770 -7575 30795 -7455
rect 30915 -7575 30960 -7455
rect 31080 -7575 31125 -7455
rect 31245 -7575 31290 -7455
rect 31410 -7575 31465 -7455
rect 31585 -7575 31630 -7455
rect 31750 -7575 31795 -7455
rect 31915 -7575 31960 -7455
rect 32080 -7575 32135 -7455
rect 32255 -7575 32300 -7455
rect 32420 -7575 32465 -7455
rect 32585 -7575 32630 -7455
rect 32750 -7575 32805 -7455
rect 32925 -7575 32970 -7455
rect 33090 -7575 33135 -7455
rect 33255 -7575 33300 -7455
rect 33420 -7575 33475 -7455
rect 33595 -7575 33640 -7455
rect 33760 -7575 33805 -7455
rect 33925 -7575 33970 -7455
rect 34090 -7575 34145 -7455
rect 34265 -7575 34310 -7455
rect 34430 -7575 34475 -7455
rect 34595 -7575 34640 -7455
rect 34760 -7575 34815 -7455
rect 34935 -7575 34980 -7455
rect 35100 -7575 35145 -7455
rect 35265 -7575 35310 -7455
rect 35430 -7575 35485 -7455
rect 35605 -7575 35650 -7455
rect 35770 -7575 35815 -7455
rect 35935 -7575 35980 -7455
rect 36100 -7575 36155 -7455
rect 36275 -7575 36485 -7455
rect 36605 -7575 36650 -7455
rect 36770 -7575 36815 -7455
rect 36935 -7575 36980 -7455
rect 37100 -7575 37155 -7455
rect 37275 -7575 37320 -7455
rect 37440 -7575 37485 -7455
rect 37605 -7575 37650 -7455
rect 37770 -7575 37825 -7455
rect 37945 -7575 37990 -7455
rect 38110 -7575 38155 -7455
rect 38275 -7575 38320 -7455
rect 38440 -7575 38495 -7455
rect 38615 -7575 38660 -7455
rect 38780 -7575 38825 -7455
rect 38945 -7575 38990 -7455
rect 39110 -7575 39165 -7455
rect 39285 -7575 39330 -7455
rect 39450 -7575 39495 -7455
rect 39615 -7575 39660 -7455
rect 39780 -7575 39835 -7455
rect 39955 -7575 40000 -7455
rect 40120 -7575 40165 -7455
rect 40285 -7575 40330 -7455
rect 40450 -7575 40505 -7455
rect 40625 -7575 40670 -7455
rect 40790 -7575 40835 -7455
rect 40955 -7575 41000 -7455
rect 41120 -7575 41175 -7455
rect 41295 -7575 41340 -7455
rect 41460 -7575 41505 -7455
rect 41625 -7575 41670 -7455
rect 41790 -7575 41845 -7455
rect 41965 -7575 42175 -7455
rect 42295 -7575 42340 -7455
rect 42460 -7575 42505 -7455
rect 42625 -7575 42670 -7455
rect 42790 -7575 42845 -7455
rect 42965 -7575 43010 -7455
rect 43130 -7575 43175 -7455
rect 43295 -7575 43340 -7455
rect 43460 -7575 43515 -7455
rect 43635 -7575 43680 -7455
rect 43800 -7575 43845 -7455
rect 43965 -7575 44010 -7455
rect 44130 -7575 44185 -7455
rect 44305 -7575 44350 -7455
rect 44470 -7575 44515 -7455
rect 44635 -7575 44680 -7455
rect 44800 -7575 44855 -7455
rect 44975 -7575 45020 -7455
rect 45140 -7575 45185 -7455
rect 45305 -7575 45350 -7455
rect 45470 -7575 45525 -7455
rect 45645 -7575 45690 -7455
rect 45810 -7575 45855 -7455
rect 45975 -7575 46020 -7455
rect 46140 -7575 46195 -7455
rect 46315 -7575 46360 -7455
rect 46480 -7575 46525 -7455
rect 46645 -7575 46690 -7455
rect 46810 -7575 46865 -7455
rect 46985 -7575 47030 -7455
rect 47150 -7575 47195 -7455
rect 47315 -7575 47360 -7455
rect 47480 -7575 47535 -7455
rect 47655 -7575 47865 -7455
rect 47985 -7575 48030 -7455
rect 48150 -7575 48195 -7455
rect 48315 -7575 48360 -7455
rect 48480 -7575 48535 -7455
rect 48655 -7575 48700 -7455
rect 48820 -7575 48865 -7455
rect 48985 -7575 49030 -7455
rect 49150 -7575 49205 -7455
rect 49325 -7575 49370 -7455
rect 49490 -7575 49535 -7455
rect 49655 -7575 49700 -7455
rect 49820 -7575 49875 -7455
rect 49995 -7575 50040 -7455
rect 50160 -7575 50205 -7455
rect 50325 -7575 50370 -7455
rect 50490 -7575 50545 -7455
rect 50665 -7575 50710 -7455
rect 50830 -7575 50875 -7455
rect 50995 -7575 51040 -7455
rect 51160 -7575 51215 -7455
rect 51335 -7575 51380 -7455
rect 51500 -7575 51545 -7455
rect 51665 -7575 51710 -7455
rect 51830 -7575 51885 -7455
rect 52005 -7575 52050 -7455
rect 52170 -7575 52215 -7455
rect 52335 -7575 52380 -7455
rect 52500 -7575 52555 -7455
rect 52675 -7575 52720 -7455
rect 52840 -7575 52885 -7455
rect 53005 -7575 53050 -7455
rect 53170 -7575 53225 -7455
rect 53345 -7575 53370 -7455
rect 30770 -7620 53370 -7575
rect 30770 -7740 30795 -7620
rect 30915 -7740 30960 -7620
rect 31080 -7740 31125 -7620
rect 31245 -7740 31290 -7620
rect 31410 -7740 31465 -7620
rect 31585 -7740 31630 -7620
rect 31750 -7740 31795 -7620
rect 31915 -7740 31960 -7620
rect 32080 -7740 32135 -7620
rect 32255 -7740 32300 -7620
rect 32420 -7740 32465 -7620
rect 32585 -7740 32630 -7620
rect 32750 -7740 32805 -7620
rect 32925 -7740 32970 -7620
rect 33090 -7740 33135 -7620
rect 33255 -7740 33300 -7620
rect 33420 -7740 33475 -7620
rect 33595 -7740 33640 -7620
rect 33760 -7740 33805 -7620
rect 33925 -7740 33970 -7620
rect 34090 -7740 34145 -7620
rect 34265 -7740 34310 -7620
rect 34430 -7740 34475 -7620
rect 34595 -7740 34640 -7620
rect 34760 -7740 34815 -7620
rect 34935 -7740 34980 -7620
rect 35100 -7740 35145 -7620
rect 35265 -7740 35310 -7620
rect 35430 -7740 35485 -7620
rect 35605 -7740 35650 -7620
rect 35770 -7740 35815 -7620
rect 35935 -7740 35980 -7620
rect 36100 -7740 36155 -7620
rect 36275 -7740 36485 -7620
rect 36605 -7740 36650 -7620
rect 36770 -7740 36815 -7620
rect 36935 -7740 36980 -7620
rect 37100 -7740 37155 -7620
rect 37275 -7740 37320 -7620
rect 37440 -7740 37485 -7620
rect 37605 -7740 37650 -7620
rect 37770 -7740 37825 -7620
rect 37945 -7740 37990 -7620
rect 38110 -7740 38155 -7620
rect 38275 -7740 38320 -7620
rect 38440 -7740 38495 -7620
rect 38615 -7740 38660 -7620
rect 38780 -7740 38825 -7620
rect 38945 -7740 38990 -7620
rect 39110 -7740 39165 -7620
rect 39285 -7740 39330 -7620
rect 39450 -7740 39495 -7620
rect 39615 -7740 39660 -7620
rect 39780 -7740 39835 -7620
rect 39955 -7740 40000 -7620
rect 40120 -7740 40165 -7620
rect 40285 -7740 40330 -7620
rect 40450 -7740 40505 -7620
rect 40625 -7740 40670 -7620
rect 40790 -7740 40835 -7620
rect 40955 -7740 41000 -7620
rect 41120 -7740 41175 -7620
rect 41295 -7740 41340 -7620
rect 41460 -7740 41505 -7620
rect 41625 -7740 41670 -7620
rect 41790 -7740 41845 -7620
rect 41965 -7740 42175 -7620
rect 42295 -7740 42340 -7620
rect 42460 -7740 42505 -7620
rect 42625 -7740 42670 -7620
rect 42790 -7740 42845 -7620
rect 42965 -7740 43010 -7620
rect 43130 -7740 43175 -7620
rect 43295 -7740 43340 -7620
rect 43460 -7740 43515 -7620
rect 43635 -7740 43680 -7620
rect 43800 -7740 43845 -7620
rect 43965 -7740 44010 -7620
rect 44130 -7740 44185 -7620
rect 44305 -7740 44350 -7620
rect 44470 -7740 44515 -7620
rect 44635 -7740 44680 -7620
rect 44800 -7740 44855 -7620
rect 44975 -7740 45020 -7620
rect 45140 -7740 45185 -7620
rect 45305 -7740 45350 -7620
rect 45470 -7740 45525 -7620
rect 45645 -7740 45690 -7620
rect 45810 -7740 45855 -7620
rect 45975 -7740 46020 -7620
rect 46140 -7740 46195 -7620
rect 46315 -7740 46360 -7620
rect 46480 -7740 46525 -7620
rect 46645 -7740 46690 -7620
rect 46810 -7740 46865 -7620
rect 46985 -7740 47030 -7620
rect 47150 -7740 47195 -7620
rect 47315 -7740 47360 -7620
rect 47480 -7740 47535 -7620
rect 47655 -7740 47865 -7620
rect 47985 -7740 48030 -7620
rect 48150 -7740 48195 -7620
rect 48315 -7740 48360 -7620
rect 48480 -7740 48535 -7620
rect 48655 -7740 48700 -7620
rect 48820 -7740 48865 -7620
rect 48985 -7740 49030 -7620
rect 49150 -7740 49205 -7620
rect 49325 -7740 49370 -7620
rect 49490 -7740 49535 -7620
rect 49655 -7740 49700 -7620
rect 49820 -7740 49875 -7620
rect 49995 -7740 50040 -7620
rect 50160 -7740 50205 -7620
rect 50325 -7740 50370 -7620
rect 50490 -7740 50545 -7620
rect 50665 -7740 50710 -7620
rect 50830 -7740 50875 -7620
rect 50995 -7740 51040 -7620
rect 51160 -7740 51215 -7620
rect 51335 -7740 51380 -7620
rect 51500 -7740 51545 -7620
rect 51665 -7740 51710 -7620
rect 51830 -7740 51885 -7620
rect 52005 -7740 52050 -7620
rect 52170 -7740 52215 -7620
rect 52335 -7740 52380 -7620
rect 52500 -7740 52555 -7620
rect 52675 -7740 52720 -7620
rect 52840 -7740 52885 -7620
rect 53005 -7740 53050 -7620
rect 53170 -7740 53225 -7620
rect 53345 -7740 53370 -7620
rect 30770 -7795 53370 -7740
rect 30770 -7915 30795 -7795
rect 30915 -7915 30960 -7795
rect 31080 -7915 31125 -7795
rect 31245 -7915 31290 -7795
rect 31410 -7915 31465 -7795
rect 31585 -7915 31630 -7795
rect 31750 -7915 31795 -7795
rect 31915 -7915 31960 -7795
rect 32080 -7915 32135 -7795
rect 32255 -7915 32300 -7795
rect 32420 -7915 32465 -7795
rect 32585 -7915 32630 -7795
rect 32750 -7915 32805 -7795
rect 32925 -7915 32970 -7795
rect 33090 -7915 33135 -7795
rect 33255 -7915 33300 -7795
rect 33420 -7915 33475 -7795
rect 33595 -7915 33640 -7795
rect 33760 -7915 33805 -7795
rect 33925 -7915 33970 -7795
rect 34090 -7915 34145 -7795
rect 34265 -7915 34310 -7795
rect 34430 -7915 34475 -7795
rect 34595 -7915 34640 -7795
rect 34760 -7915 34815 -7795
rect 34935 -7915 34980 -7795
rect 35100 -7915 35145 -7795
rect 35265 -7915 35310 -7795
rect 35430 -7915 35485 -7795
rect 35605 -7915 35650 -7795
rect 35770 -7915 35815 -7795
rect 35935 -7915 35980 -7795
rect 36100 -7915 36155 -7795
rect 36275 -7915 36485 -7795
rect 36605 -7915 36650 -7795
rect 36770 -7915 36815 -7795
rect 36935 -7915 36980 -7795
rect 37100 -7915 37155 -7795
rect 37275 -7915 37320 -7795
rect 37440 -7915 37485 -7795
rect 37605 -7915 37650 -7795
rect 37770 -7915 37825 -7795
rect 37945 -7915 37990 -7795
rect 38110 -7915 38155 -7795
rect 38275 -7915 38320 -7795
rect 38440 -7915 38495 -7795
rect 38615 -7915 38660 -7795
rect 38780 -7915 38825 -7795
rect 38945 -7915 38990 -7795
rect 39110 -7915 39165 -7795
rect 39285 -7915 39330 -7795
rect 39450 -7915 39495 -7795
rect 39615 -7915 39660 -7795
rect 39780 -7915 39835 -7795
rect 39955 -7915 40000 -7795
rect 40120 -7915 40165 -7795
rect 40285 -7915 40330 -7795
rect 40450 -7915 40505 -7795
rect 40625 -7915 40670 -7795
rect 40790 -7915 40835 -7795
rect 40955 -7915 41000 -7795
rect 41120 -7915 41175 -7795
rect 41295 -7915 41340 -7795
rect 41460 -7915 41505 -7795
rect 41625 -7915 41670 -7795
rect 41790 -7915 41845 -7795
rect 41965 -7915 42175 -7795
rect 42295 -7915 42340 -7795
rect 42460 -7915 42505 -7795
rect 42625 -7915 42670 -7795
rect 42790 -7915 42845 -7795
rect 42965 -7915 43010 -7795
rect 43130 -7915 43175 -7795
rect 43295 -7915 43340 -7795
rect 43460 -7915 43515 -7795
rect 43635 -7915 43680 -7795
rect 43800 -7915 43845 -7795
rect 43965 -7915 44010 -7795
rect 44130 -7915 44185 -7795
rect 44305 -7915 44350 -7795
rect 44470 -7915 44515 -7795
rect 44635 -7915 44680 -7795
rect 44800 -7915 44855 -7795
rect 44975 -7915 45020 -7795
rect 45140 -7915 45185 -7795
rect 45305 -7915 45350 -7795
rect 45470 -7915 45525 -7795
rect 45645 -7915 45690 -7795
rect 45810 -7915 45855 -7795
rect 45975 -7915 46020 -7795
rect 46140 -7915 46195 -7795
rect 46315 -7915 46360 -7795
rect 46480 -7915 46525 -7795
rect 46645 -7915 46690 -7795
rect 46810 -7915 46865 -7795
rect 46985 -7915 47030 -7795
rect 47150 -7915 47195 -7795
rect 47315 -7915 47360 -7795
rect 47480 -7915 47535 -7795
rect 47655 -7915 47865 -7795
rect 47985 -7915 48030 -7795
rect 48150 -7915 48195 -7795
rect 48315 -7915 48360 -7795
rect 48480 -7915 48535 -7795
rect 48655 -7915 48700 -7795
rect 48820 -7915 48865 -7795
rect 48985 -7915 49030 -7795
rect 49150 -7915 49205 -7795
rect 49325 -7915 49370 -7795
rect 49490 -7915 49535 -7795
rect 49655 -7915 49700 -7795
rect 49820 -7915 49875 -7795
rect 49995 -7915 50040 -7795
rect 50160 -7915 50205 -7795
rect 50325 -7915 50370 -7795
rect 50490 -7915 50545 -7795
rect 50665 -7915 50710 -7795
rect 50830 -7915 50875 -7795
rect 50995 -7915 51040 -7795
rect 51160 -7915 51215 -7795
rect 51335 -7915 51380 -7795
rect 51500 -7915 51545 -7795
rect 51665 -7915 51710 -7795
rect 51830 -7915 51885 -7795
rect 52005 -7915 52050 -7795
rect 52170 -7915 52215 -7795
rect 52335 -7915 52380 -7795
rect 52500 -7915 52555 -7795
rect 52675 -7915 52720 -7795
rect 52840 -7915 52885 -7795
rect 53005 -7915 53050 -7795
rect 53170 -7915 53225 -7795
rect 53345 -7915 53370 -7795
rect 30770 -7960 53370 -7915
rect 30770 -8080 30795 -7960
rect 30915 -8080 30960 -7960
rect 31080 -8080 31125 -7960
rect 31245 -8080 31290 -7960
rect 31410 -8080 31465 -7960
rect 31585 -8080 31630 -7960
rect 31750 -8080 31795 -7960
rect 31915 -8080 31960 -7960
rect 32080 -8080 32135 -7960
rect 32255 -8080 32300 -7960
rect 32420 -8080 32465 -7960
rect 32585 -8080 32630 -7960
rect 32750 -8080 32805 -7960
rect 32925 -8080 32970 -7960
rect 33090 -8080 33135 -7960
rect 33255 -8080 33300 -7960
rect 33420 -8080 33475 -7960
rect 33595 -8080 33640 -7960
rect 33760 -8080 33805 -7960
rect 33925 -8080 33970 -7960
rect 34090 -8080 34145 -7960
rect 34265 -8080 34310 -7960
rect 34430 -8080 34475 -7960
rect 34595 -8080 34640 -7960
rect 34760 -8080 34815 -7960
rect 34935 -8080 34980 -7960
rect 35100 -8080 35145 -7960
rect 35265 -8080 35310 -7960
rect 35430 -8080 35485 -7960
rect 35605 -8080 35650 -7960
rect 35770 -8080 35815 -7960
rect 35935 -8080 35980 -7960
rect 36100 -8080 36155 -7960
rect 36275 -8080 36485 -7960
rect 36605 -8080 36650 -7960
rect 36770 -8080 36815 -7960
rect 36935 -8080 36980 -7960
rect 37100 -8080 37155 -7960
rect 37275 -8080 37320 -7960
rect 37440 -8080 37485 -7960
rect 37605 -8080 37650 -7960
rect 37770 -8080 37825 -7960
rect 37945 -8080 37990 -7960
rect 38110 -8080 38155 -7960
rect 38275 -8080 38320 -7960
rect 38440 -8080 38495 -7960
rect 38615 -8080 38660 -7960
rect 38780 -8080 38825 -7960
rect 38945 -8080 38990 -7960
rect 39110 -8080 39165 -7960
rect 39285 -8080 39330 -7960
rect 39450 -8080 39495 -7960
rect 39615 -8080 39660 -7960
rect 39780 -8080 39835 -7960
rect 39955 -8080 40000 -7960
rect 40120 -8080 40165 -7960
rect 40285 -8080 40330 -7960
rect 40450 -8080 40505 -7960
rect 40625 -8080 40670 -7960
rect 40790 -8080 40835 -7960
rect 40955 -8080 41000 -7960
rect 41120 -8080 41175 -7960
rect 41295 -8080 41340 -7960
rect 41460 -8080 41505 -7960
rect 41625 -8080 41670 -7960
rect 41790 -8080 41845 -7960
rect 41965 -8080 42175 -7960
rect 42295 -8080 42340 -7960
rect 42460 -8080 42505 -7960
rect 42625 -8080 42670 -7960
rect 42790 -8080 42845 -7960
rect 42965 -8080 43010 -7960
rect 43130 -8080 43175 -7960
rect 43295 -8080 43340 -7960
rect 43460 -8080 43515 -7960
rect 43635 -8080 43680 -7960
rect 43800 -8080 43845 -7960
rect 43965 -8080 44010 -7960
rect 44130 -8080 44185 -7960
rect 44305 -8080 44350 -7960
rect 44470 -8080 44515 -7960
rect 44635 -8080 44680 -7960
rect 44800 -8080 44855 -7960
rect 44975 -8080 45020 -7960
rect 45140 -8080 45185 -7960
rect 45305 -8080 45350 -7960
rect 45470 -8080 45525 -7960
rect 45645 -8080 45690 -7960
rect 45810 -8080 45855 -7960
rect 45975 -8080 46020 -7960
rect 46140 -8080 46195 -7960
rect 46315 -8080 46360 -7960
rect 46480 -8080 46525 -7960
rect 46645 -8080 46690 -7960
rect 46810 -8080 46865 -7960
rect 46985 -8080 47030 -7960
rect 47150 -8080 47195 -7960
rect 47315 -8080 47360 -7960
rect 47480 -8080 47535 -7960
rect 47655 -8080 47865 -7960
rect 47985 -8080 48030 -7960
rect 48150 -8080 48195 -7960
rect 48315 -8080 48360 -7960
rect 48480 -8080 48535 -7960
rect 48655 -8080 48700 -7960
rect 48820 -8080 48865 -7960
rect 48985 -8080 49030 -7960
rect 49150 -8080 49205 -7960
rect 49325 -8080 49370 -7960
rect 49490 -8080 49535 -7960
rect 49655 -8080 49700 -7960
rect 49820 -8080 49875 -7960
rect 49995 -8080 50040 -7960
rect 50160 -8080 50205 -7960
rect 50325 -8080 50370 -7960
rect 50490 -8080 50545 -7960
rect 50665 -8080 50710 -7960
rect 50830 -8080 50875 -7960
rect 50995 -8080 51040 -7960
rect 51160 -8080 51215 -7960
rect 51335 -8080 51380 -7960
rect 51500 -8080 51545 -7960
rect 51665 -8080 51710 -7960
rect 51830 -8080 51885 -7960
rect 52005 -8080 52050 -7960
rect 52170 -8080 52215 -7960
rect 52335 -8080 52380 -7960
rect 52500 -8080 52555 -7960
rect 52675 -8080 52720 -7960
rect 52840 -8080 52885 -7960
rect 53005 -8080 53050 -7960
rect 53170 -8080 53225 -7960
rect 53345 -8080 53370 -7960
rect 30770 -8125 53370 -8080
rect 30770 -8245 30795 -8125
rect 30915 -8245 30960 -8125
rect 31080 -8245 31125 -8125
rect 31245 -8245 31290 -8125
rect 31410 -8245 31465 -8125
rect 31585 -8245 31630 -8125
rect 31750 -8245 31795 -8125
rect 31915 -8245 31960 -8125
rect 32080 -8245 32135 -8125
rect 32255 -8245 32300 -8125
rect 32420 -8245 32465 -8125
rect 32585 -8245 32630 -8125
rect 32750 -8245 32805 -8125
rect 32925 -8245 32970 -8125
rect 33090 -8245 33135 -8125
rect 33255 -8245 33300 -8125
rect 33420 -8245 33475 -8125
rect 33595 -8245 33640 -8125
rect 33760 -8245 33805 -8125
rect 33925 -8245 33970 -8125
rect 34090 -8245 34145 -8125
rect 34265 -8245 34310 -8125
rect 34430 -8245 34475 -8125
rect 34595 -8245 34640 -8125
rect 34760 -8245 34815 -8125
rect 34935 -8245 34980 -8125
rect 35100 -8245 35145 -8125
rect 35265 -8245 35310 -8125
rect 35430 -8245 35485 -8125
rect 35605 -8245 35650 -8125
rect 35770 -8245 35815 -8125
rect 35935 -8245 35980 -8125
rect 36100 -8245 36155 -8125
rect 36275 -8245 36485 -8125
rect 36605 -8245 36650 -8125
rect 36770 -8245 36815 -8125
rect 36935 -8245 36980 -8125
rect 37100 -8245 37155 -8125
rect 37275 -8245 37320 -8125
rect 37440 -8245 37485 -8125
rect 37605 -8245 37650 -8125
rect 37770 -8245 37825 -8125
rect 37945 -8245 37990 -8125
rect 38110 -8245 38155 -8125
rect 38275 -8245 38320 -8125
rect 38440 -8245 38495 -8125
rect 38615 -8245 38660 -8125
rect 38780 -8245 38825 -8125
rect 38945 -8245 38990 -8125
rect 39110 -8245 39165 -8125
rect 39285 -8245 39330 -8125
rect 39450 -8245 39495 -8125
rect 39615 -8245 39660 -8125
rect 39780 -8245 39835 -8125
rect 39955 -8245 40000 -8125
rect 40120 -8245 40165 -8125
rect 40285 -8245 40330 -8125
rect 40450 -8245 40505 -8125
rect 40625 -8245 40670 -8125
rect 40790 -8245 40835 -8125
rect 40955 -8245 41000 -8125
rect 41120 -8245 41175 -8125
rect 41295 -8245 41340 -8125
rect 41460 -8245 41505 -8125
rect 41625 -8245 41670 -8125
rect 41790 -8245 41845 -8125
rect 41965 -8245 42175 -8125
rect 42295 -8245 42340 -8125
rect 42460 -8245 42505 -8125
rect 42625 -8245 42670 -8125
rect 42790 -8245 42845 -8125
rect 42965 -8245 43010 -8125
rect 43130 -8245 43175 -8125
rect 43295 -8245 43340 -8125
rect 43460 -8245 43515 -8125
rect 43635 -8245 43680 -8125
rect 43800 -8245 43845 -8125
rect 43965 -8245 44010 -8125
rect 44130 -8245 44185 -8125
rect 44305 -8245 44350 -8125
rect 44470 -8245 44515 -8125
rect 44635 -8245 44680 -8125
rect 44800 -8245 44855 -8125
rect 44975 -8245 45020 -8125
rect 45140 -8245 45185 -8125
rect 45305 -8245 45350 -8125
rect 45470 -8245 45525 -8125
rect 45645 -8245 45690 -8125
rect 45810 -8245 45855 -8125
rect 45975 -8245 46020 -8125
rect 46140 -8245 46195 -8125
rect 46315 -8245 46360 -8125
rect 46480 -8245 46525 -8125
rect 46645 -8245 46690 -8125
rect 46810 -8245 46865 -8125
rect 46985 -8245 47030 -8125
rect 47150 -8245 47195 -8125
rect 47315 -8245 47360 -8125
rect 47480 -8245 47535 -8125
rect 47655 -8245 47865 -8125
rect 47985 -8245 48030 -8125
rect 48150 -8245 48195 -8125
rect 48315 -8245 48360 -8125
rect 48480 -8245 48535 -8125
rect 48655 -8245 48700 -8125
rect 48820 -8245 48865 -8125
rect 48985 -8245 49030 -8125
rect 49150 -8245 49205 -8125
rect 49325 -8245 49370 -8125
rect 49490 -8245 49535 -8125
rect 49655 -8245 49700 -8125
rect 49820 -8245 49875 -8125
rect 49995 -8245 50040 -8125
rect 50160 -8245 50205 -8125
rect 50325 -8245 50370 -8125
rect 50490 -8245 50545 -8125
rect 50665 -8245 50710 -8125
rect 50830 -8245 50875 -8125
rect 50995 -8245 51040 -8125
rect 51160 -8245 51215 -8125
rect 51335 -8245 51380 -8125
rect 51500 -8245 51545 -8125
rect 51665 -8245 51710 -8125
rect 51830 -8245 51885 -8125
rect 52005 -8245 52050 -8125
rect 52170 -8245 52215 -8125
rect 52335 -8245 52380 -8125
rect 52500 -8245 52555 -8125
rect 52675 -8245 52720 -8125
rect 52840 -8245 52885 -8125
rect 53005 -8245 53050 -8125
rect 53170 -8245 53225 -8125
rect 53345 -8245 53370 -8125
rect 30770 -8290 53370 -8245
rect 30770 -8410 30795 -8290
rect 30915 -8410 30960 -8290
rect 31080 -8410 31125 -8290
rect 31245 -8410 31290 -8290
rect 31410 -8410 31465 -8290
rect 31585 -8410 31630 -8290
rect 31750 -8410 31795 -8290
rect 31915 -8410 31960 -8290
rect 32080 -8410 32135 -8290
rect 32255 -8410 32300 -8290
rect 32420 -8410 32465 -8290
rect 32585 -8410 32630 -8290
rect 32750 -8410 32805 -8290
rect 32925 -8410 32970 -8290
rect 33090 -8410 33135 -8290
rect 33255 -8410 33300 -8290
rect 33420 -8410 33475 -8290
rect 33595 -8410 33640 -8290
rect 33760 -8410 33805 -8290
rect 33925 -8410 33970 -8290
rect 34090 -8410 34145 -8290
rect 34265 -8410 34310 -8290
rect 34430 -8410 34475 -8290
rect 34595 -8410 34640 -8290
rect 34760 -8410 34815 -8290
rect 34935 -8410 34980 -8290
rect 35100 -8410 35145 -8290
rect 35265 -8410 35310 -8290
rect 35430 -8410 35485 -8290
rect 35605 -8410 35650 -8290
rect 35770 -8410 35815 -8290
rect 35935 -8410 35980 -8290
rect 36100 -8410 36155 -8290
rect 36275 -8410 36485 -8290
rect 36605 -8410 36650 -8290
rect 36770 -8410 36815 -8290
rect 36935 -8410 36980 -8290
rect 37100 -8410 37155 -8290
rect 37275 -8410 37320 -8290
rect 37440 -8410 37485 -8290
rect 37605 -8410 37650 -8290
rect 37770 -8410 37825 -8290
rect 37945 -8410 37990 -8290
rect 38110 -8410 38155 -8290
rect 38275 -8410 38320 -8290
rect 38440 -8410 38495 -8290
rect 38615 -8410 38660 -8290
rect 38780 -8410 38825 -8290
rect 38945 -8410 38990 -8290
rect 39110 -8410 39165 -8290
rect 39285 -8410 39330 -8290
rect 39450 -8410 39495 -8290
rect 39615 -8410 39660 -8290
rect 39780 -8410 39835 -8290
rect 39955 -8410 40000 -8290
rect 40120 -8410 40165 -8290
rect 40285 -8410 40330 -8290
rect 40450 -8410 40505 -8290
rect 40625 -8410 40670 -8290
rect 40790 -8410 40835 -8290
rect 40955 -8410 41000 -8290
rect 41120 -8410 41175 -8290
rect 41295 -8410 41340 -8290
rect 41460 -8410 41505 -8290
rect 41625 -8410 41670 -8290
rect 41790 -8410 41845 -8290
rect 41965 -8410 42175 -8290
rect 42295 -8410 42340 -8290
rect 42460 -8410 42505 -8290
rect 42625 -8410 42670 -8290
rect 42790 -8410 42845 -8290
rect 42965 -8410 43010 -8290
rect 43130 -8410 43175 -8290
rect 43295 -8410 43340 -8290
rect 43460 -8410 43515 -8290
rect 43635 -8410 43680 -8290
rect 43800 -8410 43845 -8290
rect 43965 -8410 44010 -8290
rect 44130 -8410 44185 -8290
rect 44305 -8410 44350 -8290
rect 44470 -8410 44515 -8290
rect 44635 -8410 44680 -8290
rect 44800 -8410 44855 -8290
rect 44975 -8410 45020 -8290
rect 45140 -8410 45185 -8290
rect 45305 -8410 45350 -8290
rect 45470 -8410 45525 -8290
rect 45645 -8410 45690 -8290
rect 45810 -8410 45855 -8290
rect 45975 -8410 46020 -8290
rect 46140 -8410 46195 -8290
rect 46315 -8410 46360 -8290
rect 46480 -8410 46525 -8290
rect 46645 -8410 46690 -8290
rect 46810 -8410 46865 -8290
rect 46985 -8410 47030 -8290
rect 47150 -8410 47195 -8290
rect 47315 -8410 47360 -8290
rect 47480 -8410 47535 -8290
rect 47655 -8410 47865 -8290
rect 47985 -8410 48030 -8290
rect 48150 -8410 48195 -8290
rect 48315 -8410 48360 -8290
rect 48480 -8410 48535 -8290
rect 48655 -8410 48700 -8290
rect 48820 -8410 48865 -8290
rect 48985 -8410 49030 -8290
rect 49150 -8410 49205 -8290
rect 49325 -8410 49370 -8290
rect 49490 -8410 49535 -8290
rect 49655 -8410 49700 -8290
rect 49820 -8410 49875 -8290
rect 49995 -8410 50040 -8290
rect 50160 -8410 50205 -8290
rect 50325 -8410 50370 -8290
rect 50490 -8410 50545 -8290
rect 50665 -8410 50710 -8290
rect 50830 -8410 50875 -8290
rect 50995 -8410 51040 -8290
rect 51160 -8410 51215 -8290
rect 51335 -8410 51380 -8290
rect 51500 -8410 51545 -8290
rect 51665 -8410 51710 -8290
rect 51830 -8410 51885 -8290
rect 52005 -8410 52050 -8290
rect 52170 -8410 52215 -8290
rect 52335 -8410 52380 -8290
rect 52500 -8410 52555 -8290
rect 52675 -8410 52720 -8290
rect 52840 -8410 52885 -8290
rect 53005 -8410 53050 -8290
rect 53170 -8410 53225 -8290
rect 53345 -8410 53370 -8290
rect 30770 -8465 53370 -8410
rect 30770 -8585 30795 -8465
rect 30915 -8585 30960 -8465
rect 31080 -8585 31125 -8465
rect 31245 -8585 31290 -8465
rect 31410 -8585 31465 -8465
rect 31585 -8585 31630 -8465
rect 31750 -8585 31795 -8465
rect 31915 -8585 31960 -8465
rect 32080 -8585 32135 -8465
rect 32255 -8585 32300 -8465
rect 32420 -8585 32465 -8465
rect 32585 -8585 32630 -8465
rect 32750 -8585 32805 -8465
rect 32925 -8585 32970 -8465
rect 33090 -8585 33135 -8465
rect 33255 -8585 33300 -8465
rect 33420 -8585 33475 -8465
rect 33595 -8585 33640 -8465
rect 33760 -8585 33805 -8465
rect 33925 -8585 33970 -8465
rect 34090 -8585 34145 -8465
rect 34265 -8585 34310 -8465
rect 34430 -8585 34475 -8465
rect 34595 -8585 34640 -8465
rect 34760 -8585 34815 -8465
rect 34935 -8585 34980 -8465
rect 35100 -8585 35145 -8465
rect 35265 -8585 35310 -8465
rect 35430 -8585 35485 -8465
rect 35605 -8585 35650 -8465
rect 35770 -8585 35815 -8465
rect 35935 -8585 35980 -8465
rect 36100 -8585 36155 -8465
rect 36275 -8585 36485 -8465
rect 36605 -8585 36650 -8465
rect 36770 -8585 36815 -8465
rect 36935 -8585 36980 -8465
rect 37100 -8585 37155 -8465
rect 37275 -8585 37320 -8465
rect 37440 -8585 37485 -8465
rect 37605 -8585 37650 -8465
rect 37770 -8585 37825 -8465
rect 37945 -8585 37990 -8465
rect 38110 -8585 38155 -8465
rect 38275 -8585 38320 -8465
rect 38440 -8585 38495 -8465
rect 38615 -8585 38660 -8465
rect 38780 -8585 38825 -8465
rect 38945 -8585 38990 -8465
rect 39110 -8585 39165 -8465
rect 39285 -8585 39330 -8465
rect 39450 -8585 39495 -8465
rect 39615 -8585 39660 -8465
rect 39780 -8585 39835 -8465
rect 39955 -8585 40000 -8465
rect 40120 -8585 40165 -8465
rect 40285 -8585 40330 -8465
rect 40450 -8585 40505 -8465
rect 40625 -8585 40670 -8465
rect 40790 -8585 40835 -8465
rect 40955 -8585 41000 -8465
rect 41120 -8585 41175 -8465
rect 41295 -8585 41340 -8465
rect 41460 -8585 41505 -8465
rect 41625 -8585 41670 -8465
rect 41790 -8585 41845 -8465
rect 41965 -8585 42175 -8465
rect 42295 -8585 42340 -8465
rect 42460 -8585 42505 -8465
rect 42625 -8585 42670 -8465
rect 42790 -8585 42845 -8465
rect 42965 -8585 43010 -8465
rect 43130 -8585 43175 -8465
rect 43295 -8585 43340 -8465
rect 43460 -8585 43515 -8465
rect 43635 -8585 43680 -8465
rect 43800 -8585 43845 -8465
rect 43965 -8585 44010 -8465
rect 44130 -8585 44185 -8465
rect 44305 -8585 44350 -8465
rect 44470 -8585 44515 -8465
rect 44635 -8585 44680 -8465
rect 44800 -8585 44855 -8465
rect 44975 -8585 45020 -8465
rect 45140 -8585 45185 -8465
rect 45305 -8585 45350 -8465
rect 45470 -8585 45525 -8465
rect 45645 -8585 45690 -8465
rect 45810 -8585 45855 -8465
rect 45975 -8585 46020 -8465
rect 46140 -8585 46195 -8465
rect 46315 -8585 46360 -8465
rect 46480 -8585 46525 -8465
rect 46645 -8585 46690 -8465
rect 46810 -8585 46865 -8465
rect 46985 -8585 47030 -8465
rect 47150 -8585 47195 -8465
rect 47315 -8585 47360 -8465
rect 47480 -8585 47535 -8465
rect 47655 -8585 47865 -8465
rect 47985 -8585 48030 -8465
rect 48150 -8585 48195 -8465
rect 48315 -8585 48360 -8465
rect 48480 -8585 48535 -8465
rect 48655 -8585 48700 -8465
rect 48820 -8585 48865 -8465
rect 48985 -8585 49030 -8465
rect 49150 -8585 49205 -8465
rect 49325 -8585 49370 -8465
rect 49490 -8585 49535 -8465
rect 49655 -8585 49700 -8465
rect 49820 -8585 49875 -8465
rect 49995 -8585 50040 -8465
rect 50160 -8585 50205 -8465
rect 50325 -8585 50370 -8465
rect 50490 -8585 50545 -8465
rect 50665 -8585 50710 -8465
rect 50830 -8585 50875 -8465
rect 50995 -8585 51040 -8465
rect 51160 -8585 51215 -8465
rect 51335 -8585 51380 -8465
rect 51500 -8585 51545 -8465
rect 51665 -8585 51710 -8465
rect 51830 -8585 51885 -8465
rect 52005 -8585 52050 -8465
rect 52170 -8585 52215 -8465
rect 52335 -8585 52380 -8465
rect 52500 -8585 52555 -8465
rect 52675 -8585 52720 -8465
rect 52840 -8585 52885 -8465
rect 53005 -8585 53050 -8465
rect 53170 -8585 53225 -8465
rect 53345 -8585 53370 -8465
rect 30770 -8630 53370 -8585
rect 30770 -8750 30795 -8630
rect 30915 -8750 30960 -8630
rect 31080 -8750 31125 -8630
rect 31245 -8750 31290 -8630
rect 31410 -8750 31465 -8630
rect 31585 -8750 31630 -8630
rect 31750 -8750 31795 -8630
rect 31915 -8750 31960 -8630
rect 32080 -8750 32135 -8630
rect 32255 -8750 32300 -8630
rect 32420 -8750 32465 -8630
rect 32585 -8750 32630 -8630
rect 32750 -8750 32805 -8630
rect 32925 -8750 32970 -8630
rect 33090 -8750 33135 -8630
rect 33255 -8750 33300 -8630
rect 33420 -8750 33475 -8630
rect 33595 -8750 33640 -8630
rect 33760 -8750 33805 -8630
rect 33925 -8750 33970 -8630
rect 34090 -8750 34145 -8630
rect 34265 -8750 34310 -8630
rect 34430 -8750 34475 -8630
rect 34595 -8750 34640 -8630
rect 34760 -8750 34815 -8630
rect 34935 -8750 34980 -8630
rect 35100 -8750 35145 -8630
rect 35265 -8750 35310 -8630
rect 35430 -8750 35485 -8630
rect 35605 -8750 35650 -8630
rect 35770 -8750 35815 -8630
rect 35935 -8750 35980 -8630
rect 36100 -8750 36155 -8630
rect 36275 -8750 36485 -8630
rect 36605 -8750 36650 -8630
rect 36770 -8750 36815 -8630
rect 36935 -8750 36980 -8630
rect 37100 -8750 37155 -8630
rect 37275 -8750 37320 -8630
rect 37440 -8750 37485 -8630
rect 37605 -8750 37650 -8630
rect 37770 -8750 37825 -8630
rect 37945 -8750 37990 -8630
rect 38110 -8750 38155 -8630
rect 38275 -8750 38320 -8630
rect 38440 -8750 38495 -8630
rect 38615 -8750 38660 -8630
rect 38780 -8750 38825 -8630
rect 38945 -8750 38990 -8630
rect 39110 -8750 39165 -8630
rect 39285 -8750 39330 -8630
rect 39450 -8750 39495 -8630
rect 39615 -8750 39660 -8630
rect 39780 -8750 39835 -8630
rect 39955 -8750 40000 -8630
rect 40120 -8750 40165 -8630
rect 40285 -8750 40330 -8630
rect 40450 -8750 40505 -8630
rect 40625 -8750 40670 -8630
rect 40790 -8750 40835 -8630
rect 40955 -8750 41000 -8630
rect 41120 -8750 41175 -8630
rect 41295 -8750 41340 -8630
rect 41460 -8750 41505 -8630
rect 41625 -8750 41670 -8630
rect 41790 -8750 41845 -8630
rect 41965 -8750 42175 -8630
rect 42295 -8750 42340 -8630
rect 42460 -8750 42505 -8630
rect 42625 -8750 42670 -8630
rect 42790 -8750 42845 -8630
rect 42965 -8750 43010 -8630
rect 43130 -8750 43175 -8630
rect 43295 -8750 43340 -8630
rect 43460 -8750 43515 -8630
rect 43635 -8750 43680 -8630
rect 43800 -8750 43845 -8630
rect 43965 -8750 44010 -8630
rect 44130 -8750 44185 -8630
rect 44305 -8750 44350 -8630
rect 44470 -8750 44515 -8630
rect 44635 -8750 44680 -8630
rect 44800 -8750 44855 -8630
rect 44975 -8750 45020 -8630
rect 45140 -8750 45185 -8630
rect 45305 -8750 45350 -8630
rect 45470 -8750 45525 -8630
rect 45645 -8750 45690 -8630
rect 45810 -8750 45855 -8630
rect 45975 -8750 46020 -8630
rect 46140 -8750 46195 -8630
rect 46315 -8750 46360 -8630
rect 46480 -8750 46525 -8630
rect 46645 -8750 46690 -8630
rect 46810 -8750 46865 -8630
rect 46985 -8750 47030 -8630
rect 47150 -8750 47195 -8630
rect 47315 -8750 47360 -8630
rect 47480 -8750 47535 -8630
rect 47655 -8750 47865 -8630
rect 47985 -8750 48030 -8630
rect 48150 -8750 48195 -8630
rect 48315 -8750 48360 -8630
rect 48480 -8750 48535 -8630
rect 48655 -8750 48700 -8630
rect 48820 -8750 48865 -8630
rect 48985 -8750 49030 -8630
rect 49150 -8750 49205 -8630
rect 49325 -8750 49370 -8630
rect 49490 -8750 49535 -8630
rect 49655 -8750 49700 -8630
rect 49820 -8750 49875 -8630
rect 49995 -8750 50040 -8630
rect 50160 -8750 50205 -8630
rect 50325 -8750 50370 -8630
rect 50490 -8750 50545 -8630
rect 50665 -8750 50710 -8630
rect 50830 -8750 50875 -8630
rect 50995 -8750 51040 -8630
rect 51160 -8750 51215 -8630
rect 51335 -8750 51380 -8630
rect 51500 -8750 51545 -8630
rect 51665 -8750 51710 -8630
rect 51830 -8750 51885 -8630
rect 52005 -8750 52050 -8630
rect 52170 -8750 52215 -8630
rect 52335 -8750 52380 -8630
rect 52500 -8750 52555 -8630
rect 52675 -8750 52720 -8630
rect 52840 -8750 52885 -8630
rect 53005 -8750 53050 -8630
rect 53170 -8750 53225 -8630
rect 53345 -8750 53370 -8630
rect 30770 -8795 53370 -8750
rect 30770 -8915 30795 -8795
rect 30915 -8915 30960 -8795
rect 31080 -8915 31125 -8795
rect 31245 -8915 31290 -8795
rect 31410 -8915 31465 -8795
rect 31585 -8915 31630 -8795
rect 31750 -8915 31795 -8795
rect 31915 -8915 31960 -8795
rect 32080 -8915 32135 -8795
rect 32255 -8915 32300 -8795
rect 32420 -8915 32465 -8795
rect 32585 -8915 32630 -8795
rect 32750 -8915 32805 -8795
rect 32925 -8915 32970 -8795
rect 33090 -8915 33135 -8795
rect 33255 -8915 33300 -8795
rect 33420 -8915 33475 -8795
rect 33595 -8915 33640 -8795
rect 33760 -8915 33805 -8795
rect 33925 -8915 33970 -8795
rect 34090 -8915 34145 -8795
rect 34265 -8915 34310 -8795
rect 34430 -8915 34475 -8795
rect 34595 -8915 34640 -8795
rect 34760 -8915 34815 -8795
rect 34935 -8915 34980 -8795
rect 35100 -8915 35145 -8795
rect 35265 -8915 35310 -8795
rect 35430 -8915 35485 -8795
rect 35605 -8915 35650 -8795
rect 35770 -8915 35815 -8795
rect 35935 -8915 35980 -8795
rect 36100 -8915 36155 -8795
rect 36275 -8915 36485 -8795
rect 36605 -8915 36650 -8795
rect 36770 -8915 36815 -8795
rect 36935 -8915 36980 -8795
rect 37100 -8915 37155 -8795
rect 37275 -8915 37320 -8795
rect 37440 -8915 37485 -8795
rect 37605 -8915 37650 -8795
rect 37770 -8915 37825 -8795
rect 37945 -8915 37990 -8795
rect 38110 -8915 38155 -8795
rect 38275 -8915 38320 -8795
rect 38440 -8915 38495 -8795
rect 38615 -8915 38660 -8795
rect 38780 -8915 38825 -8795
rect 38945 -8915 38990 -8795
rect 39110 -8915 39165 -8795
rect 39285 -8915 39330 -8795
rect 39450 -8915 39495 -8795
rect 39615 -8915 39660 -8795
rect 39780 -8915 39835 -8795
rect 39955 -8915 40000 -8795
rect 40120 -8915 40165 -8795
rect 40285 -8915 40330 -8795
rect 40450 -8915 40505 -8795
rect 40625 -8915 40670 -8795
rect 40790 -8915 40835 -8795
rect 40955 -8915 41000 -8795
rect 41120 -8915 41175 -8795
rect 41295 -8915 41340 -8795
rect 41460 -8915 41505 -8795
rect 41625 -8915 41670 -8795
rect 41790 -8915 41845 -8795
rect 41965 -8915 42175 -8795
rect 42295 -8915 42340 -8795
rect 42460 -8915 42505 -8795
rect 42625 -8915 42670 -8795
rect 42790 -8915 42845 -8795
rect 42965 -8915 43010 -8795
rect 43130 -8915 43175 -8795
rect 43295 -8915 43340 -8795
rect 43460 -8915 43515 -8795
rect 43635 -8915 43680 -8795
rect 43800 -8915 43845 -8795
rect 43965 -8915 44010 -8795
rect 44130 -8915 44185 -8795
rect 44305 -8915 44350 -8795
rect 44470 -8915 44515 -8795
rect 44635 -8915 44680 -8795
rect 44800 -8915 44855 -8795
rect 44975 -8915 45020 -8795
rect 45140 -8915 45185 -8795
rect 45305 -8915 45350 -8795
rect 45470 -8915 45525 -8795
rect 45645 -8915 45690 -8795
rect 45810 -8915 45855 -8795
rect 45975 -8915 46020 -8795
rect 46140 -8915 46195 -8795
rect 46315 -8915 46360 -8795
rect 46480 -8915 46525 -8795
rect 46645 -8915 46690 -8795
rect 46810 -8915 46865 -8795
rect 46985 -8915 47030 -8795
rect 47150 -8915 47195 -8795
rect 47315 -8915 47360 -8795
rect 47480 -8915 47535 -8795
rect 47655 -8915 47865 -8795
rect 47985 -8915 48030 -8795
rect 48150 -8915 48195 -8795
rect 48315 -8915 48360 -8795
rect 48480 -8915 48535 -8795
rect 48655 -8915 48700 -8795
rect 48820 -8915 48865 -8795
rect 48985 -8915 49030 -8795
rect 49150 -8915 49205 -8795
rect 49325 -8915 49370 -8795
rect 49490 -8915 49535 -8795
rect 49655 -8915 49700 -8795
rect 49820 -8915 49875 -8795
rect 49995 -8915 50040 -8795
rect 50160 -8915 50205 -8795
rect 50325 -8915 50370 -8795
rect 50490 -8915 50545 -8795
rect 50665 -8915 50710 -8795
rect 50830 -8915 50875 -8795
rect 50995 -8915 51040 -8795
rect 51160 -8915 51215 -8795
rect 51335 -8915 51380 -8795
rect 51500 -8915 51545 -8795
rect 51665 -8915 51710 -8795
rect 51830 -8915 51885 -8795
rect 52005 -8915 52050 -8795
rect 52170 -8915 52215 -8795
rect 52335 -8915 52380 -8795
rect 52500 -8915 52555 -8795
rect 52675 -8915 52720 -8795
rect 52840 -8915 52885 -8795
rect 53005 -8915 53050 -8795
rect 53170 -8915 53225 -8795
rect 53345 -8915 53370 -8795
rect 30770 -8960 53370 -8915
rect 30770 -9080 30795 -8960
rect 30915 -9080 30960 -8960
rect 31080 -9080 31125 -8960
rect 31245 -9080 31290 -8960
rect 31410 -9080 31465 -8960
rect 31585 -9080 31630 -8960
rect 31750 -9080 31795 -8960
rect 31915 -9080 31960 -8960
rect 32080 -9080 32135 -8960
rect 32255 -9080 32300 -8960
rect 32420 -9080 32465 -8960
rect 32585 -9080 32630 -8960
rect 32750 -9080 32805 -8960
rect 32925 -9080 32970 -8960
rect 33090 -9080 33135 -8960
rect 33255 -9080 33300 -8960
rect 33420 -9080 33475 -8960
rect 33595 -9080 33640 -8960
rect 33760 -9080 33805 -8960
rect 33925 -9080 33970 -8960
rect 34090 -9080 34145 -8960
rect 34265 -9080 34310 -8960
rect 34430 -9080 34475 -8960
rect 34595 -9080 34640 -8960
rect 34760 -9080 34815 -8960
rect 34935 -9080 34980 -8960
rect 35100 -9080 35145 -8960
rect 35265 -9080 35310 -8960
rect 35430 -9080 35485 -8960
rect 35605 -9080 35650 -8960
rect 35770 -9080 35815 -8960
rect 35935 -9080 35980 -8960
rect 36100 -9080 36155 -8960
rect 36275 -9080 36485 -8960
rect 36605 -9080 36650 -8960
rect 36770 -9080 36815 -8960
rect 36935 -9080 36980 -8960
rect 37100 -9080 37155 -8960
rect 37275 -9080 37320 -8960
rect 37440 -9080 37485 -8960
rect 37605 -9080 37650 -8960
rect 37770 -9080 37825 -8960
rect 37945 -9080 37990 -8960
rect 38110 -9080 38155 -8960
rect 38275 -9080 38320 -8960
rect 38440 -9080 38495 -8960
rect 38615 -9080 38660 -8960
rect 38780 -9080 38825 -8960
rect 38945 -9080 38990 -8960
rect 39110 -9080 39165 -8960
rect 39285 -9080 39330 -8960
rect 39450 -9080 39495 -8960
rect 39615 -9080 39660 -8960
rect 39780 -9080 39835 -8960
rect 39955 -9080 40000 -8960
rect 40120 -9080 40165 -8960
rect 40285 -9080 40330 -8960
rect 40450 -9080 40505 -8960
rect 40625 -9080 40670 -8960
rect 40790 -9080 40835 -8960
rect 40955 -9080 41000 -8960
rect 41120 -9080 41175 -8960
rect 41295 -9080 41340 -8960
rect 41460 -9080 41505 -8960
rect 41625 -9080 41670 -8960
rect 41790 -9080 41845 -8960
rect 41965 -9080 42175 -8960
rect 42295 -9080 42340 -8960
rect 42460 -9080 42505 -8960
rect 42625 -9080 42670 -8960
rect 42790 -9080 42845 -8960
rect 42965 -9080 43010 -8960
rect 43130 -9080 43175 -8960
rect 43295 -9080 43340 -8960
rect 43460 -9080 43515 -8960
rect 43635 -9080 43680 -8960
rect 43800 -9080 43845 -8960
rect 43965 -9080 44010 -8960
rect 44130 -9080 44185 -8960
rect 44305 -9080 44350 -8960
rect 44470 -9080 44515 -8960
rect 44635 -9080 44680 -8960
rect 44800 -9080 44855 -8960
rect 44975 -9080 45020 -8960
rect 45140 -9080 45185 -8960
rect 45305 -9080 45350 -8960
rect 45470 -9080 45525 -8960
rect 45645 -9080 45690 -8960
rect 45810 -9080 45855 -8960
rect 45975 -9080 46020 -8960
rect 46140 -9080 46195 -8960
rect 46315 -9080 46360 -8960
rect 46480 -9080 46525 -8960
rect 46645 -9080 46690 -8960
rect 46810 -9080 46865 -8960
rect 46985 -9080 47030 -8960
rect 47150 -9080 47195 -8960
rect 47315 -9080 47360 -8960
rect 47480 -9080 47535 -8960
rect 47655 -9080 47865 -8960
rect 47985 -9080 48030 -8960
rect 48150 -9080 48195 -8960
rect 48315 -9080 48360 -8960
rect 48480 -9080 48535 -8960
rect 48655 -9080 48700 -8960
rect 48820 -9080 48865 -8960
rect 48985 -9080 49030 -8960
rect 49150 -9080 49205 -8960
rect 49325 -9080 49370 -8960
rect 49490 -9080 49535 -8960
rect 49655 -9080 49700 -8960
rect 49820 -9080 49875 -8960
rect 49995 -9080 50040 -8960
rect 50160 -9080 50205 -8960
rect 50325 -9080 50370 -8960
rect 50490 -9080 50545 -8960
rect 50665 -9080 50710 -8960
rect 50830 -9080 50875 -8960
rect 50995 -9080 51040 -8960
rect 51160 -9080 51215 -8960
rect 51335 -9080 51380 -8960
rect 51500 -9080 51545 -8960
rect 51665 -9080 51710 -8960
rect 51830 -9080 51885 -8960
rect 52005 -9080 52050 -8960
rect 52170 -9080 52215 -8960
rect 52335 -9080 52380 -8960
rect 52500 -9080 52555 -8960
rect 52675 -9080 52720 -8960
rect 52840 -9080 52885 -8960
rect 53005 -9080 53050 -8960
rect 53170 -9080 53225 -8960
rect 53345 -9080 53370 -8960
rect 30770 -9135 53370 -9080
rect 30770 -9255 30795 -9135
rect 30915 -9255 30960 -9135
rect 31080 -9255 31125 -9135
rect 31245 -9255 31290 -9135
rect 31410 -9255 31465 -9135
rect 31585 -9255 31630 -9135
rect 31750 -9255 31795 -9135
rect 31915 -9255 31960 -9135
rect 32080 -9255 32135 -9135
rect 32255 -9255 32300 -9135
rect 32420 -9255 32465 -9135
rect 32585 -9255 32630 -9135
rect 32750 -9255 32805 -9135
rect 32925 -9255 32970 -9135
rect 33090 -9255 33135 -9135
rect 33255 -9255 33300 -9135
rect 33420 -9255 33475 -9135
rect 33595 -9255 33640 -9135
rect 33760 -9255 33805 -9135
rect 33925 -9255 33970 -9135
rect 34090 -9255 34145 -9135
rect 34265 -9255 34310 -9135
rect 34430 -9255 34475 -9135
rect 34595 -9255 34640 -9135
rect 34760 -9255 34815 -9135
rect 34935 -9255 34980 -9135
rect 35100 -9255 35145 -9135
rect 35265 -9255 35310 -9135
rect 35430 -9255 35485 -9135
rect 35605 -9255 35650 -9135
rect 35770 -9255 35815 -9135
rect 35935 -9255 35980 -9135
rect 36100 -9255 36155 -9135
rect 36275 -9255 36485 -9135
rect 36605 -9255 36650 -9135
rect 36770 -9255 36815 -9135
rect 36935 -9255 36980 -9135
rect 37100 -9255 37155 -9135
rect 37275 -9255 37320 -9135
rect 37440 -9255 37485 -9135
rect 37605 -9255 37650 -9135
rect 37770 -9255 37825 -9135
rect 37945 -9255 37990 -9135
rect 38110 -9255 38155 -9135
rect 38275 -9255 38320 -9135
rect 38440 -9255 38495 -9135
rect 38615 -9255 38660 -9135
rect 38780 -9255 38825 -9135
rect 38945 -9255 38990 -9135
rect 39110 -9255 39165 -9135
rect 39285 -9255 39330 -9135
rect 39450 -9255 39495 -9135
rect 39615 -9255 39660 -9135
rect 39780 -9255 39835 -9135
rect 39955 -9255 40000 -9135
rect 40120 -9255 40165 -9135
rect 40285 -9255 40330 -9135
rect 40450 -9255 40505 -9135
rect 40625 -9255 40670 -9135
rect 40790 -9255 40835 -9135
rect 40955 -9255 41000 -9135
rect 41120 -9255 41175 -9135
rect 41295 -9255 41340 -9135
rect 41460 -9255 41505 -9135
rect 41625 -9255 41670 -9135
rect 41790 -9255 41845 -9135
rect 41965 -9255 42175 -9135
rect 42295 -9255 42340 -9135
rect 42460 -9255 42505 -9135
rect 42625 -9255 42670 -9135
rect 42790 -9255 42845 -9135
rect 42965 -9255 43010 -9135
rect 43130 -9255 43175 -9135
rect 43295 -9255 43340 -9135
rect 43460 -9255 43515 -9135
rect 43635 -9255 43680 -9135
rect 43800 -9255 43845 -9135
rect 43965 -9255 44010 -9135
rect 44130 -9255 44185 -9135
rect 44305 -9255 44350 -9135
rect 44470 -9255 44515 -9135
rect 44635 -9255 44680 -9135
rect 44800 -9255 44855 -9135
rect 44975 -9255 45020 -9135
rect 45140 -9255 45185 -9135
rect 45305 -9255 45350 -9135
rect 45470 -9255 45525 -9135
rect 45645 -9255 45690 -9135
rect 45810 -9255 45855 -9135
rect 45975 -9255 46020 -9135
rect 46140 -9255 46195 -9135
rect 46315 -9255 46360 -9135
rect 46480 -9255 46525 -9135
rect 46645 -9255 46690 -9135
rect 46810 -9255 46865 -9135
rect 46985 -9255 47030 -9135
rect 47150 -9255 47195 -9135
rect 47315 -9255 47360 -9135
rect 47480 -9255 47535 -9135
rect 47655 -9255 47865 -9135
rect 47985 -9255 48030 -9135
rect 48150 -9255 48195 -9135
rect 48315 -9255 48360 -9135
rect 48480 -9255 48535 -9135
rect 48655 -9255 48700 -9135
rect 48820 -9255 48865 -9135
rect 48985 -9255 49030 -9135
rect 49150 -9255 49205 -9135
rect 49325 -9255 49370 -9135
rect 49490 -9255 49535 -9135
rect 49655 -9255 49700 -9135
rect 49820 -9255 49875 -9135
rect 49995 -9255 50040 -9135
rect 50160 -9255 50205 -9135
rect 50325 -9255 50370 -9135
rect 50490 -9255 50545 -9135
rect 50665 -9255 50710 -9135
rect 50830 -9255 50875 -9135
rect 50995 -9255 51040 -9135
rect 51160 -9255 51215 -9135
rect 51335 -9255 51380 -9135
rect 51500 -9255 51545 -9135
rect 51665 -9255 51710 -9135
rect 51830 -9255 51885 -9135
rect 52005 -9255 52050 -9135
rect 52170 -9255 52215 -9135
rect 52335 -9255 52380 -9135
rect 52500 -9255 52555 -9135
rect 52675 -9255 52720 -9135
rect 52840 -9255 52885 -9135
rect 53005 -9255 53050 -9135
rect 53170 -9255 53225 -9135
rect 53345 -9255 53370 -9135
rect 30770 -9300 53370 -9255
rect 30770 -9420 30795 -9300
rect 30915 -9420 30960 -9300
rect 31080 -9420 31125 -9300
rect 31245 -9420 31290 -9300
rect 31410 -9420 31465 -9300
rect 31585 -9420 31630 -9300
rect 31750 -9420 31795 -9300
rect 31915 -9420 31960 -9300
rect 32080 -9420 32135 -9300
rect 32255 -9420 32300 -9300
rect 32420 -9420 32465 -9300
rect 32585 -9420 32630 -9300
rect 32750 -9420 32805 -9300
rect 32925 -9420 32970 -9300
rect 33090 -9420 33135 -9300
rect 33255 -9420 33300 -9300
rect 33420 -9420 33475 -9300
rect 33595 -9420 33640 -9300
rect 33760 -9420 33805 -9300
rect 33925 -9420 33970 -9300
rect 34090 -9420 34145 -9300
rect 34265 -9420 34310 -9300
rect 34430 -9420 34475 -9300
rect 34595 -9420 34640 -9300
rect 34760 -9420 34815 -9300
rect 34935 -9420 34980 -9300
rect 35100 -9420 35145 -9300
rect 35265 -9420 35310 -9300
rect 35430 -9420 35485 -9300
rect 35605 -9420 35650 -9300
rect 35770 -9420 35815 -9300
rect 35935 -9420 35980 -9300
rect 36100 -9420 36155 -9300
rect 36275 -9420 36485 -9300
rect 36605 -9420 36650 -9300
rect 36770 -9420 36815 -9300
rect 36935 -9420 36980 -9300
rect 37100 -9420 37155 -9300
rect 37275 -9420 37320 -9300
rect 37440 -9420 37485 -9300
rect 37605 -9420 37650 -9300
rect 37770 -9420 37825 -9300
rect 37945 -9420 37990 -9300
rect 38110 -9420 38155 -9300
rect 38275 -9420 38320 -9300
rect 38440 -9420 38495 -9300
rect 38615 -9420 38660 -9300
rect 38780 -9420 38825 -9300
rect 38945 -9420 38990 -9300
rect 39110 -9420 39165 -9300
rect 39285 -9420 39330 -9300
rect 39450 -9420 39495 -9300
rect 39615 -9420 39660 -9300
rect 39780 -9420 39835 -9300
rect 39955 -9420 40000 -9300
rect 40120 -9420 40165 -9300
rect 40285 -9420 40330 -9300
rect 40450 -9420 40505 -9300
rect 40625 -9420 40670 -9300
rect 40790 -9420 40835 -9300
rect 40955 -9420 41000 -9300
rect 41120 -9420 41175 -9300
rect 41295 -9420 41340 -9300
rect 41460 -9420 41505 -9300
rect 41625 -9420 41670 -9300
rect 41790 -9420 41845 -9300
rect 41965 -9420 42175 -9300
rect 42295 -9420 42340 -9300
rect 42460 -9420 42505 -9300
rect 42625 -9420 42670 -9300
rect 42790 -9420 42845 -9300
rect 42965 -9420 43010 -9300
rect 43130 -9420 43175 -9300
rect 43295 -9420 43340 -9300
rect 43460 -9420 43515 -9300
rect 43635 -9420 43680 -9300
rect 43800 -9420 43845 -9300
rect 43965 -9420 44010 -9300
rect 44130 -9420 44185 -9300
rect 44305 -9420 44350 -9300
rect 44470 -9420 44515 -9300
rect 44635 -9420 44680 -9300
rect 44800 -9420 44855 -9300
rect 44975 -9420 45020 -9300
rect 45140 -9420 45185 -9300
rect 45305 -9420 45350 -9300
rect 45470 -9420 45525 -9300
rect 45645 -9420 45690 -9300
rect 45810 -9420 45855 -9300
rect 45975 -9420 46020 -9300
rect 46140 -9420 46195 -9300
rect 46315 -9420 46360 -9300
rect 46480 -9420 46525 -9300
rect 46645 -9420 46690 -9300
rect 46810 -9420 46865 -9300
rect 46985 -9420 47030 -9300
rect 47150 -9420 47195 -9300
rect 47315 -9420 47360 -9300
rect 47480 -9420 47535 -9300
rect 47655 -9420 47865 -9300
rect 47985 -9420 48030 -9300
rect 48150 -9420 48195 -9300
rect 48315 -9420 48360 -9300
rect 48480 -9420 48535 -9300
rect 48655 -9420 48700 -9300
rect 48820 -9420 48865 -9300
rect 48985 -9420 49030 -9300
rect 49150 -9420 49205 -9300
rect 49325 -9420 49370 -9300
rect 49490 -9420 49535 -9300
rect 49655 -9420 49700 -9300
rect 49820 -9420 49875 -9300
rect 49995 -9420 50040 -9300
rect 50160 -9420 50205 -9300
rect 50325 -9420 50370 -9300
rect 50490 -9420 50545 -9300
rect 50665 -9420 50710 -9300
rect 50830 -9420 50875 -9300
rect 50995 -9420 51040 -9300
rect 51160 -9420 51215 -9300
rect 51335 -9420 51380 -9300
rect 51500 -9420 51545 -9300
rect 51665 -9420 51710 -9300
rect 51830 -9420 51885 -9300
rect 52005 -9420 52050 -9300
rect 52170 -9420 52215 -9300
rect 52335 -9420 52380 -9300
rect 52500 -9420 52555 -9300
rect 52675 -9420 52720 -9300
rect 52840 -9420 52885 -9300
rect 53005 -9420 53050 -9300
rect 53170 -9420 53225 -9300
rect 53345 -9420 53370 -9300
rect 30770 -9465 53370 -9420
rect 30770 -9585 30795 -9465
rect 30915 -9585 30960 -9465
rect 31080 -9585 31125 -9465
rect 31245 -9585 31290 -9465
rect 31410 -9585 31465 -9465
rect 31585 -9585 31630 -9465
rect 31750 -9585 31795 -9465
rect 31915 -9585 31960 -9465
rect 32080 -9585 32135 -9465
rect 32255 -9585 32300 -9465
rect 32420 -9585 32465 -9465
rect 32585 -9585 32630 -9465
rect 32750 -9585 32805 -9465
rect 32925 -9585 32970 -9465
rect 33090 -9585 33135 -9465
rect 33255 -9585 33300 -9465
rect 33420 -9585 33475 -9465
rect 33595 -9585 33640 -9465
rect 33760 -9585 33805 -9465
rect 33925 -9585 33970 -9465
rect 34090 -9585 34145 -9465
rect 34265 -9585 34310 -9465
rect 34430 -9585 34475 -9465
rect 34595 -9585 34640 -9465
rect 34760 -9585 34815 -9465
rect 34935 -9585 34980 -9465
rect 35100 -9585 35145 -9465
rect 35265 -9585 35310 -9465
rect 35430 -9585 35485 -9465
rect 35605 -9585 35650 -9465
rect 35770 -9585 35815 -9465
rect 35935 -9585 35980 -9465
rect 36100 -9585 36155 -9465
rect 36275 -9585 36485 -9465
rect 36605 -9585 36650 -9465
rect 36770 -9585 36815 -9465
rect 36935 -9585 36980 -9465
rect 37100 -9585 37155 -9465
rect 37275 -9585 37320 -9465
rect 37440 -9585 37485 -9465
rect 37605 -9585 37650 -9465
rect 37770 -9585 37825 -9465
rect 37945 -9585 37990 -9465
rect 38110 -9585 38155 -9465
rect 38275 -9585 38320 -9465
rect 38440 -9585 38495 -9465
rect 38615 -9585 38660 -9465
rect 38780 -9585 38825 -9465
rect 38945 -9585 38990 -9465
rect 39110 -9585 39165 -9465
rect 39285 -9585 39330 -9465
rect 39450 -9585 39495 -9465
rect 39615 -9585 39660 -9465
rect 39780 -9585 39835 -9465
rect 39955 -9585 40000 -9465
rect 40120 -9585 40165 -9465
rect 40285 -9585 40330 -9465
rect 40450 -9585 40505 -9465
rect 40625 -9585 40670 -9465
rect 40790 -9585 40835 -9465
rect 40955 -9585 41000 -9465
rect 41120 -9585 41175 -9465
rect 41295 -9585 41340 -9465
rect 41460 -9585 41505 -9465
rect 41625 -9585 41670 -9465
rect 41790 -9585 41845 -9465
rect 41965 -9585 42175 -9465
rect 42295 -9585 42340 -9465
rect 42460 -9585 42505 -9465
rect 42625 -9585 42670 -9465
rect 42790 -9585 42845 -9465
rect 42965 -9585 43010 -9465
rect 43130 -9585 43175 -9465
rect 43295 -9585 43340 -9465
rect 43460 -9585 43515 -9465
rect 43635 -9585 43680 -9465
rect 43800 -9585 43845 -9465
rect 43965 -9585 44010 -9465
rect 44130 -9585 44185 -9465
rect 44305 -9585 44350 -9465
rect 44470 -9585 44515 -9465
rect 44635 -9585 44680 -9465
rect 44800 -9585 44855 -9465
rect 44975 -9585 45020 -9465
rect 45140 -9585 45185 -9465
rect 45305 -9585 45350 -9465
rect 45470 -9585 45525 -9465
rect 45645 -9585 45690 -9465
rect 45810 -9585 45855 -9465
rect 45975 -9585 46020 -9465
rect 46140 -9585 46195 -9465
rect 46315 -9585 46360 -9465
rect 46480 -9585 46525 -9465
rect 46645 -9585 46690 -9465
rect 46810 -9585 46865 -9465
rect 46985 -9585 47030 -9465
rect 47150 -9585 47195 -9465
rect 47315 -9585 47360 -9465
rect 47480 -9585 47535 -9465
rect 47655 -9585 47865 -9465
rect 47985 -9585 48030 -9465
rect 48150 -9585 48195 -9465
rect 48315 -9585 48360 -9465
rect 48480 -9585 48535 -9465
rect 48655 -9585 48700 -9465
rect 48820 -9585 48865 -9465
rect 48985 -9585 49030 -9465
rect 49150 -9585 49205 -9465
rect 49325 -9585 49370 -9465
rect 49490 -9585 49535 -9465
rect 49655 -9585 49700 -9465
rect 49820 -9585 49875 -9465
rect 49995 -9585 50040 -9465
rect 50160 -9585 50205 -9465
rect 50325 -9585 50370 -9465
rect 50490 -9585 50545 -9465
rect 50665 -9585 50710 -9465
rect 50830 -9585 50875 -9465
rect 50995 -9585 51040 -9465
rect 51160 -9585 51215 -9465
rect 51335 -9585 51380 -9465
rect 51500 -9585 51545 -9465
rect 51665 -9585 51710 -9465
rect 51830 -9585 51885 -9465
rect 52005 -9585 52050 -9465
rect 52170 -9585 52215 -9465
rect 52335 -9585 52380 -9465
rect 52500 -9585 52555 -9465
rect 52675 -9585 52720 -9465
rect 52840 -9585 52885 -9465
rect 53005 -9585 53050 -9465
rect 53170 -9585 53225 -9465
rect 53345 -9585 53370 -9465
rect 30770 -9630 53370 -9585
rect 30770 -9750 30795 -9630
rect 30915 -9750 30960 -9630
rect 31080 -9750 31125 -9630
rect 31245 -9750 31290 -9630
rect 31410 -9750 31465 -9630
rect 31585 -9750 31630 -9630
rect 31750 -9750 31795 -9630
rect 31915 -9750 31960 -9630
rect 32080 -9750 32135 -9630
rect 32255 -9750 32300 -9630
rect 32420 -9750 32465 -9630
rect 32585 -9750 32630 -9630
rect 32750 -9750 32805 -9630
rect 32925 -9750 32970 -9630
rect 33090 -9750 33135 -9630
rect 33255 -9750 33300 -9630
rect 33420 -9750 33475 -9630
rect 33595 -9750 33640 -9630
rect 33760 -9750 33805 -9630
rect 33925 -9750 33970 -9630
rect 34090 -9750 34145 -9630
rect 34265 -9750 34310 -9630
rect 34430 -9750 34475 -9630
rect 34595 -9750 34640 -9630
rect 34760 -9750 34815 -9630
rect 34935 -9750 34980 -9630
rect 35100 -9750 35145 -9630
rect 35265 -9750 35310 -9630
rect 35430 -9750 35485 -9630
rect 35605 -9750 35650 -9630
rect 35770 -9750 35815 -9630
rect 35935 -9750 35980 -9630
rect 36100 -9750 36155 -9630
rect 36275 -9750 36485 -9630
rect 36605 -9750 36650 -9630
rect 36770 -9750 36815 -9630
rect 36935 -9750 36980 -9630
rect 37100 -9750 37155 -9630
rect 37275 -9750 37320 -9630
rect 37440 -9750 37485 -9630
rect 37605 -9750 37650 -9630
rect 37770 -9750 37825 -9630
rect 37945 -9750 37990 -9630
rect 38110 -9750 38155 -9630
rect 38275 -9750 38320 -9630
rect 38440 -9750 38495 -9630
rect 38615 -9750 38660 -9630
rect 38780 -9750 38825 -9630
rect 38945 -9750 38990 -9630
rect 39110 -9750 39165 -9630
rect 39285 -9750 39330 -9630
rect 39450 -9750 39495 -9630
rect 39615 -9750 39660 -9630
rect 39780 -9750 39835 -9630
rect 39955 -9750 40000 -9630
rect 40120 -9750 40165 -9630
rect 40285 -9750 40330 -9630
rect 40450 -9750 40505 -9630
rect 40625 -9750 40670 -9630
rect 40790 -9750 40835 -9630
rect 40955 -9750 41000 -9630
rect 41120 -9750 41175 -9630
rect 41295 -9750 41340 -9630
rect 41460 -9750 41505 -9630
rect 41625 -9750 41670 -9630
rect 41790 -9750 41845 -9630
rect 41965 -9750 42175 -9630
rect 42295 -9750 42340 -9630
rect 42460 -9750 42505 -9630
rect 42625 -9750 42670 -9630
rect 42790 -9750 42845 -9630
rect 42965 -9750 43010 -9630
rect 43130 -9750 43175 -9630
rect 43295 -9750 43340 -9630
rect 43460 -9750 43515 -9630
rect 43635 -9750 43680 -9630
rect 43800 -9750 43845 -9630
rect 43965 -9750 44010 -9630
rect 44130 -9750 44185 -9630
rect 44305 -9750 44350 -9630
rect 44470 -9750 44515 -9630
rect 44635 -9750 44680 -9630
rect 44800 -9750 44855 -9630
rect 44975 -9750 45020 -9630
rect 45140 -9750 45185 -9630
rect 45305 -9750 45350 -9630
rect 45470 -9750 45525 -9630
rect 45645 -9750 45690 -9630
rect 45810 -9750 45855 -9630
rect 45975 -9750 46020 -9630
rect 46140 -9750 46195 -9630
rect 46315 -9750 46360 -9630
rect 46480 -9750 46525 -9630
rect 46645 -9750 46690 -9630
rect 46810 -9750 46865 -9630
rect 46985 -9750 47030 -9630
rect 47150 -9750 47195 -9630
rect 47315 -9750 47360 -9630
rect 47480 -9750 47535 -9630
rect 47655 -9750 47865 -9630
rect 47985 -9750 48030 -9630
rect 48150 -9750 48195 -9630
rect 48315 -9750 48360 -9630
rect 48480 -9750 48535 -9630
rect 48655 -9750 48700 -9630
rect 48820 -9750 48865 -9630
rect 48985 -9750 49030 -9630
rect 49150 -9750 49205 -9630
rect 49325 -9750 49370 -9630
rect 49490 -9750 49535 -9630
rect 49655 -9750 49700 -9630
rect 49820 -9750 49875 -9630
rect 49995 -9750 50040 -9630
rect 50160 -9750 50205 -9630
rect 50325 -9750 50370 -9630
rect 50490 -9750 50545 -9630
rect 50665 -9750 50710 -9630
rect 50830 -9750 50875 -9630
rect 50995 -9750 51040 -9630
rect 51160 -9750 51215 -9630
rect 51335 -9750 51380 -9630
rect 51500 -9750 51545 -9630
rect 51665 -9750 51710 -9630
rect 51830 -9750 51885 -9630
rect 52005 -9750 52050 -9630
rect 52170 -9750 52215 -9630
rect 52335 -9750 52380 -9630
rect 52500 -9750 52555 -9630
rect 52675 -9750 52720 -9630
rect 52840 -9750 52885 -9630
rect 53005 -9750 53050 -9630
rect 53170 -9750 53225 -9630
rect 53345 -9750 53370 -9630
rect 30770 -9775 53370 -9750
rect 36300 -9825 36460 -9820
rect 41990 -9825 42150 -9820
rect 47680 -9825 47840 -9820
rect 30770 -9840 53370 -9825
rect 30770 -9960 30835 -9840
rect 30955 -9960 31000 -9840
rect 31120 -9960 31165 -9840
rect 31285 -9960 31330 -9840
rect 31450 -9960 31495 -9840
rect 31615 -9960 31660 -9840
rect 31780 -9960 31825 -9840
rect 31945 -9960 31990 -9840
rect 32110 -9960 32155 -9840
rect 32275 -9960 32320 -9840
rect 32440 -9960 32485 -9840
rect 32605 -9960 32650 -9840
rect 32770 -9960 32815 -9840
rect 32935 -9960 32980 -9840
rect 33100 -9960 33145 -9840
rect 33265 -9960 33310 -9840
rect 33430 -9960 33475 -9840
rect 33595 -9960 33640 -9840
rect 33760 -9960 33805 -9840
rect 33925 -9960 33970 -9840
rect 34090 -9960 34135 -9840
rect 34255 -9960 34300 -9840
rect 34420 -9960 34465 -9840
rect 34585 -9960 34630 -9840
rect 34750 -9960 34795 -9840
rect 34915 -9960 34960 -9840
rect 35080 -9960 35125 -9840
rect 35245 -9960 35290 -9840
rect 35410 -9960 35455 -9840
rect 35575 -9960 35620 -9840
rect 35740 -9960 35785 -9840
rect 35905 -9960 35950 -9840
rect 36070 -9960 36115 -9840
rect 36235 -9960 36525 -9840
rect 36645 -9960 36690 -9840
rect 36810 -9960 36855 -9840
rect 36975 -9960 37020 -9840
rect 37140 -9960 37185 -9840
rect 37305 -9960 37350 -9840
rect 37470 -9960 37515 -9840
rect 37635 -9960 37680 -9840
rect 37800 -9960 37845 -9840
rect 37965 -9960 38010 -9840
rect 38130 -9960 38175 -9840
rect 38295 -9960 38340 -9840
rect 38460 -9960 38505 -9840
rect 38625 -9960 38670 -9840
rect 38790 -9960 38835 -9840
rect 38955 -9960 39000 -9840
rect 39120 -9960 39165 -9840
rect 39285 -9960 39330 -9840
rect 39450 -9960 39495 -9840
rect 39615 -9960 39660 -9840
rect 39780 -9960 39825 -9840
rect 39945 -9960 39990 -9840
rect 40110 -9960 40155 -9840
rect 40275 -9960 40320 -9840
rect 40440 -9960 40485 -9840
rect 40605 -9960 40650 -9840
rect 40770 -9960 40815 -9840
rect 40935 -9960 40980 -9840
rect 41100 -9960 41145 -9840
rect 41265 -9960 41310 -9840
rect 41430 -9960 41475 -9840
rect 41595 -9960 41640 -9840
rect 41760 -9960 41805 -9840
rect 41925 -9960 42215 -9840
rect 42335 -9960 42380 -9840
rect 42500 -9960 42545 -9840
rect 42665 -9960 42710 -9840
rect 42830 -9960 42875 -9840
rect 42995 -9960 43040 -9840
rect 43160 -9960 43205 -9840
rect 43325 -9960 43370 -9840
rect 43490 -9960 43535 -9840
rect 43655 -9960 43700 -9840
rect 43820 -9960 43865 -9840
rect 43985 -9960 44030 -9840
rect 44150 -9960 44195 -9840
rect 44315 -9960 44360 -9840
rect 44480 -9960 44525 -9840
rect 44645 -9960 44690 -9840
rect 44810 -9960 44855 -9840
rect 44975 -9960 45020 -9840
rect 45140 -9960 45185 -9840
rect 45305 -9960 45350 -9840
rect 45470 -9960 45515 -9840
rect 45635 -9960 45680 -9840
rect 45800 -9960 45845 -9840
rect 45965 -9960 46010 -9840
rect 46130 -9960 46175 -9840
rect 46295 -9960 46340 -9840
rect 46460 -9960 46505 -9840
rect 46625 -9960 46670 -9840
rect 46790 -9960 46835 -9840
rect 46955 -9960 47000 -9840
rect 47120 -9960 47165 -9840
rect 47285 -9960 47330 -9840
rect 47450 -9960 47495 -9840
rect 47615 -9960 47905 -9840
rect 48025 -9960 48070 -9840
rect 48190 -9960 48235 -9840
rect 48355 -9960 48400 -9840
rect 48520 -9960 48565 -9840
rect 48685 -9960 48730 -9840
rect 48850 -9960 48895 -9840
rect 49015 -9960 49060 -9840
rect 49180 -9960 49225 -9840
rect 49345 -9960 49390 -9840
rect 49510 -9960 49555 -9840
rect 49675 -9960 49720 -9840
rect 49840 -9960 49885 -9840
rect 50005 -9960 50050 -9840
rect 50170 -9960 50215 -9840
rect 50335 -9960 50380 -9840
rect 50500 -9960 50545 -9840
rect 50665 -9960 50710 -9840
rect 50830 -9960 50875 -9840
rect 50995 -9960 51040 -9840
rect 51160 -9960 51205 -9840
rect 51325 -9960 51370 -9840
rect 51490 -9960 51535 -9840
rect 51655 -9960 51700 -9840
rect 51820 -9960 51865 -9840
rect 51985 -9960 52030 -9840
rect 52150 -9960 52195 -9840
rect 52315 -9960 52360 -9840
rect 52480 -9960 52525 -9840
rect 52645 -9960 52690 -9840
rect 52810 -9960 52855 -9840
rect 52975 -9960 53020 -9840
rect 53140 -9960 53185 -9840
rect 53305 -9960 53370 -9840
rect 30770 -9975 53370 -9960
rect 36300 -9980 36460 -9975
rect 41990 -9980 42150 -9975
rect 47680 -9980 47840 -9975
rect 30770 -10050 53370 -10025
rect 30770 -10170 30795 -10050
rect 30915 -10170 30970 -10050
rect 31090 -10170 31135 -10050
rect 31255 -10170 31300 -10050
rect 31420 -10170 31465 -10050
rect 31585 -10170 31640 -10050
rect 31760 -10170 31805 -10050
rect 31925 -10170 31970 -10050
rect 32090 -10170 32135 -10050
rect 32255 -10170 32310 -10050
rect 32430 -10170 32475 -10050
rect 32595 -10170 32640 -10050
rect 32760 -10170 32805 -10050
rect 32925 -10170 32980 -10050
rect 33100 -10170 33145 -10050
rect 33265 -10170 33310 -10050
rect 33430 -10170 33475 -10050
rect 33595 -10170 33650 -10050
rect 33770 -10170 33815 -10050
rect 33935 -10170 33980 -10050
rect 34100 -10170 34145 -10050
rect 34265 -10170 34320 -10050
rect 34440 -10170 34485 -10050
rect 34605 -10170 34650 -10050
rect 34770 -10170 34815 -10050
rect 34935 -10170 34990 -10050
rect 35110 -10170 35155 -10050
rect 35275 -10170 35320 -10050
rect 35440 -10170 35485 -10050
rect 35605 -10170 35660 -10050
rect 35780 -10170 35825 -10050
rect 35945 -10170 35990 -10050
rect 36110 -10170 36155 -10050
rect 36275 -10170 36485 -10050
rect 36605 -10170 36660 -10050
rect 36780 -10170 36825 -10050
rect 36945 -10170 36990 -10050
rect 37110 -10170 37155 -10050
rect 37275 -10170 37330 -10050
rect 37450 -10170 37495 -10050
rect 37615 -10170 37660 -10050
rect 37780 -10170 37825 -10050
rect 37945 -10170 38000 -10050
rect 38120 -10170 38165 -10050
rect 38285 -10170 38330 -10050
rect 38450 -10170 38495 -10050
rect 38615 -10170 38670 -10050
rect 38790 -10170 38835 -10050
rect 38955 -10170 39000 -10050
rect 39120 -10170 39165 -10050
rect 39285 -10170 39340 -10050
rect 39460 -10170 39505 -10050
rect 39625 -10170 39670 -10050
rect 39790 -10170 39835 -10050
rect 39955 -10170 40010 -10050
rect 40130 -10170 40175 -10050
rect 40295 -10170 40340 -10050
rect 40460 -10170 40505 -10050
rect 40625 -10170 40680 -10050
rect 40800 -10170 40845 -10050
rect 40965 -10170 41010 -10050
rect 41130 -10170 41175 -10050
rect 41295 -10170 41350 -10050
rect 41470 -10170 41515 -10050
rect 41635 -10170 41680 -10050
rect 41800 -10170 41845 -10050
rect 41965 -10170 42175 -10050
rect 42295 -10170 42350 -10050
rect 42470 -10170 42515 -10050
rect 42635 -10170 42680 -10050
rect 42800 -10170 42845 -10050
rect 42965 -10170 43020 -10050
rect 43140 -10170 43185 -10050
rect 43305 -10170 43350 -10050
rect 43470 -10170 43515 -10050
rect 43635 -10170 43690 -10050
rect 43810 -10170 43855 -10050
rect 43975 -10170 44020 -10050
rect 44140 -10170 44185 -10050
rect 44305 -10170 44360 -10050
rect 44480 -10170 44525 -10050
rect 44645 -10170 44690 -10050
rect 44810 -10170 44855 -10050
rect 44975 -10170 45030 -10050
rect 45150 -10170 45195 -10050
rect 45315 -10170 45360 -10050
rect 45480 -10170 45525 -10050
rect 45645 -10170 45700 -10050
rect 45820 -10170 45865 -10050
rect 45985 -10170 46030 -10050
rect 46150 -10170 46195 -10050
rect 46315 -10170 46370 -10050
rect 46490 -10170 46535 -10050
rect 46655 -10170 46700 -10050
rect 46820 -10170 46865 -10050
rect 46985 -10170 47040 -10050
rect 47160 -10170 47205 -10050
rect 47325 -10170 47370 -10050
rect 47490 -10170 47535 -10050
rect 47655 -10170 47865 -10050
rect 47985 -10170 48040 -10050
rect 48160 -10170 48205 -10050
rect 48325 -10170 48370 -10050
rect 48490 -10170 48535 -10050
rect 48655 -10170 48710 -10050
rect 48830 -10170 48875 -10050
rect 48995 -10170 49040 -10050
rect 49160 -10170 49205 -10050
rect 49325 -10170 49380 -10050
rect 49500 -10170 49545 -10050
rect 49665 -10170 49710 -10050
rect 49830 -10170 49875 -10050
rect 49995 -10170 50050 -10050
rect 50170 -10170 50215 -10050
rect 50335 -10170 50380 -10050
rect 50500 -10170 50545 -10050
rect 50665 -10170 50720 -10050
rect 50840 -10170 50885 -10050
rect 51005 -10170 51050 -10050
rect 51170 -10170 51215 -10050
rect 51335 -10170 51390 -10050
rect 51510 -10170 51555 -10050
rect 51675 -10170 51720 -10050
rect 51840 -10170 51885 -10050
rect 52005 -10170 52060 -10050
rect 52180 -10170 52225 -10050
rect 52345 -10170 52390 -10050
rect 52510 -10170 52555 -10050
rect 52675 -10170 52730 -10050
rect 52850 -10170 52895 -10050
rect 53015 -10170 53060 -10050
rect 53180 -10170 53225 -10050
rect 53345 -10170 53370 -10050
rect 30770 -10215 53370 -10170
rect 30770 -10335 30795 -10215
rect 30915 -10335 30970 -10215
rect 31090 -10335 31135 -10215
rect 31255 -10335 31300 -10215
rect 31420 -10335 31465 -10215
rect 31585 -10335 31640 -10215
rect 31760 -10335 31805 -10215
rect 31925 -10335 31970 -10215
rect 32090 -10335 32135 -10215
rect 32255 -10335 32310 -10215
rect 32430 -10335 32475 -10215
rect 32595 -10335 32640 -10215
rect 32760 -10335 32805 -10215
rect 32925 -10335 32980 -10215
rect 33100 -10335 33145 -10215
rect 33265 -10335 33310 -10215
rect 33430 -10335 33475 -10215
rect 33595 -10335 33650 -10215
rect 33770 -10335 33815 -10215
rect 33935 -10335 33980 -10215
rect 34100 -10335 34145 -10215
rect 34265 -10335 34320 -10215
rect 34440 -10335 34485 -10215
rect 34605 -10335 34650 -10215
rect 34770 -10335 34815 -10215
rect 34935 -10335 34990 -10215
rect 35110 -10335 35155 -10215
rect 35275 -10335 35320 -10215
rect 35440 -10335 35485 -10215
rect 35605 -10335 35660 -10215
rect 35780 -10335 35825 -10215
rect 35945 -10335 35990 -10215
rect 36110 -10335 36155 -10215
rect 36275 -10335 36485 -10215
rect 36605 -10335 36660 -10215
rect 36780 -10335 36825 -10215
rect 36945 -10335 36990 -10215
rect 37110 -10335 37155 -10215
rect 37275 -10335 37330 -10215
rect 37450 -10335 37495 -10215
rect 37615 -10335 37660 -10215
rect 37780 -10335 37825 -10215
rect 37945 -10335 38000 -10215
rect 38120 -10335 38165 -10215
rect 38285 -10335 38330 -10215
rect 38450 -10335 38495 -10215
rect 38615 -10335 38670 -10215
rect 38790 -10335 38835 -10215
rect 38955 -10335 39000 -10215
rect 39120 -10335 39165 -10215
rect 39285 -10335 39340 -10215
rect 39460 -10335 39505 -10215
rect 39625 -10335 39670 -10215
rect 39790 -10335 39835 -10215
rect 39955 -10335 40010 -10215
rect 40130 -10335 40175 -10215
rect 40295 -10335 40340 -10215
rect 40460 -10335 40505 -10215
rect 40625 -10335 40680 -10215
rect 40800 -10335 40845 -10215
rect 40965 -10335 41010 -10215
rect 41130 -10335 41175 -10215
rect 41295 -10335 41350 -10215
rect 41470 -10335 41515 -10215
rect 41635 -10335 41680 -10215
rect 41800 -10335 41845 -10215
rect 41965 -10335 42175 -10215
rect 42295 -10335 42350 -10215
rect 42470 -10335 42515 -10215
rect 42635 -10335 42680 -10215
rect 42800 -10335 42845 -10215
rect 42965 -10335 43020 -10215
rect 43140 -10335 43185 -10215
rect 43305 -10335 43350 -10215
rect 43470 -10335 43515 -10215
rect 43635 -10335 43690 -10215
rect 43810 -10335 43855 -10215
rect 43975 -10335 44020 -10215
rect 44140 -10335 44185 -10215
rect 44305 -10335 44360 -10215
rect 44480 -10335 44525 -10215
rect 44645 -10335 44690 -10215
rect 44810 -10335 44855 -10215
rect 44975 -10335 45030 -10215
rect 45150 -10335 45195 -10215
rect 45315 -10335 45360 -10215
rect 45480 -10335 45525 -10215
rect 45645 -10335 45700 -10215
rect 45820 -10335 45865 -10215
rect 45985 -10335 46030 -10215
rect 46150 -10335 46195 -10215
rect 46315 -10335 46370 -10215
rect 46490 -10335 46535 -10215
rect 46655 -10335 46700 -10215
rect 46820 -10335 46865 -10215
rect 46985 -10335 47040 -10215
rect 47160 -10335 47205 -10215
rect 47325 -10335 47370 -10215
rect 47490 -10335 47535 -10215
rect 47655 -10335 47865 -10215
rect 47985 -10335 48040 -10215
rect 48160 -10335 48205 -10215
rect 48325 -10335 48370 -10215
rect 48490 -10335 48535 -10215
rect 48655 -10335 48710 -10215
rect 48830 -10335 48875 -10215
rect 48995 -10335 49040 -10215
rect 49160 -10335 49205 -10215
rect 49325 -10335 49380 -10215
rect 49500 -10335 49545 -10215
rect 49665 -10335 49710 -10215
rect 49830 -10335 49875 -10215
rect 49995 -10335 50050 -10215
rect 50170 -10335 50215 -10215
rect 50335 -10335 50380 -10215
rect 50500 -10335 50545 -10215
rect 50665 -10335 50720 -10215
rect 50840 -10335 50885 -10215
rect 51005 -10335 51050 -10215
rect 51170 -10335 51215 -10215
rect 51335 -10335 51390 -10215
rect 51510 -10335 51555 -10215
rect 51675 -10335 51720 -10215
rect 51840 -10335 51885 -10215
rect 52005 -10335 52060 -10215
rect 52180 -10335 52225 -10215
rect 52345 -10335 52390 -10215
rect 52510 -10335 52555 -10215
rect 52675 -10335 52730 -10215
rect 52850 -10335 52895 -10215
rect 53015 -10335 53060 -10215
rect 53180 -10335 53225 -10215
rect 53345 -10335 53370 -10215
rect 30770 -10380 53370 -10335
rect 30770 -10500 30795 -10380
rect 30915 -10500 30970 -10380
rect 31090 -10500 31135 -10380
rect 31255 -10500 31300 -10380
rect 31420 -10500 31465 -10380
rect 31585 -10500 31640 -10380
rect 31760 -10500 31805 -10380
rect 31925 -10500 31970 -10380
rect 32090 -10500 32135 -10380
rect 32255 -10500 32310 -10380
rect 32430 -10500 32475 -10380
rect 32595 -10500 32640 -10380
rect 32760 -10500 32805 -10380
rect 32925 -10500 32980 -10380
rect 33100 -10500 33145 -10380
rect 33265 -10500 33310 -10380
rect 33430 -10500 33475 -10380
rect 33595 -10500 33650 -10380
rect 33770 -10500 33815 -10380
rect 33935 -10500 33980 -10380
rect 34100 -10500 34145 -10380
rect 34265 -10500 34320 -10380
rect 34440 -10500 34485 -10380
rect 34605 -10500 34650 -10380
rect 34770 -10500 34815 -10380
rect 34935 -10500 34990 -10380
rect 35110 -10500 35155 -10380
rect 35275 -10500 35320 -10380
rect 35440 -10500 35485 -10380
rect 35605 -10500 35660 -10380
rect 35780 -10500 35825 -10380
rect 35945 -10500 35990 -10380
rect 36110 -10500 36155 -10380
rect 36275 -10500 36485 -10380
rect 36605 -10500 36660 -10380
rect 36780 -10500 36825 -10380
rect 36945 -10500 36990 -10380
rect 37110 -10500 37155 -10380
rect 37275 -10500 37330 -10380
rect 37450 -10500 37495 -10380
rect 37615 -10500 37660 -10380
rect 37780 -10500 37825 -10380
rect 37945 -10500 38000 -10380
rect 38120 -10500 38165 -10380
rect 38285 -10500 38330 -10380
rect 38450 -10500 38495 -10380
rect 38615 -10500 38670 -10380
rect 38790 -10500 38835 -10380
rect 38955 -10500 39000 -10380
rect 39120 -10500 39165 -10380
rect 39285 -10500 39340 -10380
rect 39460 -10500 39505 -10380
rect 39625 -10500 39670 -10380
rect 39790 -10500 39835 -10380
rect 39955 -10500 40010 -10380
rect 40130 -10500 40175 -10380
rect 40295 -10500 40340 -10380
rect 40460 -10500 40505 -10380
rect 40625 -10500 40680 -10380
rect 40800 -10500 40845 -10380
rect 40965 -10500 41010 -10380
rect 41130 -10500 41175 -10380
rect 41295 -10500 41350 -10380
rect 41470 -10500 41515 -10380
rect 41635 -10500 41680 -10380
rect 41800 -10500 41845 -10380
rect 41965 -10500 42175 -10380
rect 42295 -10500 42350 -10380
rect 42470 -10500 42515 -10380
rect 42635 -10500 42680 -10380
rect 42800 -10500 42845 -10380
rect 42965 -10500 43020 -10380
rect 43140 -10500 43185 -10380
rect 43305 -10500 43350 -10380
rect 43470 -10500 43515 -10380
rect 43635 -10500 43690 -10380
rect 43810 -10500 43855 -10380
rect 43975 -10500 44020 -10380
rect 44140 -10500 44185 -10380
rect 44305 -10500 44360 -10380
rect 44480 -10500 44525 -10380
rect 44645 -10500 44690 -10380
rect 44810 -10500 44855 -10380
rect 44975 -10500 45030 -10380
rect 45150 -10500 45195 -10380
rect 45315 -10500 45360 -10380
rect 45480 -10500 45525 -10380
rect 45645 -10500 45700 -10380
rect 45820 -10500 45865 -10380
rect 45985 -10500 46030 -10380
rect 46150 -10500 46195 -10380
rect 46315 -10500 46370 -10380
rect 46490 -10500 46535 -10380
rect 46655 -10500 46700 -10380
rect 46820 -10500 46865 -10380
rect 46985 -10500 47040 -10380
rect 47160 -10500 47205 -10380
rect 47325 -10500 47370 -10380
rect 47490 -10500 47535 -10380
rect 47655 -10500 47865 -10380
rect 47985 -10500 48040 -10380
rect 48160 -10500 48205 -10380
rect 48325 -10500 48370 -10380
rect 48490 -10500 48535 -10380
rect 48655 -10500 48710 -10380
rect 48830 -10500 48875 -10380
rect 48995 -10500 49040 -10380
rect 49160 -10500 49205 -10380
rect 49325 -10500 49380 -10380
rect 49500 -10500 49545 -10380
rect 49665 -10500 49710 -10380
rect 49830 -10500 49875 -10380
rect 49995 -10500 50050 -10380
rect 50170 -10500 50215 -10380
rect 50335 -10500 50380 -10380
rect 50500 -10500 50545 -10380
rect 50665 -10500 50720 -10380
rect 50840 -10500 50885 -10380
rect 51005 -10500 51050 -10380
rect 51170 -10500 51215 -10380
rect 51335 -10500 51390 -10380
rect 51510 -10500 51555 -10380
rect 51675 -10500 51720 -10380
rect 51840 -10500 51885 -10380
rect 52005 -10500 52060 -10380
rect 52180 -10500 52225 -10380
rect 52345 -10500 52390 -10380
rect 52510 -10500 52555 -10380
rect 52675 -10500 52730 -10380
rect 52850 -10500 52895 -10380
rect 53015 -10500 53060 -10380
rect 53180 -10500 53225 -10380
rect 53345 -10500 53370 -10380
rect 30770 -10545 53370 -10500
rect 30770 -10665 30795 -10545
rect 30915 -10665 30970 -10545
rect 31090 -10665 31135 -10545
rect 31255 -10665 31300 -10545
rect 31420 -10665 31465 -10545
rect 31585 -10665 31640 -10545
rect 31760 -10665 31805 -10545
rect 31925 -10665 31970 -10545
rect 32090 -10665 32135 -10545
rect 32255 -10665 32310 -10545
rect 32430 -10665 32475 -10545
rect 32595 -10665 32640 -10545
rect 32760 -10665 32805 -10545
rect 32925 -10665 32980 -10545
rect 33100 -10665 33145 -10545
rect 33265 -10665 33310 -10545
rect 33430 -10665 33475 -10545
rect 33595 -10665 33650 -10545
rect 33770 -10665 33815 -10545
rect 33935 -10665 33980 -10545
rect 34100 -10665 34145 -10545
rect 34265 -10665 34320 -10545
rect 34440 -10665 34485 -10545
rect 34605 -10665 34650 -10545
rect 34770 -10665 34815 -10545
rect 34935 -10665 34990 -10545
rect 35110 -10665 35155 -10545
rect 35275 -10665 35320 -10545
rect 35440 -10665 35485 -10545
rect 35605 -10665 35660 -10545
rect 35780 -10665 35825 -10545
rect 35945 -10665 35990 -10545
rect 36110 -10665 36155 -10545
rect 36275 -10665 36485 -10545
rect 36605 -10665 36660 -10545
rect 36780 -10665 36825 -10545
rect 36945 -10665 36990 -10545
rect 37110 -10665 37155 -10545
rect 37275 -10665 37330 -10545
rect 37450 -10665 37495 -10545
rect 37615 -10665 37660 -10545
rect 37780 -10665 37825 -10545
rect 37945 -10665 38000 -10545
rect 38120 -10665 38165 -10545
rect 38285 -10665 38330 -10545
rect 38450 -10665 38495 -10545
rect 38615 -10665 38670 -10545
rect 38790 -10665 38835 -10545
rect 38955 -10665 39000 -10545
rect 39120 -10665 39165 -10545
rect 39285 -10665 39340 -10545
rect 39460 -10665 39505 -10545
rect 39625 -10665 39670 -10545
rect 39790 -10665 39835 -10545
rect 39955 -10665 40010 -10545
rect 40130 -10665 40175 -10545
rect 40295 -10665 40340 -10545
rect 40460 -10665 40505 -10545
rect 40625 -10665 40680 -10545
rect 40800 -10665 40845 -10545
rect 40965 -10665 41010 -10545
rect 41130 -10665 41175 -10545
rect 41295 -10665 41350 -10545
rect 41470 -10665 41515 -10545
rect 41635 -10665 41680 -10545
rect 41800 -10665 41845 -10545
rect 41965 -10665 42175 -10545
rect 42295 -10665 42350 -10545
rect 42470 -10665 42515 -10545
rect 42635 -10665 42680 -10545
rect 42800 -10665 42845 -10545
rect 42965 -10665 43020 -10545
rect 43140 -10665 43185 -10545
rect 43305 -10665 43350 -10545
rect 43470 -10665 43515 -10545
rect 43635 -10665 43690 -10545
rect 43810 -10665 43855 -10545
rect 43975 -10665 44020 -10545
rect 44140 -10665 44185 -10545
rect 44305 -10665 44360 -10545
rect 44480 -10665 44525 -10545
rect 44645 -10665 44690 -10545
rect 44810 -10665 44855 -10545
rect 44975 -10665 45030 -10545
rect 45150 -10665 45195 -10545
rect 45315 -10665 45360 -10545
rect 45480 -10665 45525 -10545
rect 45645 -10665 45700 -10545
rect 45820 -10665 45865 -10545
rect 45985 -10665 46030 -10545
rect 46150 -10665 46195 -10545
rect 46315 -10665 46370 -10545
rect 46490 -10665 46535 -10545
rect 46655 -10665 46700 -10545
rect 46820 -10665 46865 -10545
rect 46985 -10665 47040 -10545
rect 47160 -10665 47205 -10545
rect 47325 -10665 47370 -10545
rect 47490 -10665 47535 -10545
rect 47655 -10665 47865 -10545
rect 47985 -10665 48040 -10545
rect 48160 -10665 48205 -10545
rect 48325 -10665 48370 -10545
rect 48490 -10665 48535 -10545
rect 48655 -10665 48710 -10545
rect 48830 -10665 48875 -10545
rect 48995 -10665 49040 -10545
rect 49160 -10665 49205 -10545
rect 49325 -10665 49380 -10545
rect 49500 -10665 49545 -10545
rect 49665 -10665 49710 -10545
rect 49830 -10665 49875 -10545
rect 49995 -10665 50050 -10545
rect 50170 -10665 50215 -10545
rect 50335 -10665 50380 -10545
rect 50500 -10665 50545 -10545
rect 50665 -10665 50720 -10545
rect 50840 -10665 50885 -10545
rect 51005 -10665 51050 -10545
rect 51170 -10665 51215 -10545
rect 51335 -10665 51390 -10545
rect 51510 -10665 51555 -10545
rect 51675 -10665 51720 -10545
rect 51840 -10665 51885 -10545
rect 52005 -10665 52060 -10545
rect 52180 -10665 52225 -10545
rect 52345 -10665 52390 -10545
rect 52510 -10665 52555 -10545
rect 52675 -10665 52730 -10545
rect 52850 -10665 52895 -10545
rect 53015 -10665 53060 -10545
rect 53180 -10665 53225 -10545
rect 53345 -10665 53370 -10545
rect 30770 -10720 53370 -10665
rect 30770 -10840 30795 -10720
rect 30915 -10840 30970 -10720
rect 31090 -10840 31135 -10720
rect 31255 -10840 31300 -10720
rect 31420 -10840 31465 -10720
rect 31585 -10840 31640 -10720
rect 31760 -10840 31805 -10720
rect 31925 -10840 31970 -10720
rect 32090 -10840 32135 -10720
rect 32255 -10840 32310 -10720
rect 32430 -10840 32475 -10720
rect 32595 -10840 32640 -10720
rect 32760 -10840 32805 -10720
rect 32925 -10840 32980 -10720
rect 33100 -10840 33145 -10720
rect 33265 -10840 33310 -10720
rect 33430 -10840 33475 -10720
rect 33595 -10840 33650 -10720
rect 33770 -10840 33815 -10720
rect 33935 -10840 33980 -10720
rect 34100 -10840 34145 -10720
rect 34265 -10840 34320 -10720
rect 34440 -10840 34485 -10720
rect 34605 -10840 34650 -10720
rect 34770 -10840 34815 -10720
rect 34935 -10840 34990 -10720
rect 35110 -10840 35155 -10720
rect 35275 -10840 35320 -10720
rect 35440 -10840 35485 -10720
rect 35605 -10840 35660 -10720
rect 35780 -10840 35825 -10720
rect 35945 -10840 35990 -10720
rect 36110 -10840 36155 -10720
rect 36275 -10840 36485 -10720
rect 36605 -10840 36660 -10720
rect 36780 -10840 36825 -10720
rect 36945 -10840 36990 -10720
rect 37110 -10840 37155 -10720
rect 37275 -10840 37330 -10720
rect 37450 -10840 37495 -10720
rect 37615 -10840 37660 -10720
rect 37780 -10840 37825 -10720
rect 37945 -10840 38000 -10720
rect 38120 -10840 38165 -10720
rect 38285 -10840 38330 -10720
rect 38450 -10840 38495 -10720
rect 38615 -10840 38670 -10720
rect 38790 -10840 38835 -10720
rect 38955 -10840 39000 -10720
rect 39120 -10840 39165 -10720
rect 39285 -10840 39340 -10720
rect 39460 -10840 39505 -10720
rect 39625 -10840 39670 -10720
rect 39790 -10840 39835 -10720
rect 39955 -10840 40010 -10720
rect 40130 -10840 40175 -10720
rect 40295 -10840 40340 -10720
rect 40460 -10840 40505 -10720
rect 40625 -10840 40680 -10720
rect 40800 -10840 40845 -10720
rect 40965 -10840 41010 -10720
rect 41130 -10840 41175 -10720
rect 41295 -10840 41350 -10720
rect 41470 -10840 41515 -10720
rect 41635 -10840 41680 -10720
rect 41800 -10840 41845 -10720
rect 41965 -10840 42175 -10720
rect 42295 -10840 42350 -10720
rect 42470 -10840 42515 -10720
rect 42635 -10840 42680 -10720
rect 42800 -10840 42845 -10720
rect 42965 -10840 43020 -10720
rect 43140 -10840 43185 -10720
rect 43305 -10840 43350 -10720
rect 43470 -10840 43515 -10720
rect 43635 -10840 43690 -10720
rect 43810 -10840 43855 -10720
rect 43975 -10840 44020 -10720
rect 44140 -10840 44185 -10720
rect 44305 -10840 44360 -10720
rect 44480 -10840 44525 -10720
rect 44645 -10840 44690 -10720
rect 44810 -10840 44855 -10720
rect 44975 -10840 45030 -10720
rect 45150 -10840 45195 -10720
rect 45315 -10840 45360 -10720
rect 45480 -10840 45525 -10720
rect 45645 -10840 45700 -10720
rect 45820 -10840 45865 -10720
rect 45985 -10840 46030 -10720
rect 46150 -10840 46195 -10720
rect 46315 -10840 46370 -10720
rect 46490 -10840 46535 -10720
rect 46655 -10840 46700 -10720
rect 46820 -10840 46865 -10720
rect 46985 -10840 47040 -10720
rect 47160 -10840 47205 -10720
rect 47325 -10840 47370 -10720
rect 47490 -10840 47535 -10720
rect 47655 -10840 47865 -10720
rect 47985 -10840 48040 -10720
rect 48160 -10840 48205 -10720
rect 48325 -10840 48370 -10720
rect 48490 -10840 48535 -10720
rect 48655 -10840 48710 -10720
rect 48830 -10840 48875 -10720
rect 48995 -10840 49040 -10720
rect 49160 -10840 49205 -10720
rect 49325 -10840 49380 -10720
rect 49500 -10840 49545 -10720
rect 49665 -10840 49710 -10720
rect 49830 -10840 49875 -10720
rect 49995 -10840 50050 -10720
rect 50170 -10840 50215 -10720
rect 50335 -10840 50380 -10720
rect 50500 -10840 50545 -10720
rect 50665 -10840 50720 -10720
rect 50840 -10840 50885 -10720
rect 51005 -10840 51050 -10720
rect 51170 -10840 51215 -10720
rect 51335 -10840 51390 -10720
rect 51510 -10840 51555 -10720
rect 51675 -10840 51720 -10720
rect 51840 -10840 51885 -10720
rect 52005 -10840 52060 -10720
rect 52180 -10840 52225 -10720
rect 52345 -10840 52390 -10720
rect 52510 -10840 52555 -10720
rect 52675 -10840 52730 -10720
rect 52850 -10840 52895 -10720
rect 53015 -10840 53060 -10720
rect 53180 -10840 53225 -10720
rect 53345 -10840 53370 -10720
rect 30770 -10885 53370 -10840
rect 30770 -11005 30795 -10885
rect 30915 -11005 30970 -10885
rect 31090 -11005 31135 -10885
rect 31255 -11005 31300 -10885
rect 31420 -11005 31465 -10885
rect 31585 -11005 31640 -10885
rect 31760 -11005 31805 -10885
rect 31925 -11005 31970 -10885
rect 32090 -11005 32135 -10885
rect 32255 -11005 32310 -10885
rect 32430 -11005 32475 -10885
rect 32595 -11005 32640 -10885
rect 32760 -11005 32805 -10885
rect 32925 -11005 32980 -10885
rect 33100 -11005 33145 -10885
rect 33265 -11005 33310 -10885
rect 33430 -11005 33475 -10885
rect 33595 -11005 33650 -10885
rect 33770 -11005 33815 -10885
rect 33935 -11005 33980 -10885
rect 34100 -11005 34145 -10885
rect 34265 -11005 34320 -10885
rect 34440 -11005 34485 -10885
rect 34605 -11005 34650 -10885
rect 34770 -11005 34815 -10885
rect 34935 -11005 34990 -10885
rect 35110 -11005 35155 -10885
rect 35275 -11005 35320 -10885
rect 35440 -11005 35485 -10885
rect 35605 -11005 35660 -10885
rect 35780 -11005 35825 -10885
rect 35945 -11005 35990 -10885
rect 36110 -11005 36155 -10885
rect 36275 -11005 36485 -10885
rect 36605 -11005 36660 -10885
rect 36780 -11005 36825 -10885
rect 36945 -11005 36990 -10885
rect 37110 -11005 37155 -10885
rect 37275 -11005 37330 -10885
rect 37450 -11005 37495 -10885
rect 37615 -11005 37660 -10885
rect 37780 -11005 37825 -10885
rect 37945 -11005 38000 -10885
rect 38120 -11005 38165 -10885
rect 38285 -11005 38330 -10885
rect 38450 -11005 38495 -10885
rect 38615 -11005 38670 -10885
rect 38790 -11005 38835 -10885
rect 38955 -11005 39000 -10885
rect 39120 -11005 39165 -10885
rect 39285 -11005 39340 -10885
rect 39460 -11005 39505 -10885
rect 39625 -11005 39670 -10885
rect 39790 -11005 39835 -10885
rect 39955 -11005 40010 -10885
rect 40130 -11005 40175 -10885
rect 40295 -11005 40340 -10885
rect 40460 -11005 40505 -10885
rect 40625 -11005 40680 -10885
rect 40800 -11005 40845 -10885
rect 40965 -11005 41010 -10885
rect 41130 -11005 41175 -10885
rect 41295 -11005 41350 -10885
rect 41470 -11005 41515 -10885
rect 41635 -11005 41680 -10885
rect 41800 -11005 41845 -10885
rect 41965 -11005 42175 -10885
rect 42295 -11005 42350 -10885
rect 42470 -11005 42515 -10885
rect 42635 -11005 42680 -10885
rect 42800 -11005 42845 -10885
rect 42965 -11005 43020 -10885
rect 43140 -11005 43185 -10885
rect 43305 -11005 43350 -10885
rect 43470 -11005 43515 -10885
rect 43635 -11005 43690 -10885
rect 43810 -11005 43855 -10885
rect 43975 -11005 44020 -10885
rect 44140 -11005 44185 -10885
rect 44305 -11005 44360 -10885
rect 44480 -11005 44525 -10885
rect 44645 -11005 44690 -10885
rect 44810 -11005 44855 -10885
rect 44975 -11005 45030 -10885
rect 45150 -11005 45195 -10885
rect 45315 -11005 45360 -10885
rect 45480 -11005 45525 -10885
rect 45645 -11005 45700 -10885
rect 45820 -11005 45865 -10885
rect 45985 -11005 46030 -10885
rect 46150 -11005 46195 -10885
rect 46315 -11005 46370 -10885
rect 46490 -11005 46535 -10885
rect 46655 -11005 46700 -10885
rect 46820 -11005 46865 -10885
rect 46985 -11005 47040 -10885
rect 47160 -11005 47205 -10885
rect 47325 -11005 47370 -10885
rect 47490 -11005 47535 -10885
rect 47655 -11005 47865 -10885
rect 47985 -11005 48040 -10885
rect 48160 -11005 48205 -10885
rect 48325 -11005 48370 -10885
rect 48490 -11005 48535 -10885
rect 48655 -11005 48710 -10885
rect 48830 -11005 48875 -10885
rect 48995 -11005 49040 -10885
rect 49160 -11005 49205 -10885
rect 49325 -11005 49380 -10885
rect 49500 -11005 49545 -10885
rect 49665 -11005 49710 -10885
rect 49830 -11005 49875 -10885
rect 49995 -11005 50050 -10885
rect 50170 -11005 50215 -10885
rect 50335 -11005 50380 -10885
rect 50500 -11005 50545 -10885
rect 50665 -11005 50720 -10885
rect 50840 -11005 50885 -10885
rect 51005 -11005 51050 -10885
rect 51170 -11005 51215 -10885
rect 51335 -11005 51390 -10885
rect 51510 -11005 51555 -10885
rect 51675 -11005 51720 -10885
rect 51840 -11005 51885 -10885
rect 52005 -11005 52060 -10885
rect 52180 -11005 52225 -10885
rect 52345 -11005 52390 -10885
rect 52510 -11005 52555 -10885
rect 52675 -11005 52730 -10885
rect 52850 -11005 52895 -10885
rect 53015 -11005 53060 -10885
rect 53180 -11005 53225 -10885
rect 53345 -11005 53370 -10885
rect 30770 -11050 53370 -11005
rect 30770 -11170 30795 -11050
rect 30915 -11170 30970 -11050
rect 31090 -11170 31135 -11050
rect 31255 -11170 31300 -11050
rect 31420 -11170 31465 -11050
rect 31585 -11170 31640 -11050
rect 31760 -11170 31805 -11050
rect 31925 -11170 31970 -11050
rect 32090 -11170 32135 -11050
rect 32255 -11170 32310 -11050
rect 32430 -11170 32475 -11050
rect 32595 -11170 32640 -11050
rect 32760 -11170 32805 -11050
rect 32925 -11170 32980 -11050
rect 33100 -11170 33145 -11050
rect 33265 -11170 33310 -11050
rect 33430 -11170 33475 -11050
rect 33595 -11170 33650 -11050
rect 33770 -11170 33815 -11050
rect 33935 -11170 33980 -11050
rect 34100 -11170 34145 -11050
rect 34265 -11170 34320 -11050
rect 34440 -11170 34485 -11050
rect 34605 -11170 34650 -11050
rect 34770 -11170 34815 -11050
rect 34935 -11170 34990 -11050
rect 35110 -11170 35155 -11050
rect 35275 -11170 35320 -11050
rect 35440 -11170 35485 -11050
rect 35605 -11170 35660 -11050
rect 35780 -11170 35825 -11050
rect 35945 -11170 35990 -11050
rect 36110 -11170 36155 -11050
rect 36275 -11170 36485 -11050
rect 36605 -11170 36660 -11050
rect 36780 -11170 36825 -11050
rect 36945 -11170 36990 -11050
rect 37110 -11170 37155 -11050
rect 37275 -11170 37330 -11050
rect 37450 -11170 37495 -11050
rect 37615 -11170 37660 -11050
rect 37780 -11170 37825 -11050
rect 37945 -11170 38000 -11050
rect 38120 -11170 38165 -11050
rect 38285 -11170 38330 -11050
rect 38450 -11170 38495 -11050
rect 38615 -11170 38670 -11050
rect 38790 -11170 38835 -11050
rect 38955 -11170 39000 -11050
rect 39120 -11170 39165 -11050
rect 39285 -11170 39340 -11050
rect 39460 -11170 39505 -11050
rect 39625 -11170 39670 -11050
rect 39790 -11170 39835 -11050
rect 39955 -11170 40010 -11050
rect 40130 -11170 40175 -11050
rect 40295 -11170 40340 -11050
rect 40460 -11170 40505 -11050
rect 40625 -11170 40680 -11050
rect 40800 -11170 40845 -11050
rect 40965 -11170 41010 -11050
rect 41130 -11170 41175 -11050
rect 41295 -11170 41350 -11050
rect 41470 -11170 41515 -11050
rect 41635 -11170 41680 -11050
rect 41800 -11170 41845 -11050
rect 41965 -11170 42175 -11050
rect 42295 -11170 42350 -11050
rect 42470 -11170 42515 -11050
rect 42635 -11170 42680 -11050
rect 42800 -11170 42845 -11050
rect 42965 -11170 43020 -11050
rect 43140 -11170 43185 -11050
rect 43305 -11170 43350 -11050
rect 43470 -11170 43515 -11050
rect 43635 -11170 43690 -11050
rect 43810 -11170 43855 -11050
rect 43975 -11170 44020 -11050
rect 44140 -11170 44185 -11050
rect 44305 -11170 44360 -11050
rect 44480 -11170 44525 -11050
rect 44645 -11170 44690 -11050
rect 44810 -11170 44855 -11050
rect 44975 -11170 45030 -11050
rect 45150 -11170 45195 -11050
rect 45315 -11170 45360 -11050
rect 45480 -11170 45525 -11050
rect 45645 -11170 45700 -11050
rect 45820 -11170 45865 -11050
rect 45985 -11170 46030 -11050
rect 46150 -11170 46195 -11050
rect 46315 -11170 46370 -11050
rect 46490 -11170 46535 -11050
rect 46655 -11170 46700 -11050
rect 46820 -11170 46865 -11050
rect 46985 -11170 47040 -11050
rect 47160 -11170 47205 -11050
rect 47325 -11170 47370 -11050
rect 47490 -11170 47535 -11050
rect 47655 -11170 47865 -11050
rect 47985 -11170 48040 -11050
rect 48160 -11170 48205 -11050
rect 48325 -11170 48370 -11050
rect 48490 -11170 48535 -11050
rect 48655 -11170 48710 -11050
rect 48830 -11170 48875 -11050
rect 48995 -11170 49040 -11050
rect 49160 -11170 49205 -11050
rect 49325 -11170 49380 -11050
rect 49500 -11170 49545 -11050
rect 49665 -11170 49710 -11050
rect 49830 -11170 49875 -11050
rect 49995 -11170 50050 -11050
rect 50170 -11170 50215 -11050
rect 50335 -11170 50380 -11050
rect 50500 -11170 50545 -11050
rect 50665 -11170 50720 -11050
rect 50840 -11170 50885 -11050
rect 51005 -11170 51050 -11050
rect 51170 -11170 51215 -11050
rect 51335 -11170 51390 -11050
rect 51510 -11170 51555 -11050
rect 51675 -11170 51720 -11050
rect 51840 -11170 51885 -11050
rect 52005 -11170 52060 -11050
rect 52180 -11170 52225 -11050
rect 52345 -11170 52390 -11050
rect 52510 -11170 52555 -11050
rect 52675 -11170 52730 -11050
rect 52850 -11170 52895 -11050
rect 53015 -11170 53060 -11050
rect 53180 -11170 53225 -11050
rect 53345 -11170 53370 -11050
rect 30770 -11215 53370 -11170
rect 30770 -11335 30795 -11215
rect 30915 -11335 30970 -11215
rect 31090 -11335 31135 -11215
rect 31255 -11335 31300 -11215
rect 31420 -11335 31465 -11215
rect 31585 -11335 31640 -11215
rect 31760 -11335 31805 -11215
rect 31925 -11335 31970 -11215
rect 32090 -11335 32135 -11215
rect 32255 -11335 32310 -11215
rect 32430 -11335 32475 -11215
rect 32595 -11335 32640 -11215
rect 32760 -11335 32805 -11215
rect 32925 -11335 32980 -11215
rect 33100 -11335 33145 -11215
rect 33265 -11335 33310 -11215
rect 33430 -11335 33475 -11215
rect 33595 -11335 33650 -11215
rect 33770 -11335 33815 -11215
rect 33935 -11335 33980 -11215
rect 34100 -11335 34145 -11215
rect 34265 -11335 34320 -11215
rect 34440 -11335 34485 -11215
rect 34605 -11335 34650 -11215
rect 34770 -11335 34815 -11215
rect 34935 -11335 34990 -11215
rect 35110 -11335 35155 -11215
rect 35275 -11335 35320 -11215
rect 35440 -11335 35485 -11215
rect 35605 -11335 35660 -11215
rect 35780 -11335 35825 -11215
rect 35945 -11335 35990 -11215
rect 36110 -11335 36155 -11215
rect 36275 -11335 36485 -11215
rect 36605 -11335 36660 -11215
rect 36780 -11335 36825 -11215
rect 36945 -11335 36990 -11215
rect 37110 -11335 37155 -11215
rect 37275 -11335 37330 -11215
rect 37450 -11335 37495 -11215
rect 37615 -11335 37660 -11215
rect 37780 -11335 37825 -11215
rect 37945 -11335 38000 -11215
rect 38120 -11335 38165 -11215
rect 38285 -11335 38330 -11215
rect 38450 -11335 38495 -11215
rect 38615 -11335 38670 -11215
rect 38790 -11335 38835 -11215
rect 38955 -11335 39000 -11215
rect 39120 -11335 39165 -11215
rect 39285 -11335 39340 -11215
rect 39460 -11335 39505 -11215
rect 39625 -11335 39670 -11215
rect 39790 -11335 39835 -11215
rect 39955 -11335 40010 -11215
rect 40130 -11335 40175 -11215
rect 40295 -11335 40340 -11215
rect 40460 -11335 40505 -11215
rect 40625 -11335 40680 -11215
rect 40800 -11335 40845 -11215
rect 40965 -11335 41010 -11215
rect 41130 -11335 41175 -11215
rect 41295 -11335 41350 -11215
rect 41470 -11335 41515 -11215
rect 41635 -11335 41680 -11215
rect 41800 -11335 41845 -11215
rect 41965 -11335 42175 -11215
rect 42295 -11335 42350 -11215
rect 42470 -11335 42515 -11215
rect 42635 -11335 42680 -11215
rect 42800 -11335 42845 -11215
rect 42965 -11335 43020 -11215
rect 43140 -11335 43185 -11215
rect 43305 -11335 43350 -11215
rect 43470 -11335 43515 -11215
rect 43635 -11335 43690 -11215
rect 43810 -11335 43855 -11215
rect 43975 -11335 44020 -11215
rect 44140 -11335 44185 -11215
rect 44305 -11335 44360 -11215
rect 44480 -11335 44525 -11215
rect 44645 -11335 44690 -11215
rect 44810 -11335 44855 -11215
rect 44975 -11335 45030 -11215
rect 45150 -11335 45195 -11215
rect 45315 -11335 45360 -11215
rect 45480 -11335 45525 -11215
rect 45645 -11335 45700 -11215
rect 45820 -11335 45865 -11215
rect 45985 -11335 46030 -11215
rect 46150 -11335 46195 -11215
rect 46315 -11335 46370 -11215
rect 46490 -11335 46535 -11215
rect 46655 -11335 46700 -11215
rect 46820 -11335 46865 -11215
rect 46985 -11335 47040 -11215
rect 47160 -11335 47205 -11215
rect 47325 -11335 47370 -11215
rect 47490 -11335 47535 -11215
rect 47655 -11335 47865 -11215
rect 47985 -11335 48040 -11215
rect 48160 -11335 48205 -11215
rect 48325 -11335 48370 -11215
rect 48490 -11335 48535 -11215
rect 48655 -11335 48710 -11215
rect 48830 -11335 48875 -11215
rect 48995 -11335 49040 -11215
rect 49160 -11335 49205 -11215
rect 49325 -11335 49380 -11215
rect 49500 -11335 49545 -11215
rect 49665 -11335 49710 -11215
rect 49830 -11335 49875 -11215
rect 49995 -11335 50050 -11215
rect 50170 -11335 50215 -11215
rect 50335 -11335 50380 -11215
rect 50500 -11335 50545 -11215
rect 50665 -11335 50720 -11215
rect 50840 -11335 50885 -11215
rect 51005 -11335 51050 -11215
rect 51170 -11335 51215 -11215
rect 51335 -11335 51390 -11215
rect 51510 -11335 51555 -11215
rect 51675 -11335 51720 -11215
rect 51840 -11335 51885 -11215
rect 52005 -11335 52060 -11215
rect 52180 -11335 52225 -11215
rect 52345 -11335 52390 -11215
rect 52510 -11335 52555 -11215
rect 52675 -11335 52730 -11215
rect 52850 -11335 52895 -11215
rect 53015 -11335 53060 -11215
rect 53180 -11335 53225 -11215
rect 53345 -11335 53370 -11215
rect 30770 -11390 53370 -11335
rect 30770 -11510 30795 -11390
rect 30915 -11510 30970 -11390
rect 31090 -11510 31135 -11390
rect 31255 -11510 31300 -11390
rect 31420 -11510 31465 -11390
rect 31585 -11510 31640 -11390
rect 31760 -11510 31805 -11390
rect 31925 -11510 31970 -11390
rect 32090 -11510 32135 -11390
rect 32255 -11510 32310 -11390
rect 32430 -11510 32475 -11390
rect 32595 -11510 32640 -11390
rect 32760 -11510 32805 -11390
rect 32925 -11510 32980 -11390
rect 33100 -11510 33145 -11390
rect 33265 -11510 33310 -11390
rect 33430 -11510 33475 -11390
rect 33595 -11510 33650 -11390
rect 33770 -11510 33815 -11390
rect 33935 -11510 33980 -11390
rect 34100 -11510 34145 -11390
rect 34265 -11510 34320 -11390
rect 34440 -11510 34485 -11390
rect 34605 -11510 34650 -11390
rect 34770 -11510 34815 -11390
rect 34935 -11510 34990 -11390
rect 35110 -11510 35155 -11390
rect 35275 -11510 35320 -11390
rect 35440 -11510 35485 -11390
rect 35605 -11510 35660 -11390
rect 35780 -11510 35825 -11390
rect 35945 -11510 35990 -11390
rect 36110 -11510 36155 -11390
rect 36275 -11510 36485 -11390
rect 36605 -11510 36660 -11390
rect 36780 -11510 36825 -11390
rect 36945 -11510 36990 -11390
rect 37110 -11510 37155 -11390
rect 37275 -11510 37330 -11390
rect 37450 -11510 37495 -11390
rect 37615 -11510 37660 -11390
rect 37780 -11510 37825 -11390
rect 37945 -11510 38000 -11390
rect 38120 -11510 38165 -11390
rect 38285 -11510 38330 -11390
rect 38450 -11510 38495 -11390
rect 38615 -11510 38670 -11390
rect 38790 -11510 38835 -11390
rect 38955 -11510 39000 -11390
rect 39120 -11510 39165 -11390
rect 39285 -11510 39340 -11390
rect 39460 -11510 39505 -11390
rect 39625 -11510 39670 -11390
rect 39790 -11510 39835 -11390
rect 39955 -11510 40010 -11390
rect 40130 -11510 40175 -11390
rect 40295 -11510 40340 -11390
rect 40460 -11510 40505 -11390
rect 40625 -11510 40680 -11390
rect 40800 -11510 40845 -11390
rect 40965 -11510 41010 -11390
rect 41130 -11510 41175 -11390
rect 41295 -11510 41350 -11390
rect 41470 -11510 41515 -11390
rect 41635 -11510 41680 -11390
rect 41800 -11510 41845 -11390
rect 41965 -11510 42175 -11390
rect 42295 -11510 42350 -11390
rect 42470 -11510 42515 -11390
rect 42635 -11510 42680 -11390
rect 42800 -11510 42845 -11390
rect 42965 -11510 43020 -11390
rect 43140 -11510 43185 -11390
rect 43305 -11510 43350 -11390
rect 43470 -11510 43515 -11390
rect 43635 -11510 43690 -11390
rect 43810 -11510 43855 -11390
rect 43975 -11510 44020 -11390
rect 44140 -11510 44185 -11390
rect 44305 -11510 44360 -11390
rect 44480 -11510 44525 -11390
rect 44645 -11510 44690 -11390
rect 44810 -11510 44855 -11390
rect 44975 -11510 45030 -11390
rect 45150 -11510 45195 -11390
rect 45315 -11510 45360 -11390
rect 45480 -11510 45525 -11390
rect 45645 -11510 45700 -11390
rect 45820 -11510 45865 -11390
rect 45985 -11510 46030 -11390
rect 46150 -11510 46195 -11390
rect 46315 -11510 46370 -11390
rect 46490 -11510 46535 -11390
rect 46655 -11510 46700 -11390
rect 46820 -11510 46865 -11390
rect 46985 -11510 47040 -11390
rect 47160 -11510 47205 -11390
rect 47325 -11510 47370 -11390
rect 47490 -11510 47535 -11390
rect 47655 -11510 47865 -11390
rect 47985 -11510 48040 -11390
rect 48160 -11510 48205 -11390
rect 48325 -11510 48370 -11390
rect 48490 -11510 48535 -11390
rect 48655 -11510 48710 -11390
rect 48830 -11510 48875 -11390
rect 48995 -11510 49040 -11390
rect 49160 -11510 49205 -11390
rect 49325 -11510 49380 -11390
rect 49500 -11510 49545 -11390
rect 49665 -11510 49710 -11390
rect 49830 -11510 49875 -11390
rect 49995 -11510 50050 -11390
rect 50170 -11510 50215 -11390
rect 50335 -11510 50380 -11390
rect 50500 -11510 50545 -11390
rect 50665 -11510 50720 -11390
rect 50840 -11510 50885 -11390
rect 51005 -11510 51050 -11390
rect 51170 -11510 51215 -11390
rect 51335 -11510 51390 -11390
rect 51510 -11510 51555 -11390
rect 51675 -11510 51720 -11390
rect 51840 -11510 51885 -11390
rect 52005 -11510 52060 -11390
rect 52180 -11510 52225 -11390
rect 52345 -11510 52390 -11390
rect 52510 -11510 52555 -11390
rect 52675 -11510 52730 -11390
rect 52850 -11510 52895 -11390
rect 53015 -11510 53060 -11390
rect 53180 -11510 53225 -11390
rect 53345 -11510 53370 -11390
rect 30770 -11555 53370 -11510
rect 30770 -11675 30795 -11555
rect 30915 -11675 30970 -11555
rect 31090 -11675 31135 -11555
rect 31255 -11675 31300 -11555
rect 31420 -11675 31465 -11555
rect 31585 -11675 31640 -11555
rect 31760 -11675 31805 -11555
rect 31925 -11675 31970 -11555
rect 32090 -11675 32135 -11555
rect 32255 -11675 32310 -11555
rect 32430 -11675 32475 -11555
rect 32595 -11675 32640 -11555
rect 32760 -11675 32805 -11555
rect 32925 -11675 32980 -11555
rect 33100 -11675 33145 -11555
rect 33265 -11675 33310 -11555
rect 33430 -11675 33475 -11555
rect 33595 -11675 33650 -11555
rect 33770 -11675 33815 -11555
rect 33935 -11675 33980 -11555
rect 34100 -11675 34145 -11555
rect 34265 -11675 34320 -11555
rect 34440 -11675 34485 -11555
rect 34605 -11675 34650 -11555
rect 34770 -11675 34815 -11555
rect 34935 -11675 34990 -11555
rect 35110 -11675 35155 -11555
rect 35275 -11675 35320 -11555
rect 35440 -11675 35485 -11555
rect 35605 -11675 35660 -11555
rect 35780 -11675 35825 -11555
rect 35945 -11675 35990 -11555
rect 36110 -11675 36155 -11555
rect 36275 -11675 36485 -11555
rect 36605 -11675 36660 -11555
rect 36780 -11675 36825 -11555
rect 36945 -11675 36990 -11555
rect 37110 -11675 37155 -11555
rect 37275 -11675 37330 -11555
rect 37450 -11675 37495 -11555
rect 37615 -11675 37660 -11555
rect 37780 -11675 37825 -11555
rect 37945 -11675 38000 -11555
rect 38120 -11675 38165 -11555
rect 38285 -11675 38330 -11555
rect 38450 -11675 38495 -11555
rect 38615 -11675 38670 -11555
rect 38790 -11675 38835 -11555
rect 38955 -11675 39000 -11555
rect 39120 -11675 39165 -11555
rect 39285 -11675 39340 -11555
rect 39460 -11675 39505 -11555
rect 39625 -11675 39670 -11555
rect 39790 -11675 39835 -11555
rect 39955 -11675 40010 -11555
rect 40130 -11675 40175 -11555
rect 40295 -11675 40340 -11555
rect 40460 -11675 40505 -11555
rect 40625 -11675 40680 -11555
rect 40800 -11675 40845 -11555
rect 40965 -11675 41010 -11555
rect 41130 -11675 41175 -11555
rect 41295 -11675 41350 -11555
rect 41470 -11675 41515 -11555
rect 41635 -11675 41680 -11555
rect 41800 -11675 41845 -11555
rect 41965 -11675 42175 -11555
rect 42295 -11675 42350 -11555
rect 42470 -11675 42515 -11555
rect 42635 -11675 42680 -11555
rect 42800 -11675 42845 -11555
rect 42965 -11675 43020 -11555
rect 43140 -11675 43185 -11555
rect 43305 -11675 43350 -11555
rect 43470 -11675 43515 -11555
rect 43635 -11675 43690 -11555
rect 43810 -11675 43855 -11555
rect 43975 -11675 44020 -11555
rect 44140 -11675 44185 -11555
rect 44305 -11675 44360 -11555
rect 44480 -11675 44525 -11555
rect 44645 -11675 44690 -11555
rect 44810 -11675 44855 -11555
rect 44975 -11675 45030 -11555
rect 45150 -11675 45195 -11555
rect 45315 -11675 45360 -11555
rect 45480 -11675 45525 -11555
rect 45645 -11675 45700 -11555
rect 45820 -11675 45865 -11555
rect 45985 -11675 46030 -11555
rect 46150 -11675 46195 -11555
rect 46315 -11675 46370 -11555
rect 46490 -11675 46535 -11555
rect 46655 -11675 46700 -11555
rect 46820 -11675 46865 -11555
rect 46985 -11675 47040 -11555
rect 47160 -11675 47205 -11555
rect 47325 -11675 47370 -11555
rect 47490 -11675 47535 -11555
rect 47655 -11675 47865 -11555
rect 47985 -11675 48040 -11555
rect 48160 -11675 48205 -11555
rect 48325 -11675 48370 -11555
rect 48490 -11675 48535 -11555
rect 48655 -11675 48710 -11555
rect 48830 -11675 48875 -11555
rect 48995 -11675 49040 -11555
rect 49160 -11675 49205 -11555
rect 49325 -11675 49380 -11555
rect 49500 -11675 49545 -11555
rect 49665 -11675 49710 -11555
rect 49830 -11675 49875 -11555
rect 49995 -11675 50050 -11555
rect 50170 -11675 50215 -11555
rect 50335 -11675 50380 -11555
rect 50500 -11675 50545 -11555
rect 50665 -11675 50720 -11555
rect 50840 -11675 50885 -11555
rect 51005 -11675 51050 -11555
rect 51170 -11675 51215 -11555
rect 51335 -11675 51390 -11555
rect 51510 -11675 51555 -11555
rect 51675 -11675 51720 -11555
rect 51840 -11675 51885 -11555
rect 52005 -11675 52060 -11555
rect 52180 -11675 52225 -11555
rect 52345 -11675 52390 -11555
rect 52510 -11675 52555 -11555
rect 52675 -11675 52730 -11555
rect 52850 -11675 52895 -11555
rect 53015 -11675 53060 -11555
rect 53180 -11675 53225 -11555
rect 53345 -11675 53370 -11555
rect 30770 -11720 53370 -11675
rect 30770 -11840 30795 -11720
rect 30915 -11840 30970 -11720
rect 31090 -11840 31135 -11720
rect 31255 -11840 31300 -11720
rect 31420 -11840 31465 -11720
rect 31585 -11840 31640 -11720
rect 31760 -11840 31805 -11720
rect 31925 -11840 31970 -11720
rect 32090 -11840 32135 -11720
rect 32255 -11840 32310 -11720
rect 32430 -11840 32475 -11720
rect 32595 -11840 32640 -11720
rect 32760 -11840 32805 -11720
rect 32925 -11840 32980 -11720
rect 33100 -11840 33145 -11720
rect 33265 -11840 33310 -11720
rect 33430 -11840 33475 -11720
rect 33595 -11840 33650 -11720
rect 33770 -11840 33815 -11720
rect 33935 -11840 33980 -11720
rect 34100 -11840 34145 -11720
rect 34265 -11840 34320 -11720
rect 34440 -11840 34485 -11720
rect 34605 -11840 34650 -11720
rect 34770 -11840 34815 -11720
rect 34935 -11840 34990 -11720
rect 35110 -11840 35155 -11720
rect 35275 -11840 35320 -11720
rect 35440 -11840 35485 -11720
rect 35605 -11840 35660 -11720
rect 35780 -11840 35825 -11720
rect 35945 -11840 35990 -11720
rect 36110 -11840 36155 -11720
rect 36275 -11840 36485 -11720
rect 36605 -11840 36660 -11720
rect 36780 -11840 36825 -11720
rect 36945 -11840 36990 -11720
rect 37110 -11840 37155 -11720
rect 37275 -11840 37330 -11720
rect 37450 -11840 37495 -11720
rect 37615 -11840 37660 -11720
rect 37780 -11840 37825 -11720
rect 37945 -11840 38000 -11720
rect 38120 -11840 38165 -11720
rect 38285 -11840 38330 -11720
rect 38450 -11840 38495 -11720
rect 38615 -11840 38670 -11720
rect 38790 -11840 38835 -11720
rect 38955 -11840 39000 -11720
rect 39120 -11840 39165 -11720
rect 39285 -11840 39340 -11720
rect 39460 -11840 39505 -11720
rect 39625 -11840 39670 -11720
rect 39790 -11840 39835 -11720
rect 39955 -11840 40010 -11720
rect 40130 -11840 40175 -11720
rect 40295 -11840 40340 -11720
rect 40460 -11840 40505 -11720
rect 40625 -11840 40680 -11720
rect 40800 -11840 40845 -11720
rect 40965 -11840 41010 -11720
rect 41130 -11840 41175 -11720
rect 41295 -11840 41350 -11720
rect 41470 -11840 41515 -11720
rect 41635 -11840 41680 -11720
rect 41800 -11840 41845 -11720
rect 41965 -11840 42175 -11720
rect 42295 -11840 42350 -11720
rect 42470 -11840 42515 -11720
rect 42635 -11840 42680 -11720
rect 42800 -11840 42845 -11720
rect 42965 -11840 43020 -11720
rect 43140 -11840 43185 -11720
rect 43305 -11840 43350 -11720
rect 43470 -11840 43515 -11720
rect 43635 -11840 43690 -11720
rect 43810 -11840 43855 -11720
rect 43975 -11840 44020 -11720
rect 44140 -11840 44185 -11720
rect 44305 -11840 44360 -11720
rect 44480 -11840 44525 -11720
rect 44645 -11840 44690 -11720
rect 44810 -11840 44855 -11720
rect 44975 -11840 45030 -11720
rect 45150 -11840 45195 -11720
rect 45315 -11840 45360 -11720
rect 45480 -11840 45525 -11720
rect 45645 -11840 45700 -11720
rect 45820 -11840 45865 -11720
rect 45985 -11840 46030 -11720
rect 46150 -11840 46195 -11720
rect 46315 -11840 46370 -11720
rect 46490 -11840 46535 -11720
rect 46655 -11840 46700 -11720
rect 46820 -11840 46865 -11720
rect 46985 -11840 47040 -11720
rect 47160 -11840 47205 -11720
rect 47325 -11840 47370 -11720
rect 47490 -11840 47535 -11720
rect 47655 -11840 47865 -11720
rect 47985 -11840 48040 -11720
rect 48160 -11840 48205 -11720
rect 48325 -11840 48370 -11720
rect 48490 -11840 48535 -11720
rect 48655 -11840 48710 -11720
rect 48830 -11840 48875 -11720
rect 48995 -11840 49040 -11720
rect 49160 -11840 49205 -11720
rect 49325 -11840 49380 -11720
rect 49500 -11840 49545 -11720
rect 49665 -11840 49710 -11720
rect 49830 -11840 49875 -11720
rect 49995 -11840 50050 -11720
rect 50170 -11840 50215 -11720
rect 50335 -11840 50380 -11720
rect 50500 -11840 50545 -11720
rect 50665 -11840 50720 -11720
rect 50840 -11840 50885 -11720
rect 51005 -11840 51050 -11720
rect 51170 -11840 51215 -11720
rect 51335 -11840 51390 -11720
rect 51510 -11840 51555 -11720
rect 51675 -11840 51720 -11720
rect 51840 -11840 51885 -11720
rect 52005 -11840 52060 -11720
rect 52180 -11840 52225 -11720
rect 52345 -11840 52390 -11720
rect 52510 -11840 52555 -11720
rect 52675 -11840 52730 -11720
rect 52850 -11840 52895 -11720
rect 53015 -11840 53060 -11720
rect 53180 -11840 53225 -11720
rect 53345 -11840 53370 -11720
rect 30770 -11885 53370 -11840
rect 30770 -12005 30795 -11885
rect 30915 -12005 30970 -11885
rect 31090 -12005 31135 -11885
rect 31255 -12005 31300 -11885
rect 31420 -12005 31465 -11885
rect 31585 -12005 31640 -11885
rect 31760 -12005 31805 -11885
rect 31925 -12005 31970 -11885
rect 32090 -12005 32135 -11885
rect 32255 -12005 32310 -11885
rect 32430 -12005 32475 -11885
rect 32595 -12005 32640 -11885
rect 32760 -12005 32805 -11885
rect 32925 -12005 32980 -11885
rect 33100 -12005 33145 -11885
rect 33265 -12005 33310 -11885
rect 33430 -12005 33475 -11885
rect 33595 -12005 33650 -11885
rect 33770 -12005 33815 -11885
rect 33935 -12005 33980 -11885
rect 34100 -12005 34145 -11885
rect 34265 -12005 34320 -11885
rect 34440 -12005 34485 -11885
rect 34605 -12005 34650 -11885
rect 34770 -12005 34815 -11885
rect 34935 -12005 34990 -11885
rect 35110 -12005 35155 -11885
rect 35275 -12005 35320 -11885
rect 35440 -12005 35485 -11885
rect 35605 -12005 35660 -11885
rect 35780 -12005 35825 -11885
rect 35945 -12005 35990 -11885
rect 36110 -12005 36155 -11885
rect 36275 -12005 36485 -11885
rect 36605 -12005 36660 -11885
rect 36780 -12005 36825 -11885
rect 36945 -12005 36990 -11885
rect 37110 -12005 37155 -11885
rect 37275 -12005 37330 -11885
rect 37450 -12005 37495 -11885
rect 37615 -12005 37660 -11885
rect 37780 -12005 37825 -11885
rect 37945 -12005 38000 -11885
rect 38120 -12005 38165 -11885
rect 38285 -12005 38330 -11885
rect 38450 -12005 38495 -11885
rect 38615 -12005 38670 -11885
rect 38790 -12005 38835 -11885
rect 38955 -12005 39000 -11885
rect 39120 -12005 39165 -11885
rect 39285 -12005 39340 -11885
rect 39460 -12005 39505 -11885
rect 39625 -12005 39670 -11885
rect 39790 -12005 39835 -11885
rect 39955 -12005 40010 -11885
rect 40130 -12005 40175 -11885
rect 40295 -12005 40340 -11885
rect 40460 -12005 40505 -11885
rect 40625 -12005 40680 -11885
rect 40800 -12005 40845 -11885
rect 40965 -12005 41010 -11885
rect 41130 -12005 41175 -11885
rect 41295 -12005 41350 -11885
rect 41470 -12005 41515 -11885
rect 41635 -12005 41680 -11885
rect 41800 -12005 41845 -11885
rect 41965 -12005 42175 -11885
rect 42295 -12005 42350 -11885
rect 42470 -12005 42515 -11885
rect 42635 -12005 42680 -11885
rect 42800 -12005 42845 -11885
rect 42965 -12005 43020 -11885
rect 43140 -12005 43185 -11885
rect 43305 -12005 43350 -11885
rect 43470 -12005 43515 -11885
rect 43635 -12005 43690 -11885
rect 43810 -12005 43855 -11885
rect 43975 -12005 44020 -11885
rect 44140 -12005 44185 -11885
rect 44305 -12005 44360 -11885
rect 44480 -12005 44525 -11885
rect 44645 -12005 44690 -11885
rect 44810 -12005 44855 -11885
rect 44975 -12005 45030 -11885
rect 45150 -12005 45195 -11885
rect 45315 -12005 45360 -11885
rect 45480 -12005 45525 -11885
rect 45645 -12005 45700 -11885
rect 45820 -12005 45865 -11885
rect 45985 -12005 46030 -11885
rect 46150 -12005 46195 -11885
rect 46315 -12005 46370 -11885
rect 46490 -12005 46535 -11885
rect 46655 -12005 46700 -11885
rect 46820 -12005 46865 -11885
rect 46985 -12005 47040 -11885
rect 47160 -12005 47205 -11885
rect 47325 -12005 47370 -11885
rect 47490 -12005 47535 -11885
rect 47655 -12005 47865 -11885
rect 47985 -12005 48040 -11885
rect 48160 -12005 48205 -11885
rect 48325 -12005 48370 -11885
rect 48490 -12005 48535 -11885
rect 48655 -12005 48710 -11885
rect 48830 -12005 48875 -11885
rect 48995 -12005 49040 -11885
rect 49160 -12005 49205 -11885
rect 49325 -12005 49380 -11885
rect 49500 -12005 49545 -11885
rect 49665 -12005 49710 -11885
rect 49830 -12005 49875 -11885
rect 49995 -12005 50050 -11885
rect 50170 -12005 50215 -11885
rect 50335 -12005 50380 -11885
rect 50500 -12005 50545 -11885
rect 50665 -12005 50720 -11885
rect 50840 -12005 50885 -11885
rect 51005 -12005 51050 -11885
rect 51170 -12005 51215 -11885
rect 51335 -12005 51390 -11885
rect 51510 -12005 51555 -11885
rect 51675 -12005 51720 -11885
rect 51840 -12005 51885 -11885
rect 52005 -12005 52060 -11885
rect 52180 -12005 52225 -11885
rect 52345 -12005 52390 -11885
rect 52510 -12005 52555 -11885
rect 52675 -12005 52730 -11885
rect 52850 -12005 52895 -11885
rect 53015 -12005 53060 -11885
rect 53180 -12005 53225 -11885
rect 53345 -12005 53370 -11885
rect 30770 -12060 53370 -12005
rect 30770 -12180 30795 -12060
rect 30915 -12180 30970 -12060
rect 31090 -12180 31135 -12060
rect 31255 -12180 31300 -12060
rect 31420 -12180 31465 -12060
rect 31585 -12180 31640 -12060
rect 31760 -12180 31805 -12060
rect 31925 -12180 31970 -12060
rect 32090 -12180 32135 -12060
rect 32255 -12180 32310 -12060
rect 32430 -12180 32475 -12060
rect 32595 -12180 32640 -12060
rect 32760 -12180 32805 -12060
rect 32925 -12180 32980 -12060
rect 33100 -12180 33145 -12060
rect 33265 -12180 33310 -12060
rect 33430 -12180 33475 -12060
rect 33595 -12180 33650 -12060
rect 33770 -12180 33815 -12060
rect 33935 -12180 33980 -12060
rect 34100 -12180 34145 -12060
rect 34265 -12180 34320 -12060
rect 34440 -12180 34485 -12060
rect 34605 -12180 34650 -12060
rect 34770 -12180 34815 -12060
rect 34935 -12180 34990 -12060
rect 35110 -12180 35155 -12060
rect 35275 -12180 35320 -12060
rect 35440 -12180 35485 -12060
rect 35605 -12180 35660 -12060
rect 35780 -12180 35825 -12060
rect 35945 -12180 35990 -12060
rect 36110 -12180 36155 -12060
rect 36275 -12180 36485 -12060
rect 36605 -12180 36660 -12060
rect 36780 -12180 36825 -12060
rect 36945 -12180 36990 -12060
rect 37110 -12180 37155 -12060
rect 37275 -12180 37330 -12060
rect 37450 -12180 37495 -12060
rect 37615 -12180 37660 -12060
rect 37780 -12180 37825 -12060
rect 37945 -12180 38000 -12060
rect 38120 -12180 38165 -12060
rect 38285 -12180 38330 -12060
rect 38450 -12180 38495 -12060
rect 38615 -12180 38670 -12060
rect 38790 -12180 38835 -12060
rect 38955 -12180 39000 -12060
rect 39120 -12180 39165 -12060
rect 39285 -12180 39340 -12060
rect 39460 -12180 39505 -12060
rect 39625 -12180 39670 -12060
rect 39790 -12180 39835 -12060
rect 39955 -12180 40010 -12060
rect 40130 -12180 40175 -12060
rect 40295 -12180 40340 -12060
rect 40460 -12180 40505 -12060
rect 40625 -12180 40680 -12060
rect 40800 -12180 40845 -12060
rect 40965 -12180 41010 -12060
rect 41130 -12180 41175 -12060
rect 41295 -12180 41350 -12060
rect 41470 -12180 41515 -12060
rect 41635 -12180 41680 -12060
rect 41800 -12180 41845 -12060
rect 41965 -12180 42175 -12060
rect 42295 -12180 42350 -12060
rect 42470 -12180 42515 -12060
rect 42635 -12180 42680 -12060
rect 42800 -12180 42845 -12060
rect 42965 -12180 43020 -12060
rect 43140 -12180 43185 -12060
rect 43305 -12180 43350 -12060
rect 43470 -12180 43515 -12060
rect 43635 -12180 43690 -12060
rect 43810 -12180 43855 -12060
rect 43975 -12180 44020 -12060
rect 44140 -12180 44185 -12060
rect 44305 -12180 44360 -12060
rect 44480 -12180 44525 -12060
rect 44645 -12180 44690 -12060
rect 44810 -12180 44855 -12060
rect 44975 -12180 45030 -12060
rect 45150 -12180 45195 -12060
rect 45315 -12180 45360 -12060
rect 45480 -12180 45525 -12060
rect 45645 -12180 45700 -12060
rect 45820 -12180 45865 -12060
rect 45985 -12180 46030 -12060
rect 46150 -12180 46195 -12060
rect 46315 -12180 46370 -12060
rect 46490 -12180 46535 -12060
rect 46655 -12180 46700 -12060
rect 46820 -12180 46865 -12060
rect 46985 -12180 47040 -12060
rect 47160 -12180 47205 -12060
rect 47325 -12180 47370 -12060
rect 47490 -12180 47535 -12060
rect 47655 -12180 47865 -12060
rect 47985 -12180 48040 -12060
rect 48160 -12180 48205 -12060
rect 48325 -12180 48370 -12060
rect 48490 -12180 48535 -12060
rect 48655 -12180 48710 -12060
rect 48830 -12180 48875 -12060
rect 48995 -12180 49040 -12060
rect 49160 -12180 49205 -12060
rect 49325 -12180 49380 -12060
rect 49500 -12180 49545 -12060
rect 49665 -12180 49710 -12060
rect 49830 -12180 49875 -12060
rect 49995 -12180 50050 -12060
rect 50170 -12180 50215 -12060
rect 50335 -12180 50380 -12060
rect 50500 -12180 50545 -12060
rect 50665 -12180 50720 -12060
rect 50840 -12180 50885 -12060
rect 51005 -12180 51050 -12060
rect 51170 -12180 51215 -12060
rect 51335 -12180 51390 -12060
rect 51510 -12180 51555 -12060
rect 51675 -12180 51720 -12060
rect 51840 -12180 51885 -12060
rect 52005 -12180 52060 -12060
rect 52180 -12180 52225 -12060
rect 52345 -12180 52390 -12060
rect 52510 -12180 52555 -12060
rect 52675 -12180 52730 -12060
rect 52850 -12180 52895 -12060
rect 53015 -12180 53060 -12060
rect 53180 -12180 53225 -12060
rect 53345 -12180 53370 -12060
rect 30770 -12225 53370 -12180
rect 30770 -12345 30795 -12225
rect 30915 -12345 30970 -12225
rect 31090 -12345 31135 -12225
rect 31255 -12345 31300 -12225
rect 31420 -12345 31465 -12225
rect 31585 -12345 31640 -12225
rect 31760 -12345 31805 -12225
rect 31925 -12345 31970 -12225
rect 32090 -12345 32135 -12225
rect 32255 -12345 32310 -12225
rect 32430 -12345 32475 -12225
rect 32595 -12345 32640 -12225
rect 32760 -12345 32805 -12225
rect 32925 -12345 32980 -12225
rect 33100 -12345 33145 -12225
rect 33265 -12345 33310 -12225
rect 33430 -12345 33475 -12225
rect 33595 -12345 33650 -12225
rect 33770 -12345 33815 -12225
rect 33935 -12345 33980 -12225
rect 34100 -12345 34145 -12225
rect 34265 -12345 34320 -12225
rect 34440 -12345 34485 -12225
rect 34605 -12345 34650 -12225
rect 34770 -12345 34815 -12225
rect 34935 -12345 34990 -12225
rect 35110 -12345 35155 -12225
rect 35275 -12345 35320 -12225
rect 35440 -12345 35485 -12225
rect 35605 -12345 35660 -12225
rect 35780 -12345 35825 -12225
rect 35945 -12345 35990 -12225
rect 36110 -12345 36155 -12225
rect 36275 -12345 36485 -12225
rect 36605 -12345 36660 -12225
rect 36780 -12345 36825 -12225
rect 36945 -12345 36990 -12225
rect 37110 -12345 37155 -12225
rect 37275 -12345 37330 -12225
rect 37450 -12345 37495 -12225
rect 37615 -12345 37660 -12225
rect 37780 -12345 37825 -12225
rect 37945 -12345 38000 -12225
rect 38120 -12345 38165 -12225
rect 38285 -12345 38330 -12225
rect 38450 -12345 38495 -12225
rect 38615 -12345 38670 -12225
rect 38790 -12345 38835 -12225
rect 38955 -12345 39000 -12225
rect 39120 -12345 39165 -12225
rect 39285 -12345 39340 -12225
rect 39460 -12345 39505 -12225
rect 39625 -12345 39670 -12225
rect 39790 -12345 39835 -12225
rect 39955 -12345 40010 -12225
rect 40130 -12345 40175 -12225
rect 40295 -12345 40340 -12225
rect 40460 -12345 40505 -12225
rect 40625 -12345 40680 -12225
rect 40800 -12345 40845 -12225
rect 40965 -12345 41010 -12225
rect 41130 -12345 41175 -12225
rect 41295 -12345 41350 -12225
rect 41470 -12345 41515 -12225
rect 41635 -12345 41680 -12225
rect 41800 -12345 41845 -12225
rect 41965 -12345 42175 -12225
rect 42295 -12345 42350 -12225
rect 42470 -12345 42515 -12225
rect 42635 -12345 42680 -12225
rect 42800 -12345 42845 -12225
rect 42965 -12345 43020 -12225
rect 43140 -12345 43185 -12225
rect 43305 -12345 43350 -12225
rect 43470 -12345 43515 -12225
rect 43635 -12345 43690 -12225
rect 43810 -12345 43855 -12225
rect 43975 -12345 44020 -12225
rect 44140 -12345 44185 -12225
rect 44305 -12345 44360 -12225
rect 44480 -12345 44525 -12225
rect 44645 -12345 44690 -12225
rect 44810 -12345 44855 -12225
rect 44975 -12345 45030 -12225
rect 45150 -12345 45195 -12225
rect 45315 -12345 45360 -12225
rect 45480 -12345 45525 -12225
rect 45645 -12345 45700 -12225
rect 45820 -12345 45865 -12225
rect 45985 -12345 46030 -12225
rect 46150 -12345 46195 -12225
rect 46315 -12345 46370 -12225
rect 46490 -12345 46535 -12225
rect 46655 -12345 46700 -12225
rect 46820 -12345 46865 -12225
rect 46985 -12345 47040 -12225
rect 47160 -12345 47205 -12225
rect 47325 -12345 47370 -12225
rect 47490 -12345 47535 -12225
rect 47655 -12345 47865 -12225
rect 47985 -12345 48040 -12225
rect 48160 -12345 48205 -12225
rect 48325 -12345 48370 -12225
rect 48490 -12345 48535 -12225
rect 48655 -12345 48710 -12225
rect 48830 -12345 48875 -12225
rect 48995 -12345 49040 -12225
rect 49160 -12345 49205 -12225
rect 49325 -12345 49380 -12225
rect 49500 -12345 49545 -12225
rect 49665 -12345 49710 -12225
rect 49830 -12345 49875 -12225
rect 49995 -12345 50050 -12225
rect 50170 -12345 50215 -12225
rect 50335 -12345 50380 -12225
rect 50500 -12345 50545 -12225
rect 50665 -12345 50720 -12225
rect 50840 -12345 50885 -12225
rect 51005 -12345 51050 -12225
rect 51170 -12345 51215 -12225
rect 51335 -12345 51390 -12225
rect 51510 -12345 51555 -12225
rect 51675 -12345 51720 -12225
rect 51840 -12345 51885 -12225
rect 52005 -12345 52060 -12225
rect 52180 -12345 52225 -12225
rect 52345 -12345 52390 -12225
rect 52510 -12345 52555 -12225
rect 52675 -12345 52730 -12225
rect 52850 -12345 52895 -12225
rect 53015 -12345 53060 -12225
rect 53180 -12345 53225 -12225
rect 53345 -12345 53370 -12225
rect 30770 -12390 53370 -12345
rect 30770 -12510 30795 -12390
rect 30915 -12510 30970 -12390
rect 31090 -12510 31135 -12390
rect 31255 -12510 31300 -12390
rect 31420 -12510 31465 -12390
rect 31585 -12510 31640 -12390
rect 31760 -12510 31805 -12390
rect 31925 -12510 31970 -12390
rect 32090 -12510 32135 -12390
rect 32255 -12510 32310 -12390
rect 32430 -12510 32475 -12390
rect 32595 -12510 32640 -12390
rect 32760 -12510 32805 -12390
rect 32925 -12510 32980 -12390
rect 33100 -12510 33145 -12390
rect 33265 -12510 33310 -12390
rect 33430 -12510 33475 -12390
rect 33595 -12510 33650 -12390
rect 33770 -12510 33815 -12390
rect 33935 -12510 33980 -12390
rect 34100 -12510 34145 -12390
rect 34265 -12510 34320 -12390
rect 34440 -12510 34485 -12390
rect 34605 -12510 34650 -12390
rect 34770 -12510 34815 -12390
rect 34935 -12510 34990 -12390
rect 35110 -12510 35155 -12390
rect 35275 -12510 35320 -12390
rect 35440 -12510 35485 -12390
rect 35605 -12510 35660 -12390
rect 35780 -12510 35825 -12390
rect 35945 -12510 35990 -12390
rect 36110 -12510 36155 -12390
rect 36275 -12510 36485 -12390
rect 36605 -12510 36660 -12390
rect 36780 -12510 36825 -12390
rect 36945 -12510 36990 -12390
rect 37110 -12510 37155 -12390
rect 37275 -12510 37330 -12390
rect 37450 -12510 37495 -12390
rect 37615 -12510 37660 -12390
rect 37780 -12510 37825 -12390
rect 37945 -12510 38000 -12390
rect 38120 -12510 38165 -12390
rect 38285 -12510 38330 -12390
rect 38450 -12510 38495 -12390
rect 38615 -12510 38670 -12390
rect 38790 -12510 38835 -12390
rect 38955 -12510 39000 -12390
rect 39120 -12510 39165 -12390
rect 39285 -12510 39340 -12390
rect 39460 -12510 39505 -12390
rect 39625 -12510 39670 -12390
rect 39790 -12510 39835 -12390
rect 39955 -12510 40010 -12390
rect 40130 -12510 40175 -12390
rect 40295 -12510 40340 -12390
rect 40460 -12510 40505 -12390
rect 40625 -12510 40680 -12390
rect 40800 -12510 40845 -12390
rect 40965 -12510 41010 -12390
rect 41130 -12510 41175 -12390
rect 41295 -12510 41350 -12390
rect 41470 -12510 41515 -12390
rect 41635 -12510 41680 -12390
rect 41800 -12510 41845 -12390
rect 41965 -12510 42175 -12390
rect 42295 -12510 42350 -12390
rect 42470 -12510 42515 -12390
rect 42635 -12510 42680 -12390
rect 42800 -12510 42845 -12390
rect 42965 -12510 43020 -12390
rect 43140 -12510 43185 -12390
rect 43305 -12510 43350 -12390
rect 43470 -12510 43515 -12390
rect 43635 -12510 43690 -12390
rect 43810 -12510 43855 -12390
rect 43975 -12510 44020 -12390
rect 44140 -12510 44185 -12390
rect 44305 -12510 44360 -12390
rect 44480 -12510 44525 -12390
rect 44645 -12510 44690 -12390
rect 44810 -12510 44855 -12390
rect 44975 -12510 45030 -12390
rect 45150 -12510 45195 -12390
rect 45315 -12510 45360 -12390
rect 45480 -12510 45525 -12390
rect 45645 -12510 45700 -12390
rect 45820 -12510 45865 -12390
rect 45985 -12510 46030 -12390
rect 46150 -12510 46195 -12390
rect 46315 -12510 46370 -12390
rect 46490 -12510 46535 -12390
rect 46655 -12510 46700 -12390
rect 46820 -12510 46865 -12390
rect 46985 -12510 47040 -12390
rect 47160 -12510 47205 -12390
rect 47325 -12510 47370 -12390
rect 47490 -12510 47535 -12390
rect 47655 -12510 47865 -12390
rect 47985 -12510 48040 -12390
rect 48160 -12510 48205 -12390
rect 48325 -12510 48370 -12390
rect 48490 -12510 48535 -12390
rect 48655 -12510 48710 -12390
rect 48830 -12510 48875 -12390
rect 48995 -12510 49040 -12390
rect 49160 -12510 49205 -12390
rect 49325 -12510 49380 -12390
rect 49500 -12510 49545 -12390
rect 49665 -12510 49710 -12390
rect 49830 -12510 49875 -12390
rect 49995 -12510 50050 -12390
rect 50170 -12510 50215 -12390
rect 50335 -12510 50380 -12390
rect 50500 -12510 50545 -12390
rect 50665 -12510 50720 -12390
rect 50840 -12510 50885 -12390
rect 51005 -12510 51050 -12390
rect 51170 -12510 51215 -12390
rect 51335 -12510 51390 -12390
rect 51510 -12510 51555 -12390
rect 51675 -12510 51720 -12390
rect 51840 -12510 51885 -12390
rect 52005 -12510 52060 -12390
rect 52180 -12510 52225 -12390
rect 52345 -12510 52390 -12390
rect 52510 -12510 52555 -12390
rect 52675 -12510 52730 -12390
rect 52850 -12510 52895 -12390
rect 53015 -12510 53060 -12390
rect 53180 -12510 53225 -12390
rect 53345 -12510 53370 -12390
rect 30770 -12555 53370 -12510
rect 30770 -12675 30795 -12555
rect 30915 -12675 30970 -12555
rect 31090 -12675 31135 -12555
rect 31255 -12675 31300 -12555
rect 31420 -12675 31465 -12555
rect 31585 -12675 31640 -12555
rect 31760 -12675 31805 -12555
rect 31925 -12675 31970 -12555
rect 32090 -12675 32135 -12555
rect 32255 -12675 32310 -12555
rect 32430 -12675 32475 -12555
rect 32595 -12675 32640 -12555
rect 32760 -12675 32805 -12555
rect 32925 -12675 32980 -12555
rect 33100 -12675 33145 -12555
rect 33265 -12675 33310 -12555
rect 33430 -12675 33475 -12555
rect 33595 -12675 33650 -12555
rect 33770 -12675 33815 -12555
rect 33935 -12675 33980 -12555
rect 34100 -12675 34145 -12555
rect 34265 -12675 34320 -12555
rect 34440 -12675 34485 -12555
rect 34605 -12675 34650 -12555
rect 34770 -12675 34815 -12555
rect 34935 -12675 34990 -12555
rect 35110 -12675 35155 -12555
rect 35275 -12675 35320 -12555
rect 35440 -12675 35485 -12555
rect 35605 -12675 35660 -12555
rect 35780 -12675 35825 -12555
rect 35945 -12675 35990 -12555
rect 36110 -12675 36155 -12555
rect 36275 -12675 36485 -12555
rect 36605 -12675 36660 -12555
rect 36780 -12675 36825 -12555
rect 36945 -12675 36990 -12555
rect 37110 -12675 37155 -12555
rect 37275 -12675 37330 -12555
rect 37450 -12675 37495 -12555
rect 37615 -12675 37660 -12555
rect 37780 -12675 37825 -12555
rect 37945 -12675 38000 -12555
rect 38120 -12675 38165 -12555
rect 38285 -12675 38330 -12555
rect 38450 -12675 38495 -12555
rect 38615 -12675 38670 -12555
rect 38790 -12675 38835 -12555
rect 38955 -12675 39000 -12555
rect 39120 -12675 39165 -12555
rect 39285 -12675 39340 -12555
rect 39460 -12675 39505 -12555
rect 39625 -12675 39670 -12555
rect 39790 -12675 39835 -12555
rect 39955 -12675 40010 -12555
rect 40130 -12675 40175 -12555
rect 40295 -12675 40340 -12555
rect 40460 -12675 40505 -12555
rect 40625 -12675 40680 -12555
rect 40800 -12675 40845 -12555
rect 40965 -12675 41010 -12555
rect 41130 -12675 41175 -12555
rect 41295 -12675 41350 -12555
rect 41470 -12675 41515 -12555
rect 41635 -12675 41680 -12555
rect 41800 -12675 41845 -12555
rect 41965 -12675 42175 -12555
rect 42295 -12675 42350 -12555
rect 42470 -12675 42515 -12555
rect 42635 -12675 42680 -12555
rect 42800 -12675 42845 -12555
rect 42965 -12675 43020 -12555
rect 43140 -12675 43185 -12555
rect 43305 -12675 43350 -12555
rect 43470 -12675 43515 -12555
rect 43635 -12675 43690 -12555
rect 43810 -12675 43855 -12555
rect 43975 -12675 44020 -12555
rect 44140 -12675 44185 -12555
rect 44305 -12675 44360 -12555
rect 44480 -12675 44525 -12555
rect 44645 -12675 44690 -12555
rect 44810 -12675 44855 -12555
rect 44975 -12675 45030 -12555
rect 45150 -12675 45195 -12555
rect 45315 -12675 45360 -12555
rect 45480 -12675 45525 -12555
rect 45645 -12675 45700 -12555
rect 45820 -12675 45865 -12555
rect 45985 -12675 46030 -12555
rect 46150 -12675 46195 -12555
rect 46315 -12675 46370 -12555
rect 46490 -12675 46535 -12555
rect 46655 -12675 46700 -12555
rect 46820 -12675 46865 -12555
rect 46985 -12675 47040 -12555
rect 47160 -12675 47205 -12555
rect 47325 -12675 47370 -12555
rect 47490 -12675 47535 -12555
rect 47655 -12675 47865 -12555
rect 47985 -12675 48040 -12555
rect 48160 -12675 48205 -12555
rect 48325 -12675 48370 -12555
rect 48490 -12675 48535 -12555
rect 48655 -12675 48710 -12555
rect 48830 -12675 48875 -12555
rect 48995 -12675 49040 -12555
rect 49160 -12675 49205 -12555
rect 49325 -12675 49380 -12555
rect 49500 -12675 49545 -12555
rect 49665 -12675 49710 -12555
rect 49830 -12675 49875 -12555
rect 49995 -12675 50050 -12555
rect 50170 -12675 50215 -12555
rect 50335 -12675 50380 -12555
rect 50500 -12675 50545 -12555
rect 50665 -12675 50720 -12555
rect 50840 -12675 50885 -12555
rect 51005 -12675 51050 -12555
rect 51170 -12675 51215 -12555
rect 51335 -12675 51390 -12555
rect 51510 -12675 51555 -12555
rect 51675 -12675 51720 -12555
rect 51840 -12675 51885 -12555
rect 52005 -12675 52060 -12555
rect 52180 -12675 52225 -12555
rect 52345 -12675 52390 -12555
rect 52510 -12675 52555 -12555
rect 52675 -12675 52730 -12555
rect 52850 -12675 52895 -12555
rect 53015 -12675 53060 -12555
rect 53180 -12675 53225 -12555
rect 53345 -12675 53370 -12555
rect 30770 -12730 53370 -12675
rect 30770 -12850 30795 -12730
rect 30915 -12850 30970 -12730
rect 31090 -12850 31135 -12730
rect 31255 -12850 31300 -12730
rect 31420 -12850 31465 -12730
rect 31585 -12850 31640 -12730
rect 31760 -12850 31805 -12730
rect 31925 -12850 31970 -12730
rect 32090 -12850 32135 -12730
rect 32255 -12850 32310 -12730
rect 32430 -12850 32475 -12730
rect 32595 -12850 32640 -12730
rect 32760 -12850 32805 -12730
rect 32925 -12850 32980 -12730
rect 33100 -12850 33145 -12730
rect 33265 -12850 33310 -12730
rect 33430 -12850 33475 -12730
rect 33595 -12850 33650 -12730
rect 33770 -12850 33815 -12730
rect 33935 -12850 33980 -12730
rect 34100 -12850 34145 -12730
rect 34265 -12850 34320 -12730
rect 34440 -12850 34485 -12730
rect 34605 -12850 34650 -12730
rect 34770 -12850 34815 -12730
rect 34935 -12850 34990 -12730
rect 35110 -12850 35155 -12730
rect 35275 -12850 35320 -12730
rect 35440 -12850 35485 -12730
rect 35605 -12850 35660 -12730
rect 35780 -12850 35825 -12730
rect 35945 -12850 35990 -12730
rect 36110 -12850 36155 -12730
rect 36275 -12850 36485 -12730
rect 36605 -12850 36660 -12730
rect 36780 -12850 36825 -12730
rect 36945 -12850 36990 -12730
rect 37110 -12850 37155 -12730
rect 37275 -12850 37330 -12730
rect 37450 -12850 37495 -12730
rect 37615 -12850 37660 -12730
rect 37780 -12850 37825 -12730
rect 37945 -12850 38000 -12730
rect 38120 -12850 38165 -12730
rect 38285 -12850 38330 -12730
rect 38450 -12850 38495 -12730
rect 38615 -12850 38670 -12730
rect 38790 -12850 38835 -12730
rect 38955 -12850 39000 -12730
rect 39120 -12850 39165 -12730
rect 39285 -12850 39340 -12730
rect 39460 -12850 39505 -12730
rect 39625 -12850 39670 -12730
rect 39790 -12850 39835 -12730
rect 39955 -12850 40010 -12730
rect 40130 -12850 40175 -12730
rect 40295 -12850 40340 -12730
rect 40460 -12850 40505 -12730
rect 40625 -12850 40680 -12730
rect 40800 -12850 40845 -12730
rect 40965 -12850 41010 -12730
rect 41130 -12850 41175 -12730
rect 41295 -12850 41350 -12730
rect 41470 -12850 41515 -12730
rect 41635 -12850 41680 -12730
rect 41800 -12850 41845 -12730
rect 41965 -12850 42175 -12730
rect 42295 -12850 42350 -12730
rect 42470 -12850 42515 -12730
rect 42635 -12850 42680 -12730
rect 42800 -12850 42845 -12730
rect 42965 -12850 43020 -12730
rect 43140 -12850 43185 -12730
rect 43305 -12850 43350 -12730
rect 43470 -12850 43515 -12730
rect 43635 -12850 43690 -12730
rect 43810 -12850 43855 -12730
rect 43975 -12850 44020 -12730
rect 44140 -12850 44185 -12730
rect 44305 -12850 44360 -12730
rect 44480 -12850 44525 -12730
rect 44645 -12850 44690 -12730
rect 44810 -12850 44855 -12730
rect 44975 -12850 45030 -12730
rect 45150 -12850 45195 -12730
rect 45315 -12850 45360 -12730
rect 45480 -12850 45525 -12730
rect 45645 -12850 45700 -12730
rect 45820 -12850 45865 -12730
rect 45985 -12850 46030 -12730
rect 46150 -12850 46195 -12730
rect 46315 -12850 46370 -12730
rect 46490 -12850 46535 -12730
rect 46655 -12850 46700 -12730
rect 46820 -12850 46865 -12730
rect 46985 -12850 47040 -12730
rect 47160 -12850 47205 -12730
rect 47325 -12850 47370 -12730
rect 47490 -12850 47535 -12730
rect 47655 -12850 47865 -12730
rect 47985 -12850 48040 -12730
rect 48160 -12850 48205 -12730
rect 48325 -12850 48370 -12730
rect 48490 -12850 48535 -12730
rect 48655 -12850 48710 -12730
rect 48830 -12850 48875 -12730
rect 48995 -12850 49040 -12730
rect 49160 -12850 49205 -12730
rect 49325 -12850 49380 -12730
rect 49500 -12850 49545 -12730
rect 49665 -12850 49710 -12730
rect 49830 -12850 49875 -12730
rect 49995 -12850 50050 -12730
rect 50170 -12850 50215 -12730
rect 50335 -12850 50380 -12730
rect 50500 -12850 50545 -12730
rect 50665 -12850 50720 -12730
rect 50840 -12850 50885 -12730
rect 51005 -12850 51050 -12730
rect 51170 -12850 51215 -12730
rect 51335 -12850 51390 -12730
rect 51510 -12850 51555 -12730
rect 51675 -12850 51720 -12730
rect 51840 -12850 51885 -12730
rect 52005 -12850 52060 -12730
rect 52180 -12850 52225 -12730
rect 52345 -12850 52390 -12730
rect 52510 -12850 52555 -12730
rect 52675 -12850 52730 -12730
rect 52850 -12850 52895 -12730
rect 53015 -12850 53060 -12730
rect 53180 -12850 53225 -12730
rect 53345 -12850 53370 -12730
rect 30770 -12895 53370 -12850
rect 30770 -13015 30795 -12895
rect 30915 -13015 30970 -12895
rect 31090 -13015 31135 -12895
rect 31255 -13015 31300 -12895
rect 31420 -13015 31465 -12895
rect 31585 -13015 31640 -12895
rect 31760 -13015 31805 -12895
rect 31925 -13015 31970 -12895
rect 32090 -13015 32135 -12895
rect 32255 -13015 32310 -12895
rect 32430 -13015 32475 -12895
rect 32595 -13015 32640 -12895
rect 32760 -13015 32805 -12895
rect 32925 -13015 32980 -12895
rect 33100 -13015 33145 -12895
rect 33265 -13015 33310 -12895
rect 33430 -13015 33475 -12895
rect 33595 -13015 33650 -12895
rect 33770 -13015 33815 -12895
rect 33935 -13015 33980 -12895
rect 34100 -13015 34145 -12895
rect 34265 -13015 34320 -12895
rect 34440 -13015 34485 -12895
rect 34605 -13015 34650 -12895
rect 34770 -13015 34815 -12895
rect 34935 -13015 34990 -12895
rect 35110 -13015 35155 -12895
rect 35275 -13015 35320 -12895
rect 35440 -13015 35485 -12895
rect 35605 -13015 35660 -12895
rect 35780 -13015 35825 -12895
rect 35945 -13015 35990 -12895
rect 36110 -13015 36155 -12895
rect 36275 -13015 36485 -12895
rect 36605 -13015 36660 -12895
rect 36780 -13015 36825 -12895
rect 36945 -13015 36990 -12895
rect 37110 -13015 37155 -12895
rect 37275 -13015 37330 -12895
rect 37450 -13015 37495 -12895
rect 37615 -13015 37660 -12895
rect 37780 -13015 37825 -12895
rect 37945 -13015 38000 -12895
rect 38120 -13015 38165 -12895
rect 38285 -13015 38330 -12895
rect 38450 -13015 38495 -12895
rect 38615 -13015 38670 -12895
rect 38790 -13015 38835 -12895
rect 38955 -13015 39000 -12895
rect 39120 -13015 39165 -12895
rect 39285 -13015 39340 -12895
rect 39460 -13015 39505 -12895
rect 39625 -13015 39670 -12895
rect 39790 -13015 39835 -12895
rect 39955 -13015 40010 -12895
rect 40130 -13015 40175 -12895
rect 40295 -13015 40340 -12895
rect 40460 -13015 40505 -12895
rect 40625 -13015 40680 -12895
rect 40800 -13015 40845 -12895
rect 40965 -13015 41010 -12895
rect 41130 -13015 41175 -12895
rect 41295 -13015 41350 -12895
rect 41470 -13015 41515 -12895
rect 41635 -13015 41680 -12895
rect 41800 -13015 41845 -12895
rect 41965 -13015 42175 -12895
rect 42295 -13015 42350 -12895
rect 42470 -13015 42515 -12895
rect 42635 -13015 42680 -12895
rect 42800 -13015 42845 -12895
rect 42965 -13015 43020 -12895
rect 43140 -13015 43185 -12895
rect 43305 -13015 43350 -12895
rect 43470 -13015 43515 -12895
rect 43635 -13015 43690 -12895
rect 43810 -13015 43855 -12895
rect 43975 -13015 44020 -12895
rect 44140 -13015 44185 -12895
rect 44305 -13015 44360 -12895
rect 44480 -13015 44525 -12895
rect 44645 -13015 44690 -12895
rect 44810 -13015 44855 -12895
rect 44975 -13015 45030 -12895
rect 45150 -13015 45195 -12895
rect 45315 -13015 45360 -12895
rect 45480 -13015 45525 -12895
rect 45645 -13015 45700 -12895
rect 45820 -13015 45865 -12895
rect 45985 -13015 46030 -12895
rect 46150 -13015 46195 -12895
rect 46315 -13015 46370 -12895
rect 46490 -13015 46535 -12895
rect 46655 -13015 46700 -12895
rect 46820 -13015 46865 -12895
rect 46985 -13015 47040 -12895
rect 47160 -13015 47205 -12895
rect 47325 -13015 47370 -12895
rect 47490 -13015 47535 -12895
rect 47655 -13015 47865 -12895
rect 47985 -13015 48040 -12895
rect 48160 -13015 48205 -12895
rect 48325 -13015 48370 -12895
rect 48490 -13015 48535 -12895
rect 48655 -13015 48710 -12895
rect 48830 -13015 48875 -12895
rect 48995 -13015 49040 -12895
rect 49160 -13015 49205 -12895
rect 49325 -13015 49380 -12895
rect 49500 -13015 49545 -12895
rect 49665 -13015 49710 -12895
rect 49830 -13015 49875 -12895
rect 49995 -13015 50050 -12895
rect 50170 -13015 50215 -12895
rect 50335 -13015 50380 -12895
rect 50500 -13015 50545 -12895
rect 50665 -13015 50720 -12895
rect 50840 -13015 50885 -12895
rect 51005 -13015 51050 -12895
rect 51170 -13015 51215 -12895
rect 51335 -13015 51390 -12895
rect 51510 -13015 51555 -12895
rect 51675 -13015 51720 -12895
rect 51840 -13015 51885 -12895
rect 52005 -13015 52060 -12895
rect 52180 -13015 52225 -12895
rect 52345 -13015 52390 -12895
rect 52510 -13015 52555 -12895
rect 52675 -13015 52730 -12895
rect 52850 -13015 52895 -12895
rect 53015 -13015 53060 -12895
rect 53180 -13015 53225 -12895
rect 53345 -13015 53370 -12895
rect 30770 -13060 53370 -13015
rect 30770 -13180 30795 -13060
rect 30915 -13180 30970 -13060
rect 31090 -13180 31135 -13060
rect 31255 -13180 31300 -13060
rect 31420 -13180 31465 -13060
rect 31585 -13180 31640 -13060
rect 31760 -13180 31805 -13060
rect 31925 -13180 31970 -13060
rect 32090 -13180 32135 -13060
rect 32255 -13180 32310 -13060
rect 32430 -13180 32475 -13060
rect 32595 -13180 32640 -13060
rect 32760 -13180 32805 -13060
rect 32925 -13180 32980 -13060
rect 33100 -13180 33145 -13060
rect 33265 -13180 33310 -13060
rect 33430 -13180 33475 -13060
rect 33595 -13180 33650 -13060
rect 33770 -13180 33815 -13060
rect 33935 -13180 33980 -13060
rect 34100 -13180 34145 -13060
rect 34265 -13180 34320 -13060
rect 34440 -13180 34485 -13060
rect 34605 -13180 34650 -13060
rect 34770 -13180 34815 -13060
rect 34935 -13180 34990 -13060
rect 35110 -13180 35155 -13060
rect 35275 -13180 35320 -13060
rect 35440 -13180 35485 -13060
rect 35605 -13180 35660 -13060
rect 35780 -13180 35825 -13060
rect 35945 -13180 35990 -13060
rect 36110 -13180 36155 -13060
rect 36275 -13180 36485 -13060
rect 36605 -13180 36660 -13060
rect 36780 -13180 36825 -13060
rect 36945 -13180 36990 -13060
rect 37110 -13180 37155 -13060
rect 37275 -13180 37330 -13060
rect 37450 -13180 37495 -13060
rect 37615 -13180 37660 -13060
rect 37780 -13180 37825 -13060
rect 37945 -13180 38000 -13060
rect 38120 -13180 38165 -13060
rect 38285 -13180 38330 -13060
rect 38450 -13180 38495 -13060
rect 38615 -13180 38670 -13060
rect 38790 -13180 38835 -13060
rect 38955 -13180 39000 -13060
rect 39120 -13180 39165 -13060
rect 39285 -13180 39340 -13060
rect 39460 -13180 39505 -13060
rect 39625 -13180 39670 -13060
rect 39790 -13180 39835 -13060
rect 39955 -13180 40010 -13060
rect 40130 -13180 40175 -13060
rect 40295 -13180 40340 -13060
rect 40460 -13180 40505 -13060
rect 40625 -13180 40680 -13060
rect 40800 -13180 40845 -13060
rect 40965 -13180 41010 -13060
rect 41130 -13180 41175 -13060
rect 41295 -13180 41350 -13060
rect 41470 -13180 41515 -13060
rect 41635 -13180 41680 -13060
rect 41800 -13180 41845 -13060
rect 41965 -13180 42175 -13060
rect 42295 -13180 42350 -13060
rect 42470 -13180 42515 -13060
rect 42635 -13180 42680 -13060
rect 42800 -13180 42845 -13060
rect 42965 -13180 43020 -13060
rect 43140 -13180 43185 -13060
rect 43305 -13180 43350 -13060
rect 43470 -13180 43515 -13060
rect 43635 -13180 43690 -13060
rect 43810 -13180 43855 -13060
rect 43975 -13180 44020 -13060
rect 44140 -13180 44185 -13060
rect 44305 -13180 44360 -13060
rect 44480 -13180 44525 -13060
rect 44645 -13180 44690 -13060
rect 44810 -13180 44855 -13060
rect 44975 -13180 45030 -13060
rect 45150 -13180 45195 -13060
rect 45315 -13180 45360 -13060
rect 45480 -13180 45525 -13060
rect 45645 -13180 45700 -13060
rect 45820 -13180 45865 -13060
rect 45985 -13180 46030 -13060
rect 46150 -13180 46195 -13060
rect 46315 -13180 46370 -13060
rect 46490 -13180 46535 -13060
rect 46655 -13180 46700 -13060
rect 46820 -13180 46865 -13060
rect 46985 -13180 47040 -13060
rect 47160 -13180 47205 -13060
rect 47325 -13180 47370 -13060
rect 47490 -13180 47535 -13060
rect 47655 -13180 47865 -13060
rect 47985 -13180 48040 -13060
rect 48160 -13180 48205 -13060
rect 48325 -13180 48370 -13060
rect 48490 -13180 48535 -13060
rect 48655 -13180 48710 -13060
rect 48830 -13180 48875 -13060
rect 48995 -13180 49040 -13060
rect 49160 -13180 49205 -13060
rect 49325 -13180 49380 -13060
rect 49500 -13180 49545 -13060
rect 49665 -13180 49710 -13060
rect 49830 -13180 49875 -13060
rect 49995 -13180 50050 -13060
rect 50170 -13180 50215 -13060
rect 50335 -13180 50380 -13060
rect 50500 -13180 50545 -13060
rect 50665 -13180 50720 -13060
rect 50840 -13180 50885 -13060
rect 51005 -13180 51050 -13060
rect 51170 -13180 51215 -13060
rect 51335 -13180 51390 -13060
rect 51510 -13180 51555 -13060
rect 51675 -13180 51720 -13060
rect 51840 -13180 51885 -13060
rect 52005 -13180 52060 -13060
rect 52180 -13180 52225 -13060
rect 52345 -13180 52390 -13060
rect 52510 -13180 52555 -13060
rect 52675 -13180 52730 -13060
rect 52850 -13180 52895 -13060
rect 53015 -13180 53060 -13060
rect 53180 -13180 53225 -13060
rect 53345 -13180 53370 -13060
rect 30770 -13225 53370 -13180
rect 30770 -13345 30795 -13225
rect 30915 -13345 30970 -13225
rect 31090 -13345 31135 -13225
rect 31255 -13345 31300 -13225
rect 31420 -13345 31465 -13225
rect 31585 -13345 31640 -13225
rect 31760 -13345 31805 -13225
rect 31925 -13345 31970 -13225
rect 32090 -13345 32135 -13225
rect 32255 -13345 32310 -13225
rect 32430 -13345 32475 -13225
rect 32595 -13345 32640 -13225
rect 32760 -13345 32805 -13225
rect 32925 -13345 32980 -13225
rect 33100 -13345 33145 -13225
rect 33265 -13345 33310 -13225
rect 33430 -13345 33475 -13225
rect 33595 -13345 33650 -13225
rect 33770 -13345 33815 -13225
rect 33935 -13345 33980 -13225
rect 34100 -13345 34145 -13225
rect 34265 -13345 34320 -13225
rect 34440 -13345 34485 -13225
rect 34605 -13345 34650 -13225
rect 34770 -13345 34815 -13225
rect 34935 -13345 34990 -13225
rect 35110 -13345 35155 -13225
rect 35275 -13345 35320 -13225
rect 35440 -13345 35485 -13225
rect 35605 -13345 35660 -13225
rect 35780 -13345 35825 -13225
rect 35945 -13345 35990 -13225
rect 36110 -13345 36155 -13225
rect 36275 -13345 36485 -13225
rect 36605 -13345 36660 -13225
rect 36780 -13345 36825 -13225
rect 36945 -13345 36990 -13225
rect 37110 -13345 37155 -13225
rect 37275 -13345 37330 -13225
rect 37450 -13345 37495 -13225
rect 37615 -13345 37660 -13225
rect 37780 -13345 37825 -13225
rect 37945 -13345 38000 -13225
rect 38120 -13345 38165 -13225
rect 38285 -13345 38330 -13225
rect 38450 -13345 38495 -13225
rect 38615 -13345 38670 -13225
rect 38790 -13345 38835 -13225
rect 38955 -13345 39000 -13225
rect 39120 -13345 39165 -13225
rect 39285 -13345 39340 -13225
rect 39460 -13345 39505 -13225
rect 39625 -13345 39670 -13225
rect 39790 -13345 39835 -13225
rect 39955 -13345 40010 -13225
rect 40130 -13345 40175 -13225
rect 40295 -13345 40340 -13225
rect 40460 -13345 40505 -13225
rect 40625 -13345 40680 -13225
rect 40800 -13345 40845 -13225
rect 40965 -13345 41010 -13225
rect 41130 -13345 41175 -13225
rect 41295 -13345 41350 -13225
rect 41470 -13345 41515 -13225
rect 41635 -13345 41680 -13225
rect 41800 -13345 41845 -13225
rect 41965 -13345 42175 -13225
rect 42295 -13345 42350 -13225
rect 42470 -13345 42515 -13225
rect 42635 -13345 42680 -13225
rect 42800 -13345 42845 -13225
rect 42965 -13345 43020 -13225
rect 43140 -13345 43185 -13225
rect 43305 -13345 43350 -13225
rect 43470 -13345 43515 -13225
rect 43635 -13345 43690 -13225
rect 43810 -13345 43855 -13225
rect 43975 -13345 44020 -13225
rect 44140 -13345 44185 -13225
rect 44305 -13345 44360 -13225
rect 44480 -13345 44525 -13225
rect 44645 -13345 44690 -13225
rect 44810 -13345 44855 -13225
rect 44975 -13345 45030 -13225
rect 45150 -13345 45195 -13225
rect 45315 -13345 45360 -13225
rect 45480 -13345 45525 -13225
rect 45645 -13345 45700 -13225
rect 45820 -13345 45865 -13225
rect 45985 -13345 46030 -13225
rect 46150 -13345 46195 -13225
rect 46315 -13345 46370 -13225
rect 46490 -13345 46535 -13225
rect 46655 -13345 46700 -13225
rect 46820 -13345 46865 -13225
rect 46985 -13345 47040 -13225
rect 47160 -13345 47205 -13225
rect 47325 -13345 47370 -13225
rect 47490 -13345 47535 -13225
rect 47655 -13345 47865 -13225
rect 47985 -13345 48040 -13225
rect 48160 -13345 48205 -13225
rect 48325 -13345 48370 -13225
rect 48490 -13345 48535 -13225
rect 48655 -13345 48710 -13225
rect 48830 -13345 48875 -13225
rect 48995 -13345 49040 -13225
rect 49160 -13345 49205 -13225
rect 49325 -13345 49380 -13225
rect 49500 -13345 49545 -13225
rect 49665 -13345 49710 -13225
rect 49830 -13345 49875 -13225
rect 49995 -13345 50050 -13225
rect 50170 -13345 50215 -13225
rect 50335 -13345 50380 -13225
rect 50500 -13345 50545 -13225
rect 50665 -13345 50720 -13225
rect 50840 -13345 50885 -13225
rect 51005 -13345 51050 -13225
rect 51170 -13345 51215 -13225
rect 51335 -13345 51390 -13225
rect 51510 -13345 51555 -13225
rect 51675 -13345 51720 -13225
rect 51840 -13345 51885 -13225
rect 52005 -13345 52060 -13225
rect 52180 -13345 52225 -13225
rect 52345 -13345 52390 -13225
rect 52510 -13345 52555 -13225
rect 52675 -13345 52730 -13225
rect 52850 -13345 52895 -13225
rect 53015 -13345 53060 -13225
rect 53180 -13345 53225 -13225
rect 53345 -13345 53370 -13225
rect 30770 -13400 53370 -13345
rect 30770 -13520 30795 -13400
rect 30915 -13520 30970 -13400
rect 31090 -13520 31135 -13400
rect 31255 -13520 31300 -13400
rect 31420 -13520 31465 -13400
rect 31585 -13520 31640 -13400
rect 31760 -13520 31805 -13400
rect 31925 -13520 31970 -13400
rect 32090 -13520 32135 -13400
rect 32255 -13520 32310 -13400
rect 32430 -13520 32475 -13400
rect 32595 -13520 32640 -13400
rect 32760 -13520 32805 -13400
rect 32925 -13520 32980 -13400
rect 33100 -13520 33145 -13400
rect 33265 -13520 33310 -13400
rect 33430 -13520 33475 -13400
rect 33595 -13520 33650 -13400
rect 33770 -13520 33815 -13400
rect 33935 -13520 33980 -13400
rect 34100 -13520 34145 -13400
rect 34265 -13520 34320 -13400
rect 34440 -13520 34485 -13400
rect 34605 -13520 34650 -13400
rect 34770 -13520 34815 -13400
rect 34935 -13520 34990 -13400
rect 35110 -13520 35155 -13400
rect 35275 -13520 35320 -13400
rect 35440 -13520 35485 -13400
rect 35605 -13520 35660 -13400
rect 35780 -13520 35825 -13400
rect 35945 -13520 35990 -13400
rect 36110 -13520 36155 -13400
rect 36275 -13520 36485 -13400
rect 36605 -13520 36660 -13400
rect 36780 -13520 36825 -13400
rect 36945 -13520 36990 -13400
rect 37110 -13520 37155 -13400
rect 37275 -13520 37330 -13400
rect 37450 -13520 37495 -13400
rect 37615 -13520 37660 -13400
rect 37780 -13520 37825 -13400
rect 37945 -13520 38000 -13400
rect 38120 -13520 38165 -13400
rect 38285 -13520 38330 -13400
rect 38450 -13520 38495 -13400
rect 38615 -13520 38670 -13400
rect 38790 -13520 38835 -13400
rect 38955 -13520 39000 -13400
rect 39120 -13520 39165 -13400
rect 39285 -13520 39340 -13400
rect 39460 -13520 39505 -13400
rect 39625 -13520 39670 -13400
rect 39790 -13520 39835 -13400
rect 39955 -13520 40010 -13400
rect 40130 -13520 40175 -13400
rect 40295 -13520 40340 -13400
rect 40460 -13520 40505 -13400
rect 40625 -13520 40680 -13400
rect 40800 -13520 40845 -13400
rect 40965 -13520 41010 -13400
rect 41130 -13520 41175 -13400
rect 41295 -13520 41350 -13400
rect 41470 -13520 41515 -13400
rect 41635 -13520 41680 -13400
rect 41800 -13520 41845 -13400
rect 41965 -13520 42175 -13400
rect 42295 -13520 42350 -13400
rect 42470 -13520 42515 -13400
rect 42635 -13520 42680 -13400
rect 42800 -13520 42845 -13400
rect 42965 -13520 43020 -13400
rect 43140 -13520 43185 -13400
rect 43305 -13520 43350 -13400
rect 43470 -13520 43515 -13400
rect 43635 -13520 43690 -13400
rect 43810 -13520 43855 -13400
rect 43975 -13520 44020 -13400
rect 44140 -13520 44185 -13400
rect 44305 -13520 44360 -13400
rect 44480 -13520 44525 -13400
rect 44645 -13520 44690 -13400
rect 44810 -13520 44855 -13400
rect 44975 -13520 45030 -13400
rect 45150 -13520 45195 -13400
rect 45315 -13520 45360 -13400
rect 45480 -13520 45525 -13400
rect 45645 -13520 45700 -13400
rect 45820 -13520 45865 -13400
rect 45985 -13520 46030 -13400
rect 46150 -13520 46195 -13400
rect 46315 -13520 46370 -13400
rect 46490 -13520 46535 -13400
rect 46655 -13520 46700 -13400
rect 46820 -13520 46865 -13400
rect 46985 -13520 47040 -13400
rect 47160 -13520 47205 -13400
rect 47325 -13520 47370 -13400
rect 47490 -13520 47535 -13400
rect 47655 -13520 47865 -13400
rect 47985 -13520 48040 -13400
rect 48160 -13520 48205 -13400
rect 48325 -13520 48370 -13400
rect 48490 -13520 48535 -13400
rect 48655 -13520 48710 -13400
rect 48830 -13520 48875 -13400
rect 48995 -13520 49040 -13400
rect 49160 -13520 49205 -13400
rect 49325 -13520 49380 -13400
rect 49500 -13520 49545 -13400
rect 49665 -13520 49710 -13400
rect 49830 -13520 49875 -13400
rect 49995 -13520 50050 -13400
rect 50170 -13520 50215 -13400
rect 50335 -13520 50380 -13400
rect 50500 -13520 50545 -13400
rect 50665 -13520 50720 -13400
rect 50840 -13520 50885 -13400
rect 51005 -13520 51050 -13400
rect 51170 -13520 51215 -13400
rect 51335 -13520 51390 -13400
rect 51510 -13520 51555 -13400
rect 51675 -13520 51720 -13400
rect 51840 -13520 51885 -13400
rect 52005 -13520 52060 -13400
rect 52180 -13520 52225 -13400
rect 52345 -13520 52390 -13400
rect 52510 -13520 52555 -13400
rect 52675 -13520 52730 -13400
rect 52850 -13520 52895 -13400
rect 53015 -13520 53060 -13400
rect 53180 -13520 53225 -13400
rect 53345 -13520 53370 -13400
rect 30770 -13565 53370 -13520
rect 30770 -13685 30795 -13565
rect 30915 -13685 30970 -13565
rect 31090 -13685 31135 -13565
rect 31255 -13685 31300 -13565
rect 31420 -13685 31465 -13565
rect 31585 -13685 31640 -13565
rect 31760 -13685 31805 -13565
rect 31925 -13685 31970 -13565
rect 32090 -13685 32135 -13565
rect 32255 -13685 32310 -13565
rect 32430 -13685 32475 -13565
rect 32595 -13685 32640 -13565
rect 32760 -13685 32805 -13565
rect 32925 -13685 32980 -13565
rect 33100 -13685 33145 -13565
rect 33265 -13685 33310 -13565
rect 33430 -13685 33475 -13565
rect 33595 -13685 33650 -13565
rect 33770 -13685 33815 -13565
rect 33935 -13685 33980 -13565
rect 34100 -13685 34145 -13565
rect 34265 -13685 34320 -13565
rect 34440 -13685 34485 -13565
rect 34605 -13685 34650 -13565
rect 34770 -13685 34815 -13565
rect 34935 -13685 34990 -13565
rect 35110 -13685 35155 -13565
rect 35275 -13685 35320 -13565
rect 35440 -13685 35485 -13565
rect 35605 -13685 35660 -13565
rect 35780 -13685 35825 -13565
rect 35945 -13685 35990 -13565
rect 36110 -13685 36155 -13565
rect 36275 -13685 36485 -13565
rect 36605 -13685 36660 -13565
rect 36780 -13685 36825 -13565
rect 36945 -13685 36990 -13565
rect 37110 -13685 37155 -13565
rect 37275 -13685 37330 -13565
rect 37450 -13685 37495 -13565
rect 37615 -13685 37660 -13565
rect 37780 -13685 37825 -13565
rect 37945 -13685 38000 -13565
rect 38120 -13685 38165 -13565
rect 38285 -13685 38330 -13565
rect 38450 -13685 38495 -13565
rect 38615 -13685 38670 -13565
rect 38790 -13685 38835 -13565
rect 38955 -13685 39000 -13565
rect 39120 -13685 39165 -13565
rect 39285 -13685 39340 -13565
rect 39460 -13685 39505 -13565
rect 39625 -13685 39670 -13565
rect 39790 -13685 39835 -13565
rect 39955 -13685 40010 -13565
rect 40130 -13685 40175 -13565
rect 40295 -13685 40340 -13565
rect 40460 -13685 40505 -13565
rect 40625 -13685 40680 -13565
rect 40800 -13685 40845 -13565
rect 40965 -13685 41010 -13565
rect 41130 -13685 41175 -13565
rect 41295 -13685 41350 -13565
rect 41470 -13685 41515 -13565
rect 41635 -13685 41680 -13565
rect 41800 -13685 41845 -13565
rect 41965 -13685 42175 -13565
rect 42295 -13685 42350 -13565
rect 42470 -13685 42515 -13565
rect 42635 -13685 42680 -13565
rect 42800 -13685 42845 -13565
rect 42965 -13685 43020 -13565
rect 43140 -13685 43185 -13565
rect 43305 -13685 43350 -13565
rect 43470 -13685 43515 -13565
rect 43635 -13685 43690 -13565
rect 43810 -13685 43855 -13565
rect 43975 -13685 44020 -13565
rect 44140 -13685 44185 -13565
rect 44305 -13685 44360 -13565
rect 44480 -13685 44525 -13565
rect 44645 -13685 44690 -13565
rect 44810 -13685 44855 -13565
rect 44975 -13685 45030 -13565
rect 45150 -13685 45195 -13565
rect 45315 -13685 45360 -13565
rect 45480 -13685 45525 -13565
rect 45645 -13685 45700 -13565
rect 45820 -13685 45865 -13565
rect 45985 -13685 46030 -13565
rect 46150 -13685 46195 -13565
rect 46315 -13685 46370 -13565
rect 46490 -13685 46535 -13565
rect 46655 -13685 46700 -13565
rect 46820 -13685 46865 -13565
rect 46985 -13685 47040 -13565
rect 47160 -13685 47205 -13565
rect 47325 -13685 47370 -13565
rect 47490 -13685 47535 -13565
rect 47655 -13685 47865 -13565
rect 47985 -13685 48040 -13565
rect 48160 -13685 48205 -13565
rect 48325 -13685 48370 -13565
rect 48490 -13685 48535 -13565
rect 48655 -13685 48710 -13565
rect 48830 -13685 48875 -13565
rect 48995 -13685 49040 -13565
rect 49160 -13685 49205 -13565
rect 49325 -13685 49380 -13565
rect 49500 -13685 49545 -13565
rect 49665 -13685 49710 -13565
rect 49830 -13685 49875 -13565
rect 49995 -13685 50050 -13565
rect 50170 -13685 50215 -13565
rect 50335 -13685 50380 -13565
rect 50500 -13685 50545 -13565
rect 50665 -13685 50720 -13565
rect 50840 -13685 50885 -13565
rect 51005 -13685 51050 -13565
rect 51170 -13685 51215 -13565
rect 51335 -13685 51390 -13565
rect 51510 -13685 51555 -13565
rect 51675 -13685 51720 -13565
rect 51840 -13685 51885 -13565
rect 52005 -13685 52060 -13565
rect 52180 -13685 52225 -13565
rect 52345 -13685 52390 -13565
rect 52510 -13685 52555 -13565
rect 52675 -13685 52730 -13565
rect 52850 -13685 52895 -13565
rect 53015 -13685 53060 -13565
rect 53180 -13685 53225 -13565
rect 53345 -13685 53370 -13565
rect 30770 -13730 53370 -13685
rect 30770 -13850 30795 -13730
rect 30915 -13850 30970 -13730
rect 31090 -13850 31135 -13730
rect 31255 -13850 31300 -13730
rect 31420 -13850 31465 -13730
rect 31585 -13850 31640 -13730
rect 31760 -13850 31805 -13730
rect 31925 -13850 31970 -13730
rect 32090 -13850 32135 -13730
rect 32255 -13850 32310 -13730
rect 32430 -13850 32475 -13730
rect 32595 -13850 32640 -13730
rect 32760 -13850 32805 -13730
rect 32925 -13850 32980 -13730
rect 33100 -13850 33145 -13730
rect 33265 -13850 33310 -13730
rect 33430 -13850 33475 -13730
rect 33595 -13850 33650 -13730
rect 33770 -13850 33815 -13730
rect 33935 -13850 33980 -13730
rect 34100 -13850 34145 -13730
rect 34265 -13850 34320 -13730
rect 34440 -13850 34485 -13730
rect 34605 -13850 34650 -13730
rect 34770 -13850 34815 -13730
rect 34935 -13850 34990 -13730
rect 35110 -13850 35155 -13730
rect 35275 -13850 35320 -13730
rect 35440 -13850 35485 -13730
rect 35605 -13850 35660 -13730
rect 35780 -13850 35825 -13730
rect 35945 -13850 35990 -13730
rect 36110 -13850 36155 -13730
rect 36275 -13850 36485 -13730
rect 36605 -13850 36660 -13730
rect 36780 -13850 36825 -13730
rect 36945 -13850 36990 -13730
rect 37110 -13850 37155 -13730
rect 37275 -13850 37330 -13730
rect 37450 -13850 37495 -13730
rect 37615 -13850 37660 -13730
rect 37780 -13850 37825 -13730
rect 37945 -13850 38000 -13730
rect 38120 -13850 38165 -13730
rect 38285 -13850 38330 -13730
rect 38450 -13850 38495 -13730
rect 38615 -13850 38670 -13730
rect 38790 -13850 38835 -13730
rect 38955 -13850 39000 -13730
rect 39120 -13850 39165 -13730
rect 39285 -13850 39340 -13730
rect 39460 -13850 39505 -13730
rect 39625 -13850 39670 -13730
rect 39790 -13850 39835 -13730
rect 39955 -13850 40010 -13730
rect 40130 -13850 40175 -13730
rect 40295 -13850 40340 -13730
rect 40460 -13850 40505 -13730
rect 40625 -13850 40680 -13730
rect 40800 -13850 40845 -13730
rect 40965 -13850 41010 -13730
rect 41130 -13850 41175 -13730
rect 41295 -13850 41350 -13730
rect 41470 -13850 41515 -13730
rect 41635 -13850 41680 -13730
rect 41800 -13850 41845 -13730
rect 41965 -13850 42175 -13730
rect 42295 -13850 42350 -13730
rect 42470 -13850 42515 -13730
rect 42635 -13850 42680 -13730
rect 42800 -13850 42845 -13730
rect 42965 -13850 43020 -13730
rect 43140 -13850 43185 -13730
rect 43305 -13850 43350 -13730
rect 43470 -13850 43515 -13730
rect 43635 -13850 43690 -13730
rect 43810 -13850 43855 -13730
rect 43975 -13850 44020 -13730
rect 44140 -13850 44185 -13730
rect 44305 -13850 44360 -13730
rect 44480 -13850 44525 -13730
rect 44645 -13850 44690 -13730
rect 44810 -13850 44855 -13730
rect 44975 -13850 45030 -13730
rect 45150 -13850 45195 -13730
rect 45315 -13850 45360 -13730
rect 45480 -13850 45525 -13730
rect 45645 -13850 45700 -13730
rect 45820 -13850 45865 -13730
rect 45985 -13850 46030 -13730
rect 46150 -13850 46195 -13730
rect 46315 -13850 46370 -13730
rect 46490 -13850 46535 -13730
rect 46655 -13850 46700 -13730
rect 46820 -13850 46865 -13730
rect 46985 -13850 47040 -13730
rect 47160 -13850 47205 -13730
rect 47325 -13850 47370 -13730
rect 47490 -13850 47535 -13730
rect 47655 -13850 47865 -13730
rect 47985 -13850 48040 -13730
rect 48160 -13850 48205 -13730
rect 48325 -13850 48370 -13730
rect 48490 -13850 48535 -13730
rect 48655 -13850 48710 -13730
rect 48830 -13850 48875 -13730
rect 48995 -13850 49040 -13730
rect 49160 -13850 49205 -13730
rect 49325 -13850 49380 -13730
rect 49500 -13850 49545 -13730
rect 49665 -13850 49710 -13730
rect 49830 -13850 49875 -13730
rect 49995 -13850 50050 -13730
rect 50170 -13850 50215 -13730
rect 50335 -13850 50380 -13730
rect 50500 -13850 50545 -13730
rect 50665 -13850 50720 -13730
rect 50840 -13850 50885 -13730
rect 51005 -13850 51050 -13730
rect 51170 -13850 51215 -13730
rect 51335 -13850 51390 -13730
rect 51510 -13850 51555 -13730
rect 51675 -13850 51720 -13730
rect 51840 -13850 51885 -13730
rect 52005 -13850 52060 -13730
rect 52180 -13850 52225 -13730
rect 52345 -13850 52390 -13730
rect 52510 -13850 52555 -13730
rect 52675 -13850 52730 -13730
rect 52850 -13850 52895 -13730
rect 53015 -13850 53060 -13730
rect 53180 -13850 53225 -13730
rect 53345 -13850 53370 -13730
rect 30770 -13895 53370 -13850
rect 30770 -14015 30795 -13895
rect 30915 -14015 30970 -13895
rect 31090 -14015 31135 -13895
rect 31255 -14015 31300 -13895
rect 31420 -14015 31465 -13895
rect 31585 -14015 31640 -13895
rect 31760 -14015 31805 -13895
rect 31925 -14015 31970 -13895
rect 32090 -14015 32135 -13895
rect 32255 -14015 32310 -13895
rect 32430 -14015 32475 -13895
rect 32595 -14015 32640 -13895
rect 32760 -14015 32805 -13895
rect 32925 -14015 32980 -13895
rect 33100 -14015 33145 -13895
rect 33265 -14015 33310 -13895
rect 33430 -14015 33475 -13895
rect 33595 -14015 33650 -13895
rect 33770 -14015 33815 -13895
rect 33935 -14015 33980 -13895
rect 34100 -14015 34145 -13895
rect 34265 -14015 34320 -13895
rect 34440 -14015 34485 -13895
rect 34605 -14015 34650 -13895
rect 34770 -14015 34815 -13895
rect 34935 -14015 34990 -13895
rect 35110 -14015 35155 -13895
rect 35275 -14015 35320 -13895
rect 35440 -14015 35485 -13895
rect 35605 -14015 35660 -13895
rect 35780 -14015 35825 -13895
rect 35945 -14015 35990 -13895
rect 36110 -14015 36155 -13895
rect 36275 -14015 36485 -13895
rect 36605 -14015 36660 -13895
rect 36780 -14015 36825 -13895
rect 36945 -14015 36990 -13895
rect 37110 -14015 37155 -13895
rect 37275 -14015 37330 -13895
rect 37450 -14015 37495 -13895
rect 37615 -14015 37660 -13895
rect 37780 -14015 37825 -13895
rect 37945 -14015 38000 -13895
rect 38120 -14015 38165 -13895
rect 38285 -14015 38330 -13895
rect 38450 -14015 38495 -13895
rect 38615 -14015 38670 -13895
rect 38790 -14015 38835 -13895
rect 38955 -14015 39000 -13895
rect 39120 -14015 39165 -13895
rect 39285 -14015 39340 -13895
rect 39460 -14015 39505 -13895
rect 39625 -14015 39670 -13895
rect 39790 -14015 39835 -13895
rect 39955 -14015 40010 -13895
rect 40130 -14015 40175 -13895
rect 40295 -14015 40340 -13895
rect 40460 -14015 40505 -13895
rect 40625 -14015 40680 -13895
rect 40800 -14015 40845 -13895
rect 40965 -14015 41010 -13895
rect 41130 -14015 41175 -13895
rect 41295 -14015 41350 -13895
rect 41470 -14015 41515 -13895
rect 41635 -14015 41680 -13895
rect 41800 -14015 41845 -13895
rect 41965 -14015 42175 -13895
rect 42295 -14015 42350 -13895
rect 42470 -14015 42515 -13895
rect 42635 -14015 42680 -13895
rect 42800 -14015 42845 -13895
rect 42965 -14015 43020 -13895
rect 43140 -14015 43185 -13895
rect 43305 -14015 43350 -13895
rect 43470 -14015 43515 -13895
rect 43635 -14015 43690 -13895
rect 43810 -14015 43855 -13895
rect 43975 -14015 44020 -13895
rect 44140 -14015 44185 -13895
rect 44305 -14015 44360 -13895
rect 44480 -14015 44525 -13895
rect 44645 -14015 44690 -13895
rect 44810 -14015 44855 -13895
rect 44975 -14015 45030 -13895
rect 45150 -14015 45195 -13895
rect 45315 -14015 45360 -13895
rect 45480 -14015 45525 -13895
rect 45645 -14015 45700 -13895
rect 45820 -14015 45865 -13895
rect 45985 -14015 46030 -13895
rect 46150 -14015 46195 -13895
rect 46315 -14015 46370 -13895
rect 46490 -14015 46535 -13895
rect 46655 -14015 46700 -13895
rect 46820 -14015 46865 -13895
rect 46985 -14015 47040 -13895
rect 47160 -14015 47205 -13895
rect 47325 -14015 47370 -13895
rect 47490 -14015 47535 -13895
rect 47655 -14015 47865 -13895
rect 47985 -14015 48040 -13895
rect 48160 -14015 48205 -13895
rect 48325 -14015 48370 -13895
rect 48490 -14015 48535 -13895
rect 48655 -14015 48710 -13895
rect 48830 -14015 48875 -13895
rect 48995 -14015 49040 -13895
rect 49160 -14015 49205 -13895
rect 49325 -14015 49380 -13895
rect 49500 -14015 49545 -13895
rect 49665 -14015 49710 -13895
rect 49830 -14015 49875 -13895
rect 49995 -14015 50050 -13895
rect 50170 -14015 50215 -13895
rect 50335 -14015 50380 -13895
rect 50500 -14015 50545 -13895
rect 50665 -14015 50720 -13895
rect 50840 -14015 50885 -13895
rect 51005 -14015 51050 -13895
rect 51170 -14015 51215 -13895
rect 51335 -14015 51390 -13895
rect 51510 -14015 51555 -13895
rect 51675 -14015 51720 -13895
rect 51840 -14015 51885 -13895
rect 52005 -14015 52060 -13895
rect 52180 -14015 52225 -13895
rect 52345 -14015 52390 -13895
rect 52510 -14015 52555 -13895
rect 52675 -14015 52730 -13895
rect 52850 -14015 52895 -13895
rect 53015 -14015 53060 -13895
rect 53180 -14015 53225 -13895
rect 53345 -14015 53370 -13895
rect 30770 -14070 53370 -14015
rect 30770 -14104 30795 -14070
rect 30530 -14190 30795 -14104
rect 30915 -14190 30970 -14070
rect 31090 -14190 31135 -14070
rect 31255 -14190 31300 -14070
rect 31420 -14190 31465 -14070
rect 31585 -14190 31640 -14070
rect 31760 -14190 31805 -14070
rect 31925 -14190 31970 -14070
rect 32090 -14190 32135 -14070
rect 32255 -14190 32310 -14070
rect 32430 -14190 32475 -14070
rect 32595 -14190 32640 -14070
rect 32760 -14190 32805 -14070
rect 32925 -14190 32980 -14070
rect 33100 -14190 33145 -14070
rect 33265 -14190 33310 -14070
rect 33430 -14190 33475 -14070
rect 33595 -14190 33650 -14070
rect 33770 -14190 33815 -14070
rect 33935 -14190 33980 -14070
rect 34100 -14190 34145 -14070
rect 34265 -14190 34320 -14070
rect 34440 -14190 34485 -14070
rect 34605 -14190 34650 -14070
rect 34770 -14190 34815 -14070
rect 34935 -14190 34990 -14070
rect 35110 -14190 35155 -14070
rect 35275 -14190 35320 -14070
rect 35440 -14190 35485 -14070
rect 35605 -14190 35660 -14070
rect 35780 -14190 35825 -14070
rect 35945 -14190 35990 -14070
rect 36110 -14190 36155 -14070
rect 36275 -14190 36485 -14070
rect 36605 -14190 36660 -14070
rect 36780 -14190 36825 -14070
rect 36945 -14190 36990 -14070
rect 37110 -14190 37155 -14070
rect 37275 -14190 37330 -14070
rect 37450 -14190 37495 -14070
rect 37615 -14190 37660 -14070
rect 37780 -14190 37825 -14070
rect 37945 -14190 38000 -14070
rect 38120 -14190 38165 -14070
rect 38285 -14190 38330 -14070
rect 38450 -14190 38495 -14070
rect 38615 -14190 38670 -14070
rect 38790 -14190 38835 -14070
rect 38955 -14190 39000 -14070
rect 39120 -14190 39165 -14070
rect 39285 -14190 39340 -14070
rect 39460 -14190 39505 -14070
rect 39625 -14190 39670 -14070
rect 39790 -14190 39835 -14070
rect 39955 -14190 40010 -14070
rect 40130 -14190 40175 -14070
rect 40295 -14190 40340 -14070
rect 40460 -14190 40505 -14070
rect 40625 -14190 40680 -14070
rect 40800 -14190 40845 -14070
rect 40965 -14190 41010 -14070
rect 41130 -14190 41175 -14070
rect 41295 -14190 41350 -14070
rect 41470 -14190 41515 -14070
rect 41635 -14190 41680 -14070
rect 41800 -14190 41845 -14070
rect 41965 -14190 42175 -14070
rect 42295 -14190 42350 -14070
rect 42470 -14190 42515 -14070
rect 42635 -14190 42680 -14070
rect 42800 -14190 42845 -14070
rect 42965 -14190 43020 -14070
rect 43140 -14190 43185 -14070
rect 43305 -14190 43350 -14070
rect 43470 -14190 43515 -14070
rect 43635 -14190 43690 -14070
rect 43810 -14190 43855 -14070
rect 43975 -14190 44020 -14070
rect 44140 -14190 44185 -14070
rect 44305 -14190 44360 -14070
rect 44480 -14190 44525 -14070
rect 44645 -14190 44690 -14070
rect 44810 -14190 44855 -14070
rect 44975 -14190 45030 -14070
rect 45150 -14190 45195 -14070
rect 45315 -14190 45360 -14070
rect 45480 -14190 45525 -14070
rect 45645 -14190 45700 -14070
rect 45820 -14190 45865 -14070
rect 45985 -14190 46030 -14070
rect 46150 -14190 46195 -14070
rect 46315 -14190 46370 -14070
rect 46490 -14190 46535 -14070
rect 46655 -14190 46700 -14070
rect 46820 -14190 46865 -14070
rect 46985 -14190 47040 -14070
rect 47160 -14190 47205 -14070
rect 47325 -14190 47370 -14070
rect 47490 -14190 47535 -14070
rect 47655 -14190 47865 -14070
rect 47985 -14190 48040 -14070
rect 48160 -14190 48205 -14070
rect 48325 -14190 48370 -14070
rect 48490 -14190 48535 -14070
rect 48655 -14190 48710 -14070
rect 48830 -14190 48875 -14070
rect 48995 -14190 49040 -14070
rect 49160 -14190 49205 -14070
rect 49325 -14190 49380 -14070
rect 49500 -14190 49545 -14070
rect 49665 -14190 49710 -14070
rect 49830 -14190 49875 -14070
rect 49995 -14190 50050 -14070
rect 50170 -14190 50215 -14070
rect 50335 -14190 50380 -14070
rect 50500 -14190 50545 -14070
rect 50665 -14190 50720 -14070
rect 50840 -14190 50885 -14070
rect 51005 -14190 51050 -14070
rect 51170 -14190 51215 -14070
rect 51335 -14190 51390 -14070
rect 51510 -14190 51555 -14070
rect 51675 -14190 51720 -14070
rect 51840 -14190 51885 -14070
rect 52005 -14190 52060 -14070
rect 52180 -14190 52225 -14070
rect 52345 -14190 52390 -14070
rect 52510 -14190 52555 -14070
rect 52675 -14190 52730 -14070
rect 52850 -14190 52895 -14070
rect 53015 -14190 53060 -14070
rect 53180 -14190 53225 -14070
rect 53345 -14190 53370 -14070
rect 30530 -14235 53370 -14190
rect 30530 -14355 30795 -14235
rect 30915 -14355 30970 -14235
rect 31090 -14355 31135 -14235
rect 31255 -14355 31300 -14235
rect 31420 -14355 31465 -14235
rect 31585 -14355 31640 -14235
rect 31760 -14355 31805 -14235
rect 31925 -14355 31970 -14235
rect 32090 -14355 32135 -14235
rect 32255 -14355 32310 -14235
rect 32430 -14355 32475 -14235
rect 32595 -14355 32640 -14235
rect 32760 -14355 32805 -14235
rect 32925 -14355 32980 -14235
rect 33100 -14355 33145 -14235
rect 33265 -14355 33310 -14235
rect 33430 -14355 33475 -14235
rect 33595 -14355 33650 -14235
rect 33770 -14355 33815 -14235
rect 33935 -14355 33980 -14235
rect 34100 -14355 34145 -14235
rect 34265 -14355 34320 -14235
rect 34440 -14355 34485 -14235
rect 34605 -14355 34650 -14235
rect 34770 -14355 34815 -14235
rect 34935 -14355 34990 -14235
rect 35110 -14355 35155 -14235
rect 35275 -14355 35320 -14235
rect 35440 -14355 35485 -14235
rect 35605 -14355 35660 -14235
rect 35780 -14355 35825 -14235
rect 35945 -14355 35990 -14235
rect 36110 -14355 36155 -14235
rect 36275 -14355 36485 -14235
rect 36605 -14355 36660 -14235
rect 36780 -14355 36825 -14235
rect 36945 -14355 36990 -14235
rect 37110 -14355 37155 -14235
rect 37275 -14355 37330 -14235
rect 37450 -14355 37495 -14235
rect 37615 -14355 37660 -14235
rect 37780 -14355 37825 -14235
rect 37945 -14355 38000 -14235
rect 38120 -14355 38165 -14235
rect 38285 -14355 38330 -14235
rect 38450 -14355 38495 -14235
rect 38615 -14355 38670 -14235
rect 38790 -14355 38835 -14235
rect 38955 -14355 39000 -14235
rect 39120 -14355 39165 -14235
rect 39285 -14355 39340 -14235
rect 39460 -14355 39505 -14235
rect 39625 -14355 39670 -14235
rect 39790 -14355 39835 -14235
rect 39955 -14355 40010 -14235
rect 40130 -14355 40175 -14235
rect 40295 -14355 40340 -14235
rect 40460 -14355 40505 -14235
rect 40625 -14355 40680 -14235
rect 40800 -14355 40845 -14235
rect 40965 -14355 41010 -14235
rect 41130 -14355 41175 -14235
rect 41295 -14355 41350 -14235
rect 41470 -14355 41515 -14235
rect 41635 -14355 41680 -14235
rect 41800 -14355 41845 -14235
rect 41965 -14355 42175 -14235
rect 42295 -14355 42350 -14235
rect 42470 -14355 42515 -14235
rect 42635 -14355 42680 -14235
rect 42800 -14355 42845 -14235
rect 42965 -14355 43020 -14235
rect 43140 -14355 43185 -14235
rect 43305 -14355 43350 -14235
rect 43470 -14355 43515 -14235
rect 43635 -14355 43690 -14235
rect 43810 -14355 43855 -14235
rect 43975 -14355 44020 -14235
rect 44140 -14355 44185 -14235
rect 44305 -14355 44360 -14235
rect 44480 -14355 44525 -14235
rect 44645 -14355 44690 -14235
rect 44810 -14355 44855 -14235
rect 44975 -14355 45030 -14235
rect 45150 -14355 45195 -14235
rect 45315 -14355 45360 -14235
rect 45480 -14355 45525 -14235
rect 45645 -14355 45700 -14235
rect 45820 -14355 45865 -14235
rect 45985 -14355 46030 -14235
rect 46150 -14355 46195 -14235
rect 46315 -14355 46370 -14235
rect 46490 -14355 46535 -14235
rect 46655 -14355 46700 -14235
rect 46820 -14355 46865 -14235
rect 46985 -14355 47040 -14235
rect 47160 -14355 47205 -14235
rect 47325 -14355 47370 -14235
rect 47490 -14355 47535 -14235
rect 47655 -14355 47865 -14235
rect 47985 -14355 48040 -14235
rect 48160 -14355 48205 -14235
rect 48325 -14355 48370 -14235
rect 48490 -14355 48535 -14235
rect 48655 -14355 48710 -14235
rect 48830 -14355 48875 -14235
rect 48995 -14355 49040 -14235
rect 49160 -14355 49205 -14235
rect 49325 -14355 49380 -14235
rect 49500 -14355 49545 -14235
rect 49665 -14355 49710 -14235
rect 49830 -14355 49875 -14235
rect 49995 -14355 50050 -14235
rect 50170 -14355 50215 -14235
rect 50335 -14355 50380 -14235
rect 50500 -14355 50545 -14235
rect 50665 -14355 50720 -14235
rect 50840 -14355 50885 -14235
rect 51005 -14355 51050 -14235
rect 51170 -14355 51215 -14235
rect 51335 -14355 51390 -14235
rect 51510 -14355 51555 -14235
rect 51675 -14355 51720 -14235
rect 51840 -14355 51885 -14235
rect 52005 -14355 52060 -14235
rect 52180 -14355 52225 -14235
rect 52345 -14355 52390 -14235
rect 52510 -14355 52555 -14235
rect 52675 -14355 52730 -14235
rect 52850 -14355 52895 -14235
rect 53015 -14355 53060 -14235
rect 53180 -14355 53225 -14235
rect 53345 -14355 53370 -14235
rect 30530 -14400 53370 -14355
rect 30530 -14404 30795 -14400
rect 30770 -14520 30795 -14404
rect 30915 -14520 30970 -14400
rect 31090 -14520 31135 -14400
rect 31255 -14520 31300 -14400
rect 31420 -14520 31465 -14400
rect 31585 -14520 31640 -14400
rect 31760 -14520 31805 -14400
rect 31925 -14520 31970 -14400
rect 32090 -14520 32135 -14400
rect 32255 -14520 32310 -14400
rect 32430 -14520 32475 -14400
rect 32595 -14520 32640 -14400
rect 32760 -14520 32805 -14400
rect 32925 -14520 32980 -14400
rect 33100 -14520 33145 -14400
rect 33265 -14520 33310 -14400
rect 33430 -14520 33475 -14400
rect 33595 -14520 33650 -14400
rect 33770 -14520 33815 -14400
rect 33935 -14520 33980 -14400
rect 34100 -14520 34145 -14400
rect 34265 -14520 34320 -14400
rect 34440 -14520 34485 -14400
rect 34605 -14520 34650 -14400
rect 34770 -14520 34815 -14400
rect 34935 -14520 34990 -14400
rect 35110 -14520 35155 -14400
rect 35275 -14520 35320 -14400
rect 35440 -14520 35485 -14400
rect 35605 -14520 35660 -14400
rect 35780 -14520 35825 -14400
rect 35945 -14520 35990 -14400
rect 36110 -14520 36155 -14400
rect 36275 -14520 36485 -14400
rect 36605 -14520 36660 -14400
rect 36780 -14520 36825 -14400
rect 36945 -14520 36990 -14400
rect 37110 -14520 37155 -14400
rect 37275 -14520 37330 -14400
rect 37450 -14520 37495 -14400
rect 37615 -14520 37660 -14400
rect 37780 -14520 37825 -14400
rect 37945 -14520 38000 -14400
rect 38120 -14520 38165 -14400
rect 38285 -14520 38330 -14400
rect 38450 -14520 38495 -14400
rect 38615 -14520 38670 -14400
rect 38790 -14520 38835 -14400
rect 38955 -14520 39000 -14400
rect 39120 -14520 39165 -14400
rect 39285 -14520 39340 -14400
rect 39460 -14520 39505 -14400
rect 39625 -14520 39670 -14400
rect 39790 -14520 39835 -14400
rect 39955 -14520 40010 -14400
rect 40130 -14520 40175 -14400
rect 40295 -14520 40340 -14400
rect 40460 -14520 40505 -14400
rect 40625 -14520 40680 -14400
rect 40800 -14520 40845 -14400
rect 40965 -14520 41010 -14400
rect 41130 -14520 41175 -14400
rect 41295 -14520 41350 -14400
rect 41470 -14520 41515 -14400
rect 41635 -14520 41680 -14400
rect 41800 -14520 41845 -14400
rect 41965 -14520 42175 -14400
rect 42295 -14520 42350 -14400
rect 42470 -14520 42515 -14400
rect 42635 -14520 42680 -14400
rect 42800 -14520 42845 -14400
rect 42965 -14520 43020 -14400
rect 43140 -14520 43185 -14400
rect 43305 -14520 43350 -14400
rect 43470 -14520 43515 -14400
rect 43635 -14520 43690 -14400
rect 43810 -14520 43855 -14400
rect 43975 -14520 44020 -14400
rect 44140 -14520 44185 -14400
rect 44305 -14520 44360 -14400
rect 44480 -14520 44525 -14400
rect 44645 -14520 44690 -14400
rect 44810 -14520 44855 -14400
rect 44975 -14520 45030 -14400
rect 45150 -14520 45195 -14400
rect 45315 -14520 45360 -14400
rect 45480 -14520 45525 -14400
rect 45645 -14520 45700 -14400
rect 45820 -14520 45865 -14400
rect 45985 -14520 46030 -14400
rect 46150 -14520 46195 -14400
rect 46315 -14520 46370 -14400
rect 46490 -14520 46535 -14400
rect 46655 -14520 46700 -14400
rect 46820 -14520 46865 -14400
rect 46985 -14520 47040 -14400
rect 47160 -14520 47205 -14400
rect 47325 -14520 47370 -14400
rect 47490 -14520 47535 -14400
rect 47655 -14520 47865 -14400
rect 47985 -14520 48040 -14400
rect 48160 -14520 48205 -14400
rect 48325 -14520 48370 -14400
rect 48490 -14520 48535 -14400
rect 48655 -14520 48710 -14400
rect 48830 -14520 48875 -14400
rect 48995 -14520 49040 -14400
rect 49160 -14520 49205 -14400
rect 49325 -14520 49380 -14400
rect 49500 -14520 49545 -14400
rect 49665 -14520 49710 -14400
rect 49830 -14520 49875 -14400
rect 49995 -14520 50050 -14400
rect 50170 -14520 50215 -14400
rect 50335 -14520 50380 -14400
rect 50500 -14520 50545 -14400
rect 50665 -14520 50720 -14400
rect 50840 -14520 50885 -14400
rect 51005 -14520 51050 -14400
rect 51170 -14520 51215 -14400
rect 51335 -14520 51390 -14400
rect 51510 -14520 51555 -14400
rect 51675 -14520 51720 -14400
rect 51840 -14520 51885 -14400
rect 52005 -14520 52060 -14400
rect 52180 -14520 52225 -14400
rect 52345 -14520 52390 -14400
rect 52510 -14520 52555 -14400
rect 52675 -14520 52730 -14400
rect 52850 -14520 52895 -14400
rect 53015 -14520 53060 -14400
rect 53180 -14520 53225 -14400
rect 53345 -14520 53370 -14400
rect 30770 -14565 53370 -14520
rect 30770 -14685 30795 -14565
rect 30915 -14685 30970 -14565
rect 31090 -14685 31135 -14565
rect 31255 -14685 31300 -14565
rect 31420 -14685 31465 -14565
rect 31585 -14685 31640 -14565
rect 31760 -14685 31805 -14565
rect 31925 -14685 31970 -14565
rect 32090 -14685 32135 -14565
rect 32255 -14685 32310 -14565
rect 32430 -14685 32475 -14565
rect 32595 -14685 32640 -14565
rect 32760 -14685 32805 -14565
rect 32925 -14685 32980 -14565
rect 33100 -14685 33145 -14565
rect 33265 -14685 33310 -14565
rect 33430 -14685 33475 -14565
rect 33595 -14685 33650 -14565
rect 33770 -14685 33815 -14565
rect 33935 -14685 33980 -14565
rect 34100 -14685 34145 -14565
rect 34265 -14685 34320 -14565
rect 34440 -14685 34485 -14565
rect 34605 -14685 34650 -14565
rect 34770 -14685 34815 -14565
rect 34935 -14685 34990 -14565
rect 35110 -14685 35155 -14565
rect 35275 -14685 35320 -14565
rect 35440 -14685 35485 -14565
rect 35605 -14685 35660 -14565
rect 35780 -14685 35825 -14565
rect 35945 -14685 35990 -14565
rect 36110 -14685 36155 -14565
rect 36275 -14685 36485 -14565
rect 36605 -14685 36660 -14565
rect 36780 -14685 36825 -14565
rect 36945 -14685 36990 -14565
rect 37110 -14685 37155 -14565
rect 37275 -14685 37330 -14565
rect 37450 -14685 37495 -14565
rect 37615 -14685 37660 -14565
rect 37780 -14685 37825 -14565
rect 37945 -14685 38000 -14565
rect 38120 -14685 38165 -14565
rect 38285 -14685 38330 -14565
rect 38450 -14685 38495 -14565
rect 38615 -14685 38670 -14565
rect 38790 -14685 38835 -14565
rect 38955 -14685 39000 -14565
rect 39120 -14685 39165 -14565
rect 39285 -14685 39340 -14565
rect 39460 -14685 39505 -14565
rect 39625 -14685 39670 -14565
rect 39790 -14685 39835 -14565
rect 39955 -14685 40010 -14565
rect 40130 -14685 40175 -14565
rect 40295 -14685 40340 -14565
rect 40460 -14685 40505 -14565
rect 40625 -14685 40680 -14565
rect 40800 -14685 40845 -14565
rect 40965 -14685 41010 -14565
rect 41130 -14685 41175 -14565
rect 41295 -14685 41350 -14565
rect 41470 -14685 41515 -14565
rect 41635 -14685 41680 -14565
rect 41800 -14685 41845 -14565
rect 41965 -14685 42175 -14565
rect 42295 -14685 42350 -14565
rect 42470 -14685 42515 -14565
rect 42635 -14685 42680 -14565
rect 42800 -14685 42845 -14565
rect 42965 -14685 43020 -14565
rect 43140 -14685 43185 -14565
rect 43305 -14685 43350 -14565
rect 43470 -14685 43515 -14565
rect 43635 -14685 43690 -14565
rect 43810 -14685 43855 -14565
rect 43975 -14685 44020 -14565
rect 44140 -14685 44185 -14565
rect 44305 -14685 44360 -14565
rect 44480 -14685 44525 -14565
rect 44645 -14685 44690 -14565
rect 44810 -14685 44855 -14565
rect 44975 -14685 45030 -14565
rect 45150 -14685 45195 -14565
rect 45315 -14685 45360 -14565
rect 45480 -14685 45525 -14565
rect 45645 -14685 45700 -14565
rect 45820 -14685 45865 -14565
rect 45985 -14685 46030 -14565
rect 46150 -14685 46195 -14565
rect 46315 -14685 46370 -14565
rect 46490 -14685 46535 -14565
rect 46655 -14685 46700 -14565
rect 46820 -14685 46865 -14565
rect 46985 -14685 47040 -14565
rect 47160 -14685 47205 -14565
rect 47325 -14685 47370 -14565
rect 47490 -14685 47535 -14565
rect 47655 -14685 47865 -14565
rect 47985 -14685 48040 -14565
rect 48160 -14685 48205 -14565
rect 48325 -14685 48370 -14565
rect 48490 -14685 48535 -14565
rect 48655 -14685 48710 -14565
rect 48830 -14685 48875 -14565
rect 48995 -14685 49040 -14565
rect 49160 -14685 49205 -14565
rect 49325 -14685 49380 -14565
rect 49500 -14685 49545 -14565
rect 49665 -14685 49710 -14565
rect 49830 -14685 49875 -14565
rect 49995 -14685 50050 -14565
rect 50170 -14685 50215 -14565
rect 50335 -14685 50380 -14565
rect 50500 -14685 50545 -14565
rect 50665 -14685 50720 -14565
rect 50840 -14685 50885 -14565
rect 51005 -14685 51050 -14565
rect 51170 -14685 51215 -14565
rect 51335 -14685 51390 -14565
rect 51510 -14685 51555 -14565
rect 51675 -14685 51720 -14565
rect 51840 -14685 51885 -14565
rect 52005 -14685 52060 -14565
rect 52180 -14685 52225 -14565
rect 52345 -14685 52390 -14565
rect 52510 -14685 52555 -14565
rect 52675 -14685 52730 -14565
rect 52850 -14685 52895 -14565
rect 53015 -14685 53060 -14565
rect 53180 -14685 53225 -14565
rect 53345 -14685 53370 -14565
rect 30770 -14740 53370 -14685
rect 30770 -14860 30795 -14740
rect 30915 -14860 30970 -14740
rect 31090 -14860 31135 -14740
rect 31255 -14860 31300 -14740
rect 31420 -14860 31465 -14740
rect 31585 -14860 31640 -14740
rect 31760 -14860 31805 -14740
rect 31925 -14860 31970 -14740
rect 32090 -14860 32135 -14740
rect 32255 -14860 32310 -14740
rect 32430 -14860 32475 -14740
rect 32595 -14860 32640 -14740
rect 32760 -14860 32805 -14740
rect 32925 -14860 32980 -14740
rect 33100 -14860 33145 -14740
rect 33265 -14860 33310 -14740
rect 33430 -14860 33475 -14740
rect 33595 -14860 33650 -14740
rect 33770 -14860 33815 -14740
rect 33935 -14860 33980 -14740
rect 34100 -14860 34145 -14740
rect 34265 -14860 34320 -14740
rect 34440 -14860 34485 -14740
rect 34605 -14860 34650 -14740
rect 34770 -14860 34815 -14740
rect 34935 -14860 34990 -14740
rect 35110 -14860 35155 -14740
rect 35275 -14860 35320 -14740
rect 35440 -14860 35485 -14740
rect 35605 -14860 35660 -14740
rect 35780 -14860 35825 -14740
rect 35945 -14860 35990 -14740
rect 36110 -14860 36155 -14740
rect 36275 -14860 36485 -14740
rect 36605 -14860 36660 -14740
rect 36780 -14860 36825 -14740
rect 36945 -14860 36990 -14740
rect 37110 -14860 37155 -14740
rect 37275 -14860 37330 -14740
rect 37450 -14860 37495 -14740
rect 37615 -14860 37660 -14740
rect 37780 -14860 37825 -14740
rect 37945 -14860 38000 -14740
rect 38120 -14860 38165 -14740
rect 38285 -14860 38330 -14740
rect 38450 -14860 38495 -14740
rect 38615 -14860 38670 -14740
rect 38790 -14860 38835 -14740
rect 38955 -14860 39000 -14740
rect 39120 -14860 39165 -14740
rect 39285 -14860 39340 -14740
rect 39460 -14860 39505 -14740
rect 39625 -14860 39670 -14740
rect 39790 -14860 39835 -14740
rect 39955 -14860 40010 -14740
rect 40130 -14860 40175 -14740
rect 40295 -14860 40340 -14740
rect 40460 -14860 40505 -14740
rect 40625 -14860 40680 -14740
rect 40800 -14860 40845 -14740
rect 40965 -14860 41010 -14740
rect 41130 -14860 41175 -14740
rect 41295 -14860 41350 -14740
rect 41470 -14860 41515 -14740
rect 41635 -14860 41680 -14740
rect 41800 -14860 41845 -14740
rect 41965 -14860 42175 -14740
rect 42295 -14860 42350 -14740
rect 42470 -14860 42515 -14740
rect 42635 -14860 42680 -14740
rect 42800 -14860 42845 -14740
rect 42965 -14860 43020 -14740
rect 43140 -14860 43185 -14740
rect 43305 -14860 43350 -14740
rect 43470 -14860 43515 -14740
rect 43635 -14860 43690 -14740
rect 43810 -14860 43855 -14740
rect 43975 -14860 44020 -14740
rect 44140 -14860 44185 -14740
rect 44305 -14860 44360 -14740
rect 44480 -14860 44525 -14740
rect 44645 -14860 44690 -14740
rect 44810 -14860 44855 -14740
rect 44975 -14860 45030 -14740
rect 45150 -14860 45195 -14740
rect 45315 -14860 45360 -14740
rect 45480 -14860 45525 -14740
rect 45645 -14860 45700 -14740
rect 45820 -14860 45865 -14740
rect 45985 -14860 46030 -14740
rect 46150 -14860 46195 -14740
rect 46315 -14860 46370 -14740
rect 46490 -14860 46535 -14740
rect 46655 -14860 46700 -14740
rect 46820 -14860 46865 -14740
rect 46985 -14860 47040 -14740
rect 47160 -14860 47205 -14740
rect 47325 -14860 47370 -14740
rect 47490 -14860 47535 -14740
rect 47655 -14860 47865 -14740
rect 47985 -14860 48040 -14740
rect 48160 -14860 48205 -14740
rect 48325 -14860 48370 -14740
rect 48490 -14860 48535 -14740
rect 48655 -14860 48710 -14740
rect 48830 -14860 48875 -14740
rect 48995 -14860 49040 -14740
rect 49160 -14860 49205 -14740
rect 49325 -14860 49380 -14740
rect 49500 -14860 49545 -14740
rect 49665 -14860 49710 -14740
rect 49830 -14860 49875 -14740
rect 49995 -14860 50050 -14740
rect 50170 -14860 50215 -14740
rect 50335 -14860 50380 -14740
rect 50500 -14860 50545 -14740
rect 50665 -14860 50720 -14740
rect 50840 -14860 50885 -14740
rect 51005 -14860 51050 -14740
rect 51170 -14860 51215 -14740
rect 51335 -14860 51390 -14740
rect 51510 -14860 51555 -14740
rect 51675 -14860 51720 -14740
rect 51840 -14860 51885 -14740
rect 52005 -14860 52060 -14740
rect 52180 -14860 52225 -14740
rect 52345 -14860 52390 -14740
rect 52510 -14860 52555 -14740
rect 52675 -14860 52730 -14740
rect 52850 -14860 52895 -14740
rect 53015 -14860 53060 -14740
rect 53180 -14860 53225 -14740
rect 53345 -14860 53370 -14740
rect 30770 -14905 53370 -14860
rect 30770 -15025 30795 -14905
rect 30915 -15025 30970 -14905
rect 31090 -15025 31135 -14905
rect 31255 -15025 31300 -14905
rect 31420 -15025 31465 -14905
rect 31585 -15025 31640 -14905
rect 31760 -15025 31805 -14905
rect 31925 -15025 31970 -14905
rect 32090 -15025 32135 -14905
rect 32255 -15025 32310 -14905
rect 32430 -15025 32475 -14905
rect 32595 -15025 32640 -14905
rect 32760 -15025 32805 -14905
rect 32925 -15025 32980 -14905
rect 33100 -15025 33145 -14905
rect 33265 -15025 33310 -14905
rect 33430 -15025 33475 -14905
rect 33595 -15025 33650 -14905
rect 33770 -15025 33815 -14905
rect 33935 -15025 33980 -14905
rect 34100 -15025 34145 -14905
rect 34265 -15025 34320 -14905
rect 34440 -15025 34485 -14905
rect 34605 -15025 34650 -14905
rect 34770 -15025 34815 -14905
rect 34935 -15025 34990 -14905
rect 35110 -15025 35155 -14905
rect 35275 -15025 35320 -14905
rect 35440 -15025 35485 -14905
rect 35605 -15025 35660 -14905
rect 35780 -15025 35825 -14905
rect 35945 -15025 35990 -14905
rect 36110 -15025 36155 -14905
rect 36275 -15025 36485 -14905
rect 36605 -15025 36660 -14905
rect 36780 -15025 36825 -14905
rect 36945 -15025 36990 -14905
rect 37110 -15025 37155 -14905
rect 37275 -15025 37330 -14905
rect 37450 -15025 37495 -14905
rect 37615 -15025 37660 -14905
rect 37780 -15025 37825 -14905
rect 37945 -15025 38000 -14905
rect 38120 -15025 38165 -14905
rect 38285 -15025 38330 -14905
rect 38450 -15025 38495 -14905
rect 38615 -15025 38670 -14905
rect 38790 -15025 38835 -14905
rect 38955 -15025 39000 -14905
rect 39120 -15025 39165 -14905
rect 39285 -15025 39340 -14905
rect 39460 -15025 39505 -14905
rect 39625 -15025 39670 -14905
rect 39790 -15025 39835 -14905
rect 39955 -15025 40010 -14905
rect 40130 -15025 40175 -14905
rect 40295 -15025 40340 -14905
rect 40460 -15025 40505 -14905
rect 40625 -15025 40680 -14905
rect 40800 -15025 40845 -14905
rect 40965 -15025 41010 -14905
rect 41130 -15025 41175 -14905
rect 41295 -15025 41350 -14905
rect 41470 -15025 41515 -14905
rect 41635 -15025 41680 -14905
rect 41800 -15025 41845 -14905
rect 41965 -15025 42175 -14905
rect 42295 -15025 42350 -14905
rect 42470 -15025 42515 -14905
rect 42635 -15025 42680 -14905
rect 42800 -15025 42845 -14905
rect 42965 -15025 43020 -14905
rect 43140 -15025 43185 -14905
rect 43305 -15025 43350 -14905
rect 43470 -15025 43515 -14905
rect 43635 -15025 43690 -14905
rect 43810 -15025 43855 -14905
rect 43975 -15025 44020 -14905
rect 44140 -15025 44185 -14905
rect 44305 -15025 44360 -14905
rect 44480 -15025 44525 -14905
rect 44645 -15025 44690 -14905
rect 44810 -15025 44855 -14905
rect 44975 -15025 45030 -14905
rect 45150 -15025 45195 -14905
rect 45315 -15025 45360 -14905
rect 45480 -15025 45525 -14905
rect 45645 -15025 45700 -14905
rect 45820 -15025 45865 -14905
rect 45985 -15025 46030 -14905
rect 46150 -15025 46195 -14905
rect 46315 -15025 46370 -14905
rect 46490 -15025 46535 -14905
rect 46655 -15025 46700 -14905
rect 46820 -15025 46865 -14905
rect 46985 -15025 47040 -14905
rect 47160 -15025 47205 -14905
rect 47325 -15025 47370 -14905
rect 47490 -15025 47535 -14905
rect 47655 -15025 47865 -14905
rect 47985 -15025 48040 -14905
rect 48160 -15025 48205 -14905
rect 48325 -15025 48370 -14905
rect 48490 -15025 48535 -14905
rect 48655 -15025 48710 -14905
rect 48830 -15025 48875 -14905
rect 48995 -15025 49040 -14905
rect 49160 -15025 49205 -14905
rect 49325 -15025 49380 -14905
rect 49500 -15025 49545 -14905
rect 49665 -15025 49710 -14905
rect 49830 -15025 49875 -14905
rect 49995 -15025 50050 -14905
rect 50170 -15025 50215 -14905
rect 50335 -15025 50380 -14905
rect 50500 -15025 50545 -14905
rect 50665 -15025 50720 -14905
rect 50840 -15025 50885 -14905
rect 51005 -15025 51050 -14905
rect 51170 -15025 51215 -14905
rect 51335 -15025 51390 -14905
rect 51510 -15025 51555 -14905
rect 51675 -15025 51720 -14905
rect 51840 -15025 51885 -14905
rect 52005 -15025 52060 -14905
rect 52180 -15025 52225 -14905
rect 52345 -15025 52390 -14905
rect 52510 -15025 52555 -14905
rect 52675 -15025 52730 -14905
rect 52850 -15025 52895 -14905
rect 53015 -15025 53060 -14905
rect 53180 -15025 53225 -14905
rect 53345 -15025 53370 -14905
rect 30770 -15070 53370 -15025
rect 30770 -15190 30795 -15070
rect 30915 -15190 30970 -15070
rect 31090 -15190 31135 -15070
rect 31255 -15190 31300 -15070
rect 31420 -15190 31465 -15070
rect 31585 -15190 31640 -15070
rect 31760 -15190 31805 -15070
rect 31925 -15190 31970 -15070
rect 32090 -15190 32135 -15070
rect 32255 -15190 32310 -15070
rect 32430 -15190 32475 -15070
rect 32595 -15190 32640 -15070
rect 32760 -15190 32805 -15070
rect 32925 -15190 32980 -15070
rect 33100 -15190 33145 -15070
rect 33265 -15190 33310 -15070
rect 33430 -15190 33475 -15070
rect 33595 -15190 33650 -15070
rect 33770 -15190 33815 -15070
rect 33935 -15190 33980 -15070
rect 34100 -15190 34145 -15070
rect 34265 -15190 34320 -15070
rect 34440 -15190 34485 -15070
rect 34605 -15190 34650 -15070
rect 34770 -15190 34815 -15070
rect 34935 -15190 34990 -15070
rect 35110 -15190 35155 -15070
rect 35275 -15190 35320 -15070
rect 35440 -15190 35485 -15070
rect 35605 -15190 35660 -15070
rect 35780 -15190 35825 -15070
rect 35945 -15190 35990 -15070
rect 36110 -15190 36155 -15070
rect 36275 -15190 36485 -15070
rect 36605 -15190 36660 -15070
rect 36780 -15190 36825 -15070
rect 36945 -15190 36990 -15070
rect 37110 -15190 37155 -15070
rect 37275 -15190 37330 -15070
rect 37450 -15190 37495 -15070
rect 37615 -15190 37660 -15070
rect 37780 -15190 37825 -15070
rect 37945 -15190 38000 -15070
rect 38120 -15190 38165 -15070
rect 38285 -15190 38330 -15070
rect 38450 -15190 38495 -15070
rect 38615 -15190 38670 -15070
rect 38790 -15190 38835 -15070
rect 38955 -15190 39000 -15070
rect 39120 -15190 39165 -15070
rect 39285 -15190 39340 -15070
rect 39460 -15190 39505 -15070
rect 39625 -15190 39670 -15070
rect 39790 -15190 39835 -15070
rect 39955 -15190 40010 -15070
rect 40130 -15190 40175 -15070
rect 40295 -15190 40340 -15070
rect 40460 -15190 40505 -15070
rect 40625 -15190 40680 -15070
rect 40800 -15190 40845 -15070
rect 40965 -15190 41010 -15070
rect 41130 -15190 41175 -15070
rect 41295 -15190 41350 -15070
rect 41470 -15190 41515 -15070
rect 41635 -15190 41680 -15070
rect 41800 -15190 41845 -15070
rect 41965 -15190 42175 -15070
rect 42295 -15190 42350 -15070
rect 42470 -15190 42515 -15070
rect 42635 -15190 42680 -15070
rect 42800 -15190 42845 -15070
rect 42965 -15190 43020 -15070
rect 43140 -15190 43185 -15070
rect 43305 -15190 43350 -15070
rect 43470 -15190 43515 -15070
rect 43635 -15190 43690 -15070
rect 43810 -15190 43855 -15070
rect 43975 -15190 44020 -15070
rect 44140 -15190 44185 -15070
rect 44305 -15190 44360 -15070
rect 44480 -15190 44525 -15070
rect 44645 -15190 44690 -15070
rect 44810 -15190 44855 -15070
rect 44975 -15190 45030 -15070
rect 45150 -15190 45195 -15070
rect 45315 -15190 45360 -15070
rect 45480 -15190 45525 -15070
rect 45645 -15190 45700 -15070
rect 45820 -15190 45865 -15070
rect 45985 -15190 46030 -15070
rect 46150 -15190 46195 -15070
rect 46315 -15190 46370 -15070
rect 46490 -15190 46535 -15070
rect 46655 -15190 46700 -15070
rect 46820 -15190 46865 -15070
rect 46985 -15190 47040 -15070
rect 47160 -15190 47205 -15070
rect 47325 -15190 47370 -15070
rect 47490 -15190 47535 -15070
rect 47655 -15190 47865 -15070
rect 47985 -15190 48040 -15070
rect 48160 -15190 48205 -15070
rect 48325 -15190 48370 -15070
rect 48490 -15190 48535 -15070
rect 48655 -15190 48710 -15070
rect 48830 -15190 48875 -15070
rect 48995 -15190 49040 -15070
rect 49160 -15190 49205 -15070
rect 49325 -15190 49380 -15070
rect 49500 -15190 49545 -15070
rect 49665 -15190 49710 -15070
rect 49830 -15190 49875 -15070
rect 49995 -15190 50050 -15070
rect 50170 -15190 50215 -15070
rect 50335 -15190 50380 -15070
rect 50500 -15190 50545 -15070
rect 50665 -15190 50720 -15070
rect 50840 -15190 50885 -15070
rect 51005 -15190 51050 -15070
rect 51170 -15190 51215 -15070
rect 51335 -15190 51390 -15070
rect 51510 -15190 51555 -15070
rect 51675 -15190 51720 -15070
rect 51840 -15190 51885 -15070
rect 52005 -15190 52060 -15070
rect 52180 -15190 52225 -15070
rect 52345 -15190 52390 -15070
rect 52510 -15190 52555 -15070
rect 52675 -15190 52730 -15070
rect 52850 -15190 52895 -15070
rect 53015 -15190 53060 -15070
rect 53180 -15190 53225 -15070
rect 53345 -15190 53370 -15070
rect 30770 -15235 53370 -15190
rect 30770 -15355 30795 -15235
rect 30915 -15355 30970 -15235
rect 31090 -15355 31135 -15235
rect 31255 -15355 31300 -15235
rect 31420 -15355 31465 -15235
rect 31585 -15355 31640 -15235
rect 31760 -15355 31805 -15235
rect 31925 -15355 31970 -15235
rect 32090 -15355 32135 -15235
rect 32255 -15355 32310 -15235
rect 32430 -15355 32475 -15235
rect 32595 -15355 32640 -15235
rect 32760 -15355 32805 -15235
rect 32925 -15355 32980 -15235
rect 33100 -15355 33145 -15235
rect 33265 -15355 33310 -15235
rect 33430 -15355 33475 -15235
rect 33595 -15355 33650 -15235
rect 33770 -15355 33815 -15235
rect 33935 -15355 33980 -15235
rect 34100 -15355 34145 -15235
rect 34265 -15355 34320 -15235
rect 34440 -15355 34485 -15235
rect 34605 -15355 34650 -15235
rect 34770 -15355 34815 -15235
rect 34935 -15355 34990 -15235
rect 35110 -15355 35155 -15235
rect 35275 -15355 35320 -15235
rect 35440 -15355 35485 -15235
rect 35605 -15355 35660 -15235
rect 35780 -15355 35825 -15235
rect 35945 -15355 35990 -15235
rect 36110 -15355 36155 -15235
rect 36275 -15355 36485 -15235
rect 36605 -15355 36660 -15235
rect 36780 -15355 36825 -15235
rect 36945 -15355 36990 -15235
rect 37110 -15355 37155 -15235
rect 37275 -15355 37330 -15235
rect 37450 -15355 37495 -15235
rect 37615 -15355 37660 -15235
rect 37780 -15355 37825 -15235
rect 37945 -15355 38000 -15235
rect 38120 -15355 38165 -15235
rect 38285 -15355 38330 -15235
rect 38450 -15355 38495 -15235
rect 38615 -15355 38670 -15235
rect 38790 -15355 38835 -15235
rect 38955 -15355 39000 -15235
rect 39120 -15355 39165 -15235
rect 39285 -15355 39340 -15235
rect 39460 -15355 39505 -15235
rect 39625 -15355 39670 -15235
rect 39790 -15355 39835 -15235
rect 39955 -15355 40010 -15235
rect 40130 -15355 40175 -15235
rect 40295 -15355 40340 -15235
rect 40460 -15355 40505 -15235
rect 40625 -15355 40680 -15235
rect 40800 -15355 40845 -15235
rect 40965 -15355 41010 -15235
rect 41130 -15355 41175 -15235
rect 41295 -15355 41350 -15235
rect 41470 -15355 41515 -15235
rect 41635 -15355 41680 -15235
rect 41800 -15355 41845 -15235
rect 41965 -15355 42175 -15235
rect 42295 -15355 42350 -15235
rect 42470 -15355 42515 -15235
rect 42635 -15355 42680 -15235
rect 42800 -15355 42845 -15235
rect 42965 -15355 43020 -15235
rect 43140 -15355 43185 -15235
rect 43305 -15355 43350 -15235
rect 43470 -15355 43515 -15235
rect 43635 -15355 43690 -15235
rect 43810 -15355 43855 -15235
rect 43975 -15355 44020 -15235
rect 44140 -15355 44185 -15235
rect 44305 -15355 44360 -15235
rect 44480 -15355 44525 -15235
rect 44645 -15355 44690 -15235
rect 44810 -15355 44855 -15235
rect 44975 -15355 45030 -15235
rect 45150 -15355 45195 -15235
rect 45315 -15355 45360 -15235
rect 45480 -15355 45525 -15235
rect 45645 -15355 45700 -15235
rect 45820 -15355 45865 -15235
rect 45985 -15355 46030 -15235
rect 46150 -15355 46195 -15235
rect 46315 -15355 46370 -15235
rect 46490 -15355 46535 -15235
rect 46655 -15355 46700 -15235
rect 46820 -15355 46865 -15235
rect 46985 -15355 47040 -15235
rect 47160 -15355 47205 -15235
rect 47325 -15355 47370 -15235
rect 47490 -15355 47535 -15235
rect 47655 -15355 47865 -15235
rect 47985 -15355 48040 -15235
rect 48160 -15355 48205 -15235
rect 48325 -15355 48370 -15235
rect 48490 -15355 48535 -15235
rect 48655 -15355 48710 -15235
rect 48830 -15355 48875 -15235
rect 48995 -15355 49040 -15235
rect 49160 -15355 49205 -15235
rect 49325 -15355 49380 -15235
rect 49500 -15355 49545 -15235
rect 49665 -15355 49710 -15235
rect 49830 -15355 49875 -15235
rect 49995 -15355 50050 -15235
rect 50170 -15355 50215 -15235
rect 50335 -15355 50380 -15235
rect 50500 -15355 50545 -15235
rect 50665 -15355 50720 -15235
rect 50840 -15355 50885 -15235
rect 51005 -15355 51050 -15235
rect 51170 -15355 51215 -15235
rect 51335 -15355 51390 -15235
rect 51510 -15355 51555 -15235
rect 51675 -15355 51720 -15235
rect 51840 -15355 51885 -15235
rect 52005 -15355 52060 -15235
rect 52180 -15355 52225 -15235
rect 52345 -15355 52390 -15235
rect 52510 -15355 52555 -15235
rect 52675 -15355 52730 -15235
rect 52850 -15355 52895 -15235
rect 53015 -15355 53060 -15235
rect 53180 -15355 53225 -15235
rect 53345 -15355 53370 -15235
rect 30770 -15410 53370 -15355
rect 30770 -15530 30795 -15410
rect 30915 -15530 30970 -15410
rect 31090 -15530 31135 -15410
rect 31255 -15530 31300 -15410
rect 31420 -15530 31465 -15410
rect 31585 -15530 31640 -15410
rect 31760 -15530 31805 -15410
rect 31925 -15530 31970 -15410
rect 32090 -15530 32135 -15410
rect 32255 -15530 32310 -15410
rect 32430 -15530 32475 -15410
rect 32595 -15530 32640 -15410
rect 32760 -15530 32805 -15410
rect 32925 -15530 32980 -15410
rect 33100 -15530 33145 -15410
rect 33265 -15530 33310 -15410
rect 33430 -15530 33475 -15410
rect 33595 -15530 33650 -15410
rect 33770 -15530 33815 -15410
rect 33935 -15530 33980 -15410
rect 34100 -15530 34145 -15410
rect 34265 -15530 34320 -15410
rect 34440 -15530 34485 -15410
rect 34605 -15530 34650 -15410
rect 34770 -15530 34815 -15410
rect 34935 -15530 34990 -15410
rect 35110 -15530 35155 -15410
rect 35275 -15530 35320 -15410
rect 35440 -15530 35485 -15410
rect 35605 -15530 35660 -15410
rect 35780 -15530 35825 -15410
rect 35945 -15530 35990 -15410
rect 36110 -15530 36155 -15410
rect 36275 -15530 36485 -15410
rect 36605 -15530 36660 -15410
rect 36780 -15530 36825 -15410
rect 36945 -15530 36990 -15410
rect 37110 -15530 37155 -15410
rect 37275 -15530 37330 -15410
rect 37450 -15530 37495 -15410
rect 37615 -15530 37660 -15410
rect 37780 -15530 37825 -15410
rect 37945 -15530 38000 -15410
rect 38120 -15530 38165 -15410
rect 38285 -15530 38330 -15410
rect 38450 -15530 38495 -15410
rect 38615 -15530 38670 -15410
rect 38790 -15530 38835 -15410
rect 38955 -15530 39000 -15410
rect 39120 -15530 39165 -15410
rect 39285 -15530 39340 -15410
rect 39460 -15530 39505 -15410
rect 39625 -15530 39670 -15410
rect 39790 -15530 39835 -15410
rect 39955 -15530 40010 -15410
rect 40130 -15530 40175 -15410
rect 40295 -15530 40340 -15410
rect 40460 -15530 40505 -15410
rect 40625 -15530 40680 -15410
rect 40800 -15530 40845 -15410
rect 40965 -15530 41010 -15410
rect 41130 -15530 41175 -15410
rect 41295 -15530 41350 -15410
rect 41470 -15530 41515 -15410
rect 41635 -15530 41680 -15410
rect 41800 -15530 41845 -15410
rect 41965 -15530 42175 -15410
rect 42295 -15530 42350 -15410
rect 42470 -15530 42515 -15410
rect 42635 -15530 42680 -15410
rect 42800 -15530 42845 -15410
rect 42965 -15530 43020 -15410
rect 43140 -15530 43185 -15410
rect 43305 -15530 43350 -15410
rect 43470 -15530 43515 -15410
rect 43635 -15530 43690 -15410
rect 43810 -15530 43855 -15410
rect 43975 -15530 44020 -15410
rect 44140 -15530 44185 -15410
rect 44305 -15530 44360 -15410
rect 44480 -15530 44525 -15410
rect 44645 -15530 44690 -15410
rect 44810 -15530 44855 -15410
rect 44975 -15530 45030 -15410
rect 45150 -15530 45195 -15410
rect 45315 -15530 45360 -15410
rect 45480 -15530 45525 -15410
rect 45645 -15530 45700 -15410
rect 45820 -15530 45865 -15410
rect 45985 -15530 46030 -15410
rect 46150 -15530 46195 -15410
rect 46315 -15530 46370 -15410
rect 46490 -15530 46535 -15410
rect 46655 -15530 46700 -15410
rect 46820 -15530 46865 -15410
rect 46985 -15530 47040 -15410
rect 47160 -15530 47205 -15410
rect 47325 -15530 47370 -15410
rect 47490 -15530 47535 -15410
rect 47655 -15530 47865 -15410
rect 47985 -15530 48040 -15410
rect 48160 -15530 48205 -15410
rect 48325 -15530 48370 -15410
rect 48490 -15530 48535 -15410
rect 48655 -15530 48710 -15410
rect 48830 -15530 48875 -15410
rect 48995 -15530 49040 -15410
rect 49160 -15530 49205 -15410
rect 49325 -15530 49380 -15410
rect 49500 -15530 49545 -15410
rect 49665 -15530 49710 -15410
rect 49830 -15530 49875 -15410
rect 49995 -15530 50050 -15410
rect 50170 -15530 50215 -15410
rect 50335 -15530 50380 -15410
rect 50500 -15530 50545 -15410
rect 50665 -15530 50720 -15410
rect 50840 -15530 50885 -15410
rect 51005 -15530 51050 -15410
rect 51170 -15530 51215 -15410
rect 51335 -15530 51390 -15410
rect 51510 -15530 51555 -15410
rect 51675 -15530 51720 -15410
rect 51840 -15530 51885 -15410
rect 52005 -15530 52060 -15410
rect 52180 -15530 52225 -15410
rect 52345 -15530 52390 -15410
rect 52510 -15530 52555 -15410
rect 52675 -15530 52730 -15410
rect 52850 -15530 52895 -15410
rect 53015 -15530 53060 -15410
rect 53180 -15530 53225 -15410
rect 53345 -15530 53370 -15410
rect 30770 -15555 53370 -15530
<< via4 >>
rect 30835 1510 30955 1630
rect 31000 1510 31120 1630
rect 31165 1510 31285 1630
rect 31330 1510 31450 1630
rect 31495 1510 31615 1630
rect 31660 1510 31780 1630
rect 31825 1510 31945 1630
rect 31990 1510 32110 1630
rect 32155 1510 32275 1630
rect 32320 1510 32440 1630
rect 32485 1510 32605 1630
rect 32650 1510 32770 1630
rect 32815 1510 32935 1630
rect 32980 1510 33100 1630
rect 33145 1510 33265 1630
rect 33310 1510 33430 1630
rect 33475 1510 33595 1630
rect 33640 1510 33760 1630
rect 33805 1510 33925 1630
rect 33970 1510 34090 1630
rect 34135 1510 34255 1630
rect 34300 1510 34420 1630
rect 34465 1510 34585 1630
rect 34630 1510 34750 1630
rect 34795 1510 34915 1630
rect 34960 1510 35080 1630
rect 35125 1510 35245 1630
rect 35290 1510 35410 1630
rect 35455 1510 35575 1630
rect 35620 1510 35740 1630
rect 35785 1510 35905 1630
rect 35950 1510 36070 1630
rect 36115 1510 36235 1630
rect 36525 1510 36645 1630
rect 36690 1510 36810 1630
rect 36855 1510 36975 1630
rect 37020 1510 37140 1630
rect 37185 1510 37305 1630
rect 37350 1510 37470 1630
rect 37515 1510 37635 1630
rect 37680 1510 37800 1630
rect 37845 1510 37965 1630
rect 38010 1510 38130 1630
rect 38175 1510 38295 1630
rect 38340 1510 38460 1630
rect 38505 1510 38625 1630
rect 38670 1510 38790 1630
rect 38835 1510 38955 1630
rect 39000 1510 39120 1630
rect 39165 1510 39285 1630
rect 39330 1510 39450 1630
rect 39495 1510 39615 1630
rect 39660 1510 39780 1630
rect 39825 1510 39945 1630
rect 39990 1510 40110 1630
rect 40155 1510 40275 1630
rect 40320 1510 40440 1630
rect 40485 1510 40605 1630
rect 40650 1510 40770 1630
rect 40815 1510 40935 1630
rect 40980 1510 41100 1630
rect 41145 1510 41265 1630
rect 41310 1510 41430 1630
rect 41475 1510 41595 1630
rect 41640 1510 41760 1630
rect 41805 1510 41925 1630
rect 42215 1510 42335 1630
rect 42380 1510 42500 1630
rect 42545 1510 42665 1630
rect 42710 1510 42830 1630
rect 42875 1510 42995 1630
rect 43040 1510 43160 1630
rect 43205 1510 43325 1630
rect 43370 1510 43490 1630
rect 43535 1510 43655 1630
rect 43700 1510 43820 1630
rect 43865 1510 43985 1630
rect 44030 1510 44150 1630
rect 44195 1510 44315 1630
rect 44360 1510 44480 1630
rect 44525 1510 44645 1630
rect 44690 1510 44810 1630
rect 44855 1510 44975 1630
rect 45020 1510 45140 1630
rect 45185 1510 45305 1630
rect 45350 1510 45470 1630
rect 45515 1510 45635 1630
rect 45680 1510 45800 1630
rect 45845 1510 45965 1630
rect 46010 1510 46130 1630
rect 46175 1510 46295 1630
rect 46340 1510 46460 1630
rect 46505 1510 46625 1630
rect 46670 1510 46790 1630
rect 46835 1510 46955 1630
rect 47000 1510 47120 1630
rect 47165 1510 47285 1630
rect 47330 1510 47450 1630
rect 47495 1510 47615 1630
rect 47905 1510 48025 1630
rect 48070 1510 48190 1630
rect 48235 1510 48355 1630
rect 48400 1510 48520 1630
rect 48565 1510 48685 1630
rect 48730 1510 48850 1630
rect 48895 1510 49015 1630
rect 49060 1510 49180 1630
rect 49225 1510 49345 1630
rect 49390 1510 49510 1630
rect 49555 1510 49675 1630
rect 49720 1510 49840 1630
rect 49885 1510 50005 1630
rect 50050 1510 50170 1630
rect 50215 1510 50335 1630
rect 50380 1510 50500 1630
rect 50545 1510 50665 1630
rect 50710 1510 50830 1630
rect 50875 1510 50995 1630
rect 51040 1510 51160 1630
rect 51205 1510 51325 1630
rect 51370 1510 51490 1630
rect 51535 1510 51655 1630
rect 51700 1510 51820 1630
rect 51865 1510 51985 1630
rect 52030 1510 52150 1630
rect 52195 1510 52315 1630
rect 52360 1510 52480 1630
rect 52525 1510 52645 1630
rect 52690 1510 52810 1630
rect 52855 1510 52975 1630
rect 53020 1510 53140 1630
rect 53185 1510 53305 1630
rect 30835 -9960 30955 -9840
rect 31000 -9960 31120 -9840
rect 31165 -9960 31285 -9840
rect 31330 -9960 31450 -9840
rect 31495 -9960 31615 -9840
rect 31660 -9960 31780 -9840
rect 31825 -9960 31945 -9840
rect 31990 -9960 32110 -9840
rect 32155 -9960 32275 -9840
rect 32320 -9960 32440 -9840
rect 32485 -9960 32605 -9840
rect 32650 -9960 32770 -9840
rect 32815 -9960 32935 -9840
rect 32980 -9960 33100 -9840
rect 33145 -9960 33265 -9840
rect 33310 -9960 33430 -9840
rect 33475 -9960 33595 -9840
rect 33640 -9960 33760 -9840
rect 33805 -9960 33925 -9840
rect 33970 -9960 34090 -9840
rect 34135 -9960 34255 -9840
rect 34300 -9960 34420 -9840
rect 34465 -9960 34585 -9840
rect 34630 -9960 34750 -9840
rect 34795 -9960 34915 -9840
rect 34960 -9960 35080 -9840
rect 35125 -9960 35245 -9840
rect 35290 -9960 35410 -9840
rect 35455 -9960 35575 -9840
rect 35620 -9960 35740 -9840
rect 35785 -9960 35905 -9840
rect 35950 -9960 36070 -9840
rect 36115 -9960 36235 -9840
rect 36525 -9960 36645 -9840
rect 36690 -9960 36810 -9840
rect 36855 -9960 36975 -9840
rect 37020 -9960 37140 -9840
rect 37185 -9960 37305 -9840
rect 37350 -9960 37470 -9840
rect 37515 -9960 37635 -9840
rect 37680 -9960 37800 -9840
rect 37845 -9960 37965 -9840
rect 38010 -9960 38130 -9840
rect 38175 -9960 38295 -9840
rect 38340 -9960 38460 -9840
rect 38505 -9960 38625 -9840
rect 38670 -9960 38790 -9840
rect 38835 -9960 38955 -9840
rect 39000 -9960 39120 -9840
rect 39165 -9960 39285 -9840
rect 39330 -9960 39450 -9840
rect 39495 -9960 39615 -9840
rect 39660 -9960 39780 -9840
rect 39825 -9960 39945 -9840
rect 39990 -9960 40110 -9840
rect 40155 -9960 40275 -9840
rect 40320 -9960 40440 -9840
rect 40485 -9960 40605 -9840
rect 40650 -9960 40770 -9840
rect 40815 -9960 40935 -9840
rect 40980 -9960 41100 -9840
rect 41145 -9960 41265 -9840
rect 41310 -9960 41430 -9840
rect 41475 -9960 41595 -9840
rect 41640 -9960 41760 -9840
rect 41805 -9960 41925 -9840
rect 42215 -9960 42335 -9840
rect 42380 -9960 42500 -9840
rect 42545 -9960 42665 -9840
rect 42710 -9960 42830 -9840
rect 42875 -9960 42995 -9840
rect 43040 -9960 43160 -9840
rect 43205 -9960 43325 -9840
rect 43370 -9960 43490 -9840
rect 43535 -9960 43655 -9840
rect 43700 -9960 43820 -9840
rect 43865 -9960 43985 -9840
rect 44030 -9960 44150 -9840
rect 44195 -9960 44315 -9840
rect 44360 -9960 44480 -9840
rect 44525 -9960 44645 -9840
rect 44690 -9960 44810 -9840
rect 44855 -9960 44975 -9840
rect 45020 -9960 45140 -9840
rect 45185 -9960 45305 -9840
rect 45350 -9960 45470 -9840
rect 45515 -9960 45635 -9840
rect 45680 -9960 45800 -9840
rect 45845 -9960 45965 -9840
rect 46010 -9960 46130 -9840
rect 46175 -9960 46295 -9840
rect 46340 -9960 46460 -9840
rect 46505 -9960 46625 -9840
rect 46670 -9960 46790 -9840
rect 46835 -9960 46955 -9840
rect 47000 -9960 47120 -9840
rect 47165 -9960 47285 -9840
rect 47330 -9960 47450 -9840
rect 47495 -9960 47615 -9840
rect 47905 -9960 48025 -9840
rect 48070 -9960 48190 -9840
rect 48235 -9960 48355 -9840
rect 48400 -9960 48520 -9840
rect 48565 -9960 48685 -9840
rect 48730 -9960 48850 -9840
rect 48895 -9960 49015 -9840
rect 49060 -9960 49180 -9840
rect 49225 -9960 49345 -9840
rect 49390 -9960 49510 -9840
rect 49555 -9960 49675 -9840
rect 49720 -9960 49840 -9840
rect 49885 -9960 50005 -9840
rect 50050 -9960 50170 -9840
rect 50215 -9960 50335 -9840
rect 50380 -9960 50500 -9840
rect 50545 -9960 50665 -9840
rect 50710 -9960 50830 -9840
rect 50875 -9960 50995 -9840
rect 51040 -9960 51160 -9840
rect 51205 -9960 51325 -9840
rect 51370 -9960 51490 -9840
rect 51535 -9960 51655 -9840
rect 51700 -9960 51820 -9840
rect 51865 -9960 51985 -9840
rect 52030 -9960 52150 -9840
rect 52195 -9960 52315 -9840
rect 52360 -9960 52480 -9840
rect 52525 -9960 52645 -9840
rect 52690 -9960 52810 -9840
rect 52855 -9960 52975 -9840
rect 53020 -9960 53140 -9840
rect 53185 -9960 53305 -9840
<< mimcap2 >>
rect 30785 7200 36285 7210
rect 30785 7080 30795 7200
rect 30915 7080 30960 7200
rect 31080 7080 31125 7200
rect 31245 7080 31290 7200
rect 31410 7080 31465 7200
rect 31585 7080 31630 7200
rect 31750 7080 31795 7200
rect 31915 7080 31960 7200
rect 32080 7080 32135 7200
rect 32255 7080 32300 7200
rect 32420 7080 32465 7200
rect 32585 7080 32630 7200
rect 32750 7080 32805 7200
rect 32925 7080 32970 7200
rect 33090 7080 33135 7200
rect 33255 7080 33300 7200
rect 33420 7080 33475 7200
rect 33595 7080 33640 7200
rect 33760 7080 33805 7200
rect 33925 7080 33970 7200
rect 34090 7080 34145 7200
rect 34265 7080 34310 7200
rect 34430 7080 34475 7200
rect 34595 7080 34640 7200
rect 34760 7080 34815 7200
rect 34935 7080 34980 7200
rect 35100 7080 35145 7200
rect 35265 7080 35310 7200
rect 35430 7080 35485 7200
rect 35605 7080 35650 7200
rect 35770 7080 35815 7200
rect 35935 7080 35980 7200
rect 36100 7080 36155 7200
rect 36275 7080 36285 7200
rect 30785 7025 36285 7080
rect 30785 6905 30795 7025
rect 30915 6905 30960 7025
rect 31080 6905 31125 7025
rect 31245 6905 31290 7025
rect 31410 6905 31465 7025
rect 31585 6905 31630 7025
rect 31750 6905 31795 7025
rect 31915 6905 31960 7025
rect 32080 6905 32135 7025
rect 32255 6905 32300 7025
rect 32420 6905 32465 7025
rect 32585 6905 32630 7025
rect 32750 6905 32805 7025
rect 32925 6905 32970 7025
rect 33090 6905 33135 7025
rect 33255 6905 33300 7025
rect 33420 6905 33475 7025
rect 33595 6905 33640 7025
rect 33760 6905 33805 7025
rect 33925 6905 33970 7025
rect 34090 6905 34145 7025
rect 34265 6905 34310 7025
rect 34430 6905 34475 7025
rect 34595 6905 34640 7025
rect 34760 6905 34815 7025
rect 34935 6905 34980 7025
rect 35100 6905 35145 7025
rect 35265 6905 35310 7025
rect 35430 6905 35485 7025
rect 35605 6905 35650 7025
rect 35770 6905 35815 7025
rect 35935 6905 35980 7025
rect 36100 6905 36155 7025
rect 36275 6905 36285 7025
rect 30785 6860 36285 6905
rect 30785 6740 30795 6860
rect 30915 6740 30960 6860
rect 31080 6740 31125 6860
rect 31245 6740 31290 6860
rect 31410 6740 31465 6860
rect 31585 6740 31630 6860
rect 31750 6740 31795 6860
rect 31915 6740 31960 6860
rect 32080 6740 32135 6860
rect 32255 6740 32300 6860
rect 32420 6740 32465 6860
rect 32585 6740 32630 6860
rect 32750 6740 32805 6860
rect 32925 6740 32970 6860
rect 33090 6740 33135 6860
rect 33255 6740 33300 6860
rect 33420 6740 33475 6860
rect 33595 6740 33640 6860
rect 33760 6740 33805 6860
rect 33925 6740 33970 6860
rect 34090 6740 34145 6860
rect 34265 6740 34310 6860
rect 34430 6740 34475 6860
rect 34595 6740 34640 6860
rect 34760 6740 34815 6860
rect 34935 6740 34980 6860
rect 35100 6740 35145 6860
rect 35265 6740 35310 6860
rect 35430 6740 35485 6860
rect 35605 6740 35650 6860
rect 35770 6740 35815 6860
rect 35935 6740 35980 6860
rect 36100 6740 36155 6860
rect 36275 6740 36285 6860
rect 30785 6695 36285 6740
rect 30785 6575 30795 6695
rect 30915 6575 30960 6695
rect 31080 6575 31125 6695
rect 31245 6575 31290 6695
rect 31410 6575 31465 6695
rect 31585 6575 31630 6695
rect 31750 6575 31795 6695
rect 31915 6575 31960 6695
rect 32080 6575 32135 6695
rect 32255 6575 32300 6695
rect 32420 6575 32465 6695
rect 32585 6575 32630 6695
rect 32750 6575 32805 6695
rect 32925 6575 32970 6695
rect 33090 6575 33135 6695
rect 33255 6575 33300 6695
rect 33420 6575 33475 6695
rect 33595 6575 33640 6695
rect 33760 6575 33805 6695
rect 33925 6575 33970 6695
rect 34090 6575 34145 6695
rect 34265 6575 34310 6695
rect 34430 6575 34475 6695
rect 34595 6575 34640 6695
rect 34760 6575 34815 6695
rect 34935 6575 34980 6695
rect 35100 6575 35145 6695
rect 35265 6575 35310 6695
rect 35430 6575 35485 6695
rect 35605 6575 35650 6695
rect 35770 6575 35815 6695
rect 35935 6575 35980 6695
rect 36100 6575 36155 6695
rect 36275 6575 36285 6695
rect 30785 6530 36285 6575
rect 30785 6410 30795 6530
rect 30915 6410 30960 6530
rect 31080 6410 31125 6530
rect 31245 6410 31290 6530
rect 31410 6410 31465 6530
rect 31585 6410 31630 6530
rect 31750 6410 31795 6530
rect 31915 6410 31960 6530
rect 32080 6410 32135 6530
rect 32255 6410 32300 6530
rect 32420 6410 32465 6530
rect 32585 6410 32630 6530
rect 32750 6410 32805 6530
rect 32925 6410 32970 6530
rect 33090 6410 33135 6530
rect 33255 6410 33300 6530
rect 33420 6410 33475 6530
rect 33595 6410 33640 6530
rect 33760 6410 33805 6530
rect 33925 6410 33970 6530
rect 34090 6410 34145 6530
rect 34265 6410 34310 6530
rect 34430 6410 34475 6530
rect 34595 6410 34640 6530
rect 34760 6410 34815 6530
rect 34935 6410 34980 6530
rect 35100 6410 35145 6530
rect 35265 6410 35310 6530
rect 35430 6410 35485 6530
rect 35605 6410 35650 6530
rect 35770 6410 35815 6530
rect 35935 6410 35980 6530
rect 36100 6410 36155 6530
rect 36275 6410 36285 6530
rect 30785 6355 36285 6410
rect 30785 6235 30795 6355
rect 30915 6235 30960 6355
rect 31080 6235 31125 6355
rect 31245 6235 31290 6355
rect 31410 6235 31465 6355
rect 31585 6235 31630 6355
rect 31750 6235 31795 6355
rect 31915 6235 31960 6355
rect 32080 6235 32135 6355
rect 32255 6235 32300 6355
rect 32420 6235 32465 6355
rect 32585 6235 32630 6355
rect 32750 6235 32805 6355
rect 32925 6235 32970 6355
rect 33090 6235 33135 6355
rect 33255 6235 33300 6355
rect 33420 6235 33475 6355
rect 33595 6235 33640 6355
rect 33760 6235 33805 6355
rect 33925 6235 33970 6355
rect 34090 6235 34145 6355
rect 34265 6235 34310 6355
rect 34430 6235 34475 6355
rect 34595 6235 34640 6355
rect 34760 6235 34815 6355
rect 34935 6235 34980 6355
rect 35100 6235 35145 6355
rect 35265 6235 35310 6355
rect 35430 6235 35485 6355
rect 35605 6235 35650 6355
rect 35770 6235 35815 6355
rect 35935 6235 35980 6355
rect 36100 6235 36155 6355
rect 36275 6235 36285 6355
rect 30785 6190 36285 6235
rect 30785 6070 30795 6190
rect 30915 6070 30960 6190
rect 31080 6070 31125 6190
rect 31245 6070 31290 6190
rect 31410 6070 31465 6190
rect 31585 6070 31630 6190
rect 31750 6070 31795 6190
rect 31915 6070 31960 6190
rect 32080 6070 32135 6190
rect 32255 6070 32300 6190
rect 32420 6070 32465 6190
rect 32585 6070 32630 6190
rect 32750 6070 32805 6190
rect 32925 6070 32970 6190
rect 33090 6070 33135 6190
rect 33255 6070 33300 6190
rect 33420 6070 33475 6190
rect 33595 6070 33640 6190
rect 33760 6070 33805 6190
rect 33925 6070 33970 6190
rect 34090 6070 34145 6190
rect 34265 6070 34310 6190
rect 34430 6070 34475 6190
rect 34595 6070 34640 6190
rect 34760 6070 34815 6190
rect 34935 6070 34980 6190
rect 35100 6070 35145 6190
rect 35265 6070 35310 6190
rect 35430 6070 35485 6190
rect 35605 6070 35650 6190
rect 35770 6070 35815 6190
rect 35935 6070 35980 6190
rect 36100 6070 36155 6190
rect 36275 6070 36285 6190
rect 30785 6025 36285 6070
rect 30785 5905 30795 6025
rect 30915 5905 30960 6025
rect 31080 5905 31125 6025
rect 31245 5905 31290 6025
rect 31410 5905 31465 6025
rect 31585 5905 31630 6025
rect 31750 5905 31795 6025
rect 31915 5905 31960 6025
rect 32080 5905 32135 6025
rect 32255 5905 32300 6025
rect 32420 5905 32465 6025
rect 32585 5905 32630 6025
rect 32750 5905 32805 6025
rect 32925 5905 32970 6025
rect 33090 5905 33135 6025
rect 33255 5905 33300 6025
rect 33420 5905 33475 6025
rect 33595 5905 33640 6025
rect 33760 5905 33805 6025
rect 33925 5905 33970 6025
rect 34090 5905 34145 6025
rect 34265 5905 34310 6025
rect 34430 5905 34475 6025
rect 34595 5905 34640 6025
rect 34760 5905 34815 6025
rect 34935 5905 34980 6025
rect 35100 5905 35145 6025
rect 35265 5905 35310 6025
rect 35430 5905 35485 6025
rect 35605 5905 35650 6025
rect 35770 5905 35815 6025
rect 35935 5905 35980 6025
rect 36100 5905 36155 6025
rect 36275 5905 36285 6025
rect 30785 5860 36285 5905
rect 30785 5740 30795 5860
rect 30915 5740 30960 5860
rect 31080 5740 31125 5860
rect 31245 5740 31290 5860
rect 31410 5740 31465 5860
rect 31585 5740 31630 5860
rect 31750 5740 31795 5860
rect 31915 5740 31960 5860
rect 32080 5740 32135 5860
rect 32255 5740 32300 5860
rect 32420 5740 32465 5860
rect 32585 5740 32630 5860
rect 32750 5740 32805 5860
rect 32925 5740 32970 5860
rect 33090 5740 33135 5860
rect 33255 5740 33300 5860
rect 33420 5740 33475 5860
rect 33595 5740 33640 5860
rect 33760 5740 33805 5860
rect 33925 5740 33970 5860
rect 34090 5740 34145 5860
rect 34265 5740 34310 5860
rect 34430 5740 34475 5860
rect 34595 5740 34640 5860
rect 34760 5740 34815 5860
rect 34935 5740 34980 5860
rect 35100 5740 35145 5860
rect 35265 5740 35310 5860
rect 35430 5740 35485 5860
rect 35605 5740 35650 5860
rect 35770 5740 35815 5860
rect 35935 5740 35980 5860
rect 36100 5740 36155 5860
rect 36275 5740 36285 5860
rect 30785 5685 36285 5740
rect 30785 5565 30795 5685
rect 30915 5565 30960 5685
rect 31080 5565 31125 5685
rect 31245 5565 31290 5685
rect 31410 5565 31465 5685
rect 31585 5565 31630 5685
rect 31750 5565 31795 5685
rect 31915 5565 31960 5685
rect 32080 5565 32135 5685
rect 32255 5565 32300 5685
rect 32420 5565 32465 5685
rect 32585 5565 32630 5685
rect 32750 5565 32805 5685
rect 32925 5565 32970 5685
rect 33090 5565 33135 5685
rect 33255 5565 33300 5685
rect 33420 5565 33475 5685
rect 33595 5565 33640 5685
rect 33760 5565 33805 5685
rect 33925 5565 33970 5685
rect 34090 5565 34145 5685
rect 34265 5565 34310 5685
rect 34430 5565 34475 5685
rect 34595 5565 34640 5685
rect 34760 5565 34815 5685
rect 34935 5565 34980 5685
rect 35100 5565 35145 5685
rect 35265 5565 35310 5685
rect 35430 5565 35485 5685
rect 35605 5565 35650 5685
rect 35770 5565 35815 5685
rect 35935 5565 35980 5685
rect 36100 5565 36155 5685
rect 36275 5565 36285 5685
rect 30785 5520 36285 5565
rect 30785 5400 30795 5520
rect 30915 5400 30960 5520
rect 31080 5400 31125 5520
rect 31245 5400 31290 5520
rect 31410 5400 31465 5520
rect 31585 5400 31630 5520
rect 31750 5400 31795 5520
rect 31915 5400 31960 5520
rect 32080 5400 32135 5520
rect 32255 5400 32300 5520
rect 32420 5400 32465 5520
rect 32585 5400 32630 5520
rect 32750 5400 32805 5520
rect 32925 5400 32970 5520
rect 33090 5400 33135 5520
rect 33255 5400 33300 5520
rect 33420 5400 33475 5520
rect 33595 5400 33640 5520
rect 33760 5400 33805 5520
rect 33925 5400 33970 5520
rect 34090 5400 34145 5520
rect 34265 5400 34310 5520
rect 34430 5400 34475 5520
rect 34595 5400 34640 5520
rect 34760 5400 34815 5520
rect 34935 5400 34980 5520
rect 35100 5400 35145 5520
rect 35265 5400 35310 5520
rect 35430 5400 35485 5520
rect 35605 5400 35650 5520
rect 35770 5400 35815 5520
rect 35935 5400 35980 5520
rect 36100 5400 36155 5520
rect 36275 5400 36285 5520
rect 30785 5355 36285 5400
rect 30785 5235 30795 5355
rect 30915 5235 30960 5355
rect 31080 5235 31125 5355
rect 31245 5235 31290 5355
rect 31410 5235 31465 5355
rect 31585 5235 31630 5355
rect 31750 5235 31795 5355
rect 31915 5235 31960 5355
rect 32080 5235 32135 5355
rect 32255 5235 32300 5355
rect 32420 5235 32465 5355
rect 32585 5235 32630 5355
rect 32750 5235 32805 5355
rect 32925 5235 32970 5355
rect 33090 5235 33135 5355
rect 33255 5235 33300 5355
rect 33420 5235 33475 5355
rect 33595 5235 33640 5355
rect 33760 5235 33805 5355
rect 33925 5235 33970 5355
rect 34090 5235 34145 5355
rect 34265 5235 34310 5355
rect 34430 5235 34475 5355
rect 34595 5235 34640 5355
rect 34760 5235 34815 5355
rect 34935 5235 34980 5355
rect 35100 5235 35145 5355
rect 35265 5235 35310 5355
rect 35430 5235 35485 5355
rect 35605 5235 35650 5355
rect 35770 5235 35815 5355
rect 35935 5235 35980 5355
rect 36100 5235 36155 5355
rect 36275 5235 36285 5355
rect 30785 5190 36285 5235
rect 30785 5070 30795 5190
rect 30915 5070 30960 5190
rect 31080 5070 31125 5190
rect 31245 5070 31290 5190
rect 31410 5070 31465 5190
rect 31585 5070 31630 5190
rect 31750 5070 31795 5190
rect 31915 5070 31960 5190
rect 32080 5070 32135 5190
rect 32255 5070 32300 5190
rect 32420 5070 32465 5190
rect 32585 5070 32630 5190
rect 32750 5070 32805 5190
rect 32925 5070 32970 5190
rect 33090 5070 33135 5190
rect 33255 5070 33300 5190
rect 33420 5070 33475 5190
rect 33595 5070 33640 5190
rect 33760 5070 33805 5190
rect 33925 5070 33970 5190
rect 34090 5070 34145 5190
rect 34265 5070 34310 5190
rect 34430 5070 34475 5190
rect 34595 5070 34640 5190
rect 34760 5070 34815 5190
rect 34935 5070 34980 5190
rect 35100 5070 35145 5190
rect 35265 5070 35310 5190
rect 35430 5070 35485 5190
rect 35605 5070 35650 5190
rect 35770 5070 35815 5190
rect 35935 5070 35980 5190
rect 36100 5070 36155 5190
rect 36275 5070 36285 5190
rect 30785 5015 36285 5070
rect 30785 4895 30795 5015
rect 30915 4895 30960 5015
rect 31080 4895 31125 5015
rect 31245 4895 31290 5015
rect 31410 4895 31465 5015
rect 31585 4895 31630 5015
rect 31750 4895 31795 5015
rect 31915 4895 31960 5015
rect 32080 4895 32135 5015
rect 32255 4895 32300 5015
rect 32420 4895 32465 5015
rect 32585 4895 32630 5015
rect 32750 4895 32805 5015
rect 32925 4895 32970 5015
rect 33090 4895 33135 5015
rect 33255 4895 33300 5015
rect 33420 4895 33475 5015
rect 33595 4895 33640 5015
rect 33760 4895 33805 5015
rect 33925 4895 33970 5015
rect 34090 4895 34145 5015
rect 34265 4895 34310 5015
rect 34430 4895 34475 5015
rect 34595 4895 34640 5015
rect 34760 4895 34815 5015
rect 34935 4895 34980 5015
rect 35100 4895 35145 5015
rect 35265 4895 35310 5015
rect 35430 4895 35485 5015
rect 35605 4895 35650 5015
rect 35770 4895 35815 5015
rect 35935 4895 35980 5015
rect 36100 4895 36155 5015
rect 36275 4895 36285 5015
rect 30785 4850 36285 4895
rect 30785 4730 30795 4850
rect 30915 4730 30960 4850
rect 31080 4730 31125 4850
rect 31245 4730 31290 4850
rect 31410 4730 31465 4850
rect 31585 4730 31630 4850
rect 31750 4730 31795 4850
rect 31915 4730 31960 4850
rect 32080 4730 32135 4850
rect 32255 4730 32300 4850
rect 32420 4730 32465 4850
rect 32585 4730 32630 4850
rect 32750 4730 32805 4850
rect 32925 4730 32970 4850
rect 33090 4730 33135 4850
rect 33255 4730 33300 4850
rect 33420 4730 33475 4850
rect 33595 4730 33640 4850
rect 33760 4730 33805 4850
rect 33925 4730 33970 4850
rect 34090 4730 34145 4850
rect 34265 4730 34310 4850
rect 34430 4730 34475 4850
rect 34595 4730 34640 4850
rect 34760 4730 34815 4850
rect 34935 4730 34980 4850
rect 35100 4730 35145 4850
rect 35265 4730 35310 4850
rect 35430 4730 35485 4850
rect 35605 4730 35650 4850
rect 35770 4730 35815 4850
rect 35935 4730 35980 4850
rect 36100 4730 36155 4850
rect 36275 4730 36285 4850
rect 30785 4685 36285 4730
rect 30785 4565 30795 4685
rect 30915 4565 30960 4685
rect 31080 4565 31125 4685
rect 31245 4565 31290 4685
rect 31410 4565 31465 4685
rect 31585 4565 31630 4685
rect 31750 4565 31795 4685
rect 31915 4565 31960 4685
rect 32080 4565 32135 4685
rect 32255 4565 32300 4685
rect 32420 4565 32465 4685
rect 32585 4565 32630 4685
rect 32750 4565 32805 4685
rect 32925 4565 32970 4685
rect 33090 4565 33135 4685
rect 33255 4565 33300 4685
rect 33420 4565 33475 4685
rect 33595 4565 33640 4685
rect 33760 4565 33805 4685
rect 33925 4565 33970 4685
rect 34090 4565 34145 4685
rect 34265 4565 34310 4685
rect 34430 4565 34475 4685
rect 34595 4565 34640 4685
rect 34760 4565 34815 4685
rect 34935 4565 34980 4685
rect 35100 4565 35145 4685
rect 35265 4565 35310 4685
rect 35430 4565 35485 4685
rect 35605 4565 35650 4685
rect 35770 4565 35815 4685
rect 35935 4565 35980 4685
rect 36100 4565 36155 4685
rect 36275 4565 36285 4685
rect 30785 4520 36285 4565
rect 30785 4400 30795 4520
rect 30915 4400 30960 4520
rect 31080 4400 31125 4520
rect 31245 4400 31290 4520
rect 31410 4400 31465 4520
rect 31585 4400 31630 4520
rect 31750 4400 31795 4520
rect 31915 4400 31960 4520
rect 32080 4400 32135 4520
rect 32255 4400 32300 4520
rect 32420 4400 32465 4520
rect 32585 4400 32630 4520
rect 32750 4400 32805 4520
rect 32925 4400 32970 4520
rect 33090 4400 33135 4520
rect 33255 4400 33300 4520
rect 33420 4400 33475 4520
rect 33595 4400 33640 4520
rect 33760 4400 33805 4520
rect 33925 4400 33970 4520
rect 34090 4400 34145 4520
rect 34265 4400 34310 4520
rect 34430 4400 34475 4520
rect 34595 4400 34640 4520
rect 34760 4400 34815 4520
rect 34935 4400 34980 4520
rect 35100 4400 35145 4520
rect 35265 4400 35310 4520
rect 35430 4400 35485 4520
rect 35605 4400 35650 4520
rect 35770 4400 35815 4520
rect 35935 4400 35980 4520
rect 36100 4400 36155 4520
rect 36275 4400 36285 4520
rect 30785 4345 36285 4400
rect 30785 4225 30795 4345
rect 30915 4225 30960 4345
rect 31080 4225 31125 4345
rect 31245 4225 31290 4345
rect 31410 4225 31465 4345
rect 31585 4225 31630 4345
rect 31750 4225 31795 4345
rect 31915 4225 31960 4345
rect 32080 4225 32135 4345
rect 32255 4225 32300 4345
rect 32420 4225 32465 4345
rect 32585 4225 32630 4345
rect 32750 4225 32805 4345
rect 32925 4225 32970 4345
rect 33090 4225 33135 4345
rect 33255 4225 33300 4345
rect 33420 4225 33475 4345
rect 33595 4225 33640 4345
rect 33760 4225 33805 4345
rect 33925 4225 33970 4345
rect 34090 4225 34145 4345
rect 34265 4225 34310 4345
rect 34430 4225 34475 4345
rect 34595 4225 34640 4345
rect 34760 4225 34815 4345
rect 34935 4225 34980 4345
rect 35100 4225 35145 4345
rect 35265 4225 35310 4345
rect 35430 4225 35485 4345
rect 35605 4225 35650 4345
rect 35770 4225 35815 4345
rect 35935 4225 35980 4345
rect 36100 4225 36155 4345
rect 36275 4225 36285 4345
rect 30785 4180 36285 4225
rect 30785 4060 30795 4180
rect 30915 4060 30960 4180
rect 31080 4060 31125 4180
rect 31245 4060 31290 4180
rect 31410 4060 31465 4180
rect 31585 4060 31630 4180
rect 31750 4060 31795 4180
rect 31915 4060 31960 4180
rect 32080 4060 32135 4180
rect 32255 4060 32300 4180
rect 32420 4060 32465 4180
rect 32585 4060 32630 4180
rect 32750 4060 32805 4180
rect 32925 4060 32970 4180
rect 33090 4060 33135 4180
rect 33255 4060 33300 4180
rect 33420 4060 33475 4180
rect 33595 4060 33640 4180
rect 33760 4060 33805 4180
rect 33925 4060 33970 4180
rect 34090 4060 34145 4180
rect 34265 4060 34310 4180
rect 34430 4060 34475 4180
rect 34595 4060 34640 4180
rect 34760 4060 34815 4180
rect 34935 4060 34980 4180
rect 35100 4060 35145 4180
rect 35265 4060 35310 4180
rect 35430 4060 35485 4180
rect 35605 4060 35650 4180
rect 35770 4060 35815 4180
rect 35935 4060 35980 4180
rect 36100 4060 36155 4180
rect 36275 4060 36285 4180
rect 30785 4015 36285 4060
rect 30785 3895 30795 4015
rect 30915 3895 30960 4015
rect 31080 3895 31125 4015
rect 31245 3895 31290 4015
rect 31410 3895 31465 4015
rect 31585 3895 31630 4015
rect 31750 3895 31795 4015
rect 31915 3895 31960 4015
rect 32080 3895 32135 4015
rect 32255 3895 32300 4015
rect 32420 3895 32465 4015
rect 32585 3895 32630 4015
rect 32750 3895 32805 4015
rect 32925 3895 32970 4015
rect 33090 3895 33135 4015
rect 33255 3895 33300 4015
rect 33420 3895 33475 4015
rect 33595 3895 33640 4015
rect 33760 3895 33805 4015
rect 33925 3895 33970 4015
rect 34090 3895 34145 4015
rect 34265 3895 34310 4015
rect 34430 3895 34475 4015
rect 34595 3895 34640 4015
rect 34760 3895 34815 4015
rect 34935 3895 34980 4015
rect 35100 3895 35145 4015
rect 35265 3895 35310 4015
rect 35430 3895 35485 4015
rect 35605 3895 35650 4015
rect 35770 3895 35815 4015
rect 35935 3895 35980 4015
rect 36100 3895 36155 4015
rect 36275 3895 36285 4015
rect 30785 3850 36285 3895
rect 30785 3730 30795 3850
rect 30915 3730 30960 3850
rect 31080 3730 31125 3850
rect 31245 3730 31290 3850
rect 31410 3730 31465 3850
rect 31585 3730 31630 3850
rect 31750 3730 31795 3850
rect 31915 3730 31960 3850
rect 32080 3730 32135 3850
rect 32255 3730 32300 3850
rect 32420 3730 32465 3850
rect 32585 3730 32630 3850
rect 32750 3730 32805 3850
rect 32925 3730 32970 3850
rect 33090 3730 33135 3850
rect 33255 3730 33300 3850
rect 33420 3730 33475 3850
rect 33595 3730 33640 3850
rect 33760 3730 33805 3850
rect 33925 3730 33970 3850
rect 34090 3730 34145 3850
rect 34265 3730 34310 3850
rect 34430 3730 34475 3850
rect 34595 3730 34640 3850
rect 34760 3730 34815 3850
rect 34935 3730 34980 3850
rect 35100 3730 35145 3850
rect 35265 3730 35310 3850
rect 35430 3730 35485 3850
rect 35605 3730 35650 3850
rect 35770 3730 35815 3850
rect 35935 3730 35980 3850
rect 36100 3730 36155 3850
rect 36275 3730 36285 3850
rect 30785 3675 36285 3730
rect 30785 3555 30795 3675
rect 30915 3555 30960 3675
rect 31080 3555 31125 3675
rect 31245 3555 31290 3675
rect 31410 3555 31465 3675
rect 31585 3555 31630 3675
rect 31750 3555 31795 3675
rect 31915 3555 31960 3675
rect 32080 3555 32135 3675
rect 32255 3555 32300 3675
rect 32420 3555 32465 3675
rect 32585 3555 32630 3675
rect 32750 3555 32805 3675
rect 32925 3555 32970 3675
rect 33090 3555 33135 3675
rect 33255 3555 33300 3675
rect 33420 3555 33475 3675
rect 33595 3555 33640 3675
rect 33760 3555 33805 3675
rect 33925 3555 33970 3675
rect 34090 3555 34145 3675
rect 34265 3555 34310 3675
rect 34430 3555 34475 3675
rect 34595 3555 34640 3675
rect 34760 3555 34815 3675
rect 34935 3555 34980 3675
rect 35100 3555 35145 3675
rect 35265 3555 35310 3675
rect 35430 3555 35485 3675
rect 35605 3555 35650 3675
rect 35770 3555 35815 3675
rect 35935 3555 35980 3675
rect 36100 3555 36155 3675
rect 36275 3555 36285 3675
rect 30785 3510 36285 3555
rect 30785 3390 30795 3510
rect 30915 3390 30960 3510
rect 31080 3390 31125 3510
rect 31245 3390 31290 3510
rect 31410 3390 31465 3510
rect 31585 3390 31630 3510
rect 31750 3390 31795 3510
rect 31915 3390 31960 3510
rect 32080 3390 32135 3510
rect 32255 3390 32300 3510
rect 32420 3390 32465 3510
rect 32585 3390 32630 3510
rect 32750 3390 32805 3510
rect 32925 3390 32970 3510
rect 33090 3390 33135 3510
rect 33255 3390 33300 3510
rect 33420 3390 33475 3510
rect 33595 3390 33640 3510
rect 33760 3390 33805 3510
rect 33925 3390 33970 3510
rect 34090 3390 34145 3510
rect 34265 3390 34310 3510
rect 34430 3390 34475 3510
rect 34595 3390 34640 3510
rect 34760 3390 34815 3510
rect 34935 3390 34980 3510
rect 35100 3390 35145 3510
rect 35265 3390 35310 3510
rect 35430 3390 35485 3510
rect 35605 3390 35650 3510
rect 35770 3390 35815 3510
rect 35935 3390 35980 3510
rect 36100 3390 36155 3510
rect 36275 3390 36285 3510
rect 30785 3345 36285 3390
rect 30785 3225 30795 3345
rect 30915 3225 30960 3345
rect 31080 3225 31125 3345
rect 31245 3225 31290 3345
rect 31410 3225 31465 3345
rect 31585 3225 31630 3345
rect 31750 3225 31795 3345
rect 31915 3225 31960 3345
rect 32080 3225 32135 3345
rect 32255 3225 32300 3345
rect 32420 3225 32465 3345
rect 32585 3225 32630 3345
rect 32750 3225 32805 3345
rect 32925 3225 32970 3345
rect 33090 3225 33135 3345
rect 33255 3225 33300 3345
rect 33420 3225 33475 3345
rect 33595 3225 33640 3345
rect 33760 3225 33805 3345
rect 33925 3225 33970 3345
rect 34090 3225 34145 3345
rect 34265 3225 34310 3345
rect 34430 3225 34475 3345
rect 34595 3225 34640 3345
rect 34760 3225 34815 3345
rect 34935 3225 34980 3345
rect 35100 3225 35145 3345
rect 35265 3225 35310 3345
rect 35430 3225 35485 3345
rect 35605 3225 35650 3345
rect 35770 3225 35815 3345
rect 35935 3225 35980 3345
rect 36100 3225 36155 3345
rect 36275 3225 36285 3345
rect 30785 3180 36285 3225
rect 30785 3060 30795 3180
rect 30915 3060 30960 3180
rect 31080 3060 31125 3180
rect 31245 3060 31290 3180
rect 31410 3060 31465 3180
rect 31585 3060 31630 3180
rect 31750 3060 31795 3180
rect 31915 3060 31960 3180
rect 32080 3060 32135 3180
rect 32255 3060 32300 3180
rect 32420 3060 32465 3180
rect 32585 3060 32630 3180
rect 32750 3060 32805 3180
rect 32925 3060 32970 3180
rect 33090 3060 33135 3180
rect 33255 3060 33300 3180
rect 33420 3060 33475 3180
rect 33595 3060 33640 3180
rect 33760 3060 33805 3180
rect 33925 3060 33970 3180
rect 34090 3060 34145 3180
rect 34265 3060 34310 3180
rect 34430 3060 34475 3180
rect 34595 3060 34640 3180
rect 34760 3060 34815 3180
rect 34935 3060 34980 3180
rect 35100 3060 35145 3180
rect 35265 3060 35310 3180
rect 35430 3060 35485 3180
rect 35605 3060 35650 3180
rect 35770 3060 35815 3180
rect 35935 3060 35980 3180
rect 36100 3060 36155 3180
rect 36275 3060 36285 3180
rect 30785 3005 36285 3060
rect 30785 2885 30795 3005
rect 30915 2885 30960 3005
rect 31080 2885 31125 3005
rect 31245 2885 31290 3005
rect 31410 2885 31465 3005
rect 31585 2885 31630 3005
rect 31750 2885 31795 3005
rect 31915 2885 31960 3005
rect 32080 2885 32135 3005
rect 32255 2885 32300 3005
rect 32420 2885 32465 3005
rect 32585 2885 32630 3005
rect 32750 2885 32805 3005
rect 32925 2885 32970 3005
rect 33090 2885 33135 3005
rect 33255 2885 33300 3005
rect 33420 2885 33475 3005
rect 33595 2885 33640 3005
rect 33760 2885 33805 3005
rect 33925 2885 33970 3005
rect 34090 2885 34145 3005
rect 34265 2885 34310 3005
rect 34430 2885 34475 3005
rect 34595 2885 34640 3005
rect 34760 2885 34815 3005
rect 34935 2885 34980 3005
rect 35100 2885 35145 3005
rect 35265 2885 35310 3005
rect 35430 2885 35485 3005
rect 35605 2885 35650 3005
rect 35770 2885 35815 3005
rect 35935 2885 35980 3005
rect 36100 2885 36155 3005
rect 36275 2885 36285 3005
rect 30785 2840 36285 2885
rect 30785 2720 30795 2840
rect 30915 2720 30960 2840
rect 31080 2720 31125 2840
rect 31245 2720 31290 2840
rect 31410 2720 31465 2840
rect 31585 2720 31630 2840
rect 31750 2720 31795 2840
rect 31915 2720 31960 2840
rect 32080 2720 32135 2840
rect 32255 2720 32300 2840
rect 32420 2720 32465 2840
rect 32585 2720 32630 2840
rect 32750 2720 32805 2840
rect 32925 2720 32970 2840
rect 33090 2720 33135 2840
rect 33255 2720 33300 2840
rect 33420 2720 33475 2840
rect 33595 2720 33640 2840
rect 33760 2720 33805 2840
rect 33925 2720 33970 2840
rect 34090 2720 34145 2840
rect 34265 2720 34310 2840
rect 34430 2720 34475 2840
rect 34595 2720 34640 2840
rect 34760 2720 34815 2840
rect 34935 2720 34980 2840
rect 35100 2720 35145 2840
rect 35265 2720 35310 2840
rect 35430 2720 35485 2840
rect 35605 2720 35650 2840
rect 35770 2720 35815 2840
rect 35935 2720 35980 2840
rect 36100 2720 36155 2840
rect 36275 2720 36285 2840
rect 30785 2675 36285 2720
rect 30785 2555 30795 2675
rect 30915 2555 30960 2675
rect 31080 2555 31125 2675
rect 31245 2555 31290 2675
rect 31410 2555 31465 2675
rect 31585 2555 31630 2675
rect 31750 2555 31795 2675
rect 31915 2555 31960 2675
rect 32080 2555 32135 2675
rect 32255 2555 32300 2675
rect 32420 2555 32465 2675
rect 32585 2555 32630 2675
rect 32750 2555 32805 2675
rect 32925 2555 32970 2675
rect 33090 2555 33135 2675
rect 33255 2555 33300 2675
rect 33420 2555 33475 2675
rect 33595 2555 33640 2675
rect 33760 2555 33805 2675
rect 33925 2555 33970 2675
rect 34090 2555 34145 2675
rect 34265 2555 34310 2675
rect 34430 2555 34475 2675
rect 34595 2555 34640 2675
rect 34760 2555 34815 2675
rect 34935 2555 34980 2675
rect 35100 2555 35145 2675
rect 35265 2555 35310 2675
rect 35430 2555 35485 2675
rect 35605 2555 35650 2675
rect 35770 2555 35815 2675
rect 35935 2555 35980 2675
rect 36100 2555 36155 2675
rect 36275 2555 36285 2675
rect 30785 2510 36285 2555
rect 30785 2390 30795 2510
rect 30915 2390 30960 2510
rect 31080 2390 31125 2510
rect 31245 2390 31290 2510
rect 31410 2390 31465 2510
rect 31585 2390 31630 2510
rect 31750 2390 31795 2510
rect 31915 2390 31960 2510
rect 32080 2390 32135 2510
rect 32255 2390 32300 2510
rect 32420 2390 32465 2510
rect 32585 2390 32630 2510
rect 32750 2390 32805 2510
rect 32925 2390 32970 2510
rect 33090 2390 33135 2510
rect 33255 2390 33300 2510
rect 33420 2390 33475 2510
rect 33595 2390 33640 2510
rect 33760 2390 33805 2510
rect 33925 2390 33970 2510
rect 34090 2390 34145 2510
rect 34265 2390 34310 2510
rect 34430 2390 34475 2510
rect 34595 2390 34640 2510
rect 34760 2390 34815 2510
rect 34935 2390 34980 2510
rect 35100 2390 35145 2510
rect 35265 2390 35310 2510
rect 35430 2390 35485 2510
rect 35605 2390 35650 2510
rect 35770 2390 35815 2510
rect 35935 2390 35980 2510
rect 36100 2390 36155 2510
rect 36275 2390 36285 2510
rect 30785 2335 36285 2390
rect 30785 2215 30795 2335
rect 30915 2215 30960 2335
rect 31080 2215 31125 2335
rect 31245 2215 31290 2335
rect 31410 2215 31465 2335
rect 31585 2215 31630 2335
rect 31750 2215 31795 2335
rect 31915 2215 31960 2335
rect 32080 2215 32135 2335
rect 32255 2215 32300 2335
rect 32420 2215 32465 2335
rect 32585 2215 32630 2335
rect 32750 2215 32805 2335
rect 32925 2215 32970 2335
rect 33090 2215 33135 2335
rect 33255 2215 33300 2335
rect 33420 2215 33475 2335
rect 33595 2215 33640 2335
rect 33760 2215 33805 2335
rect 33925 2215 33970 2335
rect 34090 2215 34145 2335
rect 34265 2215 34310 2335
rect 34430 2215 34475 2335
rect 34595 2215 34640 2335
rect 34760 2215 34815 2335
rect 34935 2215 34980 2335
rect 35100 2215 35145 2335
rect 35265 2215 35310 2335
rect 35430 2215 35485 2335
rect 35605 2215 35650 2335
rect 35770 2215 35815 2335
rect 35935 2215 35980 2335
rect 36100 2215 36155 2335
rect 36275 2215 36285 2335
rect 30785 2170 36285 2215
rect 30785 2050 30795 2170
rect 30915 2050 30960 2170
rect 31080 2050 31125 2170
rect 31245 2050 31290 2170
rect 31410 2050 31465 2170
rect 31585 2050 31630 2170
rect 31750 2050 31795 2170
rect 31915 2050 31960 2170
rect 32080 2050 32135 2170
rect 32255 2050 32300 2170
rect 32420 2050 32465 2170
rect 32585 2050 32630 2170
rect 32750 2050 32805 2170
rect 32925 2050 32970 2170
rect 33090 2050 33135 2170
rect 33255 2050 33300 2170
rect 33420 2050 33475 2170
rect 33595 2050 33640 2170
rect 33760 2050 33805 2170
rect 33925 2050 33970 2170
rect 34090 2050 34145 2170
rect 34265 2050 34310 2170
rect 34430 2050 34475 2170
rect 34595 2050 34640 2170
rect 34760 2050 34815 2170
rect 34935 2050 34980 2170
rect 35100 2050 35145 2170
rect 35265 2050 35310 2170
rect 35430 2050 35485 2170
rect 35605 2050 35650 2170
rect 35770 2050 35815 2170
rect 35935 2050 35980 2170
rect 36100 2050 36155 2170
rect 36275 2050 36285 2170
rect 30785 2005 36285 2050
rect 30785 1885 30795 2005
rect 30915 1885 30960 2005
rect 31080 1885 31125 2005
rect 31245 1885 31290 2005
rect 31410 1885 31465 2005
rect 31585 1885 31630 2005
rect 31750 1885 31795 2005
rect 31915 1885 31960 2005
rect 32080 1885 32135 2005
rect 32255 1885 32300 2005
rect 32420 1885 32465 2005
rect 32585 1885 32630 2005
rect 32750 1885 32805 2005
rect 32925 1885 32970 2005
rect 33090 1885 33135 2005
rect 33255 1885 33300 2005
rect 33420 1885 33475 2005
rect 33595 1885 33640 2005
rect 33760 1885 33805 2005
rect 33925 1885 33970 2005
rect 34090 1885 34145 2005
rect 34265 1885 34310 2005
rect 34430 1885 34475 2005
rect 34595 1885 34640 2005
rect 34760 1885 34815 2005
rect 34935 1885 34980 2005
rect 35100 1885 35145 2005
rect 35265 1885 35310 2005
rect 35430 1885 35485 2005
rect 35605 1885 35650 2005
rect 35770 1885 35815 2005
rect 35935 1885 35980 2005
rect 36100 1885 36155 2005
rect 36275 1885 36285 2005
rect 30785 1840 36285 1885
rect 30785 1720 30795 1840
rect 30915 1720 30960 1840
rect 31080 1720 31125 1840
rect 31245 1720 31290 1840
rect 31410 1720 31465 1840
rect 31585 1720 31630 1840
rect 31750 1720 31795 1840
rect 31915 1720 31960 1840
rect 32080 1720 32135 1840
rect 32255 1720 32300 1840
rect 32420 1720 32465 1840
rect 32585 1720 32630 1840
rect 32750 1720 32805 1840
rect 32925 1720 32970 1840
rect 33090 1720 33135 1840
rect 33255 1720 33300 1840
rect 33420 1720 33475 1840
rect 33595 1720 33640 1840
rect 33760 1720 33805 1840
rect 33925 1720 33970 1840
rect 34090 1720 34145 1840
rect 34265 1720 34310 1840
rect 34430 1720 34475 1840
rect 34595 1720 34640 1840
rect 34760 1720 34815 1840
rect 34935 1720 34980 1840
rect 35100 1720 35145 1840
rect 35265 1720 35310 1840
rect 35430 1720 35485 1840
rect 35605 1720 35650 1840
rect 35770 1720 35815 1840
rect 35935 1720 35980 1840
rect 36100 1720 36155 1840
rect 36275 1720 36285 1840
rect 30785 1710 36285 1720
rect 36475 7200 41975 7210
rect 36475 7080 36485 7200
rect 36605 7080 36650 7200
rect 36770 7080 36815 7200
rect 36935 7080 36980 7200
rect 37100 7080 37155 7200
rect 37275 7080 37320 7200
rect 37440 7080 37485 7200
rect 37605 7080 37650 7200
rect 37770 7080 37825 7200
rect 37945 7080 37990 7200
rect 38110 7080 38155 7200
rect 38275 7080 38320 7200
rect 38440 7080 38495 7200
rect 38615 7080 38660 7200
rect 38780 7080 38825 7200
rect 38945 7080 38990 7200
rect 39110 7080 39165 7200
rect 39285 7080 39330 7200
rect 39450 7080 39495 7200
rect 39615 7080 39660 7200
rect 39780 7080 39835 7200
rect 39955 7080 40000 7200
rect 40120 7080 40165 7200
rect 40285 7080 40330 7200
rect 40450 7080 40505 7200
rect 40625 7080 40670 7200
rect 40790 7080 40835 7200
rect 40955 7080 41000 7200
rect 41120 7080 41175 7200
rect 41295 7080 41340 7200
rect 41460 7080 41505 7200
rect 41625 7080 41670 7200
rect 41790 7080 41845 7200
rect 41965 7080 41975 7200
rect 36475 7025 41975 7080
rect 36475 6905 36485 7025
rect 36605 6905 36650 7025
rect 36770 6905 36815 7025
rect 36935 6905 36980 7025
rect 37100 6905 37155 7025
rect 37275 6905 37320 7025
rect 37440 6905 37485 7025
rect 37605 6905 37650 7025
rect 37770 6905 37825 7025
rect 37945 6905 37990 7025
rect 38110 6905 38155 7025
rect 38275 6905 38320 7025
rect 38440 6905 38495 7025
rect 38615 6905 38660 7025
rect 38780 6905 38825 7025
rect 38945 6905 38990 7025
rect 39110 6905 39165 7025
rect 39285 6905 39330 7025
rect 39450 6905 39495 7025
rect 39615 6905 39660 7025
rect 39780 6905 39835 7025
rect 39955 6905 40000 7025
rect 40120 6905 40165 7025
rect 40285 6905 40330 7025
rect 40450 6905 40505 7025
rect 40625 6905 40670 7025
rect 40790 6905 40835 7025
rect 40955 6905 41000 7025
rect 41120 6905 41175 7025
rect 41295 6905 41340 7025
rect 41460 6905 41505 7025
rect 41625 6905 41670 7025
rect 41790 6905 41845 7025
rect 41965 6905 41975 7025
rect 36475 6860 41975 6905
rect 36475 6740 36485 6860
rect 36605 6740 36650 6860
rect 36770 6740 36815 6860
rect 36935 6740 36980 6860
rect 37100 6740 37155 6860
rect 37275 6740 37320 6860
rect 37440 6740 37485 6860
rect 37605 6740 37650 6860
rect 37770 6740 37825 6860
rect 37945 6740 37990 6860
rect 38110 6740 38155 6860
rect 38275 6740 38320 6860
rect 38440 6740 38495 6860
rect 38615 6740 38660 6860
rect 38780 6740 38825 6860
rect 38945 6740 38990 6860
rect 39110 6740 39165 6860
rect 39285 6740 39330 6860
rect 39450 6740 39495 6860
rect 39615 6740 39660 6860
rect 39780 6740 39835 6860
rect 39955 6740 40000 6860
rect 40120 6740 40165 6860
rect 40285 6740 40330 6860
rect 40450 6740 40505 6860
rect 40625 6740 40670 6860
rect 40790 6740 40835 6860
rect 40955 6740 41000 6860
rect 41120 6740 41175 6860
rect 41295 6740 41340 6860
rect 41460 6740 41505 6860
rect 41625 6740 41670 6860
rect 41790 6740 41845 6860
rect 41965 6740 41975 6860
rect 36475 6695 41975 6740
rect 36475 6575 36485 6695
rect 36605 6575 36650 6695
rect 36770 6575 36815 6695
rect 36935 6575 36980 6695
rect 37100 6575 37155 6695
rect 37275 6575 37320 6695
rect 37440 6575 37485 6695
rect 37605 6575 37650 6695
rect 37770 6575 37825 6695
rect 37945 6575 37990 6695
rect 38110 6575 38155 6695
rect 38275 6575 38320 6695
rect 38440 6575 38495 6695
rect 38615 6575 38660 6695
rect 38780 6575 38825 6695
rect 38945 6575 38990 6695
rect 39110 6575 39165 6695
rect 39285 6575 39330 6695
rect 39450 6575 39495 6695
rect 39615 6575 39660 6695
rect 39780 6575 39835 6695
rect 39955 6575 40000 6695
rect 40120 6575 40165 6695
rect 40285 6575 40330 6695
rect 40450 6575 40505 6695
rect 40625 6575 40670 6695
rect 40790 6575 40835 6695
rect 40955 6575 41000 6695
rect 41120 6575 41175 6695
rect 41295 6575 41340 6695
rect 41460 6575 41505 6695
rect 41625 6575 41670 6695
rect 41790 6575 41845 6695
rect 41965 6575 41975 6695
rect 36475 6530 41975 6575
rect 36475 6410 36485 6530
rect 36605 6410 36650 6530
rect 36770 6410 36815 6530
rect 36935 6410 36980 6530
rect 37100 6410 37155 6530
rect 37275 6410 37320 6530
rect 37440 6410 37485 6530
rect 37605 6410 37650 6530
rect 37770 6410 37825 6530
rect 37945 6410 37990 6530
rect 38110 6410 38155 6530
rect 38275 6410 38320 6530
rect 38440 6410 38495 6530
rect 38615 6410 38660 6530
rect 38780 6410 38825 6530
rect 38945 6410 38990 6530
rect 39110 6410 39165 6530
rect 39285 6410 39330 6530
rect 39450 6410 39495 6530
rect 39615 6410 39660 6530
rect 39780 6410 39835 6530
rect 39955 6410 40000 6530
rect 40120 6410 40165 6530
rect 40285 6410 40330 6530
rect 40450 6410 40505 6530
rect 40625 6410 40670 6530
rect 40790 6410 40835 6530
rect 40955 6410 41000 6530
rect 41120 6410 41175 6530
rect 41295 6410 41340 6530
rect 41460 6410 41505 6530
rect 41625 6410 41670 6530
rect 41790 6410 41845 6530
rect 41965 6410 41975 6530
rect 36475 6355 41975 6410
rect 36475 6235 36485 6355
rect 36605 6235 36650 6355
rect 36770 6235 36815 6355
rect 36935 6235 36980 6355
rect 37100 6235 37155 6355
rect 37275 6235 37320 6355
rect 37440 6235 37485 6355
rect 37605 6235 37650 6355
rect 37770 6235 37825 6355
rect 37945 6235 37990 6355
rect 38110 6235 38155 6355
rect 38275 6235 38320 6355
rect 38440 6235 38495 6355
rect 38615 6235 38660 6355
rect 38780 6235 38825 6355
rect 38945 6235 38990 6355
rect 39110 6235 39165 6355
rect 39285 6235 39330 6355
rect 39450 6235 39495 6355
rect 39615 6235 39660 6355
rect 39780 6235 39835 6355
rect 39955 6235 40000 6355
rect 40120 6235 40165 6355
rect 40285 6235 40330 6355
rect 40450 6235 40505 6355
rect 40625 6235 40670 6355
rect 40790 6235 40835 6355
rect 40955 6235 41000 6355
rect 41120 6235 41175 6355
rect 41295 6235 41340 6355
rect 41460 6235 41505 6355
rect 41625 6235 41670 6355
rect 41790 6235 41845 6355
rect 41965 6235 41975 6355
rect 36475 6190 41975 6235
rect 36475 6070 36485 6190
rect 36605 6070 36650 6190
rect 36770 6070 36815 6190
rect 36935 6070 36980 6190
rect 37100 6070 37155 6190
rect 37275 6070 37320 6190
rect 37440 6070 37485 6190
rect 37605 6070 37650 6190
rect 37770 6070 37825 6190
rect 37945 6070 37990 6190
rect 38110 6070 38155 6190
rect 38275 6070 38320 6190
rect 38440 6070 38495 6190
rect 38615 6070 38660 6190
rect 38780 6070 38825 6190
rect 38945 6070 38990 6190
rect 39110 6070 39165 6190
rect 39285 6070 39330 6190
rect 39450 6070 39495 6190
rect 39615 6070 39660 6190
rect 39780 6070 39835 6190
rect 39955 6070 40000 6190
rect 40120 6070 40165 6190
rect 40285 6070 40330 6190
rect 40450 6070 40505 6190
rect 40625 6070 40670 6190
rect 40790 6070 40835 6190
rect 40955 6070 41000 6190
rect 41120 6070 41175 6190
rect 41295 6070 41340 6190
rect 41460 6070 41505 6190
rect 41625 6070 41670 6190
rect 41790 6070 41845 6190
rect 41965 6070 41975 6190
rect 36475 6025 41975 6070
rect 36475 5905 36485 6025
rect 36605 5905 36650 6025
rect 36770 5905 36815 6025
rect 36935 5905 36980 6025
rect 37100 5905 37155 6025
rect 37275 5905 37320 6025
rect 37440 5905 37485 6025
rect 37605 5905 37650 6025
rect 37770 5905 37825 6025
rect 37945 5905 37990 6025
rect 38110 5905 38155 6025
rect 38275 5905 38320 6025
rect 38440 5905 38495 6025
rect 38615 5905 38660 6025
rect 38780 5905 38825 6025
rect 38945 5905 38990 6025
rect 39110 5905 39165 6025
rect 39285 5905 39330 6025
rect 39450 5905 39495 6025
rect 39615 5905 39660 6025
rect 39780 5905 39835 6025
rect 39955 5905 40000 6025
rect 40120 5905 40165 6025
rect 40285 5905 40330 6025
rect 40450 5905 40505 6025
rect 40625 5905 40670 6025
rect 40790 5905 40835 6025
rect 40955 5905 41000 6025
rect 41120 5905 41175 6025
rect 41295 5905 41340 6025
rect 41460 5905 41505 6025
rect 41625 5905 41670 6025
rect 41790 5905 41845 6025
rect 41965 5905 41975 6025
rect 36475 5860 41975 5905
rect 36475 5740 36485 5860
rect 36605 5740 36650 5860
rect 36770 5740 36815 5860
rect 36935 5740 36980 5860
rect 37100 5740 37155 5860
rect 37275 5740 37320 5860
rect 37440 5740 37485 5860
rect 37605 5740 37650 5860
rect 37770 5740 37825 5860
rect 37945 5740 37990 5860
rect 38110 5740 38155 5860
rect 38275 5740 38320 5860
rect 38440 5740 38495 5860
rect 38615 5740 38660 5860
rect 38780 5740 38825 5860
rect 38945 5740 38990 5860
rect 39110 5740 39165 5860
rect 39285 5740 39330 5860
rect 39450 5740 39495 5860
rect 39615 5740 39660 5860
rect 39780 5740 39835 5860
rect 39955 5740 40000 5860
rect 40120 5740 40165 5860
rect 40285 5740 40330 5860
rect 40450 5740 40505 5860
rect 40625 5740 40670 5860
rect 40790 5740 40835 5860
rect 40955 5740 41000 5860
rect 41120 5740 41175 5860
rect 41295 5740 41340 5860
rect 41460 5740 41505 5860
rect 41625 5740 41670 5860
rect 41790 5740 41845 5860
rect 41965 5740 41975 5860
rect 36475 5685 41975 5740
rect 36475 5565 36485 5685
rect 36605 5565 36650 5685
rect 36770 5565 36815 5685
rect 36935 5565 36980 5685
rect 37100 5565 37155 5685
rect 37275 5565 37320 5685
rect 37440 5565 37485 5685
rect 37605 5565 37650 5685
rect 37770 5565 37825 5685
rect 37945 5565 37990 5685
rect 38110 5565 38155 5685
rect 38275 5565 38320 5685
rect 38440 5565 38495 5685
rect 38615 5565 38660 5685
rect 38780 5565 38825 5685
rect 38945 5565 38990 5685
rect 39110 5565 39165 5685
rect 39285 5565 39330 5685
rect 39450 5565 39495 5685
rect 39615 5565 39660 5685
rect 39780 5565 39835 5685
rect 39955 5565 40000 5685
rect 40120 5565 40165 5685
rect 40285 5565 40330 5685
rect 40450 5565 40505 5685
rect 40625 5565 40670 5685
rect 40790 5565 40835 5685
rect 40955 5565 41000 5685
rect 41120 5565 41175 5685
rect 41295 5565 41340 5685
rect 41460 5565 41505 5685
rect 41625 5565 41670 5685
rect 41790 5565 41845 5685
rect 41965 5565 41975 5685
rect 36475 5520 41975 5565
rect 36475 5400 36485 5520
rect 36605 5400 36650 5520
rect 36770 5400 36815 5520
rect 36935 5400 36980 5520
rect 37100 5400 37155 5520
rect 37275 5400 37320 5520
rect 37440 5400 37485 5520
rect 37605 5400 37650 5520
rect 37770 5400 37825 5520
rect 37945 5400 37990 5520
rect 38110 5400 38155 5520
rect 38275 5400 38320 5520
rect 38440 5400 38495 5520
rect 38615 5400 38660 5520
rect 38780 5400 38825 5520
rect 38945 5400 38990 5520
rect 39110 5400 39165 5520
rect 39285 5400 39330 5520
rect 39450 5400 39495 5520
rect 39615 5400 39660 5520
rect 39780 5400 39835 5520
rect 39955 5400 40000 5520
rect 40120 5400 40165 5520
rect 40285 5400 40330 5520
rect 40450 5400 40505 5520
rect 40625 5400 40670 5520
rect 40790 5400 40835 5520
rect 40955 5400 41000 5520
rect 41120 5400 41175 5520
rect 41295 5400 41340 5520
rect 41460 5400 41505 5520
rect 41625 5400 41670 5520
rect 41790 5400 41845 5520
rect 41965 5400 41975 5520
rect 36475 5355 41975 5400
rect 36475 5235 36485 5355
rect 36605 5235 36650 5355
rect 36770 5235 36815 5355
rect 36935 5235 36980 5355
rect 37100 5235 37155 5355
rect 37275 5235 37320 5355
rect 37440 5235 37485 5355
rect 37605 5235 37650 5355
rect 37770 5235 37825 5355
rect 37945 5235 37990 5355
rect 38110 5235 38155 5355
rect 38275 5235 38320 5355
rect 38440 5235 38495 5355
rect 38615 5235 38660 5355
rect 38780 5235 38825 5355
rect 38945 5235 38990 5355
rect 39110 5235 39165 5355
rect 39285 5235 39330 5355
rect 39450 5235 39495 5355
rect 39615 5235 39660 5355
rect 39780 5235 39835 5355
rect 39955 5235 40000 5355
rect 40120 5235 40165 5355
rect 40285 5235 40330 5355
rect 40450 5235 40505 5355
rect 40625 5235 40670 5355
rect 40790 5235 40835 5355
rect 40955 5235 41000 5355
rect 41120 5235 41175 5355
rect 41295 5235 41340 5355
rect 41460 5235 41505 5355
rect 41625 5235 41670 5355
rect 41790 5235 41845 5355
rect 41965 5235 41975 5355
rect 36475 5190 41975 5235
rect 36475 5070 36485 5190
rect 36605 5070 36650 5190
rect 36770 5070 36815 5190
rect 36935 5070 36980 5190
rect 37100 5070 37155 5190
rect 37275 5070 37320 5190
rect 37440 5070 37485 5190
rect 37605 5070 37650 5190
rect 37770 5070 37825 5190
rect 37945 5070 37990 5190
rect 38110 5070 38155 5190
rect 38275 5070 38320 5190
rect 38440 5070 38495 5190
rect 38615 5070 38660 5190
rect 38780 5070 38825 5190
rect 38945 5070 38990 5190
rect 39110 5070 39165 5190
rect 39285 5070 39330 5190
rect 39450 5070 39495 5190
rect 39615 5070 39660 5190
rect 39780 5070 39835 5190
rect 39955 5070 40000 5190
rect 40120 5070 40165 5190
rect 40285 5070 40330 5190
rect 40450 5070 40505 5190
rect 40625 5070 40670 5190
rect 40790 5070 40835 5190
rect 40955 5070 41000 5190
rect 41120 5070 41175 5190
rect 41295 5070 41340 5190
rect 41460 5070 41505 5190
rect 41625 5070 41670 5190
rect 41790 5070 41845 5190
rect 41965 5070 41975 5190
rect 36475 5015 41975 5070
rect 36475 4895 36485 5015
rect 36605 4895 36650 5015
rect 36770 4895 36815 5015
rect 36935 4895 36980 5015
rect 37100 4895 37155 5015
rect 37275 4895 37320 5015
rect 37440 4895 37485 5015
rect 37605 4895 37650 5015
rect 37770 4895 37825 5015
rect 37945 4895 37990 5015
rect 38110 4895 38155 5015
rect 38275 4895 38320 5015
rect 38440 4895 38495 5015
rect 38615 4895 38660 5015
rect 38780 4895 38825 5015
rect 38945 4895 38990 5015
rect 39110 4895 39165 5015
rect 39285 4895 39330 5015
rect 39450 4895 39495 5015
rect 39615 4895 39660 5015
rect 39780 4895 39835 5015
rect 39955 4895 40000 5015
rect 40120 4895 40165 5015
rect 40285 4895 40330 5015
rect 40450 4895 40505 5015
rect 40625 4895 40670 5015
rect 40790 4895 40835 5015
rect 40955 4895 41000 5015
rect 41120 4895 41175 5015
rect 41295 4895 41340 5015
rect 41460 4895 41505 5015
rect 41625 4895 41670 5015
rect 41790 4895 41845 5015
rect 41965 4895 41975 5015
rect 36475 4850 41975 4895
rect 36475 4730 36485 4850
rect 36605 4730 36650 4850
rect 36770 4730 36815 4850
rect 36935 4730 36980 4850
rect 37100 4730 37155 4850
rect 37275 4730 37320 4850
rect 37440 4730 37485 4850
rect 37605 4730 37650 4850
rect 37770 4730 37825 4850
rect 37945 4730 37990 4850
rect 38110 4730 38155 4850
rect 38275 4730 38320 4850
rect 38440 4730 38495 4850
rect 38615 4730 38660 4850
rect 38780 4730 38825 4850
rect 38945 4730 38990 4850
rect 39110 4730 39165 4850
rect 39285 4730 39330 4850
rect 39450 4730 39495 4850
rect 39615 4730 39660 4850
rect 39780 4730 39835 4850
rect 39955 4730 40000 4850
rect 40120 4730 40165 4850
rect 40285 4730 40330 4850
rect 40450 4730 40505 4850
rect 40625 4730 40670 4850
rect 40790 4730 40835 4850
rect 40955 4730 41000 4850
rect 41120 4730 41175 4850
rect 41295 4730 41340 4850
rect 41460 4730 41505 4850
rect 41625 4730 41670 4850
rect 41790 4730 41845 4850
rect 41965 4730 41975 4850
rect 36475 4685 41975 4730
rect 36475 4565 36485 4685
rect 36605 4565 36650 4685
rect 36770 4565 36815 4685
rect 36935 4565 36980 4685
rect 37100 4565 37155 4685
rect 37275 4565 37320 4685
rect 37440 4565 37485 4685
rect 37605 4565 37650 4685
rect 37770 4565 37825 4685
rect 37945 4565 37990 4685
rect 38110 4565 38155 4685
rect 38275 4565 38320 4685
rect 38440 4565 38495 4685
rect 38615 4565 38660 4685
rect 38780 4565 38825 4685
rect 38945 4565 38990 4685
rect 39110 4565 39165 4685
rect 39285 4565 39330 4685
rect 39450 4565 39495 4685
rect 39615 4565 39660 4685
rect 39780 4565 39835 4685
rect 39955 4565 40000 4685
rect 40120 4565 40165 4685
rect 40285 4565 40330 4685
rect 40450 4565 40505 4685
rect 40625 4565 40670 4685
rect 40790 4565 40835 4685
rect 40955 4565 41000 4685
rect 41120 4565 41175 4685
rect 41295 4565 41340 4685
rect 41460 4565 41505 4685
rect 41625 4565 41670 4685
rect 41790 4565 41845 4685
rect 41965 4565 41975 4685
rect 36475 4520 41975 4565
rect 36475 4400 36485 4520
rect 36605 4400 36650 4520
rect 36770 4400 36815 4520
rect 36935 4400 36980 4520
rect 37100 4400 37155 4520
rect 37275 4400 37320 4520
rect 37440 4400 37485 4520
rect 37605 4400 37650 4520
rect 37770 4400 37825 4520
rect 37945 4400 37990 4520
rect 38110 4400 38155 4520
rect 38275 4400 38320 4520
rect 38440 4400 38495 4520
rect 38615 4400 38660 4520
rect 38780 4400 38825 4520
rect 38945 4400 38990 4520
rect 39110 4400 39165 4520
rect 39285 4400 39330 4520
rect 39450 4400 39495 4520
rect 39615 4400 39660 4520
rect 39780 4400 39835 4520
rect 39955 4400 40000 4520
rect 40120 4400 40165 4520
rect 40285 4400 40330 4520
rect 40450 4400 40505 4520
rect 40625 4400 40670 4520
rect 40790 4400 40835 4520
rect 40955 4400 41000 4520
rect 41120 4400 41175 4520
rect 41295 4400 41340 4520
rect 41460 4400 41505 4520
rect 41625 4400 41670 4520
rect 41790 4400 41845 4520
rect 41965 4400 41975 4520
rect 36475 4345 41975 4400
rect 36475 4225 36485 4345
rect 36605 4225 36650 4345
rect 36770 4225 36815 4345
rect 36935 4225 36980 4345
rect 37100 4225 37155 4345
rect 37275 4225 37320 4345
rect 37440 4225 37485 4345
rect 37605 4225 37650 4345
rect 37770 4225 37825 4345
rect 37945 4225 37990 4345
rect 38110 4225 38155 4345
rect 38275 4225 38320 4345
rect 38440 4225 38495 4345
rect 38615 4225 38660 4345
rect 38780 4225 38825 4345
rect 38945 4225 38990 4345
rect 39110 4225 39165 4345
rect 39285 4225 39330 4345
rect 39450 4225 39495 4345
rect 39615 4225 39660 4345
rect 39780 4225 39835 4345
rect 39955 4225 40000 4345
rect 40120 4225 40165 4345
rect 40285 4225 40330 4345
rect 40450 4225 40505 4345
rect 40625 4225 40670 4345
rect 40790 4225 40835 4345
rect 40955 4225 41000 4345
rect 41120 4225 41175 4345
rect 41295 4225 41340 4345
rect 41460 4225 41505 4345
rect 41625 4225 41670 4345
rect 41790 4225 41845 4345
rect 41965 4225 41975 4345
rect 36475 4180 41975 4225
rect 36475 4060 36485 4180
rect 36605 4060 36650 4180
rect 36770 4060 36815 4180
rect 36935 4060 36980 4180
rect 37100 4060 37155 4180
rect 37275 4060 37320 4180
rect 37440 4060 37485 4180
rect 37605 4060 37650 4180
rect 37770 4060 37825 4180
rect 37945 4060 37990 4180
rect 38110 4060 38155 4180
rect 38275 4060 38320 4180
rect 38440 4060 38495 4180
rect 38615 4060 38660 4180
rect 38780 4060 38825 4180
rect 38945 4060 38990 4180
rect 39110 4060 39165 4180
rect 39285 4060 39330 4180
rect 39450 4060 39495 4180
rect 39615 4060 39660 4180
rect 39780 4060 39835 4180
rect 39955 4060 40000 4180
rect 40120 4060 40165 4180
rect 40285 4060 40330 4180
rect 40450 4060 40505 4180
rect 40625 4060 40670 4180
rect 40790 4060 40835 4180
rect 40955 4060 41000 4180
rect 41120 4060 41175 4180
rect 41295 4060 41340 4180
rect 41460 4060 41505 4180
rect 41625 4060 41670 4180
rect 41790 4060 41845 4180
rect 41965 4060 41975 4180
rect 36475 4015 41975 4060
rect 36475 3895 36485 4015
rect 36605 3895 36650 4015
rect 36770 3895 36815 4015
rect 36935 3895 36980 4015
rect 37100 3895 37155 4015
rect 37275 3895 37320 4015
rect 37440 3895 37485 4015
rect 37605 3895 37650 4015
rect 37770 3895 37825 4015
rect 37945 3895 37990 4015
rect 38110 3895 38155 4015
rect 38275 3895 38320 4015
rect 38440 3895 38495 4015
rect 38615 3895 38660 4015
rect 38780 3895 38825 4015
rect 38945 3895 38990 4015
rect 39110 3895 39165 4015
rect 39285 3895 39330 4015
rect 39450 3895 39495 4015
rect 39615 3895 39660 4015
rect 39780 3895 39835 4015
rect 39955 3895 40000 4015
rect 40120 3895 40165 4015
rect 40285 3895 40330 4015
rect 40450 3895 40505 4015
rect 40625 3895 40670 4015
rect 40790 3895 40835 4015
rect 40955 3895 41000 4015
rect 41120 3895 41175 4015
rect 41295 3895 41340 4015
rect 41460 3895 41505 4015
rect 41625 3895 41670 4015
rect 41790 3895 41845 4015
rect 41965 3895 41975 4015
rect 36475 3850 41975 3895
rect 36475 3730 36485 3850
rect 36605 3730 36650 3850
rect 36770 3730 36815 3850
rect 36935 3730 36980 3850
rect 37100 3730 37155 3850
rect 37275 3730 37320 3850
rect 37440 3730 37485 3850
rect 37605 3730 37650 3850
rect 37770 3730 37825 3850
rect 37945 3730 37990 3850
rect 38110 3730 38155 3850
rect 38275 3730 38320 3850
rect 38440 3730 38495 3850
rect 38615 3730 38660 3850
rect 38780 3730 38825 3850
rect 38945 3730 38990 3850
rect 39110 3730 39165 3850
rect 39285 3730 39330 3850
rect 39450 3730 39495 3850
rect 39615 3730 39660 3850
rect 39780 3730 39835 3850
rect 39955 3730 40000 3850
rect 40120 3730 40165 3850
rect 40285 3730 40330 3850
rect 40450 3730 40505 3850
rect 40625 3730 40670 3850
rect 40790 3730 40835 3850
rect 40955 3730 41000 3850
rect 41120 3730 41175 3850
rect 41295 3730 41340 3850
rect 41460 3730 41505 3850
rect 41625 3730 41670 3850
rect 41790 3730 41845 3850
rect 41965 3730 41975 3850
rect 36475 3675 41975 3730
rect 36475 3555 36485 3675
rect 36605 3555 36650 3675
rect 36770 3555 36815 3675
rect 36935 3555 36980 3675
rect 37100 3555 37155 3675
rect 37275 3555 37320 3675
rect 37440 3555 37485 3675
rect 37605 3555 37650 3675
rect 37770 3555 37825 3675
rect 37945 3555 37990 3675
rect 38110 3555 38155 3675
rect 38275 3555 38320 3675
rect 38440 3555 38495 3675
rect 38615 3555 38660 3675
rect 38780 3555 38825 3675
rect 38945 3555 38990 3675
rect 39110 3555 39165 3675
rect 39285 3555 39330 3675
rect 39450 3555 39495 3675
rect 39615 3555 39660 3675
rect 39780 3555 39835 3675
rect 39955 3555 40000 3675
rect 40120 3555 40165 3675
rect 40285 3555 40330 3675
rect 40450 3555 40505 3675
rect 40625 3555 40670 3675
rect 40790 3555 40835 3675
rect 40955 3555 41000 3675
rect 41120 3555 41175 3675
rect 41295 3555 41340 3675
rect 41460 3555 41505 3675
rect 41625 3555 41670 3675
rect 41790 3555 41845 3675
rect 41965 3555 41975 3675
rect 36475 3510 41975 3555
rect 36475 3390 36485 3510
rect 36605 3390 36650 3510
rect 36770 3390 36815 3510
rect 36935 3390 36980 3510
rect 37100 3390 37155 3510
rect 37275 3390 37320 3510
rect 37440 3390 37485 3510
rect 37605 3390 37650 3510
rect 37770 3390 37825 3510
rect 37945 3390 37990 3510
rect 38110 3390 38155 3510
rect 38275 3390 38320 3510
rect 38440 3390 38495 3510
rect 38615 3390 38660 3510
rect 38780 3390 38825 3510
rect 38945 3390 38990 3510
rect 39110 3390 39165 3510
rect 39285 3390 39330 3510
rect 39450 3390 39495 3510
rect 39615 3390 39660 3510
rect 39780 3390 39835 3510
rect 39955 3390 40000 3510
rect 40120 3390 40165 3510
rect 40285 3390 40330 3510
rect 40450 3390 40505 3510
rect 40625 3390 40670 3510
rect 40790 3390 40835 3510
rect 40955 3390 41000 3510
rect 41120 3390 41175 3510
rect 41295 3390 41340 3510
rect 41460 3390 41505 3510
rect 41625 3390 41670 3510
rect 41790 3390 41845 3510
rect 41965 3390 41975 3510
rect 36475 3345 41975 3390
rect 36475 3225 36485 3345
rect 36605 3225 36650 3345
rect 36770 3225 36815 3345
rect 36935 3225 36980 3345
rect 37100 3225 37155 3345
rect 37275 3225 37320 3345
rect 37440 3225 37485 3345
rect 37605 3225 37650 3345
rect 37770 3225 37825 3345
rect 37945 3225 37990 3345
rect 38110 3225 38155 3345
rect 38275 3225 38320 3345
rect 38440 3225 38495 3345
rect 38615 3225 38660 3345
rect 38780 3225 38825 3345
rect 38945 3225 38990 3345
rect 39110 3225 39165 3345
rect 39285 3225 39330 3345
rect 39450 3225 39495 3345
rect 39615 3225 39660 3345
rect 39780 3225 39835 3345
rect 39955 3225 40000 3345
rect 40120 3225 40165 3345
rect 40285 3225 40330 3345
rect 40450 3225 40505 3345
rect 40625 3225 40670 3345
rect 40790 3225 40835 3345
rect 40955 3225 41000 3345
rect 41120 3225 41175 3345
rect 41295 3225 41340 3345
rect 41460 3225 41505 3345
rect 41625 3225 41670 3345
rect 41790 3225 41845 3345
rect 41965 3225 41975 3345
rect 36475 3180 41975 3225
rect 36475 3060 36485 3180
rect 36605 3060 36650 3180
rect 36770 3060 36815 3180
rect 36935 3060 36980 3180
rect 37100 3060 37155 3180
rect 37275 3060 37320 3180
rect 37440 3060 37485 3180
rect 37605 3060 37650 3180
rect 37770 3060 37825 3180
rect 37945 3060 37990 3180
rect 38110 3060 38155 3180
rect 38275 3060 38320 3180
rect 38440 3060 38495 3180
rect 38615 3060 38660 3180
rect 38780 3060 38825 3180
rect 38945 3060 38990 3180
rect 39110 3060 39165 3180
rect 39285 3060 39330 3180
rect 39450 3060 39495 3180
rect 39615 3060 39660 3180
rect 39780 3060 39835 3180
rect 39955 3060 40000 3180
rect 40120 3060 40165 3180
rect 40285 3060 40330 3180
rect 40450 3060 40505 3180
rect 40625 3060 40670 3180
rect 40790 3060 40835 3180
rect 40955 3060 41000 3180
rect 41120 3060 41175 3180
rect 41295 3060 41340 3180
rect 41460 3060 41505 3180
rect 41625 3060 41670 3180
rect 41790 3060 41845 3180
rect 41965 3060 41975 3180
rect 36475 3005 41975 3060
rect 36475 2885 36485 3005
rect 36605 2885 36650 3005
rect 36770 2885 36815 3005
rect 36935 2885 36980 3005
rect 37100 2885 37155 3005
rect 37275 2885 37320 3005
rect 37440 2885 37485 3005
rect 37605 2885 37650 3005
rect 37770 2885 37825 3005
rect 37945 2885 37990 3005
rect 38110 2885 38155 3005
rect 38275 2885 38320 3005
rect 38440 2885 38495 3005
rect 38615 2885 38660 3005
rect 38780 2885 38825 3005
rect 38945 2885 38990 3005
rect 39110 2885 39165 3005
rect 39285 2885 39330 3005
rect 39450 2885 39495 3005
rect 39615 2885 39660 3005
rect 39780 2885 39835 3005
rect 39955 2885 40000 3005
rect 40120 2885 40165 3005
rect 40285 2885 40330 3005
rect 40450 2885 40505 3005
rect 40625 2885 40670 3005
rect 40790 2885 40835 3005
rect 40955 2885 41000 3005
rect 41120 2885 41175 3005
rect 41295 2885 41340 3005
rect 41460 2885 41505 3005
rect 41625 2885 41670 3005
rect 41790 2885 41845 3005
rect 41965 2885 41975 3005
rect 36475 2840 41975 2885
rect 36475 2720 36485 2840
rect 36605 2720 36650 2840
rect 36770 2720 36815 2840
rect 36935 2720 36980 2840
rect 37100 2720 37155 2840
rect 37275 2720 37320 2840
rect 37440 2720 37485 2840
rect 37605 2720 37650 2840
rect 37770 2720 37825 2840
rect 37945 2720 37990 2840
rect 38110 2720 38155 2840
rect 38275 2720 38320 2840
rect 38440 2720 38495 2840
rect 38615 2720 38660 2840
rect 38780 2720 38825 2840
rect 38945 2720 38990 2840
rect 39110 2720 39165 2840
rect 39285 2720 39330 2840
rect 39450 2720 39495 2840
rect 39615 2720 39660 2840
rect 39780 2720 39835 2840
rect 39955 2720 40000 2840
rect 40120 2720 40165 2840
rect 40285 2720 40330 2840
rect 40450 2720 40505 2840
rect 40625 2720 40670 2840
rect 40790 2720 40835 2840
rect 40955 2720 41000 2840
rect 41120 2720 41175 2840
rect 41295 2720 41340 2840
rect 41460 2720 41505 2840
rect 41625 2720 41670 2840
rect 41790 2720 41845 2840
rect 41965 2720 41975 2840
rect 36475 2675 41975 2720
rect 36475 2555 36485 2675
rect 36605 2555 36650 2675
rect 36770 2555 36815 2675
rect 36935 2555 36980 2675
rect 37100 2555 37155 2675
rect 37275 2555 37320 2675
rect 37440 2555 37485 2675
rect 37605 2555 37650 2675
rect 37770 2555 37825 2675
rect 37945 2555 37990 2675
rect 38110 2555 38155 2675
rect 38275 2555 38320 2675
rect 38440 2555 38495 2675
rect 38615 2555 38660 2675
rect 38780 2555 38825 2675
rect 38945 2555 38990 2675
rect 39110 2555 39165 2675
rect 39285 2555 39330 2675
rect 39450 2555 39495 2675
rect 39615 2555 39660 2675
rect 39780 2555 39835 2675
rect 39955 2555 40000 2675
rect 40120 2555 40165 2675
rect 40285 2555 40330 2675
rect 40450 2555 40505 2675
rect 40625 2555 40670 2675
rect 40790 2555 40835 2675
rect 40955 2555 41000 2675
rect 41120 2555 41175 2675
rect 41295 2555 41340 2675
rect 41460 2555 41505 2675
rect 41625 2555 41670 2675
rect 41790 2555 41845 2675
rect 41965 2555 41975 2675
rect 36475 2510 41975 2555
rect 36475 2390 36485 2510
rect 36605 2390 36650 2510
rect 36770 2390 36815 2510
rect 36935 2390 36980 2510
rect 37100 2390 37155 2510
rect 37275 2390 37320 2510
rect 37440 2390 37485 2510
rect 37605 2390 37650 2510
rect 37770 2390 37825 2510
rect 37945 2390 37990 2510
rect 38110 2390 38155 2510
rect 38275 2390 38320 2510
rect 38440 2390 38495 2510
rect 38615 2390 38660 2510
rect 38780 2390 38825 2510
rect 38945 2390 38990 2510
rect 39110 2390 39165 2510
rect 39285 2390 39330 2510
rect 39450 2390 39495 2510
rect 39615 2390 39660 2510
rect 39780 2390 39835 2510
rect 39955 2390 40000 2510
rect 40120 2390 40165 2510
rect 40285 2390 40330 2510
rect 40450 2390 40505 2510
rect 40625 2390 40670 2510
rect 40790 2390 40835 2510
rect 40955 2390 41000 2510
rect 41120 2390 41175 2510
rect 41295 2390 41340 2510
rect 41460 2390 41505 2510
rect 41625 2390 41670 2510
rect 41790 2390 41845 2510
rect 41965 2390 41975 2510
rect 36475 2335 41975 2390
rect 36475 2215 36485 2335
rect 36605 2215 36650 2335
rect 36770 2215 36815 2335
rect 36935 2215 36980 2335
rect 37100 2215 37155 2335
rect 37275 2215 37320 2335
rect 37440 2215 37485 2335
rect 37605 2215 37650 2335
rect 37770 2215 37825 2335
rect 37945 2215 37990 2335
rect 38110 2215 38155 2335
rect 38275 2215 38320 2335
rect 38440 2215 38495 2335
rect 38615 2215 38660 2335
rect 38780 2215 38825 2335
rect 38945 2215 38990 2335
rect 39110 2215 39165 2335
rect 39285 2215 39330 2335
rect 39450 2215 39495 2335
rect 39615 2215 39660 2335
rect 39780 2215 39835 2335
rect 39955 2215 40000 2335
rect 40120 2215 40165 2335
rect 40285 2215 40330 2335
rect 40450 2215 40505 2335
rect 40625 2215 40670 2335
rect 40790 2215 40835 2335
rect 40955 2215 41000 2335
rect 41120 2215 41175 2335
rect 41295 2215 41340 2335
rect 41460 2215 41505 2335
rect 41625 2215 41670 2335
rect 41790 2215 41845 2335
rect 41965 2215 41975 2335
rect 36475 2170 41975 2215
rect 36475 2050 36485 2170
rect 36605 2050 36650 2170
rect 36770 2050 36815 2170
rect 36935 2050 36980 2170
rect 37100 2050 37155 2170
rect 37275 2050 37320 2170
rect 37440 2050 37485 2170
rect 37605 2050 37650 2170
rect 37770 2050 37825 2170
rect 37945 2050 37990 2170
rect 38110 2050 38155 2170
rect 38275 2050 38320 2170
rect 38440 2050 38495 2170
rect 38615 2050 38660 2170
rect 38780 2050 38825 2170
rect 38945 2050 38990 2170
rect 39110 2050 39165 2170
rect 39285 2050 39330 2170
rect 39450 2050 39495 2170
rect 39615 2050 39660 2170
rect 39780 2050 39835 2170
rect 39955 2050 40000 2170
rect 40120 2050 40165 2170
rect 40285 2050 40330 2170
rect 40450 2050 40505 2170
rect 40625 2050 40670 2170
rect 40790 2050 40835 2170
rect 40955 2050 41000 2170
rect 41120 2050 41175 2170
rect 41295 2050 41340 2170
rect 41460 2050 41505 2170
rect 41625 2050 41670 2170
rect 41790 2050 41845 2170
rect 41965 2050 41975 2170
rect 36475 2005 41975 2050
rect 36475 1885 36485 2005
rect 36605 1885 36650 2005
rect 36770 1885 36815 2005
rect 36935 1885 36980 2005
rect 37100 1885 37155 2005
rect 37275 1885 37320 2005
rect 37440 1885 37485 2005
rect 37605 1885 37650 2005
rect 37770 1885 37825 2005
rect 37945 1885 37990 2005
rect 38110 1885 38155 2005
rect 38275 1885 38320 2005
rect 38440 1885 38495 2005
rect 38615 1885 38660 2005
rect 38780 1885 38825 2005
rect 38945 1885 38990 2005
rect 39110 1885 39165 2005
rect 39285 1885 39330 2005
rect 39450 1885 39495 2005
rect 39615 1885 39660 2005
rect 39780 1885 39835 2005
rect 39955 1885 40000 2005
rect 40120 1885 40165 2005
rect 40285 1885 40330 2005
rect 40450 1885 40505 2005
rect 40625 1885 40670 2005
rect 40790 1885 40835 2005
rect 40955 1885 41000 2005
rect 41120 1885 41175 2005
rect 41295 1885 41340 2005
rect 41460 1885 41505 2005
rect 41625 1885 41670 2005
rect 41790 1885 41845 2005
rect 41965 1885 41975 2005
rect 36475 1840 41975 1885
rect 36475 1720 36485 1840
rect 36605 1720 36650 1840
rect 36770 1720 36815 1840
rect 36935 1720 36980 1840
rect 37100 1720 37155 1840
rect 37275 1720 37320 1840
rect 37440 1720 37485 1840
rect 37605 1720 37650 1840
rect 37770 1720 37825 1840
rect 37945 1720 37990 1840
rect 38110 1720 38155 1840
rect 38275 1720 38320 1840
rect 38440 1720 38495 1840
rect 38615 1720 38660 1840
rect 38780 1720 38825 1840
rect 38945 1720 38990 1840
rect 39110 1720 39165 1840
rect 39285 1720 39330 1840
rect 39450 1720 39495 1840
rect 39615 1720 39660 1840
rect 39780 1720 39835 1840
rect 39955 1720 40000 1840
rect 40120 1720 40165 1840
rect 40285 1720 40330 1840
rect 40450 1720 40505 1840
rect 40625 1720 40670 1840
rect 40790 1720 40835 1840
rect 40955 1720 41000 1840
rect 41120 1720 41175 1840
rect 41295 1720 41340 1840
rect 41460 1720 41505 1840
rect 41625 1720 41670 1840
rect 41790 1720 41845 1840
rect 41965 1720 41975 1840
rect 36475 1710 41975 1720
rect 42165 7200 47665 7210
rect 42165 7080 42175 7200
rect 42295 7080 42340 7200
rect 42460 7080 42505 7200
rect 42625 7080 42670 7200
rect 42790 7080 42845 7200
rect 42965 7080 43010 7200
rect 43130 7080 43175 7200
rect 43295 7080 43340 7200
rect 43460 7080 43515 7200
rect 43635 7080 43680 7200
rect 43800 7080 43845 7200
rect 43965 7080 44010 7200
rect 44130 7080 44185 7200
rect 44305 7080 44350 7200
rect 44470 7080 44515 7200
rect 44635 7080 44680 7200
rect 44800 7080 44855 7200
rect 44975 7080 45020 7200
rect 45140 7080 45185 7200
rect 45305 7080 45350 7200
rect 45470 7080 45525 7200
rect 45645 7080 45690 7200
rect 45810 7080 45855 7200
rect 45975 7080 46020 7200
rect 46140 7080 46195 7200
rect 46315 7080 46360 7200
rect 46480 7080 46525 7200
rect 46645 7080 46690 7200
rect 46810 7080 46865 7200
rect 46985 7080 47030 7200
rect 47150 7080 47195 7200
rect 47315 7080 47360 7200
rect 47480 7080 47535 7200
rect 47655 7080 47665 7200
rect 42165 7025 47665 7080
rect 42165 6905 42175 7025
rect 42295 6905 42340 7025
rect 42460 6905 42505 7025
rect 42625 6905 42670 7025
rect 42790 6905 42845 7025
rect 42965 6905 43010 7025
rect 43130 6905 43175 7025
rect 43295 6905 43340 7025
rect 43460 6905 43515 7025
rect 43635 6905 43680 7025
rect 43800 6905 43845 7025
rect 43965 6905 44010 7025
rect 44130 6905 44185 7025
rect 44305 6905 44350 7025
rect 44470 6905 44515 7025
rect 44635 6905 44680 7025
rect 44800 6905 44855 7025
rect 44975 6905 45020 7025
rect 45140 6905 45185 7025
rect 45305 6905 45350 7025
rect 45470 6905 45525 7025
rect 45645 6905 45690 7025
rect 45810 6905 45855 7025
rect 45975 6905 46020 7025
rect 46140 6905 46195 7025
rect 46315 6905 46360 7025
rect 46480 6905 46525 7025
rect 46645 6905 46690 7025
rect 46810 6905 46865 7025
rect 46985 6905 47030 7025
rect 47150 6905 47195 7025
rect 47315 6905 47360 7025
rect 47480 6905 47535 7025
rect 47655 6905 47665 7025
rect 42165 6860 47665 6905
rect 42165 6740 42175 6860
rect 42295 6740 42340 6860
rect 42460 6740 42505 6860
rect 42625 6740 42670 6860
rect 42790 6740 42845 6860
rect 42965 6740 43010 6860
rect 43130 6740 43175 6860
rect 43295 6740 43340 6860
rect 43460 6740 43515 6860
rect 43635 6740 43680 6860
rect 43800 6740 43845 6860
rect 43965 6740 44010 6860
rect 44130 6740 44185 6860
rect 44305 6740 44350 6860
rect 44470 6740 44515 6860
rect 44635 6740 44680 6860
rect 44800 6740 44855 6860
rect 44975 6740 45020 6860
rect 45140 6740 45185 6860
rect 45305 6740 45350 6860
rect 45470 6740 45525 6860
rect 45645 6740 45690 6860
rect 45810 6740 45855 6860
rect 45975 6740 46020 6860
rect 46140 6740 46195 6860
rect 46315 6740 46360 6860
rect 46480 6740 46525 6860
rect 46645 6740 46690 6860
rect 46810 6740 46865 6860
rect 46985 6740 47030 6860
rect 47150 6740 47195 6860
rect 47315 6740 47360 6860
rect 47480 6740 47535 6860
rect 47655 6740 47665 6860
rect 42165 6695 47665 6740
rect 42165 6575 42175 6695
rect 42295 6575 42340 6695
rect 42460 6575 42505 6695
rect 42625 6575 42670 6695
rect 42790 6575 42845 6695
rect 42965 6575 43010 6695
rect 43130 6575 43175 6695
rect 43295 6575 43340 6695
rect 43460 6575 43515 6695
rect 43635 6575 43680 6695
rect 43800 6575 43845 6695
rect 43965 6575 44010 6695
rect 44130 6575 44185 6695
rect 44305 6575 44350 6695
rect 44470 6575 44515 6695
rect 44635 6575 44680 6695
rect 44800 6575 44855 6695
rect 44975 6575 45020 6695
rect 45140 6575 45185 6695
rect 45305 6575 45350 6695
rect 45470 6575 45525 6695
rect 45645 6575 45690 6695
rect 45810 6575 45855 6695
rect 45975 6575 46020 6695
rect 46140 6575 46195 6695
rect 46315 6575 46360 6695
rect 46480 6575 46525 6695
rect 46645 6575 46690 6695
rect 46810 6575 46865 6695
rect 46985 6575 47030 6695
rect 47150 6575 47195 6695
rect 47315 6575 47360 6695
rect 47480 6575 47535 6695
rect 47655 6575 47665 6695
rect 42165 6530 47665 6575
rect 42165 6410 42175 6530
rect 42295 6410 42340 6530
rect 42460 6410 42505 6530
rect 42625 6410 42670 6530
rect 42790 6410 42845 6530
rect 42965 6410 43010 6530
rect 43130 6410 43175 6530
rect 43295 6410 43340 6530
rect 43460 6410 43515 6530
rect 43635 6410 43680 6530
rect 43800 6410 43845 6530
rect 43965 6410 44010 6530
rect 44130 6410 44185 6530
rect 44305 6410 44350 6530
rect 44470 6410 44515 6530
rect 44635 6410 44680 6530
rect 44800 6410 44855 6530
rect 44975 6410 45020 6530
rect 45140 6410 45185 6530
rect 45305 6410 45350 6530
rect 45470 6410 45525 6530
rect 45645 6410 45690 6530
rect 45810 6410 45855 6530
rect 45975 6410 46020 6530
rect 46140 6410 46195 6530
rect 46315 6410 46360 6530
rect 46480 6410 46525 6530
rect 46645 6410 46690 6530
rect 46810 6410 46865 6530
rect 46985 6410 47030 6530
rect 47150 6410 47195 6530
rect 47315 6410 47360 6530
rect 47480 6410 47535 6530
rect 47655 6410 47665 6530
rect 42165 6355 47665 6410
rect 42165 6235 42175 6355
rect 42295 6235 42340 6355
rect 42460 6235 42505 6355
rect 42625 6235 42670 6355
rect 42790 6235 42845 6355
rect 42965 6235 43010 6355
rect 43130 6235 43175 6355
rect 43295 6235 43340 6355
rect 43460 6235 43515 6355
rect 43635 6235 43680 6355
rect 43800 6235 43845 6355
rect 43965 6235 44010 6355
rect 44130 6235 44185 6355
rect 44305 6235 44350 6355
rect 44470 6235 44515 6355
rect 44635 6235 44680 6355
rect 44800 6235 44855 6355
rect 44975 6235 45020 6355
rect 45140 6235 45185 6355
rect 45305 6235 45350 6355
rect 45470 6235 45525 6355
rect 45645 6235 45690 6355
rect 45810 6235 45855 6355
rect 45975 6235 46020 6355
rect 46140 6235 46195 6355
rect 46315 6235 46360 6355
rect 46480 6235 46525 6355
rect 46645 6235 46690 6355
rect 46810 6235 46865 6355
rect 46985 6235 47030 6355
rect 47150 6235 47195 6355
rect 47315 6235 47360 6355
rect 47480 6235 47535 6355
rect 47655 6235 47665 6355
rect 42165 6190 47665 6235
rect 42165 6070 42175 6190
rect 42295 6070 42340 6190
rect 42460 6070 42505 6190
rect 42625 6070 42670 6190
rect 42790 6070 42845 6190
rect 42965 6070 43010 6190
rect 43130 6070 43175 6190
rect 43295 6070 43340 6190
rect 43460 6070 43515 6190
rect 43635 6070 43680 6190
rect 43800 6070 43845 6190
rect 43965 6070 44010 6190
rect 44130 6070 44185 6190
rect 44305 6070 44350 6190
rect 44470 6070 44515 6190
rect 44635 6070 44680 6190
rect 44800 6070 44855 6190
rect 44975 6070 45020 6190
rect 45140 6070 45185 6190
rect 45305 6070 45350 6190
rect 45470 6070 45525 6190
rect 45645 6070 45690 6190
rect 45810 6070 45855 6190
rect 45975 6070 46020 6190
rect 46140 6070 46195 6190
rect 46315 6070 46360 6190
rect 46480 6070 46525 6190
rect 46645 6070 46690 6190
rect 46810 6070 46865 6190
rect 46985 6070 47030 6190
rect 47150 6070 47195 6190
rect 47315 6070 47360 6190
rect 47480 6070 47535 6190
rect 47655 6070 47665 6190
rect 42165 6025 47665 6070
rect 42165 5905 42175 6025
rect 42295 5905 42340 6025
rect 42460 5905 42505 6025
rect 42625 5905 42670 6025
rect 42790 5905 42845 6025
rect 42965 5905 43010 6025
rect 43130 5905 43175 6025
rect 43295 5905 43340 6025
rect 43460 5905 43515 6025
rect 43635 5905 43680 6025
rect 43800 5905 43845 6025
rect 43965 5905 44010 6025
rect 44130 5905 44185 6025
rect 44305 5905 44350 6025
rect 44470 5905 44515 6025
rect 44635 5905 44680 6025
rect 44800 5905 44855 6025
rect 44975 5905 45020 6025
rect 45140 5905 45185 6025
rect 45305 5905 45350 6025
rect 45470 5905 45525 6025
rect 45645 5905 45690 6025
rect 45810 5905 45855 6025
rect 45975 5905 46020 6025
rect 46140 5905 46195 6025
rect 46315 5905 46360 6025
rect 46480 5905 46525 6025
rect 46645 5905 46690 6025
rect 46810 5905 46865 6025
rect 46985 5905 47030 6025
rect 47150 5905 47195 6025
rect 47315 5905 47360 6025
rect 47480 5905 47535 6025
rect 47655 5905 47665 6025
rect 42165 5860 47665 5905
rect 42165 5740 42175 5860
rect 42295 5740 42340 5860
rect 42460 5740 42505 5860
rect 42625 5740 42670 5860
rect 42790 5740 42845 5860
rect 42965 5740 43010 5860
rect 43130 5740 43175 5860
rect 43295 5740 43340 5860
rect 43460 5740 43515 5860
rect 43635 5740 43680 5860
rect 43800 5740 43845 5860
rect 43965 5740 44010 5860
rect 44130 5740 44185 5860
rect 44305 5740 44350 5860
rect 44470 5740 44515 5860
rect 44635 5740 44680 5860
rect 44800 5740 44855 5860
rect 44975 5740 45020 5860
rect 45140 5740 45185 5860
rect 45305 5740 45350 5860
rect 45470 5740 45525 5860
rect 45645 5740 45690 5860
rect 45810 5740 45855 5860
rect 45975 5740 46020 5860
rect 46140 5740 46195 5860
rect 46315 5740 46360 5860
rect 46480 5740 46525 5860
rect 46645 5740 46690 5860
rect 46810 5740 46865 5860
rect 46985 5740 47030 5860
rect 47150 5740 47195 5860
rect 47315 5740 47360 5860
rect 47480 5740 47535 5860
rect 47655 5740 47665 5860
rect 42165 5685 47665 5740
rect 42165 5565 42175 5685
rect 42295 5565 42340 5685
rect 42460 5565 42505 5685
rect 42625 5565 42670 5685
rect 42790 5565 42845 5685
rect 42965 5565 43010 5685
rect 43130 5565 43175 5685
rect 43295 5565 43340 5685
rect 43460 5565 43515 5685
rect 43635 5565 43680 5685
rect 43800 5565 43845 5685
rect 43965 5565 44010 5685
rect 44130 5565 44185 5685
rect 44305 5565 44350 5685
rect 44470 5565 44515 5685
rect 44635 5565 44680 5685
rect 44800 5565 44855 5685
rect 44975 5565 45020 5685
rect 45140 5565 45185 5685
rect 45305 5565 45350 5685
rect 45470 5565 45525 5685
rect 45645 5565 45690 5685
rect 45810 5565 45855 5685
rect 45975 5565 46020 5685
rect 46140 5565 46195 5685
rect 46315 5565 46360 5685
rect 46480 5565 46525 5685
rect 46645 5565 46690 5685
rect 46810 5565 46865 5685
rect 46985 5565 47030 5685
rect 47150 5565 47195 5685
rect 47315 5565 47360 5685
rect 47480 5565 47535 5685
rect 47655 5565 47665 5685
rect 42165 5520 47665 5565
rect 42165 5400 42175 5520
rect 42295 5400 42340 5520
rect 42460 5400 42505 5520
rect 42625 5400 42670 5520
rect 42790 5400 42845 5520
rect 42965 5400 43010 5520
rect 43130 5400 43175 5520
rect 43295 5400 43340 5520
rect 43460 5400 43515 5520
rect 43635 5400 43680 5520
rect 43800 5400 43845 5520
rect 43965 5400 44010 5520
rect 44130 5400 44185 5520
rect 44305 5400 44350 5520
rect 44470 5400 44515 5520
rect 44635 5400 44680 5520
rect 44800 5400 44855 5520
rect 44975 5400 45020 5520
rect 45140 5400 45185 5520
rect 45305 5400 45350 5520
rect 45470 5400 45525 5520
rect 45645 5400 45690 5520
rect 45810 5400 45855 5520
rect 45975 5400 46020 5520
rect 46140 5400 46195 5520
rect 46315 5400 46360 5520
rect 46480 5400 46525 5520
rect 46645 5400 46690 5520
rect 46810 5400 46865 5520
rect 46985 5400 47030 5520
rect 47150 5400 47195 5520
rect 47315 5400 47360 5520
rect 47480 5400 47535 5520
rect 47655 5400 47665 5520
rect 42165 5355 47665 5400
rect 42165 5235 42175 5355
rect 42295 5235 42340 5355
rect 42460 5235 42505 5355
rect 42625 5235 42670 5355
rect 42790 5235 42845 5355
rect 42965 5235 43010 5355
rect 43130 5235 43175 5355
rect 43295 5235 43340 5355
rect 43460 5235 43515 5355
rect 43635 5235 43680 5355
rect 43800 5235 43845 5355
rect 43965 5235 44010 5355
rect 44130 5235 44185 5355
rect 44305 5235 44350 5355
rect 44470 5235 44515 5355
rect 44635 5235 44680 5355
rect 44800 5235 44855 5355
rect 44975 5235 45020 5355
rect 45140 5235 45185 5355
rect 45305 5235 45350 5355
rect 45470 5235 45525 5355
rect 45645 5235 45690 5355
rect 45810 5235 45855 5355
rect 45975 5235 46020 5355
rect 46140 5235 46195 5355
rect 46315 5235 46360 5355
rect 46480 5235 46525 5355
rect 46645 5235 46690 5355
rect 46810 5235 46865 5355
rect 46985 5235 47030 5355
rect 47150 5235 47195 5355
rect 47315 5235 47360 5355
rect 47480 5235 47535 5355
rect 47655 5235 47665 5355
rect 42165 5190 47665 5235
rect 42165 5070 42175 5190
rect 42295 5070 42340 5190
rect 42460 5070 42505 5190
rect 42625 5070 42670 5190
rect 42790 5070 42845 5190
rect 42965 5070 43010 5190
rect 43130 5070 43175 5190
rect 43295 5070 43340 5190
rect 43460 5070 43515 5190
rect 43635 5070 43680 5190
rect 43800 5070 43845 5190
rect 43965 5070 44010 5190
rect 44130 5070 44185 5190
rect 44305 5070 44350 5190
rect 44470 5070 44515 5190
rect 44635 5070 44680 5190
rect 44800 5070 44855 5190
rect 44975 5070 45020 5190
rect 45140 5070 45185 5190
rect 45305 5070 45350 5190
rect 45470 5070 45525 5190
rect 45645 5070 45690 5190
rect 45810 5070 45855 5190
rect 45975 5070 46020 5190
rect 46140 5070 46195 5190
rect 46315 5070 46360 5190
rect 46480 5070 46525 5190
rect 46645 5070 46690 5190
rect 46810 5070 46865 5190
rect 46985 5070 47030 5190
rect 47150 5070 47195 5190
rect 47315 5070 47360 5190
rect 47480 5070 47535 5190
rect 47655 5070 47665 5190
rect 42165 5015 47665 5070
rect 42165 4895 42175 5015
rect 42295 4895 42340 5015
rect 42460 4895 42505 5015
rect 42625 4895 42670 5015
rect 42790 4895 42845 5015
rect 42965 4895 43010 5015
rect 43130 4895 43175 5015
rect 43295 4895 43340 5015
rect 43460 4895 43515 5015
rect 43635 4895 43680 5015
rect 43800 4895 43845 5015
rect 43965 4895 44010 5015
rect 44130 4895 44185 5015
rect 44305 4895 44350 5015
rect 44470 4895 44515 5015
rect 44635 4895 44680 5015
rect 44800 4895 44855 5015
rect 44975 4895 45020 5015
rect 45140 4895 45185 5015
rect 45305 4895 45350 5015
rect 45470 4895 45525 5015
rect 45645 4895 45690 5015
rect 45810 4895 45855 5015
rect 45975 4895 46020 5015
rect 46140 4895 46195 5015
rect 46315 4895 46360 5015
rect 46480 4895 46525 5015
rect 46645 4895 46690 5015
rect 46810 4895 46865 5015
rect 46985 4895 47030 5015
rect 47150 4895 47195 5015
rect 47315 4895 47360 5015
rect 47480 4895 47535 5015
rect 47655 4895 47665 5015
rect 42165 4850 47665 4895
rect 42165 4730 42175 4850
rect 42295 4730 42340 4850
rect 42460 4730 42505 4850
rect 42625 4730 42670 4850
rect 42790 4730 42845 4850
rect 42965 4730 43010 4850
rect 43130 4730 43175 4850
rect 43295 4730 43340 4850
rect 43460 4730 43515 4850
rect 43635 4730 43680 4850
rect 43800 4730 43845 4850
rect 43965 4730 44010 4850
rect 44130 4730 44185 4850
rect 44305 4730 44350 4850
rect 44470 4730 44515 4850
rect 44635 4730 44680 4850
rect 44800 4730 44855 4850
rect 44975 4730 45020 4850
rect 45140 4730 45185 4850
rect 45305 4730 45350 4850
rect 45470 4730 45525 4850
rect 45645 4730 45690 4850
rect 45810 4730 45855 4850
rect 45975 4730 46020 4850
rect 46140 4730 46195 4850
rect 46315 4730 46360 4850
rect 46480 4730 46525 4850
rect 46645 4730 46690 4850
rect 46810 4730 46865 4850
rect 46985 4730 47030 4850
rect 47150 4730 47195 4850
rect 47315 4730 47360 4850
rect 47480 4730 47535 4850
rect 47655 4730 47665 4850
rect 42165 4685 47665 4730
rect 42165 4565 42175 4685
rect 42295 4565 42340 4685
rect 42460 4565 42505 4685
rect 42625 4565 42670 4685
rect 42790 4565 42845 4685
rect 42965 4565 43010 4685
rect 43130 4565 43175 4685
rect 43295 4565 43340 4685
rect 43460 4565 43515 4685
rect 43635 4565 43680 4685
rect 43800 4565 43845 4685
rect 43965 4565 44010 4685
rect 44130 4565 44185 4685
rect 44305 4565 44350 4685
rect 44470 4565 44515 4685
rect 44635 4565 44680 4685
rect 44800 4565 44855 4685
rect 44975 4565 45020 4685
rect 45140 4565 45185 4685
rect 45305 4565 45350 4685
rect 45470 4565 45525 4685
rect 45645 4565 45690 4685
rect 45810 4565 45855 4685
rect 45975 4565 46020 4685
rect 46140 4565 46195 4685
rect 46315 4565 46360 4685
rect 46480 4565 46525 4685
rect 46645 4565 46690 4685
rect 46810 4565 46865 4685
rect 46985 4565 47030 4685
rect 47150 4565 47195 4685
rect 47315 4565 47360 4685
rect 47480 4565 47535 4685
rect 47655 4565 47665 4685
rect 42165 4520 47665 4565
rect 42165 4400 42175 4520
rect 42295 4400 42340 4520
rect 42460 4400 42505 4520
rect 42625 4400 42670 4520
rect 42790 4400 42845 4520
rect 42965 4400 43010 4520
rect 43130 4400 43175 4520
rect 43295 4400 43340 4520
rect 43460 4400 43515 4520
rect 43635 4400 43680 4520
rect 43800 4400 43845 4520
rect 43965 4400 44010 4520
rect 44130 4400 44185 4520
rect 44305 4400 44350 4520
rect 44470 4400 44515 4520
rect 44635 4400 44680 4520
rect 44800 4400 44855 4520
rect 44975 4400 45020 4520
rect 45140 4400 45185 4520
rect 45305 4400 45350 4520
rect 45470 4400 45525 4520
rect 45645 4400 45690 4520
rect 45810 4400 45855 4520
rect 45975 4400 46020 4520
rect 46140 4400 46195 4520
rect 46315 4400 46360 4520
rect 46480 4400 46525 4520
rect 46645 4400 46690 4520
rect 46810 4400 46865 4520
rect 46985 4400 47030 4520
rect 47150 4400 47195 4520
rect 47315 4400 47360 4520
rect 47480 4400 47535 4520
rect 47655 4400 47665 4520
rect 42165 4345 47665 4400
rect 42165 4225 42175 4345
rect 42295 4225 42340 4345
rect 42460 4225 42505 4345
rect 42625 4225 42670 4345
rect 42790 4225 42845 4345
rect 42965 4225 43010 4345
rect 43130 4225 43175 4345
rect 43295 4225 43340 4345
rect 43460 4225 43515 4345
rect 43635 4225 43680 4345
rect 43800 4225 43845 4345
rect 43965 4225 44010 4345
rect 44130 4225 44185 4345
rect 44305 4225 44350 4345
rect 44470 4225 44515 4345
rect 44635 4225 44680 4345
rect 44800 4225 44855 4345
rect 44975 4225 45020 4345
rect 45140 4225 45185 4345
rect 45305 4225 45350 4345
rect 45470 4225 45525 4345
rect 45645 4225 45690 4345
rect 45810 4225 45855 4345
rect 45975 4225 46020 4345
rect 46140 4225 46195 4345
rect 46315 4225 46360 4345
rect 46480 4225 46525 4345
rect 46645 4225 46690 4345
rect 46810 4225 46865 4345
rect 46985 4225 47030 4345
rect 47150 4225 47195 4345
rect 47315 4225 47360 4345
rect 47480 4225 47535 4345
rect 47655 4225 47665 4345
rect 42165 4180 47665 4225
rect 42165 4060 42175 4180
rect 42295 4060 42340 4180
rect 42460 4060 42505 4180
rect 42625 4060 42670 4180
rect 42790 4060 42845 4180
rect 42965 4060 43010 4180
rect 43130 4060 43175 4180
rect 43295 4060 43340 4180
rect 43460 4060 43515 4180
rect 43635 4060 43680 4180
rect 43800 4060 43845 4180
rect 43965 4060 44010 4180
rect 44130 4060 44185 4180
rect 44305 4060 44350 4180
rect 44470 4060 44515 4180
rect 44635 4060 44680 4180
rect 44800 4060 44855 4180
rect 44975 4060 45020 4180
rect 45140 4060 45185 4180
rect 45305 4060 45350 4180
rect 45470 4060 45525 4180
rect 45645 4060 45690 4180
rect 45810 4060 45855 4180
rect 45975 4060 46020 4180
rect 46140 4060 46195 4180
rect 46315 4060 46360 4180
rect 46480 4060 46525 4180
rect 46645 4060 46690 4180
rect 46810 4060 46865 4180
rect 46985 4060 47030 4180
rect 47150 4060 47195 4180
rect 47315 4060 47360 4180
rect 47480 4060 47535 4180
rect 47655 4060 47665 4180
rect 42165 4015 47665 4060
rect 42165 3895 42175 4015
rect 42295 3895 42340 4015
rect 42460 3895 42505 4015
rect 42625 3895 42670 4015
rect 42790 3895 42845 4015
rect 42965 3895 43010 4015
rect 43130 3895 43175 4015
rect 43295 3895 43340 4015
rect 43460 3895 43515 4015
rect 43635 3895 43680 4015
rect 43800 3895 43845 4015
rect 43965 3895 44010 4015
rect 44130 3895 44185 4015
rect 44305 3895 44350 4015
rect 44470 3895 44515 4015
rect 44635 3895 44680 4015
rect 44800 3895 44855 4015
rect 44975 3895 45020 4015
rect 45140 3895 45185 4015
rect 45305 3895 45350 4015
rect 45470 3895 45525 4015
rect 45645 3895 45690 4015
rect 45810 3895 45855 4015
rect 45975 3895 46020 4015
rect 46140 3895 46195 4015
rect 46315 3895 46360 4015
rect 46480 3895 46525 4015
rect 46645 3895 46690 4015
rect 46810 3895 46865 4015
rect 46985 3895 47030 4015
rect 47150 3895 47195 4015
rect 47315 3895 47360 4015
rect 47480 3895 47535 4015
rect 47655 3895 47665 4015
rect 42165 3850 47665 3895
rect 42165 3730 42175 3850
rect 42295 3730 42340 3850
rect 42460 3730 42505 3850
rect 42625 3730 42670 3850
rect 42790 3730 42845 3850
rect 42965 3730 43010 3850
rect 43130 3730 43175 3850
rect 43295 3730 43340 3850
rect 43460 3730 43515 3850
rect 43635 3730 43680 3850
rect 43800 3730 43845 3850
rect 43965 3730 44010 3850
rect 44130 3730 44185 3850
rect 44305 3730 44350 3850
rect 44470 3730 44515 3850
rect 44635 3730 44680 3850
rect 44800 3730 44855 3850
rect 44975 3730 45020 3850
rect 45140 3730 45185 3850
rect 45305 3730 45350 3850
rect 45470 3730 45525 3850
rect 45645 3730 45690 3850
rect 45810 3730 45855 3850
rect 45975 3730 46020 3850
rect 46140 3730 46195 3850
rect 46315 3730 46360 3850
rect 46480 3730 46525 3850
rect 46645 3730 46690 3850
rect 46810 3730 46865 3850
rect 46985 3730 47030 3850
rect 47150 3730 47195 3850
rect 47315 3730 47360 3850
rect 47480 3730 47535 3850
rect 47655 3730 47665 3850
rect 42165 3675 47665 3730
rect 42165 3555 42175 3675
rect 42295 3555 42340 3675
rect 42460 3555 42505 3675
rect 42625 3555 42670 3675
rect 42790 3555 42845 3675
rect 42965 3555 43010 3675
rect 43130 3555 43175 3675
rect 43295 3555 43340 3675
rect 43460 3555 43515 3675
rect 43635 3555 43680 3675
rect 43800 3555 43845 3675
rect 43965 3555 44010 3675
rect 44130 3555 44185 3675
rect 44305 3555 44350 3675
rect 44470 3555 44515 3675
rect 44635 3555 44680 3675
rect 44800 3555 44855 3675
rect 44975 3555 45020 3675
rect 45140 3555 45185 3675
rect 45305 3555 45350 3675
rect 45470 3555 45525 3675
rect 45645 3555 45690 3675
rect 45810 3555 45855 3675
rect 45975 3555 46020 3675
rect 46140 3555 46195 3675
rect 46315 3555 46360 3675
rect 46480 3555 46525 3675
rect 46645 3555 46690 3675
rect 46810 3555 46865 3675
rect 46985 3555 47030 3675
rect 47150 3555 47195 3675
rect 47315 3555 47360 3675
rect 47480 3555 47535 3675
rect 47655 3555 47665 3675
rect 42165 3510 47665 3555
rect 42165 3390 42175 3510
rect 42295 3390 42340 3510
rect 42460 3390 42505 3510
rect 42625 3390 42670 3510
rect 42790 3390 42845 3510
rect 42965 3390 43010 3510
rect 43130 3390 43175 3510
rect 43295 3390 43340 3510
rect 43460 3390 43515 3510
rect 43635 3390 43680 3510
rect 43800 3390 43845 3510
rect 43965 3390 44010 3510
rect 44130 3390 44185 3510
rect 44305 3390 44350 3510
rect 44470 3390 44515 3510
rect 44635 3390 44680 3510
rect 44800 3390 44855 3510
rect 44975 3390 45020 3510
rect 45140 3390 45185 3510
rect 45305 3390 45350 3510
rect 45470 3390 45525 3510
rect 45645 3390 45690 3510
rect 45810 3390 45855 3510
rect 45975 3390 46020 3510
rect 46140 3390 46195 3510
rect 46315 3390 46360 3510
rect 46480 3390 46525 3510
rect 46645 3390 46690 3510
rect 46810 3390 46865 3510
rect 46985 3390 47030 3510
rect 47150 3390 47195 3510
rect 47315 3390 47360 3510
rect 47480 3390 47535 3510
rect 47655 3390 47665 3510
rect 42165 3345 47665 3390
rect 42165 3225 42175 3345
rect 42295 3225 42340 3345
rect 42460 3225 42505 3345
rect 42625 3225 42670 3345
rect 42790 3225 42845 3345
rect 42965 3225 43010 3345
rect 43130 3225 43175 3345
rect 43295 3225 43340 3345
rect 43460 3225 43515 3345
rect 43635 3225 43680 3345
rect 43800 3225 43845 3345
rect 43965 3225 44010 3345
rect 44130 3225 44185 3345
rect 44305 3225 44350 3345
rect 44470 3225 44515 3345
rect 44635 3225 44680 3345
rect 44800 3225 44855 3345
rect 44975 3225 45020 3345
rect 45140 3225 45185 3345
rect 45305 3225 45350 3345
rect 45470 3225 45525 3345
rect 45645 3225 45690 3345
rect 45810 3225 45855 3345
rect 45975 3225 46020 3345
rect 46140 3225 46195 3345
rect 46315 3225 46360 3345
rect 46480 3225 46525 3345
rect 46645 3225 46690 3345
rect 46810 3225 46865 3345
rect 46985 3225 47030 3345
rect 47150 3225 47195 3345
rect 47315 3225 47360 3345
rect 47480 3225 47535 3345
rect 47655 3225 47665 3345
rect 42165 3180 47665 3225
rect 42165 3060 42175 3180
rect 42295 3060 42340 3180
rect 42460 3060 42505 3180
rect 42625 3060 42670 3180
rect 42790 3060 42845 3180
rect 42965 3060 43010 3180
rect 43130 3060 43175 3180
rect 43295 3060 43340 3180
rect 43460 3060 43515 3180
rect 43635 3060 43680 3180
rect 43800 3060 43845 3180
rect 43965 3060 44010 3180
rect 44130 3060 44185 3180
rect 44305 3060 44350 3180
rect 44470 3060 44515 3180
rect 44635 3060 44680 3180
rect 44800 3060 44855 3180
rect 44975 3060 45020 3180
rect 45140 3060 45185 3180
rect 45305 3060 45350 3180
rect 45470 3060 45525 3180
rect 45645 3060 45690 3180
rect 45810 3060 45855 3180
rect 45975 3060 46020 3180
rect 46140 3060 46195 3180
rect 46315 3060 46360 3180
rect 46480 3060 46525 3180
rect 46645 3060 46690 3180
rect 46810 3060 46865 3180
rect 46985 3060 47030 3180
rect 47150 3060 47195 3180
rect 47315 3060 47360 3180
rect 47480 3060 47535 3180
rect 47655 3060 47665 3180
rect 42165 3005 47665 3060
rect 42165 2885 42175 3005
rect 42295 2885 42340 3005
rect 42460 2885 42505 3005
rect 42625 2885 42670 3005
rect 42790 2885 42845 3005
rect 42965 2885 43010 3005
rect 43130 2885 43175 3005
rect 43295 2885 43340 3005
rect 43460 2885 43515 3005
rect 43635 2885 43680 3005
rect 43800 2885 43845 3005
rect 43965 2885 44010 3005
rect 44130 2885 44185 3005
rect 44305 2885 44350 3005
rect 44470 2885 44515 3005
rect 44635 2885 44680 3005
rect 44800 2885 44855 3005
rect 44975 2885 45020 3005
rect 45140 2885 45185 3005
rect 45305 2885 45350 3005
rect 45470 2885 45525 3005
rect 45645 2885 45690 3005
rect 45810 2885 45855 3005
rect 45975 2885 46020 3005
rect 46140 2885 46195 3005
rect 46315 2885 46360 3005
rect 46480 2885 46525 3005
rect 46645 2885 46690 3005
rect 46810 2885 46865 3005
rect 46985 2885 47030 3005
rect 47150 2885 47195 3005
rect 47315 2885 47360 3005
rect 47480 2885 47535 3005
rect 47655 2885 47665 3005
rect 42165 2840 47665 2885
rect 42165 2720 42175 2840
rect 42295 2720 42340 2840
rect 42460 2720 42505 2840
rect 42625 2720 42670 2840
rect 42790 2720 42845 2840
rect 42965 2720 43010 2840
rect 43130 2720 43175 2840
rect 43295 2720 43340 2840
rect 43460 2720 43515 2840
rect 43635 2720 43680 2840
rect 43800 2720 43845 2840
rect 43965 2720 44010 2840
rect 44130 2720 44185 2840
rect 44305 2720 44350 2840
rect 44470 2720 44515 2840
rect 44635 2720 44680 2840
rect 44800 2720 44855 2840
rect 44975 2720 45020 2840
rect 45140 2720 45185 2840
rect 45305 2720 45350 2840
rect 45470 2720 45525 2840
rect 45645 2720 45690 2840
rect 45810 2720 45855 2840
rect 45975 2720 46020 2840
rect 46140 2720 46195 2840
rect 46315 2720 46360 2840
rect 46480 2720 46525 2840
rect 46645 2720 46690 2840
rect 46810 2720 46865 2840
rect 46985 2720 47030 2840
rect 47150 2720 47195 2840
rect 47315 2720 47360 2840
rect 47480 2720 47535 2840
rect 47655 2720 47665 2840
rect 42165 2675 47665 2720
rect 42165 2555 42175 2675
rect 42295 2555 42340 2675
rect 42460 2555 42505 2675
rect 42625 2555 42670 2675
rect 42790 2555 42845 2675
rect 42965 2555 43010 2675
rect 43130 2555 43175 2675
rect 43295 2555 43340 2675
rect 43460 2555 43515 2675
rect 43635 2555 43680 2675
rect 43800 2555 43845 2675
rect 43965 2555 44010 2675
rect 44130 2555 44185 2675
rect 44305 2555 44350 2675
rect 44470 2555 44515 2675
rect 44635 2555 44680 2675
rect 44800 2555 44855 2675
rect 44975 2555 45020 2675
rect 45140 2555 45185 2675
rect 45305 2555 45350 2675
rect 45470 2555 45525 2675
rect 45645 2555 45690 2675
rect 45810 2555 45855 2675
rect 45975 2555 46020 2675
rect 46140 2555 46195 2675
rect 46315 2555 46360 2675
rect 46480 2555 46525 2675
rect 46645 2555 46690 2675
rect 46810 2555 46865 2675
rect 46985 2555 47030 2675
rect 47150 2555 47195 2675
rect 47315 2555 47360 2675
rect 47480 2555 47535 2675
rect 47655 2555 47665 2675
rect 42165 2510 47665 2555
rect 42165 2390 42175 2510
rect 42295 2390 42340 2510
rect 42460 2390 42505 2510
rect 42625 2390 42670 2510
rect 42790 2390 42845 2510
rect 42965 2390 43010 2510
rect 43130 2390 43175 2510
rect 43295 2390 43340 2510
rect 43460 2390 43515 2510
rect 43635 2390 43680 2510
rect 43800 2390 43845 2510
rect 43965 2390 44010 2510
rect 44130 2390 44185 2510
rect 44305 2390 44350 2510
rect 44470 2390 44515 2510
rect 44635 2390 44680 2510
rect 44800 2390 44855 2510
rect 44975 2390 45020 2510
rect 45140 2390 45185 2510
rect 45305 2390 45350 2510
rect 45470 2390 45525 2510
rect 45645 2390 45690 2510
rect 45810 2390 45855 2510
rect 45975 2390 46020 2510
rect 46140 2390 46195 2510
rect 46315 2390 46360 2510
rect 46480 2390 46525 2510
rect 46645 2390 46690 2510
rect 46810 2390 46865 2510
rect 46985 2390 47030 2510
rect 47150 2390 47195 2510
rect 47315 2390 47360 2510
rect 47480 2390 47535 2510
rect 47655 2390 47665 2510
rect 42165 2335 47665 2390
rect 42165 2215 42175 2335
rect 42295 2215 42340 2335
rect 42460 2215 42505 2335
rect 42625 2215 42670 2335
rect 42790 2215 42845 2335
rect 42965 2215 43010 2335
rect 43130 2215 43175 2335
rect 43295 2215 43340 2335
rect 43460 2215 43515 2335
rect 43635 2215 43680 2335
rect 43800 2215 43845 2335
rect 43965 2215 44010 2335
rect 44130 2215 44185 2335
rect 44305 2215 44350 2335
rect 44470 2215 44515 2335
rect 44635 2215 44680 2335
rect 44800 2215 44855 2335
rect 44975 2215 45020 2335
rect 45140 2215 45185 2335
rect 45305 2215 45350 2335
rect 45470 2215 45525 2335
rect 45645 2215 45690 2335
rect 45810 2215 45855 2335
rect 45975 2215 46020 2335
rect 46140 2215 46195 2335
rect 46315 2215 46360 2335
rect 46480 2215 46525 2335
rect 46645 2215 46690 2335
rect 46810 2215 46865 2335
rect 46985 2215 47030 2335
rect 47150 2215 47195 2335
rect 47315 2215 47360 2335
rect 47480 2215 47535 2335
rect 47655 2215 47665 2335
rect 42165 2170 47665 2215
rect 42165 2050 42175 2170
rect 42295 2050 42340 2170
rect 42460 2050 42505 2170
rect 42625 2050 42670 2170
rect 42790 2050 42845 2170
rect 42965 2050 43010 2170
rect 43130 2050 43175 2170
rect 43295 2050 43340 2170
rect 43460 2050 43515 2170
rect 43635 2050 43680 2170
rect 43800 2050 43845 2170
rect 43965 2050 44010 2170
rect 44130 2050 44185 2170
rect 44305 2050 44350 2170
rect 44470 2050 44515 2170
rect 44635 2050 44680 2170
rect 44800 2050 44855 2170
rect 44975 2050 45020 2170
rect 45140 2050 45185 2170
rect 45305 2050 45350 2170
rect 45470 2050 45525 2170
rect 45645 2050 45690 2170
rect 45810 2050 45855 2170
rect 45975 2050 46020 2170
rect 46140 2050 46195 2170
rect 46315 2050 46360 2170
rect 46480 2050 46525 2170
rect 46645 2050 46690 2170
rect 46810 2050 46865 2170
rect 46985 2050 47030 2170
rect 47150 2050 47195 2170
rect 47315 2050 47360 2170
rect 47480 2050 47535 2170
rect 47655 2050 47665 2170
rect 42165 2005 47665 2050
rect 42165 1885 42175 2005
rect 42295 1885 42340 2005
rect 42460 1885 42505 2005
rect 42625 1885 42670 2005
rect 42790 1885 42845 2005
rect 42965 1885 43010 2005
rect 43130 1885 43175 2005
rect 43295 1885 43340 2005
rect 43460 1885 43515 2005
rect 43635 1885 43680 2005
rect 43800 1885 43845 2005
rect 43965 1885 44010 2005
rect 44130 1885 44185 2005
rect 44305 1885 44350 2005
rect 44470 1885 44515 2005
rect 44635 1885 44680 2005
rect 44800 1885 44855 2005
rect 44975 1885 45020 2005
rect 45140 1885 45185 2005
rect 45305 1885 45350 2005
rect 45470 1885 45525 2005
rect 45645 1885 45690 2005
rect 45810 1885 45855 2005
rect 45975 1885 46020 2005
rect 46140 1885 46195 2005
rect 46315 1885 46360 2005
rect 46480 1885 46525 2005
rect 46645 1885 46690 2005
rect 46810 1885 46865 2005
rect 46985 1885 47030 2005
rect 47150 1885 47195 2005
rect 47315 1885 47360 2005
rect 47480 1885 47535 2005
rect 47655 1885 47665 2005
rect 42165 1840 47665 1885
rect 42165 1720 42175 1840
rect 42295 1720 42340 1840
rect 42460 1720 42505 1840
rect 42625 1720 42670 1840
rect 42790 1720 42845 1840
rect 42965 1720 43010 1840
rect 43130 1720 43175 1840
rect 43295 1720 43340 1840
rect 43460 1720 43515 1840
rect 43635 1720 43680 1840
rect 43800 1720 43845 1840
rect 43965 1720 44010 1840
rect 44130 1720 44185 1840
rect 44305 1720 44350 1840
rect 44470 1720 44515 1840
rect 44635 1720 44680 1840
rect 44800 1720 44855 1840
rect 44975 1720 45020 1840
rect 45140 1720 45185 1840
rect 45305 1720 45350 1840
rect 45470 1720 45525 1840
rect 45645 1720 45690 1840
rect 45810 1720 45855 1840
rect 45975 1720 46020 1840
rect 46140 1720 46195 1840
rect 46315 1720 46360 1840
rect 46480 1720 46525 1840
rect 46645 1720 46690 1840
rect 46810 1720 46865 1840
rect 46985 1720 47030 1840
rect 47150 1720 47195 1840
rect 47315 1720 47360 1840
rect 47480 1720 47535 1840
rect 47655 1720 47665 1840
rect 42165 1710 47665 1720
rect 47855 7200 53355 7210
rect 47855 7080 47865 7200
rect 47985 7080 48030 7200
rect 48150 7080 48195 7200
rect 48315 7080 48360 7200
rect 48480 7080 48535 7200
rect 48655 7080 48700 7200
rect 48820 7080 48865 7200
rect 48985 7080 49030 7200
rect 49150 7080 49205 7200
rect 49325 7080 49370 7200
rect 49490 7080 49535 7200
rect 49655 7080 49700 7200
rect 49820 7080 49875 7200
rect 49995 7080 50040 7200
rect 50160 7080 50205 7200
rect 50325 7080 50370 7200
rect 50490 7080 50545 7200
rect 50665 7080 50710 7200
rect 50830 7080 50875 7200
rect 50995 7080 51040 7200
rect 51160 7080 51215 7200
rect 51335 7080 51380 7200
rect 51500 7080 51545 7200
rect 51665 7080 51710 7200
rect 51830 7080 51885 7200
rect 52005 7080 52050 7200
rect 52170 7080 52215 7200
rect 52335 7080 52380 7200
rect 52500 7080 52555 7200
rect 52675 7080 52720 7200
rect 52840 7080 52885 7200
rect 53005 7080 53050 7200
rect 53170 7080 53225 7200
rect 53345 7080 53355 7200
rect 47855 7025 53355 7080
rect 47855 6905 47865 7025
rect 47985 6905 48030 7025
rect 48150 6905 48195 7025
rect 48315 6905 48360 7025
rect 48480 6905 48535 7025
rect 48655 6905 48700 7025
rect 48820 6905 48865 7025
rect 48985 6905 49030 7025
rect 49150 6905 49205 7025
rect 49325 6905 49370 7025
rect 49490 6905 49535 7025
rect 49655 6905 49700 7025
rect 49820 6905 49875 7025
rect 49995 6905 50040 7025
rect 50160 6905 50205 7025
rect 50325 6905 50370 7025
rect 50490 6905 50545 7025
rect 50665 6905 50710 7025
rect 50830 6905 50875 7025
rect 50995 6905 51040 7025
rect 51160 6905 51215 7025
rect 51335 6905 51380 7025
rect 51500 6905 51545 7025
rect 51665 6905 51710 7025
rect 51830 6905 51885 7025
rect 52005 6905 52050 7025
rect 52170 6905 52215 7025
rect 52335 6905 52380 7025
rect 52500 6905 52555 7025
rect 52675 6905 52720 7025
rect 52840 6905 52885 7025
rect 53005 6905 53050 7025
rect 53170 6905 53225 7025
rect 53345 6905 53355 7025
rect 47855 6860 53355 6905
rect 47855 6740 47865 6860
rect 47985 6740 48030 6860
rect 48150 6740 48195 6860
rect 48315 6740 48360 6860
rect 48480 6740 48535 6860
rect 48655 6740 48700 6860
rect 48820 6740 48865 6860
rect 48985 6740 49030 6860
rect 49150 6740 49205 6860
rect 49325 6740 49370 6860
rect 49490 6740 49535 6860
rect 49655 6740 49700 6860
rect 49820 6740 49875 6860
rect 49995 6740 50040 6860
rect 50160 6740 50205 6860
rect 50325 6740 50370 6860
rect 50490 6740 50545 6860
rect 50665 6740 50710 6860
rect 50830 6740 50875 6860
rect 50995 6740 51040 6860
rect 51160 6740 51215 6860
rect 51335 6740 51380 6860
rect 51500 6740 51545 6860
rect 51665 6740 51710 6860
rect 51830 6740 51885 6860
rect 52005 6740 52050 6860
rect 52170 6740 52215 6860
rect 52335 6740 52380 6860
rect 52500 6740 52555 6860
rect 52675 6740 52720 6860
rect 52840 6740 52885 6860
rect 53005 6740 53050 6860
rect 53170 6740 53225 6860
rect 53345 6740 53355 6860
rect 47855 6695 53355 6740
rect 47855 6575 47865 6695
rect 47985 6575 48030 6695
rect 48150 6575 48195 6695
rect 48315 6575 48360 6695
rect 48480 6575 48535 6695
rect 48655 6575 48700 6695
rect 48820 6575 48865 6695
rect 48985 6575 49030 6695
rect 49150 6575 49205 6695
rect 49325 6575 49370 6695
rect 49490 6575 49535 6695
rect 49655 6575 49700 6695
rect 49820 6575 49875 6695
rect 49995 6575 50040 6695
rect 50160 6575 50205 6695
rect 50325 6575 50370 6695
rect 50490 6575 50545 6695
rect 50665 6575 50710 6695
rect 50830 6575 50875 6695
rect 50995 6575 51040 6695
rect 51160 6575 51215 6695
rect 51335 6575 51380 6695
rect 51500 6575 51545 6695
rect 51665 6575 51710 6695
rect 51830 6575 51885 6695
rect 52005 6575 52050 6695
rect 52170 6575 52215 6695
rect 52335 6575 52380 6695
rect 52500 6575 52555 6695
rect 52675 6575 52720 6695
rect 52840 6575 52885 6695
rect 53005 6575 53050 6695
rect 53170 6575 53225 6695
rect 53345 6575 53355 6695
rect 47855 6530 53355 6575
rect 47855 6410 47865 6530
rect 47985 6410 48030 6530
rect 48150 6410 48195 6530
rect 48315 6410 48360 6530
rect 48480 6410 48535 6530
rect 48655 6410 48700 6530
rect 48820 6410 48865 6530
rect 48985 6410 49030 6530
rect 49150 6410 49205 6530
rect 49325 6410 49370 6530
rect 49490 6410 49535 6530
rect 49655 6410 49700 6530
rect 49820 6410 49875 6530
rect 49995 6410 50040 6530
rect 50160 6410 50205 6530
rect 50325 6410 50370 6530
rect 50490 6410 50545 6530
rect 50665 6410 50710 6530
rect 50830 6410 50875 6530
rect 50995 6410 51040 6530
rect 51160 6410 51215 6530
rect 51335 6410 51380 6530
rect 51500 6410 51545 6530
rect 51665 6410 51710 6530
rect 51830 6410 51885 6530
rect 52005 6410 52050 6530
rect 52170 6410 52215 6530
rect 52335 6410 52380 6530
rect 52500 6410 52555 6530
rect 52675 6410 52720 6530
rect 52840 6410 52885 6530
rect 53005 6410 53050 6530
rect 53170 6410 53225 6530
rect 53345 6410 53355 6530
rect 47855 6355 53355 6410
rect 47855 6235 47865 6355
rect 47985 6235 48030 6355
rect 48150 6235 48195 6355
rect 48315 6235 48360 6355
rect 48480 6235 48535 6355
rect 48655 6235 48700 6355
rect 48820 6235 48865 6355
rect 48985 6235 49030 6355
rect 49150 6235 49205 6355
rect 49325 6235 49370 6355
rect 49490 6235 49535 6355
rect 49655 6235 49700 6355
rect 49820 6235 49875 6355
rect 49995 6235 50040 6355
rect 50160 6235 50205 6355
rect 50325 6235 50370 6355
rect 50490 6235 50545 6355
rect 50665 6235 50710 6355
rect 50830 6235 50875 6355
rect 50995 6235 51040 6355
rect 51160 6235 51215 6355
rect 51335 6235 51380 6355
rect 51500 6235 51545 6355
rect 51665 6235 51710 6355
rect 51830 6235 51885 6355
rect 52005 6235 52050 6355
rect 52170 6235 52215 6355
rect 52335 6235 52380 6355
rect 52500 6235 52555 6355
rect 52675 6235 52720 6355
rect 52840 6235 52885 6355
rect 53005 6235 53050 6355
rect 53170 6235 53225 6355
rect 53345 6235 53355 6355
rect 47855 6190 53355 6235
rect 47855 6070 47865 6190
rect 47985 6070 48030 6190
rect 48150 6070 48195 6190
rect 48315 6070 48360 6190
rect 48480 6070 48535 6190
rect 48655 6070 48700 6190
rect 48820 6070 48865 6190
rect 48985 6070 49030 6190
rect 49150 6070 49205 6190
rect 49325 6070 49370 6190
rect 49490 6070 49535 6190
rect 49655 6070 49700 6190
rect 49820 6070 49875 6190
rect 49995 6070 50040 6190
rect 50160 6070 50205 6190
rect 50325 6070 50370 6190
rect 50490 6070 50545 6190
rect 50665 6070 50710 6190
rect 50830 6070 50875 6190
rect 50995 6070 51040 6190
rect 51160 6070 51215 6190
rect 51335 6070 51380 6190
rect 51500 6070 51545 6190
rect 51665 6070 51710 6190
rect 51830 6070 51885 6190
rect 52005 6070 52050 6190
rect 52170 6070 52215 6190
rect 52335 6070 52380 6190
rect 52500 6070 52555 6190
rect 52675 6070 52720 6190
rect 52840 6070 52885 6190
rect 53005 6070 53050 6190
rect 53170 6070 53225 6190
rect 53345 6070 53355 6190
rect 47855 6025 53355 6070
rect 47855 5905 47865 6025
rect 47985 5905 48030 6025
rect 48150 5905 48195 6025
rect 48315 5905 48360 6025
rect 48480 5905 48535 6025
rect 48655 5905 48700 6025
rect 48820 5905 48865 6025
rect 48985 5905 49030 6025
rect 49150 5905 49205 6025
rect 49325 5905 49370 6025
rect 49490 5905 49535 6025
rect 49655 5905 49700 6025
rect 49820 5905 49875 6025
rect 49995 5905 50040 6025
rect 50160 5905 50205 6025
rect 50325 5905 50370 6025
rect 50490 5905 50545 6025
rect 50665 5905 50710 6025
rect 50830 5905 50875 6025
rect 50995 5905 51040 6025
rect 51160 5905 51215 6025
rect 51335 5905 51380 6025
rect 51500 5905 51545 6025
rect 51665 5905 51710 6025
rect 51830 5905 51885 6025
rect 52005 5905 52050 6025
rect 52170 5905 52215 6025
rect 52335 5905 52380 6025
rect 52500 5905 52555 6025
rect 52675 5905 52720 6025
rect 52840 5905 52885 6025
rect 53005 5905 53050 6025
rect 53170 5905 53225 6025
rect 53345 5905 53355 6025
rect 47855 5860 53355 5905
rect 47855 5740 47865 5860
rect 47985 5740 48030 5860
rect 48150 5740 48195 5860
rect 48315 5740 48360 5860
rect 48480 5740 48535 5860
rect 48655 5740 48700 5860
rect 48820 5740 48865 5860
rect 48985 5740 49030 5860
rect 49150 5740 49205 5860
rect 49325 5740 49370 5860
rect 49490 5740 49535 5860
rect 49655 5740 49700 5860
rect 49820 5740 49875 5860
rect 49995 5740 50040 5860
rect 50160 5740 50205 5860
rect 50325 5740 50370 5860
rect 50490 5740 50545 5860
rect 50665 5740 50710 5860
rect 50830 5740 50875 5860
rect 50995 5740 51040 5860
rect 51160 5740 51215 5860
rect 51335 5740 51380 5860
rect 51500 5740 51545 5860
rect 51665 5740 51710 5860
rect 51830 5740 51885 5860
rect 52005 5740 52050 5860
rect 52170 5740 52215 5860
rect 52335 5740 52380 5860
rect 52500 5740 52555 5860
rect 52675 5740 52720 5860
rect 52840 5740 52885 5860
rect 53005 5740 53050 5860
rect 53170 5740 53225 5860
rect 53345 5740 53355 5860
rect 47855 5685 53355 5740
rect 47855 5565 47865 5685
rect 47985 5565 48030 5685
rect 48150 5565 48195 5685
rect 48315 5565 48360 5685
rect 48480 5565 48535 5685
rect 48655 5565 48700 5685
rect 48820 5565 48865 5685
rect 48985 5565 49030 5685
rect 49150 5565 49205 5685
rect 49325 5565 49370 5685
rect 49490 5565 49535 5685
rect 49655 5565 49700 5685
rect 49820 5565 49875 5685
rect 49995 5565 50040 5685
rect 50160 5565 50205 5685
rect 50325 5565 50370 5685
rect 50490 5565 50545 5685
rect 50665 5565 50710 5685
rect 50830 5565 50875 5685
rect 50995 5565 51040 5685
rect 51160 5565 51215 5685
rect 51335 5565 51380 5685
rect 51500 5565 51545 5685
rect 51665 5565 51710 5685
rect 51830 5565 51885 5685
rect 52005 5565 52050 5685
rect 52170 5565 52215 5685
rect 52335 5565 52380 5685
rect 52500 5565 52555 5685
rect 52675 5565 52720 5685
rect 52840 5565 52885 5685
rect 53005 5565 53050 5685
rect 53170 5565 53225 5685
rect 53345 5565 53355 5685
rect 47855 5520 53355 5565
rect 47855 5400 47865 5520
rect 47985 5400 48030 5520
rect 48150 5400 48195 5520
rect 48315 5400 48360 5520
rect 48480 5400 48535 5520
rect 48655 5400 48700 5520
rect 48820 5400 48865 5520
rect 48985 5400 49030 5520
rect 49150 5400 49205 5520
rect 49325 5400 49370 5520
rect 49490 5400 49535 5520
rect 49655 5400 49700 5520
rect 49820 5400 49875 5520
rect 49995 5400 50040 5520
rect 50160 5400 50205 5520
rect 50325 5400 50370 5520
rect 50490 5400 50545 5520
rect 50665 5400 50710 5520
rect 50830 5400 50875 5520
rect 50995 5400 51040 5520
rect 51160 5400 51215 5520
rect 51335 5400 51380 5520
rect 51500 5400 51545 5520
rect 51665 5400 51710 5520
rect 51830 5400 51885 5520
rect 52005 5400 52050 5520
rect 52170 5400 52215 5520
rect 52335 5400 52380 5520
rect 52500 5400 52555 5520
rect 52675 5400 52720 5520
rect 52840 5400 52885 5520
rect 53005 5400 53050 5520
rect 53170 5400 53225 5520
rect 53345 5400 53355 5520
rect 47855 5355 53355 5400
rect 47855 5235 47865 5355
rect 47985 5235 48030 5355
rect 48150 5235 48195 5355
rect 48315 5235 48360 5355
rect 48480 5235 48535 5355
rect 48655 5235 48700 5355
rect 48820 5235 48865 5355
rect 48985 5235 49030 5355
rect 49150 5235 49205 5355
rect 49325 5235 49370 5355
rect 49490 5235 49535 5355
rect 49655 5235 49700 5355
rect 49820 5235 49875 5355
rect 49995 5235 50040 5355
rect 50160 5235 50205 5355
rect 50325 5235 50370 5355
rect 50490 5235 50545 5355
rect 50665 5235 50710 5355
rect 50830 5235 50875 5355
rect 50995 5235 51040 5355
rect 51160 5235 51215 5355
rect 51335 5235 51380 5355
rect 51500 5235 51545 5355
rect 51665 5235 51710 5355
rect 51830 5235 51885 5355
rect 52005 5235 52050 5355
rect 52170 5235 52215 5355
rect 52335 5235 52380 5355
rect 52500 5235 52555 5355
rect 52675 5235 52720 5355
rect 52840 5235 52885 5355
rect 53005 5235 53050 5355
rect 53170 5235 53225 5355
rect 53345 5235 53355 5355
rect 47855 5190 53355 5235
rect 47855 5070 47865 5190
rect 47985 5070 48030 5190
rect 48150 5070 48195 5190
rect 48315 5070 48360 5190
rect 48480 5070 48535 5190
rect 48655 5070 48700 5190
rect 48820 5070 48865 5190
rect 48985 5070 49030 5190
rect 49150 5070 49205 5190
rect 49325 5070 49370 5190
rect 49490 5070 49535 5190
rect 49655 5070 49700 5190
rect 49820 5070 49875 5190
rect 49995 5070 50040 5190
rect 50160 5070 50205 5190
rect 50325 5070 50370 5190
rect 50490 5070 50545 5190
rect 50665 5070 50710 5190
rect 50830 5070 50875 5190
rect 50995 5070 51040 5190
rect 51160 5070 51215 5190
rect 51335 5070 51380 5190
rect 51500 5070 51545 5190
rect 51665 5070 51710 5190
rect 51830 5070 51885 5190
rect 52005 5070 52050 5190
rect 52170 5070 52215 5190
rect 52335 5070 52380 5190
rect 52500 5070 52555 5190
rect 52675 5070 52720 5190
rect 52840 5070 52885 5190
rect 53005 5070 53050 5190
rect 53170 5070 53225 5190
rect 53345 5070 53355 5190
rect 47855 5015 53355 5070
rect 47855 4895 47865 5015
rect 47985 4895 48030 5015
rect 48150 4895 48195 5015
rect 48315 4895 48360 5015
rect 48480 4895 48535 5015
rect 48655 4895 48700 5015
rect 48820 4895 48865 5015
rect 48985 4895 49030 5015
rect 49150 4895 49205 5015
rect 49325 4895 49370 5015
rect 49490 4895 49535 5015
rect 49655 4895 49700 5015
rect 49820 4895 49875 5015
rect 49995 4895 50040 5015
rect 50160 4895 50205 5015
rect 50325 4895 50370 5015
rect 50490 4895 50545 5015
rect 50665 4895 50710 5015
rect 50830 4895 50875 5015
rect 50995 4895 51040 5015
rect 51160 4895 51215 5015
rect 51335 4895 51380 5015
rect 51500 4895 51545 5015
rect 51665 4895 51710 5015
rect 51830 4895 51885 5015
rect 52005 4895 52050 5015
rect 52170 4895 52215 5015
rect 52335 4895 52380 5015
rect 52500 4895 52555 5015
rect 52675 4895 52720 5015
rect 52840 4895 52885 5015
rect 53005 4895 53050 5015
rect 53170 4895 53225 5015
rect 53345 4895 53355 5015
rect 47855 4850 53355 4895
rect 47855 4730 47865 4850
rect 47985 4730 48030 4850
rect 48150 4730 48195 4850
rect 48315 4730 48360 4850
rect 48480 4730 48535 4850
rect 48655 4730 48700 4850
rect 48820 4730 48865 4850
rect 48985 4730 49030 4850
rect 49150 4730 49205 4850
rect 49325 4730 49370 4850
rect 49490 4730 49535 4850
rect 49655 4730 49700 4850
rect 49820 4730 49875 4850
rect 49995 4730 50040 4850
rect 50160 4730 50205 4850
rect 50325 4730 50370 4850
rect 50490 4730 50545 4850
rect 50665 4730 50710 4850
rect 50830 4730 50875 4850
rect 50995 4730 51040 4850
rect 51160 4730 51215 4850
rect 51335 4730 51380 4850
rect 51500 4730 51545 4850
rect 51665 4730 51710 4850
rect 51830 4730 51885 4850
rect 52005 4730 52050 4850
rect 52170 4730 52215 4850
rect 52335 4730 52380 4850
rect 52500 4730 52555 4850
rect 52675 4730 52720 4850
rect 52840 4730 52885 4850
rect 53005 4730 53050 4850
rect 53170 4730 53225 4850
rect 53345 4730 53355 4850
rect 47855 4685 53355 4730
rect 47855 4565 47865 4685
rect 47985 4565 48030 4685
rect 48150 4565 48195 4685
rect 48315 4565 48360 4685
rect 48480 4565 48535 4685
rect 48655 4565 48700 4685
rect 48820 4565 48865 4685
rect 48985 4565 49030 4685
rect 49150 4565 49205 4685
rect 49325 4565 49370 4685
rect 49490 4565 49535 4685
rect 49655 4565 49700 4685
rect 49820 4565 49875 4685
rect 49995 4565 50040 4685
rect 50160 4565 50205 4685
rect 50325 4565 50370 4685
rect 50490 4565 50545 4685
rect 50665 4565 50710 4685
rect 50830 4565 50875 4685
rect 50995 4565 51040 4685
rect 51160 4565 51215 4685
rect 51335 4565 51380 4685
rect 51500 4565 51545 4685
rect 51665 4565 51710 4685
rect 51830 4565 51885 4685
rect 52005 4565 52050 4685
rect 52170 4565 52215 4685
rect 52335 4565 52380 4685
rect 52500 4565 52555 4685
rect 52675 4565 52720 4685
rect 52840 4565 52885 4685
rect 53005 4565 53050 4685
rect 53170 4565 53225 4685
rect 53345 4565 53355 4685
rect 47855 4520 53355 4565
rect 47855 4400 47865 4520
rect 47985 4400 48030 4520
rect 48150 4400 48195 4520
rect 48315 4400 48360 4520
rect 48480 4400 48535 4520
rect 48655 4400 48700 4520
rect 48820 4400 48865 4520
rect 48985 4400 49030 4520
rect 49150 4400 49205 4520
rect 49325 4400 49370 4520
rect 49490 4400 49535 4520
rect 49655 4400 49700 4520
rect 49820 4400 49875 4520
rect 49995 4400 50040 4520
rect 50160 4400 50205 4520
rect 50325 4400 50370 4520
rect 50490 4400 50545 4520
rect 50665 4400 50710 4520
rect 50830 4400 50875 4520
rect 50995 4400 51040 4520
rect 51160 4400 51215 4520
rect 51335 4400 51380 4520
rect 51500 4400 51545 4520
rect 51665 4400 51710 4520
rect 51830 4400 51885 4520
rect 52005 4400 52050 4520
rect 52170 4400 52215 4520
rect 52335 4400 52380 4520
rect 52500 4400 52555 4520
rect 52675 4400 52720 4520
rect 52840 4400 52885 4520
rect 53005 4400 53050 4520
rect 53170 4400 53225 4520
rect 53345 4400 53355 4520
rect 47855 4345 53355 4400
rect 47855 4225 47865 4345
rect 47985 4225 48030 4345
rect 48150 4225 48195 4345
rect 48315 4225 48360 4345
rect 48480 4225 48535 4345
rect 48655 4225 48700 4345
rect 48820 4225 48865 4345
rect 48985 4225 49030 4345
rect 49150 4225 49205 4345
rect 49325 4225 49370 4345
rect 49490 4225 49535 4345
rect 49655 4225 49700 4345
rect 49820 4225 49875 4345
rect 49995 4225 50040 4345
rect 50160 4225 50205 4345
rect 50325 4225 50370 4345
rect 50490 4225 50545 4345
rect 50665 4225 50710 4345
rect 50830 4225 50875 4345
rect 50995 4225 51040 4345
rect 51160 4225 51215 4345
rect 51335 4225 51380 4345
rect 51500 4225 51545 4345
rect 51665 4225 51710 4345
rect 51830 4225 51885 4345
rect 52005 4225 52050 4345
rect 52170 4225 52215 4345
rect 52335 4225 52380 4345
rect 52500 4225 52555 4345
rect 52675 4225 52720 4345
rect 52840 4225 52885 4345
rect 53005 4225 53050 4345
rect 53170 4225 53225 4345
rect 53345 4225 53355 4345
rect 47855 4180 53355 4225
rect 47855 4060 47865 4180
rect 47985 4060 48030 4180
rect 48150 4060 48195 4180
rect 48315 4060 48360 4180
rect 48480 4060 48535 4180
rect 48655 4060 48700 4180
rect 48820 4060 48865 4180
rect 48985 4060 49030 4180
rect 49150 4060 49205 4180
rect 49325 4060 49370 4180
rect 49490 4060 49535 4180
rect 49655 4060 49700 4180
rect 49820 4060 49875 4180
rect 49995 4060 50040 4180
rect 50160 4060 50205 4180
rect 50325 4060 50370 4180
rect 50490 4060 50545 4180
rect 50665 4060 50710 4180
rect 50830 4060 50875 4180
rect 50995 4060 51040 4180
rect 51160 4060 51215 4180
rect 51335 4060 51380 4180
rect 51500 4060 51545 4180
rect 51665 4060 51710 4180
rect 51830 4060 51885 4180
rect 52005 4060 52050 4180
rect 52170 4060 52215 4180
rect 52335 4060 52380 4180
rect 52500 4060 52555 4180
rect 52675 4060 52720 4180
rect 52840 4060 52885 4180
rect 53005 4060 53050 4180
rect 53170 4060 53225 4180
rect 53345 4060 53355 4180
rect 47855 4015 53355 4060
rect 47855 3895 47865 4015
rect 47985 3895 48030 4015
rect 48150 3895 48195 4015
rect 48315 3895 48360 4015
rect 48480 3895 48535 4015
rect 48655 3895 48700 4015
rect 48820 3895 48865 4015
rect 48985 3895 49030 4015
rect 49150 3895 49205 4015
rect 49325 3895 49370 4015
rect 49490 3895 49535 4015
rect 49655 3895 49700 4015
rect 49820 3895 49875 4015
rect 49995 3895 50040 4015
rect 50160 3895 50205 4015
rect 50325 3895 50370 4015
rect 50490 3895 50545 4015
rect 50665 3895 50710 4015
rect 50830 3895 50875 4015
rect 50995 3895 51040 4015
rect 51160 3895 51215 4015
rect 51335 3895 51380 4015
rect 51500 3895 51545 4015
rect 51665 3895 51710 4015
rect 51830 3895 51885 4015
rect 52005 3895 52050 4015
rect 52170 3895 52215 4015
rect 52335 3895 52380 4015
rect 52500 3895 52555 4015
rect 52675 3895 52720 4015
rect 52840 3895 52885 4015
rect 53005 3895 53050 4015
rect 53170 3895 53225 4015
rect 53345 3895 53355 4015
rect 47855 3850 53355 3895
rect 47855 3730 47865 3850
rect 47985 3730 48030 3850
rect 48150 3730 48195 3850
rect 48315 3730 48360 3850
rect 48480 3730 48535 3850
rect 48655 3730 48700 3850
rect 48820 3730 48865 3850
rect 48985 3730 49030 3850
rect 49150 3730 49205 3850
rect 49325 3730 49370 3850
rect 49490 3730 49535 3850
rect 49655 3730 49700 3850
rect 49820 3730 49875 3850
rect 49995 3730 50040 3850
rect 50160 3730 50205 3850
rect 50325 3730 50370 3850
rect 50490 3730 50545 3850
rect 50665 3730 50710 3850
rect 50830 3730 50875 3850
rect 50995 3730 51040 3850
rect 51160 3730 51215 3850
rect 51335 3730 51380 3850
rect 51500 3730 51545 3850
rect 51665 3730 51710 3850
rect 51830 3730 51885 3850
rect 52005 3730 52050 3850
rect 52170 3730 52215 3850
rect 52335 3730 52380 3850
rect 52500 3730 52555 3850
rect 52675 3730 52720 3850
rect 52840 3730 52885 3850
rect 53005 3730 53050 3850
rect 53170 3730 53225 3850
rect 53345 3730 53355 3850
rect 47855 3675 53355 3730
rect 47855 3555 47865 3675
rect 47985 3555 48030 3675
rect 48150 3555 48195 3675
rect 48315 3555 48360 3675
rect 48480 3555 48535 3675
rect 48655 3555 48700 3675
rect 48820 3555 48865 3675
rect 48985 3555 49030 3675
rect 49150 3555 49205 3675
rect 49325 3555 49370 3675
rect 49490 3555 49535 3675
rect 49655 3555 49700 3675
rect 49820 3555 49875 3675
rect 49995 3555 50040 3675
rect 50160 3555 50205 3675
rect 50325 3555 50370 3675
rect 50490 3555 50545 3675
rect 50665 3555 50710 3675
rect 50830 3555 50875 3675
rect 50995 3555 51040 3675
rect 51160 3555 51215 3675
rect 51335 3555 51380 3675
rect 51500 3555 51545 3675
rect 51665 3555 51710 3675
rect 51830 3555 51885 3675
rect 52005 3555 52050 3675
rect 52170 3555 52215 3675
rect 52335 3555 52380 3675
rect 52500 3555 52555 3675
rect 52675 3555 52720 3675
rect 52840 3555 52885 3675
rect 53005 3555 53050 3675
rect 53170 3555 53225 3675
rect 53345 3555 53355 3675
rect 47855 3510 53355 3555
rect 47855 3390 47865 3510
rect 47985 3390 48030 3510
rect 48150 3390 48195 3510
rect 48315 3390 48360 3510
rect 48480 3390 48535 3510
rect 48655 3390 48700 3510
rect 48820 3390 48865 3510
rect 48985 3390 49030 3510
rect 49150 3390 49205 3510
rect 49325 3390 49370 3510
rect 49490 3390 49535 3510
rect 49655 3390 49700 3510
rect 49820 3390 49875 3510
rect 49995 3390 50040 3510
rect 50160 3390 50205 3510
rect 50325 3390 50370 3510
rect 50490 3390 50545 3510
rect 50665 3390 50710 3510
rect 50830 3390 50875 3510
rect 50995 3390 51040 3510
rect 51160 3390 51215 3510
rect 51335 3390 51380 3510
rect 51500 3390 51545 3510
rect 51665 3390 51710 3510
rect 51830 3390 51885 3510
rect 52005 3390 52050 3510
rect 52170 3390 52215 3510
rect 52335 3390 52380 3510
rect 52500 3390 52555 3510
rect 52675 3390 52720 3510
rect 52840 3390 52885 3510
rect 53005 3390 53050 3510
rect 53170 3390 53225 3510
rect 53345 3390 53355 3510
rect 47855 3345 53355 3390
rect 47855 3225 47865 3345
rect 47985 3225 48030 3345
rect 48150 3225 48195 3345
rect 48315 3225 48360 3345
rect 48480 3225 48535 3345
rect 48655 3225 48700 3345
rect 48820 3225 48865 3345
rect 48985 3225 49030 3345
rect 49150 3225 49205 3345
rect 49325 3225 49370 3345
rect 49490 3225 49535 3345
rect 49655 3225 49700 3345
rect 49820 3225 49875 3345
rect 49995 3225 50040 3345
rect 50160 3225 50205 3345
rect 50325 3225 50370 3345
rect 50490 3225 50545 3345
rect 50665 3225 50710 3345
rect 50830 3225 50875 3345
rect 50995 3225 51040 3345
rect 51160 3225 51215 3345
rect 51335 3225 51380 3345
rect 51500 3225 51545 3345
rect 51665 3225 51710 3345
rect 51830 3225 51885 3345
rect 52005 3225 52050 3345
rect 52170 3225 52215 3345
rect 52335 3225 52380 3345
rect 52500 3225 52555 3345
rect 52675 3225 52720 3345
rect 52840 3225 52885 3345
rect 53005 3225 53050 3345
rect 53170 3225 53225 3345
rect 53345 3225 53355 3345
rect 47855 3180 53355 3225
rect 47855 3060 47865 3180
rect 47985 3060 48030 3180
rect 48150 3060 48195 3180
rect 48315 3060 48360 3180
rect 48480 3060 48535 3180
rect 48655 3060 48700 3180
rect 48820 3060 48865 3180
rect 48985 3060 49030 3180
rect 49150 3060 49205 3180
rect 49325 3060 49370 3180
rect 49490 3060 49535 3180
rect 49655 3060 49700 3180
rect 49820 3060 49875 3180
rect 49995 3060 50040 3180
rect 50160 3060 50205 3180
rect 50325 3060 50370 3180
rect 50490 3060 50545 3180
rect 50665 3060 50710 3180
rect 50830 3060 50875 3180
rect 50995 3060 51040 3180
rect 51160 3060 51215 3180
rect 51335 3060 51380 3180
rect 51500 3060 51545 3180
rect 51665 3060 51710 3180
rect 51830 3060 51885 3180
rect 52005 3060 52050 3180
rect 52170 3060 52215 3180
rect 52335 3060 52380 3180
rect 52500 3060 52555 3180
rect 52675 3060 52720 3180
rect 52840 3060 52885 3180
rect 53005 3060 53050 3180
rect 53170 3060 53225 3180
rect 53345 3060 53355 3180
rect 47855 3005 53355 3060
rect 47855 2885 47865 3005
rect 47985 2885 48030 3005
rect 48150 2885 48195 3005
rect 48315 2885 48360 3005
rect 48480 2885 48535 3005
rect 48655 2885 48700 3005
rect 48820 2885 48865 3005
rect 48985 2885 49030 3005
rect 49150 2885 49205 3005
rect 49325 2885 49370 3005
rect 49490 2885 49535 3005
rect 49655 2885 49700 3005
rect 49820 2885 49875 3005
rect 49995 2885 50040 3005
rect 50160 2885 50205 3005
rect 50325 2885 50370 3005
rect 50490 2885 50545 3005
rect 50665 2885 50710 3005
rect 50830 2885 50875 3005
rect 50995 2885 51040 3005
rect 51160 2885 51215 3005
rect 51335 2885 51380 3005
rect 51500 2885 51545 3005
rect 51665 2885 51710 3005
rect 51830 2885 51885 3005
rect 52005 2885 52050 3005
rect 52170 2885 52215 3005
rect 52335 2885 52380 3005
rect 52500 2885 52555 3005
rect 52675 2885 52720 3005
rect 52840 2885 52885 3005
rect 53005 2885 53050 3005
rect 53170 2885 53225 3005
rect 53345 2885 53355 3005
rect 47855 2840 53355 2885
rect 47855 2720 47865 2840
rect 47985 2720 48030 2840
rect 48150 2720 48195 2840
rect 48315 2720 48360 2840
rect 48480 2720 48535 2840
rect 48655 2720 48700 2840
rect 48820 2720 48865 2840
rect 48985 2720 49030 2840
rect 49150 2720 49205 2840
rect 49325 2720 49370 2840
rect 49490 2720 49535 2840
rect 49655 2720 49700 2840
rect 49820 2720 49875 2840
rect 49995 2720 50040 2840
rect 50160 2720 50205 2840
rect 50325 2720 50370 2840
rect 50490 2720 50545 2840
rect 50665 2720 50710 2840
rect 50830 2720 50875 2840
rect 50995 2720 51040 2840
rect 51160 2720 51215 2840
rect 51335 2720 51380 2840
rect 51500 2720 51545 2840
rect 51665 2720 51710 2840
rect 51830 2720 51885 2840
rect 52005 2720 52050 2840
rect 52170 2720 52215 2840
rect 52335 2720 52380 2840
rect 52500 2720 52555 2840
rect 52675 2720 52720 2840
rect 52840 2720 52885 2840
rect 53005 2720 53050 2840
rect 53170 2720 53225 2840
rect 53345 2720 53355 2840
rect 47855 2675 53355 2720
rect 47855 2555 47865 2675
rect 47985 2555 48030 2675
rect 48150 2555 48195 2675
rect 48315 2555 48360 2675
rect 48480 2555 48535 2675
rect 48655 2555 48700 2675
rect 48820 2555 48865 2675
rect 48985 2555 49030 2675
rect 49150 2555 49205 2675
rect 49325 2555 49370 2675
rect 49490 2555 49535 2675
rect 49655 2555 49700 2675
rect 49820 2555 49875 2675
rect 49995 2555 50040 2675
rect 50160 2555 50205 2675
rect 50325 2555 50370 2675
rect 50490 2555 50545 2675
rect 50665 2555 50710 2675
rect 50830 2555 50875 2675
rect 50995 2555 51040 2675
rect 51160 2555 51215 2675
rect 51335 2555 51380 2675
rect 51500 2555 51545 2675
rect 51665 2555 51710 2675
rect 51830 2555 51885 2675
rect 52005 2555 52050 2675
rect 52170 2555 52215 2675
rect 52335 2555 52380 2675
rect 52500 2555 52555 2675
rect 52675 2555 52720 2675
rect 52840 2555 52885 2675
rect 53005 2555 53050 2675
rect 53170 2555 53225 2675
rect 53345 2555 53355 2675
rect 47855 2510 53355 2555
rect 47855 2390 47865 2510
rect 47985 2390 48030 2510
rect 48150 2390 48195 2510
rect 48315 2390 48360 2510
rect 48480 2390 48535 2510
rect 48655 2390 48700 2510
rect 48820 2390 48865 2510
rect 48985 2390 49030 2510
rect 49150 2390 49205 2510
rect 49325 2390 49370 2510
rect 49490 2390 49535 2510
rect 49655 2390 49700 2510
rect 49820 2390 49875 2510
rect 49995 2390 50040 2510
rect 50160 2390 50205 2510
rect 50325 2390 50370 2510
rect 50490 2390 50545 2510
rect 50665 2390 50710 2510
rect 50830 2390 50875 2510
rect 50995 2390 51040 2510
rect 51160 2390 51215 2510
rect 51335 2390 51380 2510
rect 51500 2390 51545 2510
rect 51665 2390 51710 2510
rect 51830 2390 51885 2510
rect 52005 2390 52050 2510
rect 52170 2390 52215 2510
rect 52335 2390 52380 2510
rect 52500 2390 52555 2510
rect 52675 2390 52720 2510
rect 52840 2390 52885 2510
rect 53005 2390 53050 2510
rect 53170 2390 53225 2510
rect 53345 2390 53355 2510
rect 47855 2335 53355 2390
rect 47855 2215 47865 2335
rect 47985 2215 48030 2335
rect 48150 2215 48195 2335
rect 48315 2215 48360 2335
rect 48480 2215 48535 2335
rect 48655 2215 48700 2335
rect 48820 2215 48865 2335
rect 48985 2215 49030 2335
rect 49150 2215 49205 2335
rect 49325 2215 49370 2335
rect 49490 2215 49535 2335
rect 49655 2215 49700 2335
rect 49820 2215 49875 2335
rect 49995 2215 50040 2335
rect 50160 2215 50205 2335
rect 50325 2215 50370 2335
rect 50490 2215 50545 2335
rect 50665 2215 50710 2335
rect 50830 2215 50875 2335
rect 50995 2215 51040 2335
rect 51160 2215 51215 2335
rect 51335 2215 51380 2335
rect 51500 2215 51545 2335
rect 51665 2215 51710 2335
rect 51830 2215 51885 2335
rect 52005 2215 52050 2335
rect 52170 2215 52215 2335
rect 52335 2215 52380 2335
rect 52500 2215 52555 2335
rect 52675 2215 52720 2335
rect 52840 2215 52885 2335
rect 53005 2215 53050 2335
rect 53170 2215 53225 2335
rect 53345 2215 53355 2335
rect 47855 2170 53355 2215
rect 47855 2050 47865 2170
rect 47985 2050 48030 2170
rect 48150 2050 48195 2170
rect 48315 2050 48360 2170
rect 48480 2050 48535 2170
rect 48655 2050 48700 2170
rect 48820 2050 48865 2170
rect 48985 2050 49030 2170
rect 49150 2050 49205 2170
rect 49325 2050 49370 2170
rect 49490 2050 49535 2170
rect 49655 2050 49700 2170
rect 49820 2050 49875 2170
rect 49995 2050 50040 2170
rect 50160 2050 50205 2170
rect 50325 2050 50370 2170
rect 50490 2050 50545 2170
rect 50665 2050 50710 2170
rect 50830 2050 50875 2170
rect 50995 2050 51040 2170
rect 51160 2050 51215 2170
rect 51335 2050 51380 2170
rect 51500 2050 51545 2170
rect 51665 2050 51710 2170
rect 51830 2050 51885 2170
rect 52005 2050 52050 2170
rect 52170 2050 52215 2170
rect 52335 2050 52380 2170
rect 52500 2050 52555 2170
rect 52675 2050 52720 2170
rect 52840 2050 52885 2170
rect 53005 2050 53050 2170
rect 53170 2050 53225 2170
rect 53345 2050 53355 2170
rect 47855 2005 53355 2050
rect 47855 1885 47865 2005
rect 47985 1885 48030 2005
rect 48150 1885 48195 2005
rect 48315 1885 48360 2005
rect 48480 1885 48535 2005
rect 48655 1885 48700 2005
rect 48820 1885 48865 2005
rect 48985 1885 49030 2005
rect 49150 1885 49205 2005
rect 49325 1885 49370 2005
rect 49490 1885 49535 2005
rect 49655 1885 49700 2005
rect 49820 1885 49875 2005
rect 49995 1885 50040 2005
rect 50160 1885 50205 2005
rect 50325 1885 50370 2005
rect 50490 1885 50545 2005
rect 50665 1885 50710 2005
rect 50830 1885 50875 2005
rect 50995 1885 51040 2005
rect 51160 1885 51215 2005
rect 51335 1885 51380 2005
rect 51500 1885 51545 2005
rect 51665 1885 51710 2005
rect 51830 1885 51885 2005
rect 52005 1885 52050 2005
rect 52170 1885 52215 2005
rect 52335 1885 52380 2005
rect 52500 1885 52555 2005
rect 52675 1885 52720 2005
rect 52840 1885 52885 2005
rect 53005 1885 53050 2005
rect 53170 1885 53225 2005
rect 53345 1885 53355 2005
rect 47855 1840 53355 1885
rect 47855 1720 47865 1840
rect 47985 1720 48030 1840
rect 48150 1720 48195 1840
rect 48315 1720 48360 1840
rect 48480 1720 48535 1840
rect 48655 1720 48700 1840
rect 48820 1720 48865 1840
rect 48985 1720 49030 1840
rect 49150 1720 49205 1840
rect 49325 1720 49370 1840
rect 49490 1720 49535 1840
rect 49655 1720 49700 1840
rect 49820 1720 49875 1840
rect 49995 1720 50040 1840
rect 50160 1720 50205 1840
rect 50325 1720 50370 1840
rect 50490 1720 50545 1840
rect 50665 1720 50710 1840
rect 50830 1720 50875 1840
rect 50995 1720 51040 1840
rect 51160 1720 51215 1840
rect 51335 1720 51380 1840
rect 51500 1720 51545 1840
rect 51665 1720 51710 1840
rect 51830 1720 51885 1840
rect 52005 1720 52050 1840
rect 52170 1720 52215 1840
rect 52335 1720 52380 1840
rect 52500 1720 52555 1840
rect 52675 1720 52720 1840
rect 52840 1720 52885 1840
rect 53005 1720 53050 1840
rect 53170 1720 53225 1840
rect 53345 1720 53355 1840
rect 47855 1710 53355 1720
rect 30785 1420 36285 1430
rect 30785 1300 30795 1420
rect 30915 1300 30970 1420
rect 31090 1300 31135 1420
rect 31255 1300 31300 1420
rect 31420 1300 31465 1420
rect 31585 1300 31640 1420
rect 31760 1300 31805 1420
rect 31925 1300 31970 1420
rect 32090 1300 32135 1420
rect 32255 1300 32310 1420
rect 32430 1300 32475 1420
rect 32595 1300 32640 1420
rect 32760 1300 32805 1420
rect 32925 1300 32980 1420
rect 33100 1300 33145 1420
rect 33265 1300 33310 1420
rect 33430 1300 33475 1420
rect 33595 1300 33650 1420
rect 33770 1300 33815 1420
rect 33935 1300 33980 1420
rect 34100 1300 34145 1420
rect 34265 1300 34320 1420
rect 34440 1300 34485 1420
rect 34605 1300 34650 1420
rect 34770 1300 34815 1420
rect 34935 1300 34990 1420
rect 35110 1300 35155 1420
rect 35275 1300 35320 1420
rect 35440 1300 35485 1420
rect 35605 1300 35660 1420
rect 35780 1300 35825 1420
rect 35945 1300 35990 1420
rect 36110 1300 36155 1420
rect 36275 1300 36285 1420
rect 30785 1255 36285 1300
rect 30785 1135 30795 1255
rect 30915 1135 30970 1255
rect 31090 1135 31135 1255
rect 31255 1135 31300 1255
rect 31420 1135 31465 1255
rect 31585 1135 31640 1255
rect 31760 1135 31805 1255
rect 31925 1135 31970 1255
rect 32090 1135 32135 1255
rect 32255 1135 32310 1255
rect 32430 1135 32475 1255
rect 32595 1135 32640 1255
rect 32760 1135 32805 1255
rect 32925 1135 32980 1255
rect 33100 1135 33145 1255
rect 33265 1135 33310 1255
rect 33430 1135 33475 1255
rect 33595 1135 33650 1255
rect 33770 1135 33815 1255
rect 33935 1135 33980 1255
rect 34100 1135 34145 1255
rect 34265 1135 34320 1255
rect 34440 1135 34485 1255
rect 34605 1135 34650 1255
rect 34770 1135 34815 1255
rect 34935 1135 34990 1255
rect 35110 1135 35155 1255
rect 35275 1135 35320 1255
rect 35440 1135 35485 1255
rect 35605 1135 35660 1255
rect 35780 1135 35825 1255
rect 35945 1135 35990 1255
rect 36110 1135 36155 1255
rect 36275 1135 36285 1255
rect 30785 1090 36285 1135
rect 30785 970 30795 1090
rect 30915 970 30970 1090
rect 31090 970 31135 1090
rect 31255 970 31300 1090
rect 31420 970 31465 1090
rect 31585 970 31640 1090
rect 31760 970 31805 1090
rect 31925 970 31970 1090
rect 32090 970 32135 1090
rect 32255 970 32310 1090
rect 32430 970 32475 1090
rect 32595 970 32640 1090
rect 32760 970 32805 1090
rect 32925 970 32980 1090
rect 33100 970 33145 1090
rect 33265 970 33310 1090
rect 33430 970 33475 1090
rect 33595 970 33650 1090
rect 33770 970 33815 1090
rect 33935 970 33980 1090
rect 34100 970 34145 1090
rect 34265 970 34320 1090
rect 34440 970 34485 1090
rect 34605 970 34650 1090
rect 34770 970 34815 1090
rect 34935 970 34990 1090
rect 35110 970 35155 1090
rect 35275 970 35320 1090
rect 35440 970 35485 1090
rect 35605 970 35660 1090
rect 35780 970 35825 1090
rect 35945 970 35990 1090
rect 36110 970 36155 1090
rect 36275 970 36285 1090
rect 30785 925 36285 970
rect 30785 805 30795 925
rect 30915 805 30970 925
rect 31090 805 31135 925
rect 31255 805 31300 925
rect 31420 805 31465 925
rect 31585 805 31640 925
rect 31760 805 31805 925
rect 31925 805 31970 925
rect 32090 805 32135 925
rect 32255 805 32310 925
rect 32430 805 32475 925
rect 32595 805 32640 925
rect 32760 805 32805 925
rect 32925 805 32980 925
rect 33100 805 33145 925
rect 33265 805 33310 925
rect 33430 805 33475 925
rect 33595 805 33650 925
rect 33770 805 33815 925
rect 33935 805 33980 925
rect 34100 805 34145 925
rect 34265 805 34320 925
rect 34440 805 34485 925
rect 34605 805 34650 925
rect 34770 805 34815 925
rect 34935 805 34990 925
rect 35110 805 35155 925
rect 35275 805 35320 925
rect 35440 805 35485 925
rect 35605 805 35660 925
rect 35780 805 35825 925
rect 35945 805 35990 925
rect 36110 805 36155 925
rect 36275 805 36285 925
rect 30785 750 36285 805
rect 30785 630 30795 750
rect 30915 630 30970 750
rect 31090 630 31135 750
rect 31255 630 31300 750
rect 31420 630 31465 750
rect 31585 630 31640 750
rect 31760 630 31805 750
rect 31925 630 31970 750
rect 32090 630 32135 750
rect 32255 630 32310 750
rect 32430 630 32475 750
rect 32595 630 32640 750
rect 32760 630 32805 750
rect 32925 630 32980 750
rect 33100 630 33145 750
rect 33265 630 33310 750
rect 33430 630 33475 750
rect 33595 630 33650 750
rect 33770 630 33815 750
rect 33935 630 33980 750
rect 34100 630 34145 750
rect 34265 630 34320 750
rect 34440 630 34485 750
rect 34605 630 34650 750
rect 34770 630 34815 750
rect 34935 630 34990 750
rect 35110 630 35155 750
rect 35275 630 35320 750
rect 35440 630 35485 750
rect 35605 630 35660 750
rect 35780 630 35825 750
rect 35945 630 35990 750
rect 36110 630 36155 750
rect 36275 630 36285 750
rect 30785 585 36285 630
rect 30785 465 30795 585
rect 30915 465 30970 585
rect 31090 465 31135 585
rect 31255 465 31300 585
rect 31420 465 31465 585
rect 31585 465 31640 585
rect 31760 465 31805 585
rect 31925 465 31970 585
rect 32090 465 32135 585
rect 32255 465 32310 585
rect 32430 465 32475 585
rect 32595 465 32640 585
rect 32760 465 32805 585
rect 32925 465 32980 585
rect 33100 465 33145 585
rect 33265 465 33310 585
rect 33430 465 33475 585
rect 33595 465 33650 585
rect 33770 465 33815 585
rect 33935 465 33980 585
rect 34100 465 34145 585
rect 34265 465 34320 585
rect 34440 465 34485 585
rect 34605 465 34650 585
rect 34770 465 34815 585
rect 34935 465 34990 585
rect 35110 465 35155 585
rect 35275 465 35320 585
rect 35440 465 35485 585
rect 35605 465 35660 585
rect 35780 465 35825 585
rect 35945 465 35990 585
rect 36110 465 36155 585
rect 36275 465 36285 585
rect 30785 420 36285 465
rect 30785 300 30795 420
rect 30915 300 30970 420
rect 31090 300 31135 420
rect 31255 300 31300 420
rect 31420 300 31465 420
rect 31585 300 31640 420
rect 31760 300 31805 420
rect 31925 300 31970 420
rect 32090 300 32135 420
rect 32255 300 32310 420
rect 32430 300 32475 420
rect 32595 300 32640 420
rect 32760 300 32805 420
rect 32925 300 32980 420
rect 33100 300 33145 420
rect 33265 300 33310 420
rect 33430 300 33475 420
rect 33595 300 33650 420
rect 33770 300 33815 420
rect 33935 300 33980 420
rect 34100 300 34145 420
rect 34265 300 34320 420
rect 34440 300 34485 420
rect 34605 300 34650 420
rect 34770 300 34815 420
rect 34935 300 34990 420
rect 35110 300 35155 420
rect 35275 300 35320 420
rect 35440 300 35485 420
rect 35605 300 35660 420
rect 35780 300 35825 420
rect 35945 300 35990 420
rect 36110 300 36155 420
rect 36275 300 36285 420
rect 30785 255 36285 300
rect 30785 135 30795 255
rect 30915 135 30970 255
rect 31090 135 31135 255
rect 31255 135 31300 255
rect 31420 135 31465 255
rect 31585 135 31640 255
rect 31760 135 31805 255
rect 31925 135 31970 255
rect 32090 135 32135 255
rect 32255 135 32310 255
rect 32430 135 32475 255
rect 32595 135 32640 255
rect 32760 135 32805 255
rect 32925 135 32980 255
rect 33100 135 33145 255
rect 33265 135 33310 255
rect 33430 135 33475 255
rect 33595 135 33650 255
rect 33770 135 33815 255
rect 33935 135 33980 255
rect 34100 135 34145 255
rect 34265 135 34320 255
rect 34440 135 34485 255
rect 34605 135 34650 255
rect 34770 135 34815 255
rect 34935 135 34990 255
rect 35110 135 35155 255
rect 35275 135 35320 255
rect 35440 135 35485 255
rect 35605 135 35660 255
rect 35780 135 35825 255
rect 35945 135 35990 255
rect 36110 135 36155 255
rect 36275 135 36285 255
rect 30785 80 36285 135
rect 30785 -40 30795 80
rect 30915 -40 30970 80
rect 31090 -40 31135 80
rect 31255 -40 31300 80
rect 31420 -40 31465 80
rect 31585 -40 31640 80
rect 31760 -40 31805 80
rect 31925 -40 31970 80
rect 32090 -40 32135 80
rect 32255 -40 32310 80
rect 32430 -40 32475 80
rect 32595 -40 32640 80
rect 32760 -40 32805 80
rect 32925 -40 32980 80
rect 33100 -40 33145 80
rect 33265 -40 33310 80
rect 33430 -40 33475 80
rect 33595 -40 33650 80
rect 33770 -40 33815 80
rect 33935 -40 33980 80
rect 34100 -40 34145 80
rect 34265 -40 34320 80
rect 34440 -40 34485 80
rect 34605 -40 34650 80
rect 34770 -40 34815 80
rect 34935 -40 34990 80
rect 35110 -40 35155 80
rect 35275 -40 35320 80
rect 35440 -40 35485 80
rect 35605 -40 35660 80
rect 35780 -40 35825 80
rect 35945 -40 35990 80
rect 36110 -40 36155 80
rect 36275 -40 36285 80
rect 30785 -85 36285 -40
rect 30785 -205 30795 -85
rect 30915 -205 30970 -85
rect 31090 -205 31135 -85
rect 31255 -205 31300 -85
rect 31420 -205 31465 -85
rect 31585 -205 31640 -85
rect 31760 -205 31805 -85
rect 31925 -205 31970 -85
rect 32090 -205 32135 -85
rect 32255 -205 32310 -85
rect 32430 -205 32475 -85
rect 32595 -205 32640 -85
rect 32760 -205 32805 -85
rect 32925 -205 32980 -85
rect 33100 -205 33145 -85
rect 33265 -205 33310 -85
rect 33430 -205 33475 -85
rect 33595 -205 33650 -85
rect 33770 -205 33815 -85
rect 33935 -205 33980 -85
rect 34100 -205 34145 -85
rect 34265 -205 34320 -85
rect 34440 -205 34485 -85
rect 34605 -205 34650 -85
rect 34770 -205 34815 -85
rect 34935 -205 34990 -85
rect 35110 -205 35155 -85
rect 35275 -205 35320 -85
rect 35440 -205 35485 -85
rect 35605 -205 35660 -85
rect 35780 -205 35825 -85
rect 35945 -205 35990 -85
rect 36110 -205 36155 -85
rect 36275 -205 36285 -85
rect 30785 -250 36285 -205
rect 30785 -370 30795 -250
rect 30915 -370 30970 -250
rect 31090 -370 31135 -250
rect 31255 -370 31300 -250
rect 31420 -370 31465 -250
rect 31585 -370 31640 -250
rect 31760 -370 31805 -250
rect 31925 -370 31970 -250
rect 32090 -370 32135 -250
rect 32255 -370 32310 -250
rect 32430 -370 32475 -250
rect 32595 -370 32640 -250
rect 32760 -370 32805 -250
rect 32925 -370 32980 -250
rect 33100 -370 33145 -250
rect 33265 -370 33310 -250
rect 33430 -370 33475 -250
rect 33595 -370 33650 -250
rect 33770 -370 33815 -250
rect 33935 -370 33980 -250
rect 34100 -370 34145 -250
rect 34265 -370 34320 -250
rect 34440 -370 34485 -250
rect 34605 -370 34650 -250
rect 34770 -370 34815 -250
rect 34935 -370 34990 -250
rect 35110 -370 35155 -250
rect 35275 -370 35320 -250
rect 35440 -370 35485 -250
rect 35605 -370 35660 -250
rect 35780 -370 35825 -250
rect 35945 -370 35990 -250
rect 36110 -370 36155 -250
rect 36275 -370 36285 -250
rect 30785 -415 36285 -370
rect 30785 -535 30795 -415
rect 30915 -535 30970 -415
rect 31090 -535 31135 -415
rect 31255 -535 31300 -415
rect 31420 -535 31465 -415
rect 31585 -535 31640 -415
rect 31760 -535 31805 -415
rect 31925 -535 31970 -415
rect 32090 -535 32135 -415
rect 32255 -535 32310 -415
rect 32430 -535 32475 -415
rect 32595 -535 32640 -415
rect 32760 -535 32805 -415
rect 32925 -535 32980 -415
rect 33100 -535 33145 -415
rect 33265 -535 33310 -415
rect 33430 -535 33475 -415
rect 33595 -535 33650 -415
rect 33770 -535 33815 -415
rect 33935 -535 33980 -415
rect 34100 -535 34145 -415
rect 34265 -535 34320 -415
rect 34440 -535 34485 -415
rect 34605 -535 34650 -415
rect 34770 -535 34815 -415
rect 34935 -535 34990 -415
rect 35110 -535 35155 -415
rect 35275 -535 35320 -415
rect 35440 -535 35485 -415
rect 35605 -535 35660 -415
rect 35780 -535 35825 -415
rect 35945 -535 35990 -415
rect 36110 -535 36155 -415
rect 36275 -535 36285 -415
rect 30785 -590 36285 -535
rect 30785 -710 30795 -590
rect 30915 -710 30970 -590
rect 31090 -710 31135 -590
rect 31255 -710 31300 -590
rect 31420 -710 31465 -590
rect 31585 -710 31640 -590
rect 31760 -710 31805 -590
rect 31925 -710 31970 -590
rect 32090 -710 32135 -590
rect 32255 -710 32310 -590
rect 32430 -710 32475 -590
rect 32595 -710 32640 -590
rect 32760 -710 32805 -590
rect 32925 -710 32980 -590
rect 33100 -710 33145 -590
rect 33265 -710 33310 -590
rect 33430 -710 33475 -590
rect 33595 -710 33650 -590
rect 33770 -710 33815 -590
rect 33935 -710 33980 -590
rect 34100 -710 34145 -590
rect 34265 -710 34320 -590
rect 34440 -710 34485 -590
rect 34605 -710 34650 -590
rect 34770 -710 34815 -590
rect 34935 -710 34990 -590
rect 35110 -710 35155 -590
rect 35275 -710 35320 -590
rect 35440 -710 35485 -590
rect 35605 -710 35660 -590
rect 35780 -710 35825 -590
rect 35945 -710 35990 -590
rect 36110 -710 36155 -590
rect 36275 -710 36285 -590
rect 30785 -755 36285 -710
rect 30785 -875 30795 -755
rect 30915 -875 30970 -755
rect 31090 -875 31135 -755
rect 31255 -875 31300 -755
rect 31420 -875 31465 -755
rect 31585 -875 31640 -755
rect 31760 -875 31805 -755
rect 31925 -875 31970 -755
rect 32090 -875 32135 -755
rect 32255 -875 32310 -755
rect 32430 -875 32475 -755
rect 32595 -875 32640 -755
rect 32760 -875 32805 -755
rect 32925 -875 32980 -755
rect 33100 -875 33145 -755
rect 33265 -875 33310 -755
rect 33430 -875 33475 -755
rect 33595 -875 33650 -755
rect 33770 -875 33815 -755
rect 33935 -875 33980 -755
rect 34100 -875 34145 -755
rect 34265 -875 34320 -755
rect 34440 -875 34485 -755
rect 34605 -875 34650 -755
rect 34770 -875 34815 -755
rect 34935 -875 34990 -755
rect 35110 -875 35155 -755
rect 35275 -875 35320 -755
rect 35440 -875 35485 -755
rect 35605 -875 35660 -755
rect 35780 -875 35825 -755
rect 35945 -875 35990 -755
rect 36110 -875 36155 -755
rect 36275 -875 36285 -755
rect 30785 -920 36285 -875
rect 30785 -1040 30795 -920
rect 30915 -1040 30970 -920
rect 31090 -1040 31135 -920
rect 31255 -1040 31300 -920
rect 31420 -1040 31465 -920
rect 31585 -1040 31640 -920
rect 31760 -1040 31805 -920
rect 31925 -1040 31970 -920
rect 32090 -1040 32135 -920
rect 32255 -1040 32310 -920
rect 32430 -1040 32475 -920
rect 32595 -1040 32640 -920
rect 32760 -1040 32805 -920
rect 32925 -1040 32980 -920
rect 33100 -1040 33145 -920
rect 33265 -1040 33310 -920
rect 33430 -1040 33475 -920
rect 33595 -1040 33650 -920
rect 33770 -1040 33815 -920
rect 33935 -1040 33980 -920
rect 34100 -1040 34145 -920
rect 34265 -1040 34320 -920
rect 34440 -1040 34485 -920
rect 34605 -1040 34650 -920
rect 34770 -1040 34815 -920
rect 34935 -1040 34990 -920
rect 35110 -1040 35155 -920
rect 35275 -1040 35320 -920
rect 35440 -1040 35485 -920
rect 35605 -1040 35660 -920
rect 35780 -1040 35825 -920
rect 35945 -1040 35990 -920
rect 36110 -1040 36155 -920
rect 36275 -1040 36285 -920
rect 30785 -1085 36285 -1040
rect 30785 -1205 30795 -1085
rect 30915 -1205 30970 -1085
rect 31090 -1205 31135 -1085
rect 31255 -1205 31300 -1085
rect 31420 -1205 31465 -1085
rect 31585 -1205 31640 -1085
rect 31760 -1205 31805 -1085
rect 31925 -1205 31970 -1085
rect 32090 -1205 32135 -1085
rect 32255 -1205 32310 -1085
rect 32430 -1205 32475 -1085
rect 32595 -1205 32640 -1085
rect 32760 -1205 32805 -1085
rect 32925 -1205 32980 -1085
rect 33100 -1205 33145 -1085
rect 33265 -1205 33310 -1085
rect 33430 -1205 33475 -1085
rect 33595 -1205 33650 -1085
rect 33770 -1205 33815 -1085
rect 33935 -1205 33980 -1085
rect 34100 -1205 34145 -1085
rect 34265 -1205 34320 -1085
rect 34440 -1205 34485 -1085
rect 34605 -1205 34650 -1085
rect 34770 -1205 34815 -1085
rect 34935 -1205 34990 -1085
rect 35110 -1205 35155 -1085
rect 35275 -1205 35320 -1085
rect 35440 -1205 35485 -1085
rect 35605 -1205 35660 -1085
rect 35780 -1205 35825 -1085
rect 35945 -1205 35990 -1085
rect 36110 -1205 36155 -1085
rect 36275 -1205 36285 -1085
rect 30785 -1260 36285 -1205
rect 30785 -1380 30795 -1260
rect 30915 -1380 30970 -1260
rect 31090 -1380 31135 -1260
rect 31255 -1380 31300 -1260
rect 31420 -1380 31465 -1260
rect 31585 -1380 31640 -1260
rect 31760 -1380 31805 -1260
rect 31925 -1380 31970 -1260
rect 32090 -1380 32135 -1260
rect 32255 -1380 32310 -1260
rect 32430 -1380 32475 -1260
rect 32595 -1380 32640 -1260
rect 32760 -1380 32805 -1260
rect 32925 -1380 32980 -1260
rect 33100 -1380 33145 -1260
rect 33265 -1380 33310 -1260
rect 33430 -1380 33475 -1260
rect 33595 -1380 33650 -1260
rect 33770 -1380 33815 -1260
rect 33935 -1380 33980 -1260
rect 34100 -1380 34145 -1260
rect 34265 -1380 34320 -1260
rect 34440 -1380 34485 -1260
rect 34605 -1380 34650 -1260
rect 34770 -1380 34815 -1260
rect 34935 -1380 34990 -1260
rect 35110 -1380 35155 -1260
rect 35275 -1380 35320 -1260
rect 35440 -1380 35485 -1260
rect 35605 -1380 35660 -1260
rect 35780 -1380 35825 -1260
rect 35945 -1380 35990 -1260
rect 36110 -1380 36155 -1260
rect 36275 -1380 36285 -1260
rect 30785 -1425 36285 -1380
rect 30785 -1545 30795 -1425
rect 30915 -1545 30970 -1425
rect 31090 -1545 31135 -1425
rect 31255 -1545 31300 -1425
rect 31420 -1545 31465 -1425
rect 31585 -1545 31640 -1425
rect 31760 -1545 31805 -1425
rect 31925 -1545 31970 -1425
rect 32090 -1545 32135 -1425
rect 32255 -1545 32310 -1425
rect 32430 -1545 32475 -1425
rect 32595 -1545 32640 -1425
rect 32760 -1545 32805 -1425
rect 32925 -1545 32980 -1425
rect 33100 -1545 33145 -1425
rect 33265 -1545 33310 -1425
rect 33430 -1545 33475 -1425
rect 33595 -1545 33650 -1425
rect 33770 -1545 33815 -1425
rect 33935 -1545 33980 -1425
rect 34100 -1545 34145 -1425
rect 34265 -1545 34320 -1425
rect 34440 -1545 34485 -1425
rect 34605 -1545 34650 -1425
rect 34770 -1545 34815 -1425
rect 34935 -1545 34990 -1425
rect 35110 -1545 35155 -1425
rect 35275 -1545 35320 -1425
rect 35440 -1545 35485 -1425
rect 35605 -1545 35660 -1425
rect 35780 -1545 35825 -1425
rect 35945 -1545 35990 -1425
rect 36110 -1545 36155 -1425
rect 36275 -1545 36285 -1425
rect 30785 -1590 36285 -1545
rect 30785 -1710 30795 -1590
rect 30915 -1710 30970 -1590
rect 31090 -1710 31135 -1590
rect 31255 -1710 31300 -1590
rect 31420 -1710 31465 -1590
rect 31585 -1710 31640 -1590
rect 31760 -1710 31805 -1590
rect 31925 -1710 31970 -1590
rect 32090 -1710 32135 -1590
rect 32255 -1710 32310 -1590
rect 32430 -1710 32475 -1590
rect 32595 -1710 32640 -1590
rect 32760 -1710 32805 -1590
rect 32925 -1710 32980 -1590
rect 33100 -1710 33145 -1590
rect 33265 -1710 33310 -1590
rect 33430 -1710 33475 -1590
rect 33595 -1710 33650 -1590
rect 33770 -1710 33815 -1590
rect 33935 -1710 33980 -1590
rect 34100 -1710 34145 -1590
rect 34265 -1710 34320 -1590
rect 34440 -1710 34485 -1590
rect 34605 -1710 34650 -1590
rect 34770 -1710 34815 -1590
rect 34935 -1710 34990 -1590
rect 35110 -1710 35155 -1590
rect 35275 -1710 35320 -1590
rect 35440 -1710 35485 -1590
rect 35605 -1710 35660 -1590
rect 35780 -1710 35825 -1590
rect 35945 -1710 35990 -1590
rect 36110 -1710 36155 -1590
rect 36275 -1710 36285 -1590
rect 30785 -1755 36285 -1710
rect 30785 -1875 30795 -1755
rect 30915 -1875 30970 -1755
rect 31090 -1875 31135 -1755
rect 31255 -1875 31300 -1755
rect 31420 -1875 31465 -1755
rect 31585 -1875 31640 -1755
rect 31760 -1875 31805 -1755
rect 31925 -1875 31970 -1755
rect 32090 -1875 32135 -1755
rect 32255 -1875 32310 -1755
rect 32430 -1875 32475 -1755
rect 32595 -1875 32640 -1755
rect 32760 -1875 32805 -1755
rect 32925 -1875 32980 -1755
rect 33100 -1875 33145 -1755
rect 33265 -1875 33310 -1755
rect 33430 -1875 33475 -1755
rect 33595 -1875 33650 -1755
rect 33770 -1875 33815 -1755
rect 33935 -1875 33980 -1755
rect 34100 -1875 34145 -1755
rect 34265 -1875 34320 -1755
rect 34440 -1875 34485 -1755
rect 34605 -1875 34650 -1755
rect 34770 -1875 34815 -1755
rect 34935 -1875 34990 -1755
rect 35110 -1875 35155 -1755
rect 35275 -1875 35320 -1755
rect 35440 -1875 35485 -1755
rect 35605 -1875 35660 -1755
rect 35780 -1875 35825 -1755
rect 35945 -1875 35990 -1755
rect 36110 -1875 36155 -1755
rect 36275 -1875 36285 -1755
rect 30785 -1930 36285 -1875
rect 30785 -2050 30795 -1930
rect 30915 -2050 30970 -1930
rect 31090 -2050 31135 -1930
rect 31255 -2050 31300 -1930
rect 31420 -2050 31465 -1930
rect 31585 -2050 31640 -1930
rect 31760 -2050 31805 -1930
rect 31925 -2050 31970 -1930
rect 32090 -2050 32135 -1930
rect 32255 -2050 32310 -1930
rect 32430 -2050 32475 -1930
rect 32595 -2050 32640 -1930
rect 32760 -2050 32805 -1930
rect 32925 -2050 32980 -1930
rect 33100 -2050 33145 -1930
rect 33265 -2050 33310 -1930
rect 33430 -2050 33475 -1930
rect 33595 -2050 33650 -1930
rect 33770 -2050 33815 -1930
rect 33935 -2050 33980 -1930
rect 34100 -2050 34145 -1930
rect 34265 -2050 34320 -1930
rect 34440 -2050 34485 -1930
rect 34605 -2050 34650 -1930
rect 34770 -2050 34815 -1930
rect 34935 -2050 34990 -1930
rect 35110 -2050 35155 -1930
rect 35275 -2050 35320 -1930
rect 35440 -2050 35485 -1930
rect 35605 -2050 35660 -1930
rect 35780 -2050 35825 -1930
rect 35945 -2050 35990 -1930
rect 36110 -2050 36155 -1930
rect 36275 -2050 36285 -1930
rect 30785 -2095 36285 -2050
rect 30785 -2215 30795 -2095
rect 30915 -2215 30970 -2095
rect 31090 -2215 31135 -2095
rect 31255 -2215 31300 -2095
rect 31420 -2215 31465 -2095
rect 31585 -2215 31640 -2095
rect 31760 -2215 31805 -2095
rect 31925 -2215 31970 -2095
rect 32090 -2215 32135 -2095
rect 32255 -2215 32310 -2095
rect 32430 -2215 32475 -2095
rect 32595 -2215 32640 -2095
rect 32760 -2215 32805 -2095
rect 32925 -2215 32980 -2095
rect 33100 -2215 33145 -2095
rect 33265 -2215 33310 -2095
rect 33430 -2215 33475 -2095
rect 33595 -2215 33650 -2095
rect 33770 -2215 33815 -2095
rect 33935 -2215 33980 -2095
rect 34100 -2215 34145 -2095
rect 34265 -2215 34320 -2095
rect 34440 -2215 34485 -2095
rect 34605 -2215 34650 -2095
rect 34770 -2215 34815 -2095
rect 34935 -2215 34990 -2095
rect 35110 -2215 35155 -2095
rect 35275 -2215 35320 -2095
rect 35440 -2215 35485 -2095
rect 35605 -2215 35660 -2095
rect 35780 -2215 35825 -2095
rect 35945 -2215 35990 -2095
rect 36110 -2215 36155 -2095
rect 36275 -2215 36285 -2095
rect 30785 -2260 36285 -2215
rect 30785 -2380 30795 -2260
rect 30915 -2380 30970 -2260
rect 31090 -2380 31135 -2260
rect 31255 -2380 31300 -2260
rect 31420 -2380 31465 -2260
rect 31585 -2380 31640 -2260
rect 31760 -2380 31805 -2260
rect 31925 -2380 31970 -2260
rect 32090 -2380 32135 -2260
rect 32255 -2380 32310 -2260
rect 32430 -2380 32475 -2260
rect 32595 -2380 32640 -2260
rect 32760 -2380 32805 -2260
rect 32925 -2380 32980 -2260
rect 33100 -2380 33145 -2260
rect 33265 -2380 33310 -2260
rect 33430 -2380 33475 -2260
rect 33595 -2380 33650 -2260
rect 33770 -2380 33815 -2260
rect 33935 -2380 33980 -2260
rect 34100 -2380 34145 -2260
rect 34265 -2380 34320 -2260
rect 34440 -2380 34485 -2260
rect 34605 -2380 34650 -2260
rect 34770 -2380 34815 -2260
rect 34935 -2380 34990 -2260
rect 35110 -2380 35155 -2260
rect 35275 -2380 35320 -2260
rect 35440 -2380 35485 -2260
rect 35605 -2380 35660 -2260
rect 35780 -2380 35825 -2260
rect 35945 -2380 35990 -2260
rect 36110 -2380 36155 -2260
rect 36275 -2380 36285 -2260
rect 30785 -2425 36285 -2380
rect 30785 -2545 30795 -2425
rect 30915 -2545 30970 -2425
rect 31090 -2545 31135 -2425
rect 31255 -2545 31300 -2425
rect 31420 -2545 31465 -2425
rect 31585 -2545 31640 -2425
rect 31760 -2545 31805 -2425
rect 31925 -2545 31970 -2425
rect 32090 -2545 32135 -2425
rect 32255 -2545 32310 -2425
rect 32430 -2545 32475 -2425
rect 32595 -2545 32640 -2425
rect 32760 -2545 32805 -2425
rect 32925 -2545 32980 -2425
rect 33100 -2545 33145 -2425
rect 33265 -2545 33310 -2425
rect 33430 -2545 33475 -2425
rect 33595 -2545 33650 -2425
rect 33770 -2545 33815 -2425
rect 33935 -2545 33980 -2425
rect 34100 -2545 34145 -2425
rect 34265 -2545 34320 -2425
rect 34440 -2545 34485 -2425
rect 34605 -2545 34650 -2425
rect 34770 -2545 34815 -2425
rect 34935 -2545 34990 -2425
rect 35110 -2545 35155 -2425
rect 35275 -2545 35320 -2425
rect 35440 -2545 35485 -2425
rect 35605 -2545 35660 -2425
rect 35780 -2545 35825 -2425
rect 35945 -2545 35990 -2425
rect 36110 -2545 36155 -2425
rect 36275 -2545 36285 -2425
rect 30785 -2600 36285 -2545
rect 30785 -2720 30795 -2600
rect 30915 -2720 30970 -2600
rect 31090 -2720 31135 -2600
rect 31255 -2720 31300 -2600
rect 31420 -2720 31465 -2600
rect 31585 -2720 31640 -2600
rect 31760 -2720 31805 -2600
rect 31925 -2720 31970 -2600
rect 32090 -2720 32135 -2600
rect 32255 -2720 32310 -2600
rect 32430 -2720 32475 -2600
rect 32595 -2720 32640 -2600
rect 32760 -2720 32805 -2600
rect 32925 -2720 32980 -2600
rect 33100 -2720 33145 -2600
rect 33265 -2720 33310 -2600
rect 33430 -2720 33475 -2600
rect 33595 -2720 33650 -2600
rect 33770 -2720 33815 -2600
rect 33935 -2720 33980 -2600
rect 34100 -2720 34145 -2600
rect 34265 -2720 34320 -2600
rect 34440 -2720 34485 -2600
rect 34605 -2720 34650 -2600
rect 34770 -2720 34815 -2600
rect 34935 -2720 34990 -2600
rect 35110 -2720 35155 -2600
rect 35275 -2720 35320 -2600
rect 35440 -2720 35485 -2600
rect 35605 -2720 35660 -2600
rect 35780 -2720 35825 -2600
rect 35945 -2720 35990 -2600
rect 36110 -2720 36155 -2600
rect 36275 -2720 36285 -2600
rect 30785 -2765 36285 -2720
rect 30785 -2885 30795 -2765
rect 30915 -2885 30970 -2765
rect 31090 -2885 31135 -2765
rect 31255 -2885 31300 -2765
rect 31420 -2885 31465 -2765
rect 31585 -2885 31640 -2765
rect 31760 -2885 31805 -2765
rect 31925 -2885 31970 -2765
rect 32090 -2885 32135 -2765
rect 32255 -2885 32310 -2765
rect 32430 -2885 32475 -2765
rect 32595 -2885 32640 -2765
rect 32760 -2885 32805 -2765
rect 32925 -2885 32980 -2765
rect 33100 -2885 33145 -2765
rect 33265 -2885 33310 -2765
rect 33430 -2885 33475 -2765
rect 33595 -2885 33650 -2765
rect 33770 -2885 33815 -2765
rect 33935 -2885 33980 -2765
rect 34100 -2885 34145 -2765
rect 34265 -2885 34320 -2765
rect 34440 -2885 34485 -2765
rect 34605 -2885 34650 -2765
rect 34770 -2885 34815 -2765
rect 34935 -2885 34990 -2765
rect 35110 -2885 35155 -2765
rect 35275 -2885 35320 -2765
rect 35440 -2885 35485 -2765
rect 35605 -2885 35660 -2765
rect 35780 -2885 35825 -2765
rect 35945 -2885 35990 -2765
rect 36110 -2885 36155 -2765
rect 36275 -2885 36285 -2765
rect 30785 -2930 36285 -2885
rect 30785 -3050 30795 -2930
rect 30915 -3050 30970 -2930
rect 31090 -3050 31135 -2930
rect 31255 -3050 31300 -2930
rect 31420 -3050 31465 -2930
rect 31585 -3050 31640 -2930
rect 31760 -3050 31805 -2930
rect 31925 -3050 31970 -2930
rect 32090 -3050 32135 -2930
rect 32255 -3050 32310 -2930
rect 32430 -3050 32475 -2930
rect 32595 -3050 32640 -2930
rect 32760 -3050 32805 -2930
rect 32925 -3050 32980 -2930
rect 33100 -3050 33145 -2930
rect 33265 -3050 33310 -2930
rect 33430 -3050 33475 -2930
rect 33595 -3050 33650 -2930
rect 33770 -3050 33815 -2930
rect 33935 -3050 33980 -2930
rect 34100 -3050 34145 -2930
rect 34265 -3050 34320 -2930
rect 34440 -3050 34485 -2930
rect 34605 -3050 34650 -2930
rect 34770 -3050 34815 -2930
rect 34935 -3050 34990 -2930
rect 35110 -3050 35155 -2930
rect 35275 -3050 35320 -2930
rect 35440 -3050 35485 -2930
rect 35605 -3050 35660 -2930
rect 35780 -3050 35825 -2930
rect 35945 -3050 35990 -2930
rect 36110 -3050 36155 -2930
rect 36275 -3050 36285 -2930
rect 30785 -3095 36285 -3050
rect 30785 -3215 30795 -3095
rect 30915 -3215 30970 -3095
rect 31090 -3215 31135 -3095
rect 31255 -3215 31300 -3095
rect 31420 -3215 31465 -3095
rect 31585 -3215 31640 -3095
rect 31760 -3215 31805 -3095
rect 31925 -3215 31970 -3095
rect 32090 -3215 32135 -3095
rect 32255 -3215 32310 -3095
rect 32430 -3215 32475 -3095
rect 32595 -3215 32640 -3095
rect 32760 -3215 32805 -3095
rect 32925 -3215 32980 -3095
rect 33100 -3215 33145 -3095
rect 33265 -3215 33310 -3095
rect 33430 -3215 33475 -3095
rect 33595 -3215 33650 -3095
rect 33770 -3215 33815 -3095
rect 33935 -3215 33980 -3095
rect 34100 -3215 34145 -3095
rect 34265 -3215 34320 -3095
rect 34440 -3215 34485 -3095
rect 34605 -3215 34650 -3095
rect 34770 -3215 34815 -3095
rect 34935 -3215 34990 -3095
rect 35110 -3215 35155 -3095
rect 35275 -3215 35320 -3095
rect 35440 -3215 35485 -3095
rect 35605 -3215 35660 -3095
rect 35780 -3215 35825 -3095
rect 35945 -3215 35990 -3095
rect 36110 -3215 36155 -3095
rect 36275 -3215 36285 -3095
rect 30785 -3270 36285 -3215
rect 30785 -3390 30795 -3270
rect 30915 -3390 30970 -3270
rect 31090 -3390 31135 -3270
rect 31255 -3390 31300 -3270
rect 31420 -3390 31465 -3270
rect 31585 -3390 31640 -3270
rect 31760 -3390 31805 -3270
rect 31925 -3390 31970 -3270
rect 32090 -3390 32135 -3270
rect 32255 -3390 32310 -3270
rect 32430 -3390 32475 -3270
rect 32595 -3390 32640 -3270
rect 32760 -3390 32805 -3270
rect 32925 -3390 32980 -3270
rect 33100 -3390 33145 -3270
rect 33265 -3390 33310 -3270
rect 33430 -3390 33475 -3270
rect 33595 -3390 33650 -3270
rect 33770 -3390 33815 -3270
rect 33935 -3390 33980 -3270
rect 34100 -3390 34145 -3270
rect 34265 -3390 34320 -3270
rect 34440 -3390 34485 -3270
rect 34605 -3390 34650 -3270
rect 34770 -3390 34815 -3270
rect 34935 -3390 34990 -3270
rect 35110 -3390 35155 -3270
rect 35275 -3390 35320 -3270
rect 35440 -3390 35485 -3270
rect 35605 -3390 35660 -3270
rect 35780 -3390 35825 -3270
rect 35945 -3390 35990 -3270
rect 36110 -3390 36155 -3270
rect 36275 -3390 36285 -3270
rect 30785 -3435 36285 -3390
rect 30785 -3555 30795 -3435
rect 30915 -3555 30970 -3435
rect 31090 -3555 31135 -3435
rect 31255 -3555 31300 -3435
rect 31420 -3555 31465 -3435
rect 31585 -3555 31640 -3435
rect 31760 -3555 31805 -3435
rect 31925 -3555 31970 -3435
rect 32090 -3555 32135 -3435
rect 32255 -3555 32310 -3435
rect 32430 -3555 32475 -3435
rect 32595 -3555 32640 -3435
rect 32760 -3555 32805 -3435
rect 32925 -3555 32980 -3435
rect 33100 -3555 33145 -3435
rect 33265 -3555 33310 -3435
rect 33430 -3555 33475 -3435
rect 33595 -3555 33650 -3435
rect 33770 -3555 33815 -3435
rect 33935 -3555 33980 -3435
rect 34100 -3555 34145 -3435
rect 34265 -3555 34320 -3435
rect 34440 -3555 34485 -3435
rect 34605 -3555 34650 -3435
rect 34770 -3555 34815 -3435
rect 34935 -3555 34990 -3435
rect 35110 -3555 35155 -3435
rect 35275 -3555 35320 -3435
rect 35440 -3555 35485 -3435
rect 35605 -3555 35660 -3435
rect 35780 -3555 35825 -3435
rect 35945 -3555 35990 -3435
rect 36110 -3555 36155 -3435
rect 36275 -3555 36285 -3435
rect 30785 -3600 36285 -3555
rect 30785 -3720 30795 -3600
rect 30915 -3720 30970 -3600
rect 31090 -3720 31135 -3600
rect 31255 -3720 31300 -3600
rect 31420 -3720 31465 -3600
rect 31585 -3720 31640 -3600
rect 31760 -3720 31805 -3600
rect 31925 -3720 31970 -3600
rect 32090 -3720 32135 -3600
rect 32255 -3720 32310 -3600
rect 32430 -3720 32475 -3600
rect 32595 -3720 32640 -3600
rect 32760 -3720 32805 -3600
rect 32925 -3720 32980 -3600
rect 33100 -3720 33145 -3600
rect 33265 -3720 33310 -3600
rect 33430 -3720 33475 -3600
rect 33595 -3720 33650 -3600
rect 33770 -3720 33815 -3600
rect 33935 -3720 33980 -3600
rect 34100 -3720 34145 -3600
rect 34265 -3720 34320 -3600
rect 34440 -3720 34485 -3600
rect 34605 -3720 34650 -3600
rect 34770 -3720 34815 -3600
rect 34935 -3720 34990 -3600
rect 35110 -3720 35155 -3600
rect 35275 -3720 35320 -3600
rect 35440 -3720 35485 -3600
rect 35605 -3720 35660 -3600
rect 35780 -3720 35825 -3600
rect 35945 -3720 35990 -3600
rect 36110 -3720 36155 -3600
rect 36275 -3720 36285 -3600
rect 30785 -3765 36285 -3720
rect 30785 -3885 30795 -3765
rect 30915 -3885 30970 -3765
rect 31090 -3885 31135 -3765
rect 31255 -3885 31300 -3765
rect 31420 -3885 31465 -3765
rect 31585 -3885 31640 -3765
rect 31760 -3885 31805 -3765
rect 31925 -3885 31970 -3765
rect 32090 -3885 32135 -3765
rect 32255 -3885 32310 -3765
rect 32430 -3885 32475 -3765
rect 32595 -3885 32640 -3765
rect 32760 -3885 32805 -3765
rect 32925 -3885 32980 -3765
rect 33100 -3885 33145 -3765
rect 33265 -3885 33310 -3765
rect 33430 -3885 33475 -3765
rect 33595 -3885 33650 -3765
rect 33770 -3885 33815 -3765
rect 33935 -3885 33980 -3765
rect 34100 -3885 34145 -3765
rect 34265 -3885 34320 -3765
rect 34440 -3885 34485 -3765
rect 34605 -3885 34650 -3765
rect 34770 -3885 34815 -3765
rect 34935 -3885 34990 -3765
rect 35110 -3885 35155 -3765
rect 35275 -3885 35320 -3765
rect 35440 -3885 35485 -3765
rect 35605 -3885 35660 -3765
rect 35780 -3885 35825 -3765
rect 35945 -3885 35990 -3765
rect 36110 -3885 36155 -3765
rect 36275 -3885 36285 -3765
rect 30785 -3940 36285 -3885
rect 30785 -4060 30795 -3940
rect 30915 -4060 30970 -3940
rect 31090 -4060 31135 -3940
rect 31255 -4060 31300 -3940
rect 31420 -4060 31465 -3940
rect 31585 -4060 31640 -3940
rect 31760 -4060 31805 -3940
rect 31925 -4060 31970 -3940
rect 32090 -4060 32135 -3940
rect 32255 -4060 32310 -3940
rect 32430 -4060 32475 -3940
rect 32595 -4060 32640 -3940
rect 32760 -4060 32805 -3940
rect 32925 -4060 32980 -3940
rect 33100 -4060 33145 -3940
rect 33265 -4060 33310 -3940
rect 33430 -4060 33475 -3940
rect 33595 -4060 33650 -3940
rect 33770 -4060 33815 -3940
rect 33935 -4060 33980 -3940
rect 34100 -4060 34145 -3940
rect 34265 -4060 34320 -3940
rect 34440 -4060 34485 -3940
rect 34605 -4060 34650 -3940
rect 34770 -4060 34815 -3940
rect 34935 -4060 34990 -3940
rect 35110 -4060 35155 -3940
rect 35275 -4060 35320 -3940
rect 35440 -4060 35485 -3940
rect 35605 -4060 35660 -3940
rect 35780 -4060 35825 -3940
rect 35945 -4060 35990 -3940
rect 36110 -4060 36155 -3940
rect 36275 -4060 36285 -3940
rect 30785 -4070 36285 -4060
rect 36475 1420 41975 1430
rect 36475 1300 36485 1420
rect 36605 1300 36660 1420
rect 36780 1300 36825 1420
rect 36945 1300 36990 1420
rect 37110 1300 37155 1420
rect 37275 1300 37330 1420
rect 37450 1300 37495 1420
rect 37615 1300 37660 1420
rect 37780 1300 37825 1420
rect 37945 1300 38000 1420
rect 38120 1300 38165 1420
rect 38285 1300 38330 1420
rect 38450 1300 38495 1420
rect 38615 1300 38670 1420
rect 38790 1300 38835 1420
rect 38955 1300 39000 1420
rect 39120 1300 39165 1420
rect 39285 1300 39340 1420
rect 39460 1300 39505 1420
rect 39625 1300 39670 1420
rect 39790 1300 39835 1420
rect 39955 1300 40010 1420
rect 40130 1300 40175 1420
rect 40295 1300 40340 1420
rect 40460 1300 40505 1420
rect 40625 1300 40680 1420
rect 40800 1300 40845 1420
rect 40965 1300 41010 1420
rect 41130 1300 41175 1420
rect 41295 1300 41350 1420
rect 41470 1300 41515 1420
rect 41635 1300 41680 1420
rect 41800 1300 41845 1420
rect 41965 1300 41975 1420
rect 36475 1255 41975 1300
rect 36475 1135 36485 1255
rect 36605 1135 36660 1255
rect 36780 1135 36825 1255
rect 36945 1135 36990 1255
rect 37110 1135 37155 1255
rect 37275 1135 37330 1255
rect 37450 1135 37495 1255
rect 37615 1135 37660 1255
rect 37780 1135 37825 1255
rect 37945 1135 38000 1255
rect 38120 1135 38165 1255
rect 38285 1135 38330 1255
rect 38450 1135 38495 1255
rect 38615 1135 38670 1255
rect 38790 1135 38835 1255
rect 38955 1135 39000 1255
rect 39120 1135 39165 1255
rect 39285 1135 39340 1255
rect 39460 1135 39505 1255
rect 39625 1135 39670 1255
rect 39790 1135 39835 1255
rect 39955 1135 40010 1255
rect 40130 1135 40175 1255
rect 40295 1135 40340 1255
rect 40460 1135 40505 1255
rect 40625 1135 40680 1255
rect 40800 1135 40845 1255
rect 40965 1135 41010 1255
rect 41130 1135 41175 1255
rect 41295 1135 41350 1255
rect 41470 1135 41515 1255
rect 41635 1135 41680 1255
rect 41800 1135 41845 1255
rect 41965 1135 41975 1255
rect 36475 1090 41975 1135
rect 36475 970 36485 1090
rect 36605 970 36660 1090
rect 36780 970 36825 1090
rect 36945 970 36990 1090
rect 37110 970 37155 1090
rect 37275 970 37330 1090
rect 37450 970 37495 1090
rect 37615 970 37660 1090
rect 37780 970 37825 1090
rect 37945 970 38000 1090
rect 38120 970 38165 1090
rect 38285 970 38330 1090
rect 38450 970 38495 1090
rect 38615 970 38670 1090
rect 38790 970 38835 1090
rect 38955 970 39000 1090
rect 39120 970 39165 1090
rect 39285 970 39340 1090
rect 39460 970 39505 1090
rect 39625 970 39670 1090
rect 39790 970 39835 1090
rect 39955 970 40010 1090
rect 40130 970 40175 1090
rect 40295 970 40340 1090
rect 40460 970 40505 1090
rect 40625 970 40680 1090
rect 40800 970 40845 1090
rect 40965 970 41010 1090
rect 41130 970 41175 1090
rect 41295 970 41350 1090
rect 41470 970 41515 1090
rect 41635 970 41680 1090
rect 41800 970 41845 1090
rect 41965 970 41975 1090
rect 36475 925 41975 970
rect 36475 805 36485 925
rect 36605 805 36660 925
rect 36780 805 36825 925
rect 36945 805 36990 925
rect 37110 805 37155 925
rect 37275 805 37330 925
rect 37450 805 37495 925
rect 37615 805 37660 925
rect 37780 805 37825 925
rect 37945 805 38000 925
rect 38120 805 38165 925
rect 38285 805 38330 925
rect 38450 805 38495 925
rect 38615 805 38670 925
rect 38790 805 38835 925
rect 38955 805 39000 925
rect 39120 805 39165 925
rect 39285 805 39340 925
rect 39460 805 39505 925
rect 39625 805 39670 925
rect 39790 805 39835 925
rect 39955 805 40010 925
rect 40130 805 40175 925
rect 40295 805 40340 925
rect 40460 805 40505 925
rect 40625 805 40680 925
rect 40800 805 40845 925
rect 40965 805 41010 925
rect 41130 805 41175 925
rect 41295 805 41350 925
rect 41470 805 41515 925
rect 41635 805 41680 925
rect 41800 805 41845 925
rect 41965 805 41975 925
rect 36475 750 41975 805
rect 36475 630 36485 750
rect 36605 630 36660 750
rect 36780 630 36825 750
rect 36945 630 36990 750
rect 37110 630 37155 750
rect 37275 630 37330 750
rect 37450 630 37495 750
rect 37615 630 37660 750
rect 37780 630 37825 750
rect 37945 630 38000 750
rect 38120 630 38165 750
rect 38285 630 38330 750
rect 38450 630 38495 750
rect 38615 630 38670 750
rect 38790 630 38835 750
rect 38955 630 39000 750
rect 39120 630 39165 750
rect 39285 630 39340 750
rect 39460 630 39505 750
rect 39625 630 39670 750
rect 39790 630 39835 750
rect 39955 630 40010 750
rect 40130 630 40175 750
rect 40295 630 40340 750
rect 40460 630 40505 750
rect 40625 630 40680 750
rect 40800 630 40845 750
rect 40965 630 41010 750
rect 41130 630 41175 750
rect 41295 630 41350 750
rect 41470 630 41515 750
rect 41635 630 41680 750
rect 41800 630 41845 750
rect 41965 630 41975 750
rect 36475 585 41975 630
rect 36475 465 36485 585
rect 36605 465 36660 585
rect 36780 465 36825 585
rect 36945 465 36990 585
rect 37110 465 37155 585
rect 37275 465 37330 585
rect 37450 465 37495 585
rect 37615 465 37660 585
rect 37780 465 37825 585
rect 37945 465 38000 585
rect 38120 465 38165 585
rect 38285 465 38330 585
rect 38450 465 38495 585
rect 38615 465 38670 585
rect 38790 465 38835 585
rect 38955 465 39000 585
rect 39120 465 39165 585
rect 39285 465 39340 585
rect 39460 465 39505 585
rect 39625 465 39670 585
rect 39790 465 39835 585
rect 39955 465 40010 585
rect 40130 465 40175 585
rect 40295 465 40340 585
rect 40460 465 40505 585
rect 40625 465 40680 585
rect 40800 465 40845 585
rect 40965 465 41010 585
rect 41130 465 41175 585
rect 41295 465 41350 585
rect 41470 465 41515 585
rect 41635 465 41680 585
rect 41800 465 41845 585
rect 41965 465 41975 585
rect 36475 420 41975 465
rect 36475 300 36485 420
rect 36605 300 36660 420
rect 36780 300 36825 420
rect 36945 300 36990 420
rect 37110 300 37155 420
rect 37275 300 37330 420
rect 37450 300 37495 420
rect 37615 300 37660 420
rect 37780 300 37825 420
rect 37945 300 38000 420
rect 38120 300 38165 420
rect 38285 300 38330 420
rect 38450 300 38495 420
rect 38615 300 38670 420
rect 38790 300 38835 420
rect 38955 300 39000 420
rect 39120 300 39165 420
rect 39285 300 39340 420
rect 39460 300 39505 420
rect 39625 300 39670 420
rect 39790 300 39835 420
rect 39955 300 40010 420
rect 40130 300 40175 420
rect 40295 300 40340 420
rect 40460 300 40505 420
rect 40625 300 40680 420
rect 40800 300 40845 420
rect 40965 300 41010 420
rect 41130 300 41175 420
rect 41295 300 41350 420
rect 41470 300 41515 420
rect 41635 300 41680 420
rect 41800 300 41845 420
rect 41965 300 41975 420
rect 36475 255 41975 300
rect 36475 135 36485 255
rect 36605 135 36660 255
rect 36780 135 36825 255
rect 36945 135 36990 255
rect 37110 135 37155 255
rect 37275 135 37330 255
rect 37450 135 37495 255
rect 37615 135 37660 255
rect 37780 135 37825 255
rect 37945 135 38000 255
rect 38120 135 38165 255
rect 38285 135 38330 255
rect 38450 135 38495 255
rect 38615 135 38670 255
rect 38790 135 38835 255
rect 38955 135 39000 255
rect 39120 135 39165 255
rect 39285 135 39340 255
rect 39460 135 39505 255
rect 39625 135 39670 255
rect 39790 135 39835 255
rect 39955 135 40010 255
rect 40130 135 40175 255
rect 40295 135 40340 255
rect 40460 135 40505 255
rect 40625 135 40680 255
rect 40800 135 40845 255
rect 40965 135 41010 255
rect 41130 135 41175 255
rect 41295 135 41350 255
rect 41470 135 41515 255
rect 41635 135 41680 255
rect 41800 135 41845 255
rect 41965 135 41975 255
rect 36475 80 41975 135
rect 36475 -40 36485 80
rect 36605 -40 36660 80
rect 36780 -40 36825 80
rect 36945 -40 36990 80
rect 37110 -40 37155 80
rect 37275 -40 37330 80
rect 37450 -40 37495 80
rect 37615 -40 37660 80
rect 37780 -40 37825 80
rect 37945 -40 38000 80
rect 38120 -40 38165 80
rect 38285 -40 38330 80
rect 38450 -40 38495 80
rect 38615 -40 38670 80
rect 38790 -40 38835 80
rect 38955 -40 39000 80
rect 39120 -40 39165 80
rect 39285 -40 39340 80
rect 39460 -40 39505 80
rect 39625 -40 39670 80
rect 39790 -40 39835 80
rect 39955 -40 40010 80
rect 40130 -40 40175 80
rect 40295 -40 40340 80
rect 40460 -40 40505 80
rect 40625 -40 40680 80
rect 40800 -40 40845 80
rect 40965 -40 41010 80
rect 41130 -40 41175 80
rect 41295 -40 41350 80
rect 41470 -40 41515 80
rect 41635 -40 41680 80
rect 41800 -40 41845 80
rect 41965 -40 41975 80
rect 36475 -85 41975 -40
rect 36475 -205 36485 -85
rect 36605 -205 36660 -85
rect 36780 -205 36825 -85
rect 36945 -205 36990 -85
rect 37110 -205 37155 -85
rect 37275 -205 37330 -85
rect 37450 -205 37495 -85
rect 37615 -205 37660 -85
rect 37780 -205 37825 -85
rect 37945 -205 38000 -85
rect 38120 -205 38165 -85
rect 38285 -205 38330 -85
rect 38450 -205 38495 -85
rect 38615 -205 38670 -85
rect 38790 -205 38835 -85
rect 38955 -205 39000 -85
rect 39120 -205 39165 -85
rect 39285 -205 39340 -85
rect 39460 -205 39505 -85
rect 39625 -205 39670 -85
rect 39790 -205 39835 -85
rect 39955 -205 40010 -85
rect 40130 -205 40175 -85
rect 40295 -205 40340 -85
rect 40460 -205 40505 -85
rect 40625 -205 40680 -85
rect 40800 -205 40845 -85
rect 40965 -205 41010 -85
rect 41130 -205 41175 -85
rect 41295 -205 41350 -85
rect 41470 -205 41515 -85
rect 41635 -205 41680 -85
rect 41800 -205 41845 -85
rect 41965 -205 41975 -85
rect 36475 -250 41975 -205
rect 36475 -370 36485 -250
rect 36605 -370 36660 -250
rect 36780 -370 36825 -250
rect 36945 -370 36990 -250
rect 37110 -370 37155 -250
rect 37275 -370 37330 -250
rect 37450 -370 37495 -250
rect 37615 -370 37660 -250
rect 37780 -370 37825 -250
rect 37945 -370 38000 -250
rect 38120 -370 38165 -250
rect 38285 -370 38330 -250
rect 38450 -370 38495 -250
rect 38615 -370 38670 -250
rect 38790 -370 38835 -250
rect 38955 -370 39000 -250
rect 39120 -370 39165 -250
rect 39285 -370 39340 -250
rect 39460 -370 39505 -250
rect 39625 -370 39670 -250
rect 39790 -370 39835 -250
rect 39955 -370 40010 -250
rect 40130 -370 40175 -250
rect 40295 -370 40340 -250
rect 40460 -370 40505 -250
rect 40625 -370 40680 -250
rect 40800 -370 40845 -250
rect 40965 -370 41010 -250
rect 41130 -370 41175 -250
rect 41295 -370 41350 -250
rect 41470 -370 41515 -250
rect 41635 -370 41680 -250
rect 41800 -370 41845 -250
rect 41965 -370 41975 -250
rect 36475 -415 41975 -370
rect 36475 -535 36485 -415
rect 36605 -535 36660 -415
rect 36780 -535 36825 -415
rect 36945 -535 36990 -415
rect 37110 -535 37155 -415
rect 37275 -535 37330 -415
rect 37450 -535 37495 -415
rect 37615 -535 37660 -415
rect 37780 -535 37825 -415
rect 37945 -535 38000 -415
rect 38120 -535 38165 -415
rect 38285 -535 38330 -415
rect 38450 -535 38495 -415
rect 38615 -535 38670 -415
rect 38790 -535 38835 -415
rect 38955 -535 39000 -415
rect 39120 -535 39165 -415
rect 39285 -535 39340 -415
rect 39460 -535 39505 -415
rect 39625 -535 39670 -415
rect 39790 -535 39835 -415
rect 39955 -535 40010 -415
rect 40130 -535 40175 -415
rect 40295 -535 40340 -415
rect 40460 -535 40505 -415
rect 40625 -535 40680 -415
rect 40800 -535 40845 -415
rect 40965 -535 41010 -415
rect 41130 -535 41175 -415
rect 41295 -535 41350 -415
rect 41470 -535 41515 -415
rect 41635 -535 41680 -415
rect 41800 -535 41845 -415
rect 41965 -535 41975 -415
rect 36475 -590 41975 -535
rect 36475 -710 36485 -590
rect 36605 -710 36660 -590
rect 36780 -710 36825 -590
rect 36945 -710 36990 -590
rect 37110 -710 37155 -590
rect 37275 -710 37330 -590
rect 37450 -710 37495 -590
rect 37615 -710 37660 -590
rect 37780 -710 37825 -590
rect 37945 -710 38000 -590
rect 38120 -710 38165 -590
rect 38285 -710 38330 -590
rect 38450 -710 38495 -590
rect 38615 -710 38670 -590
rect 38790 -710 38835 -590
rect 38955 -710 39000 -590
rect 39120 -710 39165 -590
rect 39285 -710 39340 -590
rect 39460 -710 39505 -590
rect 39625 -710 39670 -590
rect 39790 -710 39835 -590
rect 39955 -710 40010 -590
rect 40130 -710 40175 -590
rect 40295 -710 40340 -590
rect 40460 -710 40505 -590
rect 40625 -710 40680 -590
rect 40800 -710 40845 -590
rect 40965 -710 41010 -590
rect 41130 -710 41175 -590
rect 41295 -710 41350 -590
rect 41470 -710 41515 -590
rect 41635 -710 41680 -590
rect 41800 -710 41845 -590
rect 41965 -710 41975 -590
rect 36475 -755 41975 -710
rect 36475 -875 36485 -755
rect 36605 -875 36660 -755
rect 36780 -875 36825 -755
rect 36945 -875 36990 -755
rect 37110 -875 37155 -755
rect 37275 -875 37330 -755
rect 37450 -875 37495 -755
rect 37615 -875 37660 -755
rect 37780 -875 37825 -755
rect 37945 -875 38000 -755
rect 38120 -875 38165 -755
rect 38285 -875 38330 -755
rect 38450 -875 38495 -755
rect 38615 -875 38670 -755
rect 38790 -875 38835 -755
rect 38955 -875 39000 -755
rect 39120 -875 39165 -755
rect 39285 -875 39340 -755
rect 39460 -875 39505 -755
rect 39625 -875 39670 -755
rect 39790 -875 39835 -755
rect 39955 -875 40010 -755
rect 40130 -875 40175 -755
rect 40295 -875 40340 -755
rect 40460 -875 40505 -755
rect 40625 -875 40680 -755
rect 40800 -875 40845 -755
rect 40965 -875 41010 -755
rect 41130 -875 41175 -755
rect 41295 -875 41350 -755
rect 41470 -875 41515 -755
rect 41635 -875 41680 -755
rect 41800 -875 41845 -755
rect 41965 -875 41975 -755
rect 36475 -920 41975 -875
rect 36475 -1040 36485 -920
rect 36605 -1040 36660 -920
rect 36780 -1040 36825 -920
rect 36945 -1040 36990 -920
rect 37110 -1040 37155 -920
rect 37275 -1040 37330 -920
rect 37450 -1040 37495 -920
rect 37615 -1040 37660 -920
rect 37780 -1040 37825 -920
rect 37945 -1040 38000 -920
rect 38120 -1040 38165 -920
rect 38285 -1040 38330 -920
rect 38450 -1040 38495 -920
rect 38615 -1040 38670 -920
rect 38790 -1040 38835 -920
rect 38955 -1040 39000 -920
rect 39120 -1040 39165 -920
rect 39285 -1040 39340 -920
rect 39460 -1040 39505 -920
rect 39625 -1040 39670 -920
rect 39790 -1040 39835 -920
rect 39955 -1040 40010 -920
rect 40130 -1040 40175 -920
rect 40295 -1040 40340 -920
rect 40460 -1040 40505 -920
rect 40625 -1040 40680 -920
rect 40800 -1040 40845 -920
rect 40965 -1040 41010 -920
rect 41130 -1040 41175 -920
rect 41295 -1040 41350 -920
rect 41470 -1040 41515 -920
rect 41635 -1040 41680 -920
rect 41800 -1040 41845 -920
rect 41965 -1040 41975 -920
rect 36475 -1085 41975 -1040
rect 36475 -1205 36485 -1085
rect 36605 -1205 36660 -1085
rect 36780 -1205 36825 -1085
rect 36945 -1205 36990 -1085
rect 37110 -1205 37155 -1085
rect 37275 -1205 37330 -1085
rect 37450 -1205 37495 -1085
rect 37615 -1205 37660 -1085
rect 37780 -1205 37825 -1085
rect 37945 -1205 38000 -1085
rect 38120 -1205 38165 -1085
rect 38285 -1205 38330 -1085
rect 38450 -1205 38495 -1085
rect 38615 -1205 38670 -1085
rect 38790 -1205 38835 -1085
rect 38955 -1205 39000 -1085
rect 39120 -1205 39165 -1085
rect 39285 -1205 39340 -1085
rect 39460 -1205 39505 -1085
rect 39625 -1205 39670 -1085
rect 39790 -1205 39835 -1085
rect 39955 -1205 40010 -1085
rect 40130 -1205 40175 -1085
rect 40295 -1205 40340 -1085
rect 40460 -1205 40505 -1085
rect 40625 -1205 40680 -1085
rect 40800 -1205 40845 -1085
rect 40965 -1205 41010 -1085
rect 41130 -1205 41175 -1085
rect 41295 -1205 41350 -1085
rect 41470 -1205 41515 -1085
rect 41635 -1205 41680 -1085
rect 41800 -1205 41845 -1085
rect 41965 -1205 41975 -1085
rect 36475 -1260 41975 -1205
rect 36475 -1380 36485 -1260
rect 36605 -1380 36660 -1260
rect 36780 -1380 36825 -1260
rect 36945 -1380 36990 -1260
rect 37110 -1380 37155 -1260
rect 37275 -1380 37330 -1260
rect 37450 -1380 37495 -1260
rect 37615 -1380 37660 -1260
rect 37780 -1380 37825 -1260
rect 37945 -1380 38000 -1260
rect 38120 -1380 38165 -1260
rect 38285 -1380 38330 -1260
rect 38450 -1380 38495 -1260
rect 38615 -1380 38670 -1260
rect 38790 -1380 38835 -1260
rect 38955 -1380 39000 -1260
rect 39120 -1380 39165 -1260
rect 39285 -1380 39340 -1260
rect 39460 -1380 39505 -1260
rect 39625 -1380 39670 -1260
rect 39790 -1380 39835 -1260
rect 39955 -1380 40010 -1260
rect 40130 -1380 40175 -1260
rect 40295 -1380 40340 -1260
rect 40460 -1380 40505 -1260
rect 40625 -1380 40680 -1260
rect 40800 -1380 40845 -1260
rect 40965 -1380 41010 -1260
rect 41130 -1380 41175 -1260
rect 41295 -1380 41350 -1260
rect 41470 -1380 41515 -1260
rect 41635 -1380 41680 -1260
rect 41800 -1380 41845 -1260
rect 41965 -1380 41975 -1260
rect 36475 -1425 41975 -1380
rect 36475 -1545 36485 -1425
rect 36605 -1545 36660 -1425
rect 36780 -1545 36825 -1425
rect 36945 -1545 36990 -1425
rect 37110 -1545 37155 -1425
rect 37275 -1545 37330 -1425
rect 37450 -1545 37495 -1425
rect 37615 -1545 37660 -1425
rect 37780 -1545 37825 -1425
rect 37945 -1545 38000 -1425
rect 38120 -1545 38165 -1425
rect 38285 -1545 38330 -1425
rect 38450 -1545 38495 -1425
rect 38615 -1545 38670 -1425
rect 38790 -1545 38835 -1425
rect 38955 -1545 39000 -1425
rect 39120 -1545 39165 -1425
rect 39285 -1545 39340 -1425
rect 39460 -1545 39505 -1425
rect 39625 -1545 39670 -1425
rect 39790 -1545 39835 -1425
rect 39955 -1545 40010 -1425
rect 40130 -1545 40175 -1425
rect 40295 -1545 40340 -1425
rect 40460 -1545 40505 -1425
rect 40625 -1545 40680 -1425
rect 40800 -1545 40845 -1425
rect 40965 -1545 41010 -1425
rect 41130 -1545 41175 -1425
rect 41295 -1545 41350 -1425
rect 41470 -1545 41515 -1425
rect 41635 -1545 41680 -1425
rect 41800 -1545 41845 -1425
rect 41965 -1545 41975 -1425
rect 36475 -1590 41975 -1545
rect 36475 -1710 36485 -1590
rect 36605 -1710 36660 -1590
rect 36780 -1710 36825 -1590
rect 36945 -1710 36990 -1590
rect 37110 -1710 37155 -1590
rect 37275 -1710 37330 -1590
rect 37450 -1710 37495 -1590
rect 37615 -1710 37660 -1590
rect 37780 -1710 37825 -1590
rect 37945 -1710 38000 -1590
rect 38120 -1710 38165 -1590
rect 38285 -1710 38330 -1590
rect 38450 -1710 38495 -1590
rect 38615 -1710 38670 -1590
rect 38790 -1710 38835 -1590
rect 38955 -1710 39000 -1590
rect 39120 -1710 39165 -1590
rect 39285 -1710 39340 -1590
rect 39460 -1710 39505 -1590
rect 39625 -1710 39670 -1590
rect 39790 -1710 39835 -1590
rect 39955 -1710 40010 -1590
rect 40130 -1710 40175 -1590
rect 40295 -1710 40340 -1590
rect 40460 -1710 40505 -1590
rect 40625 -1710 40680 -1590
rect 40800 -1710 40845 -1590
rect 40965 -1710 41010 -1590
rect 41130 -1710 41175 -1590
rect 41295 -1710 41350 -1590
rect 41470 -1710 41515 -1590
rect 41635 -1710 41680 -1590
rect 41800 -1710 41845 -1590
rect 41965 -1710 41975 -1590
rect 36475 -1755 41975 -1710
rect 36475 -1875 36485 -1755
rect 36605 -1875 36660 -1755
rect 36780 -1875 36825 -1755
rect 36945 -1875 36990 -1755
rect 37110 -1875 37155 -1755
rect 37275 -1875 37330 -1755
rect 37450 -1875 37495 -1755
rect 37615 -1875 37660 -1755
rect 37780 -1875 37825 -1755
rect 37945 -1875 38000 -1755
rect 38120 -1875 38165 -1755
rect 38285 -1875 38330 -1755
rect 38450 -1875 38495 -1755
rect 38615 -1875 38670 -1755
rect 38790 -1875 38835 -1755
rect 38955 -1875 39000 -1755
rect 39120 -1875 39165 -1755
rect 39285 -1875 39340 -1755
rect 39460 -1875 39505 -1755
rect 39625 -1875 39670 -1755
rect 39790 -1875 39835 -1755
rect 39955 -1875 40010 -1755
rect 40130 -1875 40175 -1755
rect 40295 -1875 40340 -1755
rect 40460 -1875 40505 -1755
rect 40625 -1875 40680 -1755
rect 40800 -1875 40845 -1755
rect 40965 -1875 41010 -1755
rect 41130 -1875 41175 -1755
rect 41295 -1875 41350 -1755
rect 41470 -1875 41515 -1755
rect 41635 -1875 41680 -1755
rect 41800 -1875 41845 -1755
rect 41965 -1875 41975 -1755
rect 36475 -1930 41975 -1875
rect 36475 -2050 36485 -1930
rect 36605 -2050 36660 -1930
rect 36780 -2050 36825 -1930
rect 36945 -2050 36990 -1930
rect 37110 -2050 37155 -1930
rect 37275 -2050 37330 -1930
rect 37450 -2050 37495 -1930
rect 37615 -2050 37660 -1930
rect 37780 -2050 37825 -1930
rect 37945 -2050 38000 -1930
rect 38120 -2050 38165 -1930
rect 38285 -2050 38330 -1930
rect 38450 -2050 38495 -1930
rect 38615 -2050 38670 -1930
rect 38790 -2050 38835 -1930
rect 38955 -2050 39000 -1930
rect 39120 -2050 39165 -1930
rect 39285 -2050 39340 -1930
rect 39460 -2050 39505 -1930
rect 39625 -2050 39670 -1930
rect 39790 -2050 39835 -1930
rect 39955 -2050 40010 -1930
rect 40130 -2050 40175 -1930
rect 40295 -2050 40340 -1930
rect 40460 -2050 40505 -1930
rect 40625 -2050 40680 -1930
rect 40800 -2050 40845 -1930
rect 40965 -2050 41010 -1930
rect 41130 -2050 41175 -1930
rect 41295 -2050 41350 -1930
rect 41470 -2050 41515 -1930
rect 41635 -2050 41680 -1930
rect 41800 -2050 41845 -1930
rect 41965 -2050 41975 -1930
rect 36475 -2095 41975 -2050
rect 36475 -2215 36485 -2095
rect 36605 -2215 36660 -2095
rect 36780 -2215 36825 -2095
rect 36945 -2215 36990 -2095
rect 37110 -2215 37155 -2095
rect 37275 -2215 37330 -2095
rect 37450 -2215 37495 -2095
rect 37615 -2215 37660 -2095
rect 37780 -2215 37825 -2095
rect 37945 -2215 38000 -2095
rect 38120 -2215 38165 -2095
rect 38285 -2215 38330 -2095
rect 38450 -2215 38495 -2095
rect 38615 -2215 38670 -2095
rect 38790 -2215 38835 -2095
rect 38955 -2215 39000 -2095
rect 39120 -2215 39165 -2095
rect 39285 -2215 39340 -2095
rect 39460 -2215 39505 -2095
rect 39625 -2215 39670 -2095
rect 39790 -2215 39835 -2095
rect 39955 -2215 40010 -2095
rect 40130 -2215 40175 -2095
rect 40295 -2215 40340 -2095
rect 40460 -2215 40505 -2095
rect 40625 -2215 40680 -2095
rect 40800 -2215 40845 -2095
rect 40965 -2215 41010 -2095
rect 41130 -2215 41175 -2095
rect 41295 -2215 41350 -2095
rect 41470 -2215 41515 -2095
rect 41635 -2215 41680 -2095
rect 41800 -2215 41845 -2095
rect 41965 -2215 41975 -2095
rect 36475 -2260 41975 -2215
rect 36475 -2380 36485 -2260
rect 36605 -2380 36660 -2260
rect 36780 -2380 36825 -2260
rect 36945 -2380 36990 -2260
rect 37110 -2380 37155 -2260
rect 37275 -2380 37330 -2260
rect 37450 -2380 37495 -2260
rect 37615 -2380 37660 -2260
rect 37780 -2380 37825 -2260
rect 37945 -2380 38000 -2260
rect 38120 -2380 38165 -2260
rect 38285 -2380 38330 -2260
rect 38450 -2380 38495 -2260
rect 38615 -2380 38670 -2260
rect 38790 -2380 38835 -2260
rect 38955 -2380 39000 -2260
rect 39120 -2380 39165 -2260
rect 39285 -2380 39340 -2260
rect 39460 -2380 39505 -2260
rect 39625 -2380 39670 -2260
rect 39790 -2380 39835 -2260
rect 39955 -2380 40010 -2260
rect 40130 -2380 40175 -2260
rect 40295 -2380 40340 -2260
rect 40460 -2380 40505 -2260
rect 40625 -2380 40680 -2260
rect 40800 -2380 40845 -2260
rect 40965 -2380 41010 -2260
rect 41130 -2380 41175 -2260
rect 41295 -2380 41350 -2260
rect 41470 -2380 41515 -2260
rect 41635 -2380 41680 -2260
rect 41800 -2380 41845 -2260
rect 41965 -2380 41975 -2260
rect 36475 -2425 41975 -2380
rect 36475 -2545 36485 -2425
rect 36605 -2545 36660 -2425
rect 36780 -2545 36825 -2425
rect 36945 -2545 36990 -2425
rect 37110 -2545 37155 -2425
rect 37275 -2545 37330 -2425
rect 37450 -2545 37495 -2425
rect 37615 -2545 37660 -2425
rect 37780 -2545 37825 -2425
rect 37945 -2545 38000 -2425
rect 38120 -2545 38165 -2425
rect 38285 -2545 38330 -2425
rect 38450 -2545 38495 -2425
rect 38615 -2545 38670 -2425
rect 38790 -2545 38835 -2425
rect 38955 -2545 39000 -2425
rect 39120 -2545 39165 -2425
rect 39285 -2545 39340 -2425
rect 39460 -2545 39505 -2425
rect 39625 -2545 39670 -2425
rect 39790 -2545 39835 -2425
rect 39955 -2545 40010 -2425
rect 40130 -2545 40175 -2425
rect 40295 -2545 40340 -2425
rect 40460 -2545 40505 -2425
rect 40625 -2545 40680 -2425
rect 40800 -2545 40845 -2425
rect 40965 -2545 41010 -2425
rect 41130 -2545 41175 -2425
rect 41295 -2545 41350 -2425
rect 41470 -2545 41515 -2425
rect 41635 -2545 41680 -2425
rect 41800 -2545 41845 -2425
rect 41965 -2545 41975 -2425
rect 36475 -2600 41975 -2545
rect 36475 -2720 36485 -2600
rect 36605 -2720 36660 -2600
rect 36780 -2720 36825 -2600
rect 36945 -2720 36990 -2600
rect 37110 -2720 37155 -2600
rect 37275 -2720 37330 -2600
rect 37450 -2720 37495 -2600
rect 37615 -2720 37660 -2600
rect 37780 -2720 37825 -2600
rect 37945 -2720 38000 -2600
rect 38120 -2720 38165 -2600
rect 38285 -2720 38330 -2600
rect 38450 -2720 38495 -2600
rect 38615 -2720 38670 -2600
rect 38790 -2720 38835 -2600
rect 38955 -2720 39000 -2600
rect 39120 -2720 39165 -2600
rect 39285 -2720 39340 -2600
rect 39460 -2720 39505 -2600
rect 39625 -2720 39670 -2600
rect 39790 -2720 39835 -2600
rect 39955 -2720 40010 -2600
rect 40130 -2720 40175 -2600
rect 40295 -2720 40340 -2600
rect 40460 -2720 40505 -2600
rect 40625 -2720 40680 -2600
rect 40800 -2720 40845 -2600
rect 40965 -2720 41010 -2600
rect 41130 -2720 41175 -2600
rect 41295 -2720 41350 -2600
rect 41470 -2720 41515 -2600
rect 41635 -2720 41680 -2600
rect 41800 -2720 41845 -2600
rect 41965 -2720 41975 -2600
rect 36475 -2765 41975 -2720
rect 36475 -2885 36485 -2765
rect 36605 -2885 36660 -2765
rect 36780 -2885 36825 -2765
rect 36945 -2885 36990 -2765
rect 37110 -2885 37155 -2765
rect 37275 -2885 37330 -2765
rect 37450 -2885 37495 -2765
rect 37615 -2885 37660 -2765
rect 37780 -2885 37825 -2765
rect 37945 -2885 38000 -2765
rect 38120 -2885 38165 -2765
rect 38285 -2885 38330 -2765
rect 38450 -2885 38495 -2765
rect 38615 -2885 38670 -2765
rect 38790 -2885 38835 -2765
rect 38955 -2885 39000 -2765
rect 39120 -2885 39165 -2765
rect 39285 -2885 39340 -2765
rect 39460 -2885 39505 -2765
rect 39625 -2885 39670 -2765
rect 39790 -2885 39835 -2765
rect 39955 -2885 40010 -2765
rect 40130 -2885 40175 -2765
rect 40295 -2885 40340 -2765
rect 40460 -2885 40505 -2765
rect 40625 -2885 40680 -2765
rect 40800 -2885 40845 -2765
rect 40965 -2885 41010 -2765
rect 41130 -2885 41175 -2765
rect 41295 -2885 41350 -2765
rect 41470 -2885 41515 -2765
rect 41635 -2885 41680 -2765
rect 41800 -2885 41845 -2765
rect 41965 -2885 41975 -2765
rect 36475 -2930 41975 -2885
rect 36475 -3050 36485 -2930
rect 36605 -3050 36660 -2930
rect 36780 -3050 36825 -2930
rect 36945 -3050 36990 -2930
rect 37110 -3050 37155 -2930
rect 37275 -3050 37330 -2930
rect 37450 -3050 37495 -2930
rect 37615 -3050 37660 -2930
rect 37780 -3050 37825 -2930
rect 37945 -3050 38000 -2930
rect 38120 -3050 38165 -2930
rect 38285 -3050 38330 -2930
rect 38450 -3050 38495 -2930
rect 38615 -3050 38670 -2930
rect 38790 -3050 38835 -2930
rect 38955 -3050 39000 -2930
rect 39120 -3050 39165 -2930
rect 39285 -3050 39340 -2930
rect 39460 -3050 39505 -2930
rect 39625 -3050 39670 -2930
rect 39790 -3050 39835 -2930
rect 39955 -3050 40010 -2930
rect 40130 -3050 40175 -2930
rect 40295 -3050 40340 -2930
rect 40460 -3050 40505 -2930
rect 40625 -3050 40680 -2930
rect 40800 -3050 40845 -2930
rect 40965 -3050 41010 -2930
rect 41130 -3050 41175 -2930
rect 41295 -3050 41350 -2930
rect 41470 -3050 41515 -2930
rect 41635 -3050 41680 -2930
rect 41800 -3050 41845 -2930
rect 41965 -3050 41975 -2930
rect 36475 -3095 41975 -3050
rect 36475 -3215 36485 -3095
rect 36605 -3215 36660 -3095
rect 36780 -3215 36825 -3095
rect 36945 -3215 36990 -3095
rect 37110 -3215 37155 -3095
rect 37275 -3215 37330 -3095
rect 37450 -3215 37495 -3095
rect 37615 -3215 37660 -3095
rect 37780 -3215 37825 -3095
rect 37945 -3215 38000 -3095
rect 38120 -3215 38165 -3095
rect 38285 -3215 38330 -3095
rect 38450 -3215 38495 -3095
rect 38615 -3215 38670 -3095
rect 38790 -3215 38835 -3095
rect 38955 -3215 39000 -3095
rect 39120 -3215 39165 -3095
rect 39285 -3215 39340 -3095
rect 39460 -3215 39505 -3095
rect 39625 -3215 39670 -3095
rect 39790 -3215 39835 -3095
rect 39955 -3215 40010 -3095
rect 40130 -3215 40175 -3095
rect 40295 -3215 40340 -3095
rect 40460 -3215 40505 -3095
rect 40625 -3215 40680 -3095
rect 40800 -3215 40845 -3095
rect 40965 -3215 41010 -3095
rect 41130 -3215 41175 -3095
rect 41295 -3215 41350 -3095
rect 41470 -3215 41515 -3095
rect 41635 -3215 41680 -3095
rect 41800 -3215 41845 -3095
rect 41965 -3215 41975 -3095
rect 36475 -3270 41975 -3215
rect 36475 -3390 36485 -3270
rect 36605 -3390 36660 -3270
rect 36780 -3390 36825 -3270
rect 36945 -3390 36990 -3270
rect 37110 -3390 37155 -3270
rect 37275 -3390 37330 -3270
rect 37450 -3390 37495 -3270
rect 37615 -3390 37660 -3270
rect 37780 -3390 37825 -3270
rect 37945 -3390 38000 -3270
rect 38120 -3390 38165 -3270
rect 38285 -3390 38330 -3270
rect 38450 -3390 38495 -3270
rect 38615 -3390 38670 -3270
rect 38790 -3390 38835 -3270
rect 38955 -3390 39000 -3270
rect 39120 -3390 39165 -3270
rect 39285 -3390 39340 -3270
rect 39460 -3390 39505 -3270
rect 39625 -3390 39670 -3270
rect 39790 -3390 39835 -3270
rect 39955 -3390 40010 -3270
rect 40130 -3390 40175 -3270
rect 40295 -3390 40340 -3270
rect 40460 -3390 40505 -3270
rect 40625 -3390 40680 -3270
rect 40800 -3390 40845 -3270
rect 40965 -3390 41010 -3270
rect 41130 -3390 41175 -3270
rect 41295 -3390 41350 -3270
rect 41470 -3390 41515 -3270
rect 41635 -3390 41680 -3270
rect 41800 -3390 41845 -3270
rect 41965 -3390 41975 -3270
rect 36475 -3435 41975 -3390
rect 36475 -3555 36485 -3435
rect 36605 -3555 36660 -3435
rect 36780 -3555 36825 -3435
rect 36945 -3555 36990 -3435
rect 37110 -3555 37155 -3435
rect 37275 -3555 37330 -3435
rect 37450 -3555 37495 -3435
rect 37615 -3555 37660 -3435
rect 37780 -3555 37825 -3435
rect 37945 -3555 38000 -3435
rect 38120 -3555 38165 -3435
rect 38285 -3555 38330 -3435
rect 38450 -3555 38495 -3435
rect 38615 -3555 38670 -3435
rect 38790 -3555 38835 -3435
rect 38955 -3555 39000 -3435
rect 39120 -3555 39165 -3435
rect 39285 -3555 39340 -3435
rect 39460 -3555 39505 -3435
rect 39625 -3555 39670 -3435
rect 39790 -3555 39835 -3435
rect 39955 -3555 40010 -3435
rect 40130 -3555 40175 -3435
rect 40295 -3555 40340 -3435
rect 40460 -3555 40505 -3435
rect 40625 -3555 40680 -3435
rect 40800 -3555 40845 -3435
rect 40965 -3555 41010 -3435
rect 41130 -3555 41175 -3435
rect 41295 -3555 41350 -3435
rect 41470 -3555 41515 -3435
rect 41635 -3555 41680 -3435
rect 41800 -3555 41845 -3435
rect 41965 -3555 41975 -3435
rect 36475 -3600 41975 -3555
rect 36475 -3720 36485 -3600
rect 36605 -3720 36660 -3600
rect 36780 -3720 36825 -3600
rect 36945 -3720 36990 -3600
rect 37110 -3720 37155 -3600
rect 37275 -3720 37330 -3600
rect 37450 -3720 37495 -3600
rect 37615 -3720 37660 -3600
rect 37780 -3720 37825 -3600
rect 37945 -3720 38000 -3600
rect 38120 -3720 38165 -3600
rect 38285 -3720 38330 -3600
rect 38450 -3720 38495 -3600
rect 38615 -3720 38670 -3600
rect 38790 -3720 38835 -3600
rect 38955 -3720 39000 -3600
rect 39120 -3720 39165 -3600
rect 39285 -3720 39340 -3600
rect 39460 -3720 39505 -3600
rect 39625 -3720 39670 -3600
rect 39790 -3720 39835 -3600
rect 39955 -3720 40010 -3600
rect 40130 -3720 40175 -3600
rect 40295 -3720 40340 -3600
rect 40460 -3720 40505 -3600
rect 40625 -3720 40680 -3600
rect 40800 -3720 40845 -3600
rect 40965 -3720 41010 -3600
rect 41130 -3720 41175 -3600
rect 41295 -3720 41350 -3600
rect 41470 -3720 41515 -3600
rect 41635 -3720 41680 -3600
rect 41800 -3720 41845 -3600
rect 41965 -3720 41975 -3600
rect 36475 -3765 41975 -3720
rect 36475 -3885 36485 -3765
rect 36605 -3885 36660 -3765
rect 36780 -3885 36825 -3765
rect 36945 -3885 36990 -3765
rect 37110 -3885 37155 -3765
rect 37275 -3885 37330 -3765
rect 37450 -3885 37495 -3765
rect 37615 -3885 37660 -3765
rect 37780 -3885 37825 -3765
rect 37945 -3885 38000 -3765
rect 38120 -3885 38165 -3765
rect 38285 -3885 38330 -3765
rect 38450 -3885 38495 -3765
rect 38615 -3885 38670 -3765
rect 38790 -3885 38835 -3765
rect 38955 -3885 39000 -3765
rect 39120 -3885 39165 -3765
rect 39285 -3885 39340 -3765
rect 39460 -3885 39505 -3765
rect 39625 -3885 39670 -3765
rect 39790 -3885 39835 -3765
rect 39955 -3885 40010 -3765
rect 40130 -3885 40175 -3765
rect 40295 -3885 40340 -3765
rect 40460 -3885 40505 -3765
rect 40625 -3885 40680 -3765
rect 40800 -3885 40845 -3765
rect 40965 -3885 41010 -3765
rect 41130 -3885 41175 -3765
rect 41295 -3885 41350 -3765
rect 41470 -3885 41515 -3765
rect 41635 -3885 41680 -3765
rect 41800 -3885 41845 -3765
rect 41965 -3885 41975 -3765
rect 36475 -3940 41975 -3885
rect 36475 -4060 36485 -3940
rect 36605 -4060 36660 -3940
rect 36780 -4060 36825 -3940
rect 36945 -4060 36990 -3940
rect 37110 -4060 37155 -3940
rect 37275 -4060 37330 -3940
rect 37450 -4060 37495 -3940
rect 37615 -4060 37660 -3940
rect 37780 -4060 37825 -3940
rect 37945 -4060 38000 -3940
rect 38120 -4060 38165 -3940
rect 38285 -4060 38330 -3940
rect 38450 -4060 38495 -3940
rect 38615 -4060 38670 -3940
rect 38790 -4060 38835 -3940
rect 38955 -4060 39000 -3940
rect 39120 -4060 39165 -3940
rect 39285 -4060 39340 -3940
rect 39460 -4060 39505 -3940
rect 39625 -4060 39670 -3940
rect 39790 -4060 39835 -3940
rect 39955 -4060 40010 -3940
rect 40130 -4060 40175 -3940
rect 40295 -4060 40340 -3940
rect 40460 -4060 40505 -3940
rect 40625 -4060 40680 -3940
rect 40800 -4060 40845 -3940
rect 40965 -4060 41010 -3940
rect 41130 -4060 41175 -3940
rect 41295 -4060 41350 -3940
rect 41470 -4060 41515 -3940
rect 41635 -4060 41680 -3940
rect 41800 -4060 41845 -3940
rect 41965 -4060 41975 -3940
rect 36475 -4070 41975 -4060
rect 42165 1420 47665 1430
rect 42165 1300 42175 1420
rect 42295 1300 42350 1420
rect 42470 1300 42515 1420
rect 42635 1300 42680 1420
rect 42800 1300 42845 1420
rect 42965 1300 43020 1420
rect 43140 1300 43185 1420
rect 43305 1300 43350 1420
rect 43470 1300 43515 1420
rect 43635 1300 43690 1420
rect 43810 1300 43855 1420
rect 43975 1300 44020 1420
rect 44140 1300 44185 1420
rect 44305 1300 44360 1420
rect 44480 1300 44525 1420
rect 44645 1300 44690 1420
rect 44810 1300 44855 1420
rect 44975 1300 45030 1420
rect 45150 1300 45195 1420
rect 45315 1300 45360 1420
rect 45480 1300 45525 1420
rect 45645 1300 45700 1420
rect 45820 1300 45865 1420
rect 45985 1300 46030 1420
rect 46150 1300 46195 1420
rect 46315 1300 46370 1420
rect 46490 1300 46535 1420
rect 46655 1300 46700 1420
rect 46820 1300 46865 1420
rect 46985 1300 47040 1420
rect 47160 1300 47205 1420
rect 47325 1300 47370 1420
rect 47490 1300 47535 1420
rect 47655 1300 47665 1420
rect 42165 1255 47665 1300
rect 42165 1135 42175 1255
rect 42295 1135 42350 1255
rect 42470 1135 42515 1255
rect 42635 1135 42680 1255
rect 42800 1135 42845 1255
rect 42965 1135 43020 1255
rect 43140 1135 43185 1255
rect 43305 1135 43350 1255
rect 43470 1135 43515 1255
rect 43635 1135 43690 1255
rect 43810 1135 43855 1255
rect 43975 1135 44020 1255
rect 44140 1135 44185 1255
rect 44305 1135 44360 1255
rect 44480 1135 44525 1255
rect 44645 1135 44690 1255
rect 44810 1135 44855 1255
rect 44975 1135 45030 1255
rect 45150 1135 45195 1255
rect 45315 1135 45360 1255
rect 45480 1135 45525 1255
rect 45645 1135 45700 1255
rect 45820 1135 45865 1255
rect 45985 1135 46030 1255
rect 46150 1135 46195 1255
rect 46315 1135 46370 1255
rect 46490 1135 46535 1255
rect 46655 1135 46700 1255
rect 46820 1135 46865 1255
rect 46985 1135 47040 1255
rect 47160 1135 47205 1255
rect 47325 1135 47370 1255
rect 47490 1135 47535 1255
rect 47655 1135 47665 1255
rect 42165 1090 47665 1135
rect 42165 970 42175 1090
rect 42295 970 42350 1090
rect 42470 970 42515 1090
rect 42635 970 42680 1090
rect 42800 970 42845 1090
rect 42965 970 43020 1090
rect 43140 970 43185 1090
rect 43305 970 43350 1090
rect 43470 970 43515 1090
rect 43635 970 43690 1090
rect 43810 970 43855 1090
rect 43975 970 44020 1090
rect 44140 970 44185 1090
rect 44305 970 44360 1090
rect 44480 970 44525 1090
rect 44645 970 44690 1090
rect 44810 970 44855 1090
rect 44975 970 45030 1090
rect 45150 970 45195 1090
rect 45315 970 45360 1090
rect 45480 970 45525 1090
rect 45645 970 45700 1090
rect 45820 970 45865 1090
rect 45985 970 46030 1090
rect 46150 970 46195 1090
rect 46315 970 46370 1090
rect 46490 970 46535 1090
rect 46655 970 46700 1090
rect 46820 970 46865 1090
rect 46985 970 47040 1090
rect 47160 970 47205 1090
rect 47325 970 47370 1090
rect 47490 970 47535 1090
rect 47655 970 47665 1090
rect 42165 925 47665 970
rect 42165 805 42175 925
rect 42295 805 42350 925
rect 42470 805 42515 925
rect 42635 805 42680 925
rect 42800 805 42845 925
rect 42965 805 43020 925
rect 43140 805 43185 925
rect 43305 805 43350 925
rect 43470 805 43515 925
rect 43635 805 43690 925
rect 43810 805 43855 925
rect 43975 805 44020 925
rect 44140 805 44185 925
rect 44305 805 44360 925
rect 44480 805 44525 925
rect 44645 805 44690 925
rect 44810 805 44855 925
rect 44975 805 45030 925
rect 45150 805 45195 925
rect 45315 805 45360 925
rect 45480 805 45525 925
rect 45645 805 45700 925
rect 45820 805 45865 925
rect 45985 805 46030 925
rect 46150 805 46195 925
rect 46315 805 46370 925
rect 46490 805 46535 925
rect 46655 805 46700 925
rect 46820 805 46865 925
rect 46985 805 47040 925
rect 47160 805 47205 925
rect 47325 805 47370 925
rect 47490 805 47535 925
rect 47655 805 47665 925
rect 42165 750 47665 805
rect 42165 630 42175 750
rect 42295 630 42350 750
rect 42470 630 42515 750
rect 42635 630 42680 750
rect 42800 630 42845 750
rect 42965 630 43020 750
rect 43140 630 43185 750
rect 43305 630 43350 750
rect 43470 630 43515 750
rect 43635 630 43690 750
rect 43810 630 43855 750
rect 43975 630 44020 750
rect 44140 630 44185 750
rect 44305 630 44360 750
rect 44480 630 44525 750
rect 44645 630 44690 750
rect 44810 630 44855 750
rect 44975 630 45030 750
rect 45150 630 45195 750
rect 45315 630 45360 750
rect 45480 630 45525 750
rect 45645 630 45700 750
rect 45820 630 45865 750
rect 45985 630 46030 750
rect 46150 630 46195 750
rect 46315 630 46370 750
rect 46490 630 46535 750
rect 46655 630 46700 750
rect 46820 630 46865 750
rect 46985 630 47040 750
rect 47160 630 47205 750
rect 47325 630 47370 750
rect 47490 630 47535 750
rect 47655 630 47665 750
rect 42165 585 47665 630
rect 42165 465 42175 585
rect 42295 465 42350 585
rect 42470 465 42515 585
rect 42635 465 42680 585
rect 42800 465 42845 585
rect 42965 465 43020 585
rect 43140 465 43185 585
rect 43305 465 43350 585
rect 43470 465 43515 585
rect 43635 465 43690 585
rect 43810 465 43855 585
rect 43975 465 44020 585
rect 44140 465 44185 585
rect 44305 465 44360 585
rect 44480 465 44525 585
rect 44645 465 44690 585
rect 44810 465 44855 585
rect 44975 465 45030 585
rect 45150 465 45195 585
rect 45315 465 45360 585
rect 45480 465 45525 585
rect 45645 465 45700 585
rect 45820 465 45865 585
rect 45985 465 46030 585
rect 46150 465 46195 585
rect 46315 465 46370 585
rect 46490 465 46535 585
rect 46655 465 46700 585
rect 46820 465 46865 585
rect 46985 465 47040 585
rect 47160 465 47205 585
rect 47325 465 47370 585
rect 47490 465 47535 585
rect 47655 465 47665 585
rect 42165 420 47665 465
rect 42165 300 42175 420
rect 42295 300 42350 420
rect 42470 300 42515 420
rect 42635 300 42680 420
rect 42800 300 42845 420
rect 42965 300 43020 420
rect 43140 300 43185 420
rect 43305 300 43350 420
rect 43470 300 43515 420
rect 43635 300 43690 420
rect 43810 300 43855 420
rect 43975 300 44020 420
rect 44140 300 44185 420
rect 44305 300 44360 420
rect 44480 300 44525 420
rect 44645 300 44690 420
rect 44810 300 44855 420
rect 44975 300 45030 420
rect 45150 300 45195 420
rect 45315 300 45360 420
rect 45480 300 45525 420
rect 45645 300 45700 420
rect 45820 300 45865 420
rect 45985 300 46030 420
rect 46150 300 46195 420
rect 46315 300 46370 420
rect 46490 300 46535 420
rect 46655 300 46700 420
rect 46820 300 46865 420
rect 46985 300 47040 420
rect 47160 300 47205 420
rect 47325 300 47370 420
rect 47490 300 47535 420
rect 47655 300 47665 420
rect 42165 255 47665 300
rect 42165 135 42175 255
rect 42295 135 42350 255
rect 42470 135 42515 255
rect 42635 135 42680 255
rect 42800 135 42845 255
rect 42965 135 43020 255
rect 43140 135 43185 255
rect 43305 135 43350 255
rect 43470 135 43515 255
rect 43635 135 43690 255
rect 43810 135 43855 255
rect 43975 135 44020 255
rect 44140 135 44185 255
rect 44305 135 44360 255
rect 44480 135 44525 255
rect 44645 135 44690 255
rect 44810 135 44855 255
rect 44975 135 45030 255
rect 45150 135 45195 255
rect 45315 135 45360 255
rect 45480 135 45525 255
rect 45645 135 45700 255
rect 45820 135 45865 255
rect 45985 135 46030 255
rect 46150 135 46195 255
rect 46315 135 46370 255
rect 46490 135 46535 255
rect 46655 135 46700 255
rect 46820 135 46865 255
rect 46985 135 47040 255
rect 47160 135 47205 255
rect 47325 135 47370 255
rect 47490 135 47535 255
rect 47655 135 47665 255
rect 42165 80 47665 135
rect 42165 -40 42175 80
rect 42295 -40 42350 80
rect 42470 -40 42515 80
rect 42635 -40 42680 80
rect 42800 -40 42845 80
rect 42965 -40 43020 80
rect 43140 -40 43185 80
rect 43305 -40 43350 80
rect 43470 -40 43515 80
rect 43635 -40 43690 80
rect 43810 -40 43855 80
rect 43975 -40 44020 80
rect 44140 -40 44185 80
rect 44305 -40 44360 80
rect 44480 -40 44525 80
rect 44645 -40 44690 80
rect 44810 -40 44855 80
rect 44975 -40 45030 80
rect 45150 -40 45195 80
rect 45315 -40 45360 80
rect 45480 -40 45525 80
rect 45645 -40 45700 80
rect 45820 -40 45865 80
rect 45985 -40 46030 80
rect 46150 -40 46195 80
rect 46315 -40 46370 80
rect 46490 -40 46535 80
rect 46655 -40 46700 80
rect 46820 -40 46865 80
rect 46985 -40 47040 80
rect 47160 -40 47205 80
rect 47325 -40 47370 80
rect 47490 -40 47535 80
rect 47655 -40 47665 80
rect 42165 -85 47665 -40
rect 42165 -205 42175 -85
rect 42295 -205 42350 -85
rect 42470 -205 42515 -85
rect 42635 -205 42680 -85
rect 42800 -205 42845 -85
rect 42965 -205 43020 -85
rect 43140 -205 43185 -85
rect 43305 -205 43350 -85
rect 43470 -205 43515 -85
rect 43635 -205 43690 -85
rect 43810 -205 43855 -85
rect 43975 -205 44020 -85
rect 44140 -205 44185 -85
rect 44305 -205 44360 -85
rect 44480 -205 44525 -85
rect 44645 -205 44690 -85
rect 44810 -205 44855 -85
rect 44975 -205 45030 -85
rect 45150 -205 45195 -85
rect 45315 -205 45360 -85
rect 45480 -205 45525 -85
rect 45645 -205 45700 -85
rect 45820 -205 45865 -85
rect 45985 -205 46030 -85
rect 46150 -205 46195 -85
rect 46315 -205 46370 -85
rect 46490 -205 46535 -85
rect 46655 -205 46700 -85
rect 46820 -205 46865 -85
rect 46985 -205 47040 -85
rect 47160 -205 47205 -85
rect 47325 -205 47370 -85
rect 47490 -205 47535 -85
rect 47655 -205 47665 -85
rect 42165 -250 47665 -205
rect 42165 -370 42175 -250
rect 42295 -370 42350 -250
rect 42470 -370 42515 -250
rect 42635 -370 42680 -250
rect 42800 -370 42845 -250
rect 42965 -370 43020 -250
rect 43140 -370 43185 -250
rect 43305 -370 43350 -250
rect 43470 -370 43515 -250
rect 43635 -370 43690 -250
rect 43810 -370 43855 -250
rect 43975 -370 44020 -250
rect 44140 -370 44185 -250
rect 44305 -370 44360 -250
rect 44480 -370 44525 -250
rect 44645 -370 44690 -250
rect 44810 -370 44855 -250
rect 44975 -370 45030 -250
rect 45150 -370 45195 -250
rect 45315 -370 45360 -250
rect 45480 -370 45525 -250
rect 45645 -370 45700 -250
rect 45820 -370 45865 -250
rect 45985 -370 46030 -250
rect 46150 -370 46195 -250
rect 46315 -370 46370 -250
rect 46490 -370 46535 -250
rect 46655 -370 46700 -250
rect 46820 -370 46865 -250
rect 46985 -370 47040 -250
rect 47160 -370 47205 -250
rect 47325 -370 47370 -250
rect 47490 -370 47535 -250
rect 47655 -370 47665 -250
rect 42165 -415 47665 -370
rect 42165 -535 42175 -415
rect 42295 -535 42350 -415
rect 42470 -535 42515 -415
rect 42635 -535 42680 -415
rect 42800 -535 42845 -415
rect 42965 -535 43020 -415
rect 43140 -535 43185 -415
rect 43305 -535 43350 -415
rect 43470 -535 43515 -415
rect 43635 -535 43690 -415
rect 43810 -535 43855 -415
rect 43975 -535 44020 -415
rect 44140 -535 44185 -415
rect 44305 -535 44360 -415
rect 44480 -535 44525 -415
rect 44645 -535 44690 -415
rect 44810 -535 44855 -415
rect 44975 -535 45030 -415
rect 45150 -535 45195 -415
rect 45315 -535 45360 -415
rect 45480 -535 45525 -415
rect 45645 -535 45700 -415
rect 45820 -535 45865 -415
rect 45985 -535 46030 -415
rect 46150 -535 46195 -415
rect 46315 -535 46370 -415
rect 46490 -535 46535 -415
rect 46655 -535 46700 -415
rect 46820 -535 46865 -415
rect 46985 -535 47040 -415
rect 47160 -535 47205 -415
rect 47325 -535 47370 -415
rect 47490 -535 47535 -415
rect 47655 -535 47665 -415
rect 42165 -590 47665 -535
rect 42165 -710 42175 -590
rect 42295 -710 42350 -590
rect 42470 -710 42515 -590
rect 42635 -710 42680 -590
rect 42800 -710 42845 -590
rect 42965 -710 43020 -590
rect 43140 -710 43185 -590
rect 43305 -710 43350 -590
rect 43470 -710 43515 -590
rect 43635 -710 43690 -590
rect 43810 -710 43855 -590
rect 43975 -710 44020 -590
rect 44140 -710 44185 -590
rect 44305 -710 44360 -590
rect 44480 -710 44525 -590
rect 44645 -710 44690 -590
rect 44810 -710 44855 -590
rect 44975 -710 45030 -590
rect 45150 -710 45195 -590
rect 45315 -710 45360 -590
rect 45480 -710 45525 -590
rect 45645 -710 45700 -590
rect 45820 -710 45865 -590
rect 45985 -710 46030 -590
rect 46150 -710 46195 -590
rect 46315 -710 46370 -590
rect 46490 -710 46535 -590
rect 46655 -710 46700 -590
rect 46820 -710 46865 -590
rect 46985 -710 47040 -590
rect 47160 -710 47205 -590
rect 47325 -710 47370 -590
rect 47490 -710 47535 -590
rect 47655 -710 47665 -590
rect 42165 -755 47665 -710
rect 42165 -875 42175 -755
rect 42295 -875 42350 -755
rect 42470 -875 42515 -755
rect 42635 -875 42680 -755
rect 42800 -875 42845 -755
rect 42965 -875 43020 -755
rect 43140 -875 43185 -755
rect 43305 -875 43350 -755
rect 43470 -875 43515 -755
rect 43635 -875 43690 -755
rect 43810 -875 43855 -755
rect 43975 -875 44020 -755
rect 44140 -875 44185 -755
rect 44305 -875 44360 -755
rect 44480 -875 44525 -755
rect 44645 -875 44690 -755
rect 44810 -875 44855 -755
rect 44975 -875 45030 -755
rect 45150 -875 45195 -755
rect 45315 -875 45360 -755
rect 45480 -875 45525 -755
rect 45645 -875 45700 -755
rect 45820 -875 45865 -755
rect 45985 -875 46030 -755
rect 46150 -875 46195 -755
rect 46315 -875 46370 -755
rect 46490 -875 46535 -755
rect 46655 -875 46700 -755
rect 46820 -875 46865 -755
rect 46985 -875 47040 -755
rect 47160 -875 47205 -755
rect 47325 -875 47370 -755
rect 47490 -875 47535 -755
rect 47655 -875 47665 -755
rect 42165 -920 47665 -875
rect 42165 -1040 42175 -920
rect 42295 -1040 42350 -920
rect 42470 -1040 42515 -920
rect 42635 -1040 42680 -920
rect 42800 -1040 42845 -920
rect 42965 -1040 43020 -920
rect 43140 -1040 43185 -920
rect 43305 -1040 43350 -920
rect 43470 -1040 43515 -920
rect 43635 -1040 43690 -920
rect 43810 -1040 43855 -920
rect 43975 -1040 44020 -920
rect 44140 -1040 44185 -920
rect 44305 -1040 44360 -920
rect 44480 -1040 44525 -920
rect 44645 -1040 44690 -920
rect 44810 -1040 44855 -920
rect 44975 -1040 45030 -920
rect 45150 -1040 45195 -920
rect 45315 -1040 45360 -920
rect 45480 -1040 45525 -920
rect 45645 -1040 45700 -920
rect 45820 -1040 45865 -920
rect 45985 -1040 46030 -920
rect 46150 -1040 46195 -920
rect 46315 -1040 46370 -920
rect 46490 -1040 46535 -920
rect 46655 -1040 46700 -920
rect 46820 -1040 46865 -920
rect 46985 -1040 47040 -920
rect 47160 -1040 47205 -920
rect 47325 -1040 47370 -920
rect 47490 -1040 47535 -920
rect 47655 -1040 47665 -920
rect 42165 -1085 47665 -1040
rect 42165 -1205 42175 -1085
rect 42295 -1205 42350 -1085
rect 42470 -1205 42515 -1085
rect 42635 -1205 42680 -1085
rect 42800 -1205 42845 -1085
rect 42965 -1205 43020 -1085
rect 43140 -1205 43185 -1085
rect 43305 -1205 43350 -1085
rect 43470 -1205 43515 -1085
rect 43635 -1205 43690 -1085
rect 43810 -1205 43855 -1085
rect 43975 -1205 44020 -1085
rect 44140 -1205 44185 -1085
rect 44305 -1205 44360 -1085
rect 44480 -1205 44525 -1085
rect 44645 -1205 44690 -1085
rect 44810 -1205 44855 -1085
rect 44975 -1205 45030 -1085
rect 45150 -1205 45195 -1085
rect 45315 -1205 45360 -1085
rect 45480 -1205 45525 -1085
rect 45645 -1205 45700 -1085
rect 45820 -1205 45865 -1085
rect 45985 -1205 46030 -1085
rect 46150 -1205 46195 -1085
rect 46315 -1205 46370 -1085
rect 46490 -1205 46535 -1085
rect 46655 -1205 46700 -1085
rect 46820 -1205 46865 -1085
rect 46985 -1205 47040 -1085
rect 47160 -1205 47205 -1085
rect 47325 -1205 47370 -1085
rect 47490 -1205 47535 -1085
rect 47655 -1205 47665 -1085
rect 42165 -1260 47665 -1205
rect 42165 -1380 42175 -1260
rect 42295 -1380 42350 -1260
rect 42470 -1380 42515 -1260
rect 42635 -1380 42680 -1260
rect 42800 -1380 42845 -1260
rect 42965 -1380 43020 -1260
rect 43140 -1380 43185 -1260
rect 43305 -1380 43350 -1260
rect 43470 -1380 43515 -1260
rect 43635 -1380 43690 -1260
rect 43810 -1380 43855 -1260
rect 43975 -1380 44020 -1260
rect 44140 -1380 44185 -1260
rect 44305 -1380 44360 -1260
rect 44480 -1380 44525 -1260
rect 44645 -1380 44690 -1260
rect 44810 -1380 44855 -1260
rect 44975 -1380 45030 -1260
rect 45150 -1380 45195 -1260
rect 45315 -1380 45360 -1260
rect 45480 -1380 45525 -1260
rect 45645 -1380 45700 -1260
rect 45820 -1380 45865 -1260
rect 45985 -1380 46030 -1260
rect 46150 -1380 46195 -1260
rect 46315 -1380 46370 -1260
rect 46490 -1380 46535 -1260
rect 46655 -1380 46700 -1260
rect 46820 -1380 46865 -1260
rect 46985 -1380 47040 -1260
rect 47160 -1380 47205 -1260
rect 47325 -1380 47370 -1260
rect 47490 -1380 47535 -1260
rect 47655 -1380 47665 -1260
rect 42165 -1425 47665 -1380
rect 42165 -1545 42175 -1425
rect 42295 -1545 42350 -1425
rect 42470 -1545 42515 -1425
rect 42635 -1545 42680 -1425
rect 42800 -1545 42845 -1425
rect 42965 -1545 43020 -1425
rect 43140 -1545 43185 -1425
rect 43305 -1545 43350 -1425
rect 43470 -1545 43515 -1425
rect 43635 -1545 43690 -1425
rect 43810 -1545 43855 -1425
rect 43975 -1545 44020 -1425
rect 44140 -1545 44185 -1425
rect 44305 -1545 44360 -1425
rect 44480 -1545 44525 -1425
rect 44645 -1545 44690 -1425
rect 44810 -1545 44855 -1425
rect 44975 -1545 45030 -1425
rect 45150 -1545 45195 -1425
rect 45315 -1545 45360 -1425
rect 45480 -1545 45525 -1425
rect 45645 -1545 45700 -1425
rect 45820 -1545 45865 -1425
rect 45985 -1545 46030 -1425
rect 46150 -1545 46195 -1425
rect 46315 -1545 46370 -1425
rect 46490 -1545 46535 -1425
rect 46655 -1545 46700 -1425
rect 46820 -1545 46865 -1425
rect 46985 -1545 47040 -1425
rect 47160 -1545 47205 -1425
rect 47325 -1545 47370 -1425
rect 47490 -1545 47535 -1425
rect 47655 -1545 47665 -1425
rect 42165 -1590 47665 -1545
rect 42165 -1710 42175 -1590
rect 42295 -1710 42350 -1590
rect 42470 -1710 42515 -1590
rect 42635 -1710 42680 -1590
rect 42800 -1710 42845 -1590
rect 42965 -1710 43020 -1590
rect 43140 -1710 43185 -1590
rect 43305 -1710 43350 -1590
rect 43470 -1710 43515 -1590
rect 43635 -1710 43690 -1590
rect 43810 -1710 43855 -1590
rect 43975 -1710 44020 -1590
rect 44140 -1710 44185 -1590
rect 44305 -1710 44360 -1590
rect 44480 -1710 44525 -1590
rect 44645 -1710 44690 -1590
rect 44810 -1710 44855 -1590
rect 44975 -1710 45030 -1590
rect 45150 -1710 45195 -1590
rect 45315 -1710 45360 -1590
rect 45480 -1710 45525 -1590
rect 45645 -1710 45700 -1590
rect 45820 -1710 45865 -1590
rect 45985 -1710 46030 -1590
rect 46150 -1710 46195 -1590
rect 46315 -1710 46370 -1590
rect 46490 -1710 46535 -1590
rect 46655 -1710 46700 -1590
rect 46820 -1710 46865 -1590
rect 46985 -1710 47040 -1590
rect 47160 -1710 47205 -1590
rect 47325 -1710 47370 -1590
rect 47490 -1710 47535 -1590
rect 47655 -1710 47665 -1590
rect 42165 -1755 47665 -1710
rect 42165 -1875 42175 -1755
rect 42295 -1875 42350 -1755
rect 42470 -1875 42515 -1755
rect 42635 -1875 42680 -1755
rect 42800 -1875 42845 -1755
rect 42965 -1875 43020 -1755
rect 43140 -1875 43185 -1755
rect 43305 -1875 43350 -1755
rect 43470 -1875 43515 -1755
rect 43635 -1875 43690 -1755
rect 43810 -1875 43855 -1755
rect 43975 -1875 44020 -1755
rect 44140 -1875 44185 -1755
rect 44305 -1875 44360 -1755
rect 44480 -1875 44525 -1755
rect 44645 -1875 44690 -1755
rect 44810 -1875 44855 -1755
rect 44975 -1875 45030 -1755
rect 45150 -1875 45195 -1755
rect 45315 -1875 45360 -1755
rect 45480 -1875 45525 -1755
rect 45645 -1875 45700 -1755
rect 45820 -1875 45865 -1755
rect 45985 -1875 46030 -1755
rect 46150 -1875 46195 -1755
rect 46315 -1875 46370 -1755
rect 46490 -1875 46535 -1755
rect 46655 -1875 46700 -1755
rect 46820 -1875 46865 -1755
rect 46985 -1875 47040 -1755
rect 47160 -1875 47205 -1755
rect 47325 -1875 47370 -1755
rect 47490 -1875 47535 -1755
rect 47655 -1875 47665 -1755
rect 42165 -1930 47665 -1875
rect 42165 -2050 42175 -1930
rect 42295 -2050 42350 -1930
rect 42470 -2050 42515 -1930
rect 42635 -2050 42680 -1930
rect 42800 -2050 42845 -1930
rect 42965 -2050 43020 -1930
rect 43140 -2050 43185 -1930
rect 43305 -2050 43350 -1930
rect 43470 -2050 43515 -1930
rect 43635 -2050 43690 -1930
rect 43810 -2050 43855 -1930
rect 43975 -2050 44020 -1930
rect 44140 -2050 44185 -1930
rect 44305 -2050 44360 -1930
rect 44480 -2050 44525 -1930
rect 44645 -2050 44690 -1930
rect 44810 -2050 44855 -1930
rect 44975 -2050 45030 -1930
rect 45150 -2050 45195 -1930
rect 45315 -2050 45360 -1930
rect 45480 -2050 45525 -1930
rect 45645 -2050 45700 -1930
rect 45820 -2050 45865 -1930
rect 45985 -2050 46030 -1930
rect 46150 -2050 46195 -1930
rect 46315 -2050 46370 -1930
rect 46490 -2050 46535 -1930
rect 46655 -2050 46700 -1930
rect 46820 -2050 46865 -1930
rect 46985 -2050 47040 -1930
rect 47160 -2050 47205 -1930
rect 47325 -2050 47370 -1930
rect 47490 -2050 47535 -1930
rect 47655 -2050 47665 -1930
rect 42165 -2095 47665 -2050
rect 42165 -2215 42175 -2095
rect 42295 -2215 42350 -2095
rect 42470 -2215 42515 -2095
rect 42635 -2215 42680 -2095
rect 42800 -2215 42845 -2095
rect 42965 -2215 43020 -2095
rect 43140 -2215 43185 -2095
rect 43305 -2215 43350 -2095
rect 43470 -2215 43515 -2095
rect 43635 -2215 43690 -2095
rect 43810 -2215 43855 -2095
rect 43975 -2215 44020 -2095
rect 44140 -2215 44185 -2095
rect 44305 -2215 44360 -2095
rect 44480 -2215 44525 -2095
rect 44645 -2215 44690 -2095
rect 44810 -2215 44855 -2095
rect 44975 -2215 45030 -2095
rect 45150 -2215 45195 -2095
rect 45315 -2215 45360 -2095
rect 45480 -2215 45525 -2095
rect 45645 -2215 45700 -2095
rect 45820 -2215 45865 -2095
rect 45985 -2215 46030 -2095
rect 46150 -2215 46195 -2095
rect 46315 -2215 46370 -2095
rect 46490 -2215 46535 -2095
rect 46655 -2215 46700 -2095
rect 46820 -2215 46865 -2095
rect 46985 -2215 47040 -2095
rect 47160 -2215 47205 -2095
rect 47325 -2215 47370 -2095
rect 47490 -2215 47535 -2095
rect 47655 -2215 47665 -2095
rect 42165 -2260 47665 -2215
rect 42165 -2380 42175 -2260
rect 42295 -2380 42350 -2260
rect 42470 -2380 42515 -2260
rect 42635 -2380 42680 -2260
rect 42800 -2380 42845 -2260
rect 42965 -2380 43020 -2260
rect 43140 -2380 43185 -2260
rect 43305 -2380 43350 -2260
rect 43470 -2380 43515 -2260
rect 43635 -2380 43690 -2260
rect 43810 -2380 43855 -2260
rect 43975 -2380 44020 -2260
rect 44140 -2380 44185 -2260
rect 44305 -2380 44360 -2260
rect 44480 -2380 44525 -2260
rect 44645 -2380 44690 -2260
rect 44810 -2380 44855 -2260
rect 44975 -2380 45030 -2260
rect 45150 -2380 45195 -2260
rect 45315 -2380 45360 -2260
rect 45480 -2380 45525 -2260
rect 45645 -2380 45700 -2260
rect 45820 -2380 45865 -2260
rect 45985 -2380 46030 -2260
rect 46150 -2380 46195 -2260
rect 46315 -2380 46370 -2260
rect 46490 -2380 46535 -2260
rect 46655 -2380 46700 -2260
rect 46820 -2380 46865 -2260
rect 46985 -2380 47040 -2260
rect 47160 -2380 47205 -2260
rect 47325 -2380 47370 -2260
rect 47490 -2380 47535 -2260
rect 47655 -2380 47665 -2260
rect 42165 -2425 47665 -2380
rect 42165 -2545 42175 -2425
rect 42295 -2545 42350 -2425
rect 42470 -2545 42515 -2425
rect 42635 -2545 42680 -2425
rect 42800 -2545 42845 -2425
rect 42965 -2545 43020 -2425
rect 43140 -2545 43185 -2425
rect 43305 -2545 43350 -2425
rect 43470 -2545 43515 -2425
rect 43635 -2545 43690 -2425
rect 43810 -2545 43855 -2425
rect 43975 -2545 44020 -2425
rect 44140 -2545 44185 -2425
rect 44305 -2545 44360 -2425
rect 44480 -2545 44525 -2425
rect 44645 -2545 44690 -2425
rect 44810 -2545 44855 -2425
rect 44975 -2545 45030 -2425
rect 45150 -2545 45195 -2425
rect 45315 -2545 45360 -2425
rect 45480 -2545 45525 -2425
rect 45645 -2545 45700 -2425
rect 45820 -2545 45865 -2425
rect 45985 -2545 46030 -2425
rect 46150 -2545 46195 -2425
rect 46315 -2545 46370 -2425
rect 46490 -2545 46535 -2425
rect 46655 -2545 46700 -2425
rect 46820 -2545 46865 -2425
rect 46985 -2545 47040 -2425
rect 47160 -2545 47205 -2425
rect 47325 -2545 47370 -2425
rect 47490 -2545 47535 -2425
rect 47655 -2545 47665 -2425
rect 42165 -2600 47665 -2545
rect 42165 -2720 42175 -2600
rect 42295 -2720 42350 -2600
rect 42470 -2720 42515 -2600
rect 42635 -2720 42680 -2600
rect 42800 -2720 42845 -2600
rect 42965 -2720 43020 -2600
rect 43140 -2720 43185 -2600
rect 43305 -2720 43350 -2600
rect 43470 -2720 43515 -2600
rect 43635 -2720 43690 -2600
rect 43810 -2720 43855 -2600
rect 43975 -2720 44020 -2600
rect 44140 -2720 44185 -2600
rect 44305 -2720 44360 -2600
rect 44480 -2720 44525 -2600
rect 44645 -2720 44690 -2600
rect 44810 -2720 44855 -2600
rect 44975 -2720 45030 -2600
rect 45150 -2720 45195 -2600
rect 45315 -2720 45360 -2600
rect 45480 -2720 45525 -2600
rect 45645 -2720 45700 -2600
rect 45820 -2720 45865 -2600
rect 45985 -2720 46030 -2600
rect 46150 -2720 46195 -2600
rect 46315 -2720 46370 -2600
rect 46490 -2720 46535 -2600
rect 46655 -2720 46700 -2600
rect 46820 -2720 46865 -2600
rect 46985 -2720 47040 -2600
rect 47160 -2720 47205 -2600
rect 47325 -2720 47370 -2600
rect 47490 -2720 47535 -2600
rect 47655 -2720 47665 -2600
rect 42165 -2765 47665 -2720
rect 42165 -2885 42175 -2765
rect 42295 -2885 42350 -2765
rect 42470 -2885 42515 -2765
rect 42635 -2885 42680 -2765
rect 42800 -2885 42845 -2765
rect 42965 -2885 43020 -2765
rect 43140 -2885 43185 -2765
rect 43305 -2885 43350 -2765
rect 43470 -2885 43515 -2765
rect 43635 -2885 43690 -2765
rect 43810 -2885 43855 -2765
rect 43975 -2885 44020 -2765
rect 44140 -2885 44185 -2765
rect 44305 -2885 44360 -2765
rect 44480 -2885 44525 -2765
rect 44645 -2885 44690 -2765
rect 44810 -2885 44855 -2765
rect 44975 -2885 45030 -2765
rect 45150 -2885 45195 -2765
rect 45315 -2885 45360 -2765
rect 45480 -2885 45525 -2765
rect 45645 -2885 45700 -2765
rect 45820 -2885 45865 -2765
rect 45985 -2885 46030 -2765
rect 46150 -2885 46195 -2765
rect 46315 -2885 46370 -2765
rect 46490 -2885 46535 -2765
rect 46655 -2885 46700 -2765
rect 46820 -2885 46865 -2765
rect 46985 -2885 47040 -2765
rect 47160 -2885 47205 -2765
rect 47325 -2885 47370 -2765
rect 47490 -2885 47535 -2765
rect 47655 -2885 47665 -2765
rect 42165 -2930 47665 -2885
rect 42165 -3050 42175 -2930
rect 42295 -3050 42350 -2930
rect 42470 -3050 42515 -2930
rect 42635 -3050 42680 -2930
rect 42800 -3050 42845 -2930
rect 42965 -3050 43020 -2930
rect 43140 -3050 43185 -2930
rect 43305 -3050 43350 -2930
rect 43470 -3050 43515 -2930
rect 43635 -3050 43690 -2930
rect 43810 -3050 43855 -2930
rect 43975 -3050 44020 -2930
rect 44140 -3050 44185 -2930
rect 44305 -3050 44360 -2930
rect 44480 -3050 44525 -2930
rect 44645 -3050 44690 -2930
rect 44810 -3050 44855 -2930
rect 44975 -3050 45030 -2930
rect 45150 -3050 45195 -2930
rect 45315 -3050 45360 -2930
rect 45480 -3050 45525 -2930
rect 45645 -3050 45700 -2930
rect 45820 -3050 45865 -2930
rect 45985 -3050 46030 -2930
rect 46150 -3050 46195 -2930
rect 46315 -3050 46370 -2930
rect 46490 -3050 46535 -2930
rect 46655 -3050 46700 -2930
rect 46820 -3050 46865 -2930
rect 46985 -3050 47040 -2930
rect 47160 -3050 47205 -2930
rect 47325 -3050 47370 -2930
rect 47490 -3050 47535 -2930
rect 47655 -3050 47665 -2930
rect 42165 -3095 47665 -3050
rect 42165 -3215 42175 -3095
rect 42295 -3215 42350 -3095
rect 42470 -3215 42515 -3095
rect 42635 -3215 42680 -3095
rect 42800 -3215 42845 -3095
rect 42965 -3215 43020 -3095
rect 43140 -3215 43185 -3095
rect 43305 -3215 43350 -3095
rect 43470 -3215 43515 -3095
rect 43635 -3215 43690 -3095
rect 43810 -3215 43855 -3095
rect 43975 -3215 44020 -3095
rect 44140 -3215 44185 -3095
rect 44305 -3215 44360 -3095
rect 44480 -3215 44525 -3095
rect 44645 -3215 44690 -3095
rect 44810 -3215 44855 -3095
rect 44975 -3215 45030 -3095
rect 45150 -3215 45195 -3095
rect 45315 -3215 45360 -3095
rect 45480 -3215 45525 -3095
rect 45645 -3215 45700 -3095
rect 45820 -3215 45865 -3095
rect 45985 -3215 46030 -3095
rect 46150 -3215 46195 -3095
rect 46315 -3215 46370 -3095
rect 46490 -3215 46535 -3095
rect 46655 -3215 46700 -3095
rect 46820 -3215 46865 -3095
rect 46985 -3215 47040 -3095
rect 47160 -3215 47205 -3095
rect 47325 -3215 47370 -3095
rect 47490 -3215 47535 -3095
rect 47655 -3215 47665 -3095
rect 42165 -3270 47665 -3215
rect 42165 -3390 42175 -3270
rect 42295 -3390 42350 -3270
rect 42470 -3390 42515 -3270
rect 42635 -3390 42680 -3270
rect 42800 -3390 42845 -3270
rect 42965 -3390 43020 -3270
rect 43140 -3390 43185 -3270
rect 43305 -3390 43350 -3270
rect 43470 -3390 43515 -3270
rect 43635 -3390 43690 -3270
rect 43810 -3390 43855 -3270
rect 43975 -3390 44020 -3270
rect 44140 -3390 44185 -3270
rect 44305 -3390 44360 -3270
rect 44480 -3390 44525 -3270
rect 44645 -3390 44690 -3270
rect 44810 -3390 44855 -3270
rect 44975 -3390 45030 -3270
rect 45150 -3390 45195 -3270
rect 45315 -3390 45360 -3270
rect 45480 -3390 45525 -3270
rect 45645 -3390 45700 -3270
rect 45820 -3390 45865 -3270
rect 45985 -3390 46030 -3270
rect 46150 -3390 46195 -3270
rect 46315 -3390 46370 -3270
rect 46490 -3390 46535 -3270
rect 46655 -3390 46700 -3270
rect 46820 -3390 46865 -3270
rect 46985 -3390 47040 -3270
rect 47160 -3390 47205 -3270
rect 47325 -3390 47370 -3270
rect 47490 -3390 47535 -3270
rect 47655 -3390 47665 -3270
rect 42165 -3435 47665 -3390
rect 42165 -3555 42175 -3435
rect 42295 -3555 42350 -3435
rect 42470 -3555 42515 -3435
rect 42635 -3555 42680 -3435
rect 42800 -3555 42845 -3435
rect 42965 -3555 43020 -3435
rect 43140 -3555 43185 -3435
rect 43305 -3555 43350 -3435
rect 43470 -3555 43515 -3435
rect 43635 -3555 43690 -3435
rect 43810 -3555 43855 -3435
rect 43975 -3555 44020 -3435
rect 44140 -3555 44185 -3435
rect 44305 -3555 44360 -3435
rect 44480 -3555 44525 -3435
rect 44645 -3555 44690 -3435
rect 44810 -3555 44855 -3435
rect 44975 -3555 45030 -3435
rect 45150 -3555 45195 -3435
rect 45315 -3555 45360 -3435
rect 45480 -3555 45525 -3435
rect 45645 -3555 45700 -3435
rect 45820 -3555 45865 -3435
rect 45985 -3555 46030 -3435
rect 46150 -3555 46195 -3435
rect 46315 -3555 46370 -3435
rect 46490 -3555 46535 -3435
rect 46655 -3555 46700 -3435
rect 46820 -3555 46865 -3435
rect 46985 -3555 47040 -3435
rect 47160 -3555 47205 -3435
rect 47325 -3555 47370 -3435
rect 47490 -3555 47535 -3435
rect 47655 -3555 47665 -3435
rect 42165 -3600 47665 -3555
rect 42165 -3720 42175 -3600
rect 42295 -3720 42350 -3600
rect 42470 -3720 42515 -3600
rect 42635 -3720 42680 -3600
rect 42800 -3720 42845 -3600
rect 42965 -3720 43020 -3600
rect 43140 -3720 43185 -3600
rect 43305 -3720 43350 -3600
rect 43470 -3720 43515 -3600
rect 43635 -3720 43690 -3600
rect 43810 -3720 43855 -3600
rect 43975 -3720 44020 -3600
rect 44140 -3720 44185 -3600
rect 44305 -3720 44360 -3600
rect 44480 -3720 44525 -3600
rect 44645 -3720 44690 -3600
rect 44810 -3720 44855 -3600
rect 44975 -3720 45030 -3600
rect 45150 -3720 45195 -3600
rect 45315 -3720 45360 -3600
rect 45480 -3720 45525 -3600
rect 45645 -3720 45700 -3600
rect 45820 -3720 45865 -3600
rect 45985 -3720 46030 -3600
rect 46150 -3720 46195 -3600
rect 46315 -3720 46370 -3600
rect 46490 -3720 46535 -3600
rect 46655 -3720 46700 -3600
rect 46820 -3720 46865 -3600
rect 46985 -3720 47040 -3600
rect 47160 -3720 47205 -3600
rect 47325 -3720 47370 -3600
rect 47490 -3720 47535 -3600
rect 47655 -3720 47665 -3600
rect 42165 -3765 47665 -3720
rect 42165 -3885 42175 -3765
rect 42295 -3885 42350 -3765
rect 42470 -3885 42515 -3765
rect 42635 -3885 42680 -3765
rect 42800 -3885 42845 -3765
rect 42965 -3885 43020 -3765
rect 43140 -3885 43185 -3765
rect 43305 -3885 43350 -3765
rect 43470 -3885 43515 -3765
rect 43635 -3885 43690 -3765
rect 43810 -3885 43855 -3765
rect 43975 -3885 44020 -3765
rect 44140 -3885 44185 -3765
rect 44305 -3885 44360 -3765
rect 44480 -3885 44525 -3765
rect 44645 -3885 44690 -3765
rect 44810 -3885 44855 -3765
rect 44975 -3885 45030 -3765
rect 45150 -3885 45195 -3765
rect 45315 -3885 45360 -3765
rect 45480 -3885 45525 -3765
rect 45645 -3885 45700 -3765
rect 45820 -3885 45865 -3765
rect 45985 -3885 46030 -3765
rect 46150 -3885 46195 -3765
rect 46315 -3885 46370 -3765
rect 46490 -3885 46535 -3765
rect 46655 -3885 46700 -3765
rect 46820 -3885 46865 -3765
rect 46985 -3885 47040 -3765
rect 47160 -3885 47205 -3765
rect 47325 -3885 47370 -3765
rect 47490 -3885 47535 -3765
rect 47655 -3885 47665 -3765
rect 42165 -3940 47665 -3885
rect 42165 -4060 42175 -3940
rect 42295 -4060 42350 -3940
rect 42470 -4060 42515 -3940
rect 42635 -4060 42680 -3940
rect 42800 -4060 42845 -3940
rect 42965 -4060 43020 -3940
rect 43140 -4060 43185 -3940
rect 43305 -4060 43350 -3940
rect 43470 -4060 43515 -3940
rect 43635 -4060 43690 -3940
rect 43810 -4060 43855 -3940
rect 43975 -4060 44020 -3940
rect 44140 -4060 44185 -3940
rect 44305 -4060 44360 -3940
rect 44480 -4060 44525 -3940
rect 44645 -4060 44690 -3940
rect 44810 -4060 44855 -3940
rect 44975 -4060 45030 -3940
rect 45150 -4060 45195 -3940
rect 45315 -4060 45360 -3940
rect 45480 -4060 45525 -3940
rect 45645 -4060 45700 -3940
rect 45820 -4060 45865 -3940
rect 45985 -4060 46030 -3940
rect 46150 -4060 46195 -3940
rect 46315 -4060 46370 -3940
rect 46490 -4060 46535 -3940
rect 46655 -4060 46700 -3940
rect 46820 -4060 46865 -3940
rect 46985 -4060 47040 -3940
rect 47160 -4060 47205 -3940
rect 47325 -4060 47370 -3940
rect 47490 -4060 47535 -3940
rect 47655 -4060 47665 -3940
rect 42165 -4070 47665 -4060
rect 47855 1420 53355 1430
rect 47855 1300 47865 1420
rect 47985 1300 48040 1420
rect 48160 1300 48205 1420
rect 48325 1300 48370 1420
rect 48490 1300 48535 1420
rect 48655 1300 48710 1420
rect 48830 1300 48875 1420
rect 48995 1300 49040 1420
rect 49160 1300 49205 1420
rect 49325 1300 49380 1420
rect 49500 1300 49545 1420
rect 49665 1300 49710 1420
rect 49830 1300 49875 1420
rect 49995 1300 50050 1420
rect 50170 1300 50215 1420
rect 50335 1300 50380 1420
rect 50500 1300 50545 1420
rect 50665 1300 50720 1420
rect 50840 1300 50885 1420
rect 51005 1300 51050 1420
rect 51170 1300 51215 1420
rect 51335 1300 51390 1420
rect 51510 1300 51555 1420
rect 51675 1300 51720 1420
rect 51840 1300 51885 1420
rect 52005 1300 52060 1420
rect 52180 1300 52225 1420
rect 52345 1300 52390 1420
rect 52510 1300 52555 1420
rect 52675 1300 52730 1420
rect 52850 1300 52895 1420
rect 53015 1300 53060 1420
rect 53180 1300 53225 1420
rect 53345 1300 53355 1420
rect 47855 1255 53355 1300
rect 47855 1135 47865 1255
rect 47985 1135 48040 1255
rect 48160 1135 48205 1255
rect 48325 1135 48370 1255
rect 48490 1135 48535 1255
rect 48655 1135 48710 1255
rect 48830 1135 48875 1255
rect 48995 1135 49040 1255
rect 49160 1135 49205 1255
rect 49325 1135 49380 1255
rect 49500 1135 49545 1255
rect 49665 1135 49710 1255
rect 49830 1135 49875 1255
rect 49995 1135 50050 1255
rect 50170 1135 50215 1255
rect 50335 1135 50380 1255
rect 50500 1135 50545 1255
rect 50665 1135 50720 1255
rect 50840 1135 50885 1255
rect 51005 1135 51050 1255
rect 51170 1135 51215 1255
rect 51335 1135 51390 1255
rect 51510 1135 51555 1255
rect 51675 1135 51720 1255
rect 51840 1135 51885 1255
rect 52005 1135 52060 1255
rect 52180 1135 52225 1255
rect 52345 1135 52390 1255
rect 52510 1135 52555 1255
rect 52675 1135 52730 1255
rect 52850 1135 52895 1255
rect 53015 1135 53060 1255
rect 53180 1135 53225 1255
rect 53345 1135 53355 1255
rect 47855 1090 53355 1135
rect 47855 970 47865 1090
rect 47985 970 48040 1090
rect 48160 970 48205 1090
rect 48325 970 48370 1090
rect 48490 970 48535 1090
rect 48655 970 48710 1090
rect 48830 970 48875 1090
rect 48995 970 49040 1090
rect 49160 970 49205 1090
rect 49325 970 49380 1090
rect 49500 970 49545 1090
rect 49665 970 49710 1090
rect 49830 970 49875 1090
rect 49995 970 50050 1090
rect 50170 970 50215 1090
rect 50335 970 50380 1090
rect 50500 970 50545 1090
rect 50665 970 50720 1090
rect 50840 970 50885 1090
rect 51005 970 51050 1090
rect 51170 970 51215 1090
rect 51335 970 51390 1090
rect 51510 970 51555 1090
rect 51675 970 51720 1090
rect 51840 970 51885 1090
rect 52005 970 52060 1090
rect 52180 970 52225 1090
rect 52345 970 52390 1090
rect 52510 970 52555 1090
rect 52675 970 52730 1090
rect 52850 970 52895 1090
rect 53015 970 53060 1090
rect 53180 970 53225 1090
rect 53345 970 53355 1090
rect 47855 925 53355 970
rect 47855 805 47865 925
rect 47985 805 48040 925
rect 48160 805 48205 925
rect 48325 805 48370 925
rect 48490 805 48535 925
rect 48655 805 48710 925
rect 48830 805 48875 925
rect 48995 805 49040 925
rect 49160 805 49205 925
rect 49325 805 49380 925
rect 49500 805 49545 925
rect 49665 805 49710 925
rect 49830 805 49875 925
rect 49995 805 50050 925
rect 50170 805 50215 925
rect 50335 805 50380 925
rect 50500 805 50545 925
rect 50665 805 50720 925
rect 50840 805 50885 925
rect 51005 805 51050 925
rect 51170 805 51215 925
rect 51335 805 51390 925
rect 51510 805 51555 925
rect 51675 805 51720 925
rect 51840 805 51885 925
rect 52005 805 52060 925
rect 52180 805 52225 925
rect 52345 805 52390 925
rect 52510 805 52555 925
rect 52675 805 52730 925
rect 52850 805 52895 925
rect 53015 805 53060 925
rect 53180 805 53225 925
rect 53345 805 53355 925
rect 47855 750 53355 805
rect 47855 630 47865 750
rect 47985 630 48040 750
rect 48160 630 48205 750
rect 48325 630 48370 750
rect 48490 630 48535 750
rect 48655 630 48710 750
rect 48830 630 48875 750
rect 48995 630 49040 750
rect 49160 630 49205 750
rect 49325 630 49380 750
rect 49500 630 49545 750
rect 49665 630 49710 750
rect 49830 630 49875 750
rect 49995 630 50050 750
rect 50170 630 50215 750
rect 50335 630 50380 750
rect 50500 630 50545 750
rect 50665 630 50720 750
rect 50840 630 50885 750
rect 51005 630 51050 750
rect 51170 630 51215 750
rect 51335 630 51390 750
rect 51510 630 51555 750
rect 51675 630 51720 750
rect 51840 630 51885 750
rect 52005 630 52060 750
rect 52180 630 52225 750
rect 52345 630 52390 750
rect 52510 630 52555 750
rect 52675 630 52730 750
rect 52850 630 52895 750
rect 53015 630 53060 750
rect 53180 630 53225 750
rect 53345 630 53355 750
rect 47855 585 53355 630
rect 47855 465 47865 585
rect 47985 465 48040 585
rect 48160 465 48205 585
rect 48325 465 48370 585
rect 48490 465 48535 585
rect 48655 465 48710 585
rect 48830 465 48875 585
rect 48995 465 49040 585
rect 49160 465 49205 585
rect 49325 465 49380 585
rect 49500 465 49545 585
rect 49665 465 49710 585
rect 49830 465 49875 585
rect 49995 465 50050 585
rect 50170 465 50215 585
rect 50335 465 50380 585
rect 50500 465 50545 585
rect 50665 465 50720 585
rect 50840 465 50885 585
rect 51005 465 51050 585
rect 51170 465 51215 585
rect 51335 465 51390 585
rect 51510 465 51555 585
rect 51675 465 51720 585
rect 51840 465 51885 585
rect 52005 465 52060 585
rect 52180 465 52225 585
rect 52345 465 52390 585
rect 52510 465 52555 585
rect 52675 465 52730 585
rect 52850 465 52895 585
rect 53015 465 53060 585
rect 53180 465 53225 585
rect 53345 465 53355 585
rect 47855 420 53355 465
rect 47855 300 47865 420
rect 47985 300 48040 420
rect 48160 300 48205 420
rect 48325 300 48370 420
rect 48490 300 48535 420
rect 48655 300 48710 420
rect 48830 300 48875 420
rect 48995 300 49040 420
rect 49160 300 49205 420
rect 49325 300 49380 420
rect 49500 300 49545 420
rect 49665 300 49710 420
rect 49830 300 49875 420
rect 49995 300 50050 420
rect 50170 300 50215 420
rect 50335 300 50380 420
rect 50500 300 50545 420
rect 50665 300 50720 420
rect 50840 300 50885 420
rect 51005 300 51050 420
rect 51170 300 51215 420
rect 51335 300 51390 420
rect 51510 300 51555 420
rect 51675 300 51720 420
rect 51840 300 51885 420
rect 52005 300 52060 420
rect 52180 300 52225 420
rect 52345 300 52390 420
rect 52510 300 52555 420
rect 52675 300 52730 420
rect 52850 300 52895 420
rect 53015 300 53060 420
rect 53180 300 53225 420
rect 53345 300 53355 420
rect 47855 255 53355 300
rect 47855 135 47865 255
rect 47985 135 48040 255
rect 48160 135 48205 255
rect 48325 135 48370 255
rect 48490 135 48535 255
rect 48655 135 48710 255
rect 48830 135 48875 255
rect 48995 135 49040 255
rect 49160 135 49205 255
rect 49325 135 49380 255
rect 49500 135 49545 255
rect 49665 135 49710 255
rect 49830 135 49875 255
rect 49995 135 50050 255
rect 50170 135 50215 255
rect 50335 135 50380 255
rect 50500 135 50545 255
rect 50665 135 50720 255
rect 50840 135 50885 255
rect 51005 135 51050 255
rect 51170 135 51215 255
rect 51335 135 51390 255
rect 51510 135 51555 255
rect 51675 135 51720 255
rect 51840 135 51885 255
rect 52005 135 52060 255
rect 52180 135 52225 255
rect 52345 135 52390 255
rect 52510 135 52555 255
rect 52675 135 52730 255
rect 52850 135 52895 255
rect 53015 135 53060 255
rect 53180 135 53225 255
rect 53345 135 53355 255
rect 47855 80 53355 135
rect 47855 -40 47865 80
rect 47985 -40 48040 80
rect 48160 -40 48205 80
rect 48325 -40 48370 80
rect 48490 -40 48535 80
rect 48655 -40 48710 80
rect 48830 -40 48875 80
rect 48995 -40 49040 80
rect 49160 -40 49205 80
rect 49325 -40 49380 80
rect 49500 -40 49545 80
rect 49665 -40 49710 80
rect 49830 -40 49875 80
rect 49995 -40 50050 80
rect 50170 -40 50215 80
rect 50335 -40 50380 80
rect 50500 -40 50545 80
rect 50665 -40 50720 80
rect 50840 -40 50885 80
rect 51005 -40 51050 80
rect 51170 -40 51215 80
rect 51335 -40 51390 80
rect 51510 -40 51555 80
rect 51675 -40 51720 80
rect 51840 -40 51885 80
rect 52005 -40 52060 80
rect 52180 -40 52225 80
rect 52345 -40 52390 80
rect 52510 -40 52555 80
rect 52675 -40 52730 80
rect 52850 -40 52895 80
rect 53015 -40 53060 80
rect 53180 -40 53225 80
rect 53345 -40 53355 80
rect 47855 -85 53355 -40
rect 47855 -205 47865 -85
rect 47985 -205 48040 -85
rect 48160 -205 48205 -85
rect 48325 -205 48370 -85
rect 48490 -205 48535 -85
rect 48655 -205 48710 -85
rect 48830 -205 48875 -85
rect 48995 -205 49040 -85
rect 49160 -205 49205 -85
rect 49325 -205 49380 -85
rect 49500 -205 49545 -85
rect 49665 -205 49710 -85
rect 49830 -205 49875 -85
rect 49995 -205 50050 -85
rect 50170 -205 50215 -85
rect 50335 -205 50380 -85
rect 50500 -205 50545 -85
rect 50665 -205 50720 -85
rect 50840 -205 50885 -85
rect 51005 -205 51050 -85
rect 51170 -205 51215 -85
rect 51335 -205 51390 -85
rect 51510 -205 51555 -85
rect 51675 -205 51720 -85
rect 51840 -205 51885 -85
rect 52005 -205 52060 -85
rect 52180 -205 52225 -85
rect 52345 -205 52390 -85
rect 52510 -205 52555 -85
rect 52675 -205 52730 -85
rect 52850 -205 52895 -85
rect 53015 -205 53060 -85
rect 53180 -205 53225 -85
rect 53345 -205 53355 -85
rect 47855 -250 53355 -205
rect 47855 -370 47865 -250
rect 47985 -370 48040 -250
rect 48160 -370 48205 -250
rect 48325 -370 48370 -250
rect 48490 -370 48535 -250
rect 48655 -370 48710 -250
rect 48830 -370 48875 -250
rect 48995 -370 49040 -250
rect 49160 -370 49205 -250
rect 49325 -370 49380 -250
rect 49500 -370 49545 -250
rect 49665 -370 49710 -250
rect 49830 -370 49875 -250
rect 49995 -370 50050 -250
rect 50170 -370 50215 -250
rect 50335 -370 50380 -250
rect 50500 -370 50545 -250
rect 50665 -370 50720 -250
rect 50840 -370 50885 -250
rect 51005 -370 51050 -250
rect 51170 -370 51215 -250
rect 51335 -370 51390 -250
rect 51510 -370 51555 -250
rect 51675 -370 51720 -250
rect 51840 -370 51885 -250
rect 52005 -370 52060 -250
rect 52180 -370 52225 -250
rect 52345 -370 52390 -250
rect 52510 -370 52555 -250
rect 52675 -370 52730 -250
rect 52850 -370 52895 -250
rect 53015 -370 53060 -250
rect 53180 -370 53225 -250
rect 53345 -370 53355 -250
rect 47855 -415 53355 -370
rect 47855 -535 47865 -415
rect 47985 -535 48040 -415
rect 48160 -535 48205 -415
rect 48325 -535 48370 -415
rect 48490 -535 48535 -415
rect 48655 -535 48710 -415
rect 48830 -535 48875 -415
rect 48995 -535 49040 -415
rect 49160 -535 49205 -415
rect 49325 -535 49380 -415
rect 49500 -535 49545 -415
rect 49665 -535 49710 -415
rect 49830 -535 49875 -415
rect 49995 -535 50050 -415
rect 50170 -535 50215 -415
rect 50335 -535 50380 -415
rect 50500 -535 50545 -415
rect 50665 -535 50720 -415
rect 50840 -535 50885 -415
rect 51005 -535 51050 -415
rect 51170 -535 51215 -415
rect 51335 -535 51390 -415
rect 51510 -535 51555 -415
rect 51675 -535 51720 -415
rect 51840 -535 51885 -415
rect 52005 -535 52060 -415
rect 52180 -535 52225 -415
rect 52345 -535 52390 -415
rect 52510 -535 52555 -415
rect 52675 -535 52730 -415
rect 52850 -535 52895 -415
rect 53015 -535 53060 -415
rect 53180 -535 53225 -415
rect 53345 -535 53355 -415
rect 47855 -590 53355 -535
rect 47855 -710 47865 -590
rect 47985 -710 48040 -590
rect 48160 -710 48205 -590
rect 48325 -710 48370 -590
rect 48490 -710 48535 -590
rect 48655 -710 48710 -590
rect 48830 -710 48875 -590
rect 48995 -710 49040 -590
rect 49160 -710 49205 -590
rect 49325 -710 49380 -590
rect 49500 -710 49545 -590
rect 49665 -710 49710 -590
rect 49830 -710 49875 -590
rect 49995 -710 50050 -590
rect 50170 -710 50215 -590
rect 50335 -710 50380 -590
rect 50500 -710 50545 -590
rect 50665 -710 50720 -590
rect 50840 -710 50885 -590
rect 51005 -710 51050 -590
rect 51170 -710 51215 -590
rect 51335 -710 51390 -590
rect 51510 -710 51555 -590
rect 51675 -710 51720 -590
rect 51840 -710 51885 -590
rect 52005 -710 52060 -590
rect 52180 -710 52225 -590
rect 52345 -710 52390 -590
rect 52510 -710 52555 -590
rect 52675 -710 52730 -590
rect 52850 -710 52895 -590
rect 53015 -710 53060 -590
rect 53180 -710 53225 -590
rect 53345 -710 53355 -590
rect 47855 -755 53355 -710
rect 47855 -875 47865 -755
rect 47985 -875 48040 -755
rect 48160 -875 48205 -755
rect 48325 -875 48370 -755
rect 48490 -875 48535 -755
rect 48655 -875 48710 -755
rect 48830 -875 48875 -755
rect 48995 -875 49040 -755
rect 49160 -875 49205 -755
rect 49325 -875 49380 -755
rect 49500 -875 49545 -755
rect 49665 -875 49710 -755
rect 49830 -875 49875 -755
rect 49995 -875 50050 -755
rect 50170 -875 50215 -755
rect 50335 -875 50380 -755
rect 50500 -875 50545 -755
rect 50665 -875 50720 -755
rect 50840 -875 50885 -755
rect 51005 -875 51050 -755
rect 51170 -875 51215 -755
rect 51335 -875 51390 -755
rect 51510 -875 51555 -755
rect 51675 -875 51720 -755
rect 51840 -875 51885 -755
rect 52005 -875 52060 -755
rect 52180 -875 52225 -755
rect 52345 -875 52390 -755
rect 52510 -875 52555 -755
rect 52675 -875 52730 -755
rect 52850 -875 52895 -755
rect 53015 -875 53060 -755
rect 53180 -875 53225 -755
rect 53345 -875 53355 -755
rect 47855 -920 53355 -875
rect 47855 -1040 47865 -920
rect 47985 -1040 48040 -920
rect 48160 -1040 48205 -920
rect 48325 -1040 48370 -920
rect 48490 -1040 48535 -920
rect 48655 -1040 48710 -920
rect 48830 -1040 48875 -920
rect 48995 -1040 49040 -920
rect 49160 -1040 49205 -920
rect 49325 -1040 49380 -920
rect 49500 -1040 49545 -920
rect 49665 -1040 49710 -920
rect 49830 -1040 49875 -920
rect 49995 -1040 50050 -920
rect 50170 -1040 50215 -920
rect 50335 -1040 50380 -920
rect 50500 -1040 50545 -920
rect 50665 -1040 50720 -920
rect 50840 -1040 50885 -920
rect 51005 -1040 51050 -920
rect 51170 -1040 51215 -920
rect 51335 -1040 51390 -920
rect 51510 -1040 51555 -920
rect 51675 -1040 51720 -920
rect 51840 -1040 51885 -920
rect 52005 -1040 52060 -920
rect 52180 -1040 52225 -920
rect 52345 -1040 52390 -920
rect 52510 -1040 52555 -920
rect 52675 -1040 52730 -920
rect 52850 -1040 52895 -920
rect 53015 -1040 53060 -920
rect 53180 -1040 53225 -920
rect 53345 -1040 53355 -920
rect 47855 -1085 53355 -1040
rect 47855 -1205 47865 -1085
rect 47985 -1205 48040 -1085
rect 48160 -1205 48205 -1085
rect 48325 -1205 48370 -1085
rect 48490 -1205 48535 -1085
rect 48655 -1205 48710 -1085
rect 48830 -1205 48875 -1085
rect 48995 -1205 49040 -1085
rect 49160 -1205 49205 -1085
rect 49325 -1205 49380 -1085
rect 49500 -1205 49545 -1085
rect 49665 -1205 49710 -1085
rect 49830 -1205 49875 -1085
rect 49995 -1205 50050 -1085
rect 50170 -1205 50215 -1085
rect 50335 -1205 50380 -1085
rect 50500 -1205 50545 -1085
rect 50665 -1205 50720 -1085
rect 50840 -1205 50885 -1085
rect 51005 -1205 51050 -1085
rect 51170 -1205 51215 -1085
rect 51335 -1205 51390 -1085
rect 51510 -1205 51555 -1085
rect 51675 -1205 51720 -1085
rect 51840 -1205 51885 -1085
rect 52005 -1205 52060 -1085
rect 52180 -1205 52225 -1085
rect 52345 -1205 52390 -1085
rect 52510 -1205 52555 -1085
rect 52675 -1205 52730 -1085
rect 52850 -1205 52895 -1085
rect 53015 -1205 53060 -1085
rect 53180 -1205 53225 -1085
rect 53345 -1205 53355 -1085
rect 47855 -1260 53355 -1205
rect 47855 -1380 47865 -1260
rect 47985 -1380 48040 -1260
rect 48160 -1380 48205 -1260
rect 48325 -1380 48370 -1260
rect 48490 -1380 48535 -1260
rect 48655 -1380 48710 -1260
rect 48830 -1380 48875 -1260
rect 48995 -1380 49040 -1260
rect 49160 -1380 49205 -1260
rect 49325 -1380 49380 -1260
rect 49500 -1380 49545 -1260
rect 49665 -1380 49710 -1260
rect 49830 -1380 49875 -1260
rect 49995 -1380 50050 -1260
rect 50170 -1380 50215 -1260
rect 50335 -1380 50380 -1260
rect 50500 -1380 50545 -1260
rect 50665 -1380 50720 -1260
rect 50840 -1380 50885 -1260
rect 51005 -1380 51050 -1260
rect 51170 -1380 51215 -1260
rect 51335 -1380 51390 -1260
rect 51510 -1380 51555 -1260
rect 51675 -1380 51720 -1260
rect 51840 -1380 51885 -1260
rect 52005 -1380 52060 -1260
rect 52180 -1380 52225 -1260
rect 52345 -1380 52390 -1260
rect 52510 -1380 52555 -1260
rect 52675 -1380 52730 -1260
rect 52850 -1380 52895 -1260
rect 53015 -1380 53060 -1260
rect 53180 -1380 53225 -1260
rect 53345 -1380 53355 -1260
rect 47855 -1425 53355 -1380
rect 47855 -1545 47865 -1425
rect 47985 -1545 48040 -1425
rect 48160 -1545 48205 -1425
rect 48325 -1545 48370 -1425
rect 48490 -1545 48535 -1425
rect 48655 -1545 48710 -1425
rect 48830 -1545 48875 -1425
rect 48995 -1545 49040 -1425
rect 49160 -1545 49205 -1425
rect 49325 -1545 49380 -1425
rect 49500 -1545 49545 -1425
rect 49665 -1545 49710 -1425
rect 49830 -1545 49875 -1425
rect 49995 -1545 50050 -1425
rect 50170 -1545 50215 -1425
rect 50335 -1545 50380 -1425
rect 50500 -1545 50545 -1425
rect 50665 -1545 50720 -1425
rect 50840 -1545 50885 -1425
rect 51005 -1545 51050 -1425
rect 51170 -1545 51215 -1425
rect 51335 -1545 51390 -1425
rect 51510 -1545 51555 -1425
rect 51675 -1545 51720 -1425
rect 51840 -1545 51885 -1425
rect 52005 -1545 52060 -1425
rect 52180 -1545 52225 -1425
rect 52345 -1545 52390 -1425
rect 52510 -1545 52555 -1425
rect 52675 -1545 52730 -1425
rect 52850 -1545 52895 -1425
rect 53015 -1545 53060 -1425
rect 53180 -1545 53225 -1425
rect 53345 -1545 53355 -1425
rect 47855 -1590 53355 -1545
rect 47855 -1710 47865 -1590
rect 47985 -1710 48040 -1590
rect 48160 -1710 48205 -1590
rect 48325 -1710 48370 -1590
rect 48490 -1710 48535 -1590
rect 48655 -1710 48710 -1590
rect 48830 -1710 48875 -1590
rect 48995 -1710 49040 -1590
rect 49160 -1710 49205 -1590
rect 49325 -1710 49380 -1590
rect 49500 -1710 49545 -1590
rect 49665 -1710 49710 -1590
rect 49830 -1710 49875 -1590
rect 49995 -1710 50050 -1590
rect 50170 -1710 50215 -1590
rect 50335 -1710 50380 -1590
rect 50500 -1710 50545 -1590
rect 50665 -1710 50720 -1590
rect 50840 -1710 50885 -1590
rect 51005 -1710 51050 -1590
rect 51170 -1710 51215 -1590
rect 51335 -1710 51390 -1590
rect 51510 -1710 51555 -1590
rect 51675 -1710 51720 -1590
rect 51840 -1710 51885 -1590
rect 52005 -1710 52060 -1590
rect 52180 -1710 52225 -1590
rect 52345 -1710 52390 -1590
rect 52510 -1710 52555 -1590
rect 52675 -1710 52730 -1590
rect 52850 -1710 52895 -1590
rect 53015 -1710 53060 -1590
rect 53180 -1710 53225 -1590
rect 53345 -1710 53355 -1590
rect 47855 -1755 53355 -1710
rect 47855 -1875 47865 -1755
rect 47985 -1875 48040 -1755
rect 48160 -1875 48205 -1755
rect 48325 -1875 48370 -1755
rect 48490 -1875 48535 -1755
rect 48655 -1875 48710 -1755
rect 48830 -1875 48875 -1755
rect 48995 -1875 49040 -1755
rect 49160 -1875 49205 -1755
rect 49325 -1875 49380 -1755
rect 49500 -1875 49545 -1755
rect 49665 -1875 49710 -1755
rect 49830 -1875 49875 -1755
rect 49995 -1875 50050 -1755
rect 50170 -1875 50215 -1755
rect 50335 -1875 50380 -1755
rect 50500 -1875 50545 -1755
rect 50665 -1875 50720 -1755
rect 50840 -1875 50885 -1755
rect 51005 -1875 51050 -1755
rect 51170 -1875 51215 -1755
rect 51335 -1875 51390 -1755
rect 51510 -1875 51555 -1755
rect 51675 -1875 51720 -1755
rect 51840 -1875 51885 -1755
rect 52005 -1875 52060 -1755
rect 52180 -1875 52225 -1755
rect 52345 -1875 52390 -1755
rect 52510 -1875 52555 -1755
rect 52675 -1875 52730 -1755
rect 52850 -1875 52895 -1755
rect 53015 -1875 53060 -1755
rect 53180 -1875 53225 -1755
rect 53345 -1875 53355 -1755
rect 47855 -1930 53355 -1875
rect 47855 -2050 47865 -1930
rect 47985 -2050 48040 -1930
rect 48160 -2050 48205 -1930
rect 48325 -2050 48370 -1930
rect 48490 -2050 48535 -1930
rect 48655 -2050 48710 -1930
rect 48830 -2050 48875 -1930
rect 48995 -2050 49040 -1930
rect 49160 -2050 49205 -1930
rect 49325 -2050 49380 -1930
rect 49500 -2050 49545 -1930
rect 49665 -2050 49710 -1930
rect 49830 -2050 49875 -1930
rect 49995 -2050 50050 -1930
rect 50170 -2050 50215 -1930
rect 50335 -2050 50380 -1930
rect 50500 -2050 50545 -1930
rect 50665 -2050 50720 -1930
rect 50840 -2050 50885 -1930
rect 51005 -2050 51050 -1930
rect 51170 -2050 51215 -1930
rect 51335 -2050 51390 -1930
rect 51510 -2050 51555 -1930
rect 51675 -2050 51720 -1930
rect 51840 -2050 51885 -1930
rect 52005 -2050 52060 -1930
rect 52180 -2050 52225 -1930
rect 52345 -2050 52390 -1930
rect 52510 -2050 52555 -1930
rect 52675 -2050 52730 -1930
rect 52850 -2050 52895 -1930
rect 53015 -2050 53060 -1930
rect 53180 -2050 53225 -1930
rect 53345 -2050 53355 -1930
rect 47855 -2095 53355 -2050
rect 47855 -2215 47865 -2095
rect 47985 -2215 48040 -2095
rect 48160 -2215 48205 -2095
rect 48325 -2215 48370 -2095
rect 48490 -2215 48535 -2095
rect 48655 -2215 48710 -2095
rect 48830 -2215 48875 -2095
rect 48995 -2215 49040 -2095
rect 49160 -2215 49205 -2095
rect 49325 -2215 49380 -2095
rect 49500 -2215 49545 -2095
rect 49665 -2215 49710 -2095
rect 49830 -2215 49875 -2095
rect 49995 -2215 50050 -2095
rect 50170 -2215 50215 -2095
rect 50335 -2215 50380 -2095
rect 50500 -2215 50545 -2095
rect 50665 -2215 50720 -2095
rect 50840 -2215 50885 -2095
rect 51005 -2215 51050 -2095
rect 51170 -2215 51215 -2095
rect 51335 -2215 51390 -2095
rect 51510 -2215 51555 -2095
rect 51675 -2215 51720 -2095
rect 51840 -2215 51885 -2095
rect 52005 -2215 52060 -2095
rect 52180 -2215 52225 -2095
rect 52345 -2215 52390 -2095
rect 52510 -2215 52555 -2095
rect 52675 -2215 52730 -2095
rect 52850 -2215 52895 -2095
rect 53015 -2215 53060 -2095
rect 53180 -2215 53225 -2095
rect 53345 -2215 53355 -2095
rect 47855 -2260 53355 -2215
rect 47855 -2380 47865 -2260
rect 47985 -2380 48040 -2260
rect 48160 -2380 48205 -2260
rect 48325 -2380 48370 -2260
rect 48490 -2380 48535 -2260
rect 48655 -2380 48710 -2260
rect 48830 -2380 48875 -2260
rect 48995 -2380 49040 -2260
rect 49160 -2380 49205 -2260
rect 49325 -2380 49380 -2260
rect 49500 -2380 49545 -2260
rect 49665 -2380 49710 -2260
rect 49830 -2380 49875 -2260
rect 49995 -2380 50050 -2260
rect 50170 -2380 50215 -2260
rect 50335 -2380 50380 -2260
rect 50500 -2380 50545 -2260
rect 50665 -2380 50720 -2260
rect 50840 -2380 50885 -2260
rect 51005 -2380 51050 -2260
rect 51170 -2380 51215 -2260
rect 51335 -2380 51390 -2260
rect 51510 -2380 51555 -2260
rect 51675 -2380 51720 -2260
rect 51840 -2380 51885 -2260
rect 52005 -2380 52060 -2260
rect 52180 -2380 52225 -2260
rect 52345 -2380 52390 -2260
rect 52510 -2380 52555 -2260
rect 52675 -2380 52730 -2260
rect 52850 -2380 52895 -2260
rect 53015 -2380 53060 -2260
rect 53180 -2380 53225 -2260
rect 53345 -2380 53355 -2260
rect 47855 -2425 53355 -2380
rect 47855 -2545 47865 -2425
rect 47985 -2545 48040 -2425
rect 48160 -2545 48205 -2425
rect 48325 -2545 48370 -2425
rect 48490 -2545 48535 -2425
rect 48655 -2545 48710 -2425
rect 48830 -2545 48875 -2425
rect 48995 -2545 49040 -2425
rect 49160 -2545 49205 -2425
rect 49325 -2545 49380 -2425
rect 49500 -2545 49545 -2425
rect 49665 -2545 49710 -2425
rect 49830 -2545 49875 -2425
rect 49995 -2545 50050 -2425
rect 50170 -2545 50215 -2425
rect 50335 -2545 50380 -2425
rect 50500 -2545 50545 -2425
rect 50665 -2545 50720 -2425
rect 50840 -2545 50885 -2425
rect 51005 -2545 51050 -2425
rect 51170 -2545 51215 -2425
rect 51335 -2545 51390 -2425
rect 51510 -2545 51555 -2425
rect 51675 -2545 51720 -2425
rect 51840 -2545 51885 -2425
rect 52005 -2545 52060 -2425
rect 52180 -2545 52225 -2425
rect 52345 -2545 52390 -2425
rect 52510 -2545 52555 -2425
rect 52675 -2545 52730 -2425
rect 52850 -2545 52895 -2425
rect 53015 -2545 53060 -2425
rect 53180 -2545 53225 -2425
rect 53345 -2545 53355 -2425
rect 47855 -2600 53355 -2545
rect 47855 -2720 47865 -2600
rect 47985 -2720 48040 -2600
rect 48160 -2720 48205 -2600
rect 48325 -2720 48370 -2600
rect 48490 -2720 48535 -2600
rect 48655 -2720 48710 -2600
rect 48830 -2720 48875 -2600
rect 48995 -2720 49040 -2600
rect 49160 -2720 49205 -2600
rect 49325 -2720 49380 -2600
rect 49500 -2720 49545 -2600
rect 49665 -2720 49710 -2600
rect 49830 -2720 49875 -2600
rect 49995 -2720 50050 -2600
rect 50170 -2720 50215 -2600
rect 50335 -2720 50380 -2600
rect 50500 -2720 50545 -2600
rect 50665 -2720 50720 -2600
rect 50840 -2720 50885 -2600
rect 51005 -2720 51050 -2600
rect 51170 -2720 51215 -2600
rect 51335 -2720 51390 -2600
rect 51510 -2720 51555 -2600
rect 51675 -2720 51720 -2600
rect 51840 -2720 51885 -2600
rect 52005 -2720 52060 -2600
rect 52180 -2720 52225 -2600
rect 52345 -2720 52390 -2600
rect 52510 -2720 52555 -2600
rect 52675 -2720 52730 -2600
rect 52850 -2720 52895 -2600
rect 53015 -2720 53060 -2600
rect 53180 -2720 53225 -2600
rect 53345 -2720 53355 -2600
rect 47855 -2765 53355 -2720
rect 47855 -2885 47865 -2765
rect 47985 -2885 48040 -2765
rect 48160 -2885 48205 -2765
rect 48325 -2885 48370 -2765
rect 48490 -2885 48535 -2765
rect 48655 -2885 48710 -2765
rect 48830 -2885 48875 -2765
rect 48995 -2885 49040 -2765
rect 49160 -2885 49205 -2765
rect 49325 -2885 49380 -2765
rect 49500 -2885 49545 -2765
rect 49665 -2885 49710 -2765
rect 49830 -2885 49875 -2765
rect 49995 -2885 50050 -2765
rect 50170 -2885 50215 -2765
rect 50335 -2885 50380 -2765
rect 50500 -2885 50545 -2765
rect 50665 -2885 50720 -2765
rect 50840 -2885 50885 -2765
rect 51005 -2885 51050 -2765
rect 51170 -2885 51215 -2765
rect 51335 -2885 51390 -2765
rect 51510 -2885 51555 -2765
rect 51675 -2885 51720 -2765
rect 51840 -2885 51885 -2765
rect 52005 -2885 52060 -2765
rect 52180 -2885 52225 -2765
rect 52345 -2885 52390 -2765
rect 52510 -2885 52555 -2765
rect 52675 -2885 52730 -2765
rect 52850 -2885 52895 -2765
rect 53015 -2885 53060 -2765
rect 53180 -2885 53225 -2765
rect 53345 -2885 53355 -2765
rect 47855 -2930 53355 -2885
rect 47855 -3050 47865 -2930
rect 47985 -3050 48040 -2930
rect 48160 -3050 48205 -2930
rect 48325 -3050 48370 -2930
rect 48490 -3050 48535 -2930
rect 48655 -3050 48710 -2930
rect 48830 -3050 48875 -2930
rect 48995 -3050 49040 -2930
rect 49160 -3050 49205 -2930
rect 49325 -3050 49380 -2930
rect 49500 -3050 49545 -2930
rect 49665 -3050 49710 -2930
rect 49830 -3050 49875 -2930
rect 49995 -3050 50050 -2930
rect 50170 -3050 50215 -2930
rect 50335 -3050 50380 -2930
rect 50500 -3050 50545 -2930
rect 50665 -3050 50720 -2930
rect 50840 -3050 50885 -2930
rect 51005 -3050 51050 -2930
rect 51170 -3050 51215 -2930
rect 51335 -3050 51390 -2930
rect 51510 -3050 51555 -2930
rect 51675 -3050 51720 -2930
rect 51840 -3050 51885 -2930
rect 52005 -3050 52060 -2930
rect 52180 -3050 52225 -2930
rect 52345 -3050 52390 -2930
rect 52510 -3050 52555 -2930
rect 52675 -3050 52730 -2930
rect 52850 -3050 52895 -2930
rect 53015 -3050 53060 -2930
rect 53180 -3050 53225 -2930
rect 53345 -3050 53355 -2930
rect 47855 -3095 53355 -3050
rect 47855 -3215 47865 -3095
rect 47985 -3215 48040 -3095
rect 48160 -3215 48205 -3095
rect 48325 -3215 48370 -3095
rect 48490 -3215 48535 -3095
rect 48655 -3215 48710 -3095
rect 48830 -3215 48875 -3095
rect 48995 -3215 49040 -3095
rect 49160 -3215 49205 -3095
rect 49325 -3215 49380 -3095
rect 49500 -3215 49545 -3095
rect 49665 -3215 49710 -3095
rect 49830 -3215 49875 -3095
rect 49995 -3215 50050 -3095
rect 50170 -3215 50215 -3095
rect 50335 -3215 50380 -3095
rect 50500 -3215 50545 -3095
rect 50665 -3215 50720 -3095
rect 50840 -3215 50885 -3095
rect 51005 -3215 51050 -3095
rect 51170 -3215 51215 -3095
rect 51335 -3215 51390 -3095
rect 51510 -3215 51555 -3095
rect 51675 -3215 51720 -3095
rect 51840 -3215 51885 -3095
rect 52005 -3215 52060 -3095
rect 52180 -3215 52225 -3095
rect 52345 -3215 52390 -3095
rect 52510 -3215 52555 -3095
rect 52675 -3215 52730 -3095
rect 52850 -3215 52895 -3095
rect 53015 -3215 53060 -3095
rect 53180 -3215 53225 -3095
rect 53345 -3215 53355 -3095
rect 47855 -3270 53355 -3215
rect 47855 -3390 47865 -3270
rect 47985 -3390 48040 -3270
rect 48160 -3390 48205 -3270
rect 48325 -3390 48370 -3270
rect 48490 -3390 48535 -3270
rect 48655 -3390 48710 -3270
rect 48830 -3390 48875 -3270
rect 48995 -3390 49040 -3270
rect 49160 -3390 49205 -3270
rect 49325 -3390 49380 -3270
rect 49500 -3390 49545 -3270
rect 49665 -3390 49710 -3270
rect 49830 -3390 49875 -3270
rect 49995 -3390 50050 -3270
rect 50170 -3390 50215 -3270
rect 50335 -3390 50380 -3270
rect 50500 -3390 50545 -3270
rect 50665 -3390 50720 -3270
rect 50840 -3390 50885 -3270
rect 51005 -3390 51050 -3270
rect 51170 -3390 51215 -3270
rect 51335 -3390 51390 -3270
rect 51510 -3390 51555 -3270
rect 51675 -3390 51720 -3270
rect 51840 -3390 51885 -3270
rect 52005 -3390 52060 -3270
rect 52180 -3390 52225 -3270
rect 52345 -3390 52390 -3270
rect 52510 -3390 52555 -3270
rect 52675 -3390 52730 -3270
rect 52850 -3390 52895 -3270
rect 53015 -3390 53060 -3270
rect 53180 -3390 53225 -3270
rect 53345 -3390 53355 -3270
rect 47855 -3435 53355 -3390
rect 47855 -3555 47865 -3435
rect 47985 -3555 48040 -3435
rect 48160 -3555 48205 -3435
rect 48325 -3555 48370 -3435
rect 48490 -3555 48535 -3435
rect 48655 -3555 48710 -3435
rect 48830 -3555 48875 -3435
rect 48995 -3555 49040 -3435
rect 49160 -3555 49205 -3435
rect 49325 -3555 49380 -3435
rect 49500 -3555 49545 -3435
rect 49665 -3555 49710 -3435
rect 49830 -3555 49875 -3435
rect 49995 -3555 50050 -3435
rect 50170 -3555 50215 -3435
rect 50335 -3555 50380 -3435
rect 50500 -3555 50545 -3435
rect 50665 -3555 50720 -3435
rect 50840 -3555 50885 -3435
rect 51005 -3555 51050 -3435
rect 51170 -3555 51215 -3435
rect 51335 -3555 51390 -3435
rect 51510 -3555 51555 -3435
rect 51675 -3555 51720 -3435
rect 51840 -3555 51885 -3435
rect 52005 -3555 52060 -3435
rect 52180 -3555 52225 -3435
rect 52345 -3555 52390 -3435
rect 52510 -3555 52555 -3435
rect 52675 -3555 52730 -3435
rect 52850 -3555 52895 -3435
rect 53015 -3555 53060 -3435
rect 53180 -3555 53225 -3435
rect 53345 -3555 53355 -3435
rect 47855 -3600 53355 -3555
rect 47855 -3720 47865 -3600
rect 47985 -3720 48040 -3600
rect 48160 -3720 48205 -3600
rect 48325 -3720 48370 -3600
rect 48490 -3720 48535 -3600
rect 48655 -3720 48710 -3600
rect 48830 -3720 48875 -3600
rect 48995 -3720 49040 -3600
rect 49160 -3720 49205 -3600
rect 49325 -3720 49380 -3600
rect 49500 -3720 49545 -3600
rect 49665 -3720 49710 -3600
rect 49830 -3720 49875 -3600
rect 49995 -3720 50050 -3600
rect 50170 -3720 50215 -3600
rect 50335 -3720 50380 -3600
rect 50500 -3720 50545 -3600
rect 50665 -3720 50720 -3600
rect 50840 -3720 50885 -3600
rect 51005 -3720 51050 -3600
rect 51170 -3720 51215 -3600
rect 51335 -3720 51390 -3600
rect 51510 -3720 51555 -3600
rect 51675 -3720 51720 -3600
rect 51840 -3720 51885 -3600
rect 52005 -3720 52060 -3600
rect 52180 -3720 52225 -3600
rect 52345 -3720 52390 -3600
rect 52510 -3720 52555 -3600
rect 52675 -3720 52730 -3600
rect 52850 -3720 52895 -3600
rect 53015 -3720 53060 -3600
rect 53180 -3720 53225 -3600
rect 53345 -3720 53355 -3600
rect 47855 -3765 53355 -3720
rect 47855 -3885 47865 -3765
rect 47985 -3885 48040 -3765
rect 48160 -3885 48205 -3765
rect 48325 -3885 48370 -3765
rect 48490 -3885 48535 -3765
rect 48655 -3885 48710 -3765
rect 48830 -3885 48875 -3765
rect 48995 -3885 49040 -3765
rect 49160 -3885 49205 -3765
rect 49325 -3885 49380 -3765
rect 49500 -3885 49545 -3765
rect 49665 -3885 49710 -3765
rect 49830 -3885 49875 -3765
rect 49995 -3885 50050 -3765
rect 50170 -3885 50215 -3765
rect 50335 -3885 50380 -3765
rect 50500 -3885 50545 -3765
rect 50665 -3885 50720 -3765
rect 50840 -3885 50885 -3765
rect 51005 -3885 51050 -3765
rect 51170 -3885 51215 -3765
rect 51335 -3885 51390 -3765
rect 51510 -3885 51555 -3765
rect 51675 -3885 51720 -3765
rect 51840 -3885 51885 -3765
rect 52005 -3885 52060 -3765
rect 52180 -3885 52225 -3765
rect 52345 -3885 52390 -3765
rect 52510 -3885 52555 -3765
rect 52675 -3885 52730 -3765
rect 52850 -3885 52895 -3765
rect 53015 -3885 53060 -3765
rect 53180 -3885 53225 -3765
rect 53345 -3885 53355 -3765
rect 47855 -3940 53355 -3885
rect 47855 -4060 47865 -3940
rect 47985 -4060 48040 -3940
rect 48160 -4060 48205 -3940
rect 48325 -4060 48370 -3940
rect 48490 -4060 48535 -3940
rect 48655 -4060 48710 -3940
rect 48830 -4060 48875 -3940
rect 48995 -4060 49040 -3940
rect 49160 -4060 49205 -3940
rect 49325 -4060 49380 -3940
rect 49500 -4060 49545 -3940
rect 49665 -4060 49710 -3940
rect 49830 -4060 49875 -3940
rect 49995 -4060 50050 -3940
rect 50170 -4060 50215 -3940
rect 50335 -4060 50380 -3940
rect 50500 -4060 50545 -3940
rect 50665 -4060 50720 -3940
rect 50840 -4060 50885 -3940
rect 51005 -4060 51050 -3940
rect 51170 -4060 51215 -3940
rect 51335 -4060 51390 -3940
rect 51510 -4060 51555 -3940
rect 51675 -4060 51720 -3940
rect 51840 -4060 51885 -3940
rect 52005 -4060 52060 -3940
rect 52180 -4060 52225 -3940
rect 52345 -4060 52390 -3940
rect 52510 -4060 52555 -3940
rect 52675 -4060 52730 -3940
rect 52850 -4060 52895 -3940
rect 53015 -4060 53060 -3940
rect 53180 -4060 53225 -3940
rect 53345 -4060 53355 -3940
rect 47855 -4070 53355 -4060
rect 30785 -4270 36285 -4260
rect 30785 -4390 30795 -4270
rect 30915 -4390 30960 -4270
rect 31080 -4390 31125 -4270
rect 31245 -4390 31290 -4270
rect 31410 -4390 31465 -4270
rect 31585 -4390 31630 -4270
rect 31750 -4390 31795 -4270
rect 31915 -4390 31960 -4270
rect 32080 -4390 32135 -4270
rect 32255 -4390 32300 -4270
rect 32420 -4390 32465 -4270
rect 32585 -4390 32630 -4270
rect 32750 -4390 32805 -4270
rect 32925 -4390 32970 -4270
rect 33090 -4390 33135 -4270
rect 33255 -4390 33300 -4270
rect 33420 -4390 33475 -4270
rect 33595 -4390 33640 -4270
rect 33760 -4390 33805 -4270
rect 33925 -4390 33970 -4270
rect 34090 -4390 34145 -4270
rect 34265 -4390 34310 -4270
rect 34430 -4390 34475 -4270
rect 34595 -4390 34640 -4270
rect 34760 -4390 34815 -4270
rect 34935 -4390 34980 -4270
rect 35100 -4390 35145 -4270
rect 35265 -4390 35310 -4270
rect 35430 -4390 35485 -4270
rect 35605 -4390 35650 -4270
rect 35770 -4390 35815 -4270
rect 35935 -4390 35980 -4270
rect 36100 -4390 36155 -4270
rect 36275 -4390 36285 -4270
rect 30785 -4445 36285 -4390
rect 30785 -4565 30795 -4445
rect 30915 -4565 30960 -4445
rect 31080 -4565 31125 -4445
rect 31245 -4565 31290 -4445
rect 31410 -4565 31465 -4445
rect 31585 -4565 31630 -4445
rect 31750 -4565 31795 -4445
rect 31915 -4565 31960 -4445
rect 32080 -4565 32135 -4445
rect 32255 -4565 32300 -4445
rect 32420 -4565 32465 -4445
rect 32585 -4565 32630 -4445
rect 32750 -4565 32805 -4445
rect 32925 -4565 32970 -4445
rect 33090 -4565 33135 -4445
rect 33255 -4565 33300 -4445
rect 33420 -4565 33475 -4445
rect 33595 -4565 33640 -4445
rect 33760 -4565 33805 -4445
rect 33925 -4565 33970 -4445
rect 34090 -4565 34145 -4445
rect 34265 -4565 34310 -4445
rect 34430 -4565 34475 -4445
rect 34595 -4565 34640 -4445
rect 34760 -4565 34815 -4445
rect 34935 -4565 34980 -4445
rect 35100 -4565 35145 -4445
rect 35265 -4565 35310 -4445
rect 35430 -4565 35485 -4445
rect 35605 -4565 35650 -4445
rect 35770 -4565 35815 -4445
rect 35935 -4565 35980 -4445
rect 36100 -4565 36155 -4445
rect 36275 -4565 36285 -4445
rect 30785 -4610 36285 -4565
rect 30785 -4730 30795 -4610
rect 30915 -4730 30960 -4610
rect 31080 -4730 31125 -4610
rect 31245 -4730 31290 -4610
rect 31410 -4730 31465 -4610
rect 31585 -4730 31630 -4610
rect 31750 -4730 31795 -4610
rect 31915 -4730 31960 -4610
rect 32080 -4730 32135 -4610
rect 32255 -4730 32300 -4610
rect 32420 -4730 32465 -4610
rect 32585 -4730 32630 -4610
rect 32750 -4730 32805 -4610
rect 32925 -4730 32970 -4610
rect 33090 -4730 33135 -4610
rect 33255 -4730 33300 -4610
rect 33420 -4730 33475 -4610
rect 33595 -4730 33640 -4610
rect 33760 -4730 33805 -4610
rect 33925 -4730 33970 -4610
rect 34090 -4730 34145 -4610
rect 34265 -4730 34310 -4610
rect 34430 -4730 34475 -4610
rect 34595 -4730 34640 -4610
rect 34760 -4730 34815 -4610
rect 34935 -4730 34980 -4610
rect 35100 -4730 35145 -4610
rect 35265 -4730 35310 -4610
rect 35430 -4730 35485 -4610
rect 35605 -4730 35650 -4610
rect 35770 -4730 35815 -4610
rect 35935 -4730 35980 -4610
rect 36100 -4730 36155 -4610
rect 36275 -4730 36285 -4610
rect 30785 -4775 36285 -4730
rect 30785 -4895 30795 -4775
rect 30915 -4895 30960 -4775
rect 31080 -4895 31125 -4775
rect 31245 -4895 31290 -4775
rect 31410 -4895 31465 -4775
rect 31585 -4895 31630 -4775
rect 31750 -4895 31795 -4775
rect 31915 -4895 31960 -4775
rect 32080 -4895 32135 -4775
rect 32255 -4895 32300 -4775
rect 32420 -4895 32465 -4775
rect 32585 -4895 32630 -4775
rect 32750 -4895 32805 -4775
rect 32925 -4895 32970 -4775
rect 33090 -4895 33135 -4775
rect 33255 -4895 33300 -4775
rect 33420 -4895 33475 -4775
rect 33595 -4895 33640 -4775
rect 33760 -4895 33805 -4775
rect 33925 -4895 33970 -4775
rect 34090 -4895 34145 -4775
rect 34265 -4895 34310 -4775
rect 34430 -4895 34475 -4775
rect 34595 -4895 34640 -4775
rect 34760 -4895 34815 -4775
rect 34935 -4895 34980 -4775
rect 35100 -4895 35145 -4775
rect 35265 -4895 35310 -4775
rect 35430 -4895 35485 -4775
rect 35605 -4895 35650 -4775
rect 35770 -4895 35815 -4775
rect 35935 -4895 35980 -4775
rect 36100 -4895 36155 -4775
rect 36275 -4895 36285 -4775
rect 30785 -4940 36285 -4895
rect 30785 -5060 30795 -4940
rect 30915 -5060 30960 -4940
rect 31080 -5060 31125 -4940
rect 31245 -5060 31290 -4940
rect 31410 -5060 31465 -4940
rect 31585 -5060 31630 -4940
rect 31750 -5060 31795 -4940
rect 31915 -5060 31960 -4940
rect 32080 -5060 32135 -4940
rect 32255 -5060 32300 -4940
rect 32420 -5060 32465 -4940
rect 32585 -5060 32630 -4940
rect 32750 -5060 32805 -4940
rect 32925 -5060 32970 -4940
rect 33090 -5060 33135 -4940
rect 33255 -5060 33300 -4940
rect 33420 -5060 33475 -4940
rect 33595 -5060 33640 -4940
rect 33760 -5060 33805 -4940
rect 33925 -5060 33970 -4940
rect 34090 -5060 34145 -4940
rect 34265 -5060 34310 -4940
rect 34430 -5060 34475 -4940
rect 34595 -5060 34640 -4940
rect 34760 -5060 34815 -4940
rect 34935 -5060 34980 -4940
rect 35100 -5060 35145 -4940
rect 35265 -5060 35310 -4940
rect 35430 -5060 35485 -4940
rect 35605 -5060 35650 -4940
rect 35770 -5060 35815 -4940
rect 35935 -5060 35980 -4940
rect 36100 -5060 36155 -4940
rect 36275 -5060 36285 -4940
rect 30785 -5115 36285 -5060
rect 30785 -5235 30795 -5115
rect 30915 -5235 30960 -5115
rect 31080 -5235 31125 -5115
rect 31245 -5235 31290 -5115
rect 31410 -5235 31465 -5115
rect 31585 -5235 31630 -5115
rect 31750 -5235 31795 -5115
rect 31915 -5235 31960 -5115
rect 32080 -5235 32135 -5115
rect 32255 -5235 32300 -5115
rect 32420 -5235 32465 -5115
rect 32585 -5235 32630 -5115
rect 32750 -5235 32805 -5115
rect 32925 -5235 32970 -5115
rect 33090 -5235 33135 -5115
rect 33255 -5235 33300 -5115
rect 33420 -5235 33475 -5115
rect 33595 -5235 33640 -5115
rect 33760 -5235 33805 -5115
rect 33925 -5235 33970 -5115
rect 34090 -5235 34145 -5115
rect 34265 -5235 34310 -5115
rect 34430 -5235 34475 -5115
rect 34595 -5235 34640 -5115
rect 34760 -5235 34815 -5115
rect 34935 -5235 34980 -5115
rect 35100 -5235 35145 -5115
rect 35265 -5235 35310 -5115
rect 35430 -5235 35485 -5115
rect 35605 -5235 35650 -5115
rect 35770 -5235 35815 -5115
rect 35935 -5235 35980 -5115
rect 36100 -5235 36155 -5115
rect 36275 -5235 36285 -5115
rect 30785 -5280 36285 -5235
rect 30785 -5400 30795 -5280
rect 30915 -5400 30960 -5280
rect 31080 -5400 31125 -5280
rect 31245 -5400 31290 -5280
rect 31410 -5400 31465 -5280
rect 31585 -5400 31630 -5280
rect 31750 -5400 31795 -5280
rect 31915 -5400 31960 -5280
rect 32080 -5400 32135 -5280
rect 32255 -5400 32300 -5280
rect 32420 -5400 32465 -5280
rect 32585 -5400 32630 -5280
rect 32750 -5400 32805 -5280
rect 32925 -5400 32970 -5280
rect 33090 -5400 33135 -5280
rect 33255 -5400 33300 -5280
rect 33420 -5400 33475 -5280
rect 33595 -5400 33640 -5280
rect 33760 -5400 33805 -5280
rect 33925 -5400 33970 -5280
rect 34090 -5400 34145 -5280
rect 34265 -5400 34310 -5280
rect 34430 -5400 34475 -5280
rect 34595 -5400 34640 -5280
rect 34760 -5400 34815 -5280
rect 34935 -5400 34980 -5280
rect 35100 -5400 35145 -5280
rect 35265 -5400 35310 -5280
rect 35430 -5400 35485 -5280
rect 35605 -5400 35650 -5280
rect 35770 -5400 35815 -5280
rect 35935 -5400 35980 -5280
rect 36100 -5400 36155 -5280
rect 36275 -5400 36285 -5280
rect 30785 -5445 36285 -5400
rect 30785 -5565 30795 -5445
rect 30915 -5565 30960 -5445
rect 31080 -5565 31125 -5445
rect 31245 -5565 31290 -5445
rect 31410 -5565 31465 -5445
rect 31585 -5565 31630 -5445
rect 31750 -5565 31795 -5445
rect 31915 -5565 31960 -5445
rect 32080 -5565 32135 -5445
rect 32255 -5565 32300 -5445
rect 32420 -5565 32465 -5445
rect 32585 -5565 32630 -5445
rect 32750 -5565 32805 -5445
rect 32925 -5565 32970 -5445
rect 33090 -5565 33135 -5445
rect 33255 -5565 33300 -5445
rect 33420 -5565 33475 -5445
rect 33595 -5565 33640 -5445
rect 33760 -5565 33805 -5445
rect 33925 -5565 33970 -5445
rect 34090 -5565 34145 -5445
rect 34265 -5565 34310 -5445
rect 34430 -5565 34475 -5445
rect 34595 -5565 34640 -5445
rect 34760 -5565 34815 -5445
rect 34935 -5565 34980 -5445
rect 35100 -5565 35145 -5445
rect 35265 -5565 35310 -5445
rect 35430 -5565 35485 -5445
rect 35605 -5565 35650 -5445
rect 35770 -5565 35815 -5445
rect 35935 -5565 35980 -5445
rect 36100 -5565 36155 -5445
rect 36275 -5565 36285 -5445
rect 30785 -5610 36285 -5565
rect 30785 -5730 30795 -5610
rect 30915 -5730 30960 -5610
rect 31080 -5730 31125 -5610
rect 31245 -5730 31290 -5610
rect 31410 -5730 31465 -5610
rect 31585 -5730 31630 -5610
rect 31750 -5730 31795 -5610
rect 31915 -5730 31960 -5610
rect 32080 -5730 32135 -5610
rect 32255 -5730 32300 -5610
rect 32420 -5730 32465 -5610
rect 32585 -5730 32630 -5610
rect 32750 -5730 32805 -5610
rect 32925 -5730 32970 -5610
rect 33090 -5730 33135 -5610
rect 33255 -5730 33300 -5610
rect 33420 -5730 33475 -5610
rect 33595 -5730 33640 -5610
rect 33760 -5730 33805 -5610
rect 33925 -5730 33970 -5610
rect 34090 -5730 34145 -5610
rect 34265 -5730 34310 -5610
rect 34430 -5730 34475 -5610
rect 34595 -5730 34640 -5610
rect 34760 -5730 34815 -5610
rect 34935 -5730 34980 -5610
rect 35100 -5730 35145 -5610
rect 35265 -5730 35310 -5610
rect 35430 -5730 35485 -5610
rect 35605 -5730 35650 -5610
rect 35770 -5730 35815 -5610
rect 35935 -5730 35980 -5610
rect 36100 -5730 36155 -5610
rect 36275 -5730 36285 -5610
rect 30785 -5785 36285 -5730
rect 30785 -5905 30795 -5785
rect 30915 -5905 30960 -5785
rect 31080 -5905 31125 -5785
rect 31245 -5905 31290 -5785
rect 31410 -5905 31465 -5785
rect 31585 -5905 31630 -5785
rect 31750 -5905 31795 -5785
rect 31915 -5905 31960 -5785
rect 32080 -5905 32135 -5785
rect 32255 -5905 32300 -5785
rect 32420 -5905 32465 -5785
rect 32585 -5905 32630 -5785
rect 32750 -5905 32805 -5785
rect 32925 -5905 32970 -5785
rect 33090 -5905 33135 -5785
rect 33255 -5905 33300 -5785
rect 33420 -5905 33475 -5785
rect 33595 -5905 33640 -5785
rect 33760 -5905 33805 -5785
rect 33925 -5905 33970 -5785
rect 34090 -5905 34145 -5785
rect 34265 -5905 34310 -5785
rect 34430 -5905 34475 -5785
rect 34595 -5905 34640 -5785
rect 34760 -5905 34815 -5785
rect 34935 -5905 34980 -5785
rect 35100 -5905 35145 -5785
rect 35265 -5905 35310 -5785
rect 35430 -5905 35485 -5785
rect 35605 -5905 35650 -5785
rect 35770 -5905 35815 -5785
rect 35935 -5905 35980 -5785
rect 36100 -5905 36155 -5785
rect 36275 -5905 36285 -5785
rect 30785 -5950 36285 -5905
rect 30785 -6070 30795 -5950
rect 30915 -6070 30960 -5950
rect 31080 -6070 31125 -5950
rect 31245 -6070 31290 -5950
rect 31410 -6070 31465 -5950
rect 31585 -6070 31630 -5950
rect 31750 -6070 31795 -5950
rect 31915 -6070 31960 -5950
rect 32080 -6070 32135 -5950
rect 32255 -6070 32300 -5950
rect 32420 -6070 32465 -5950
rect 32585 -6070 32630 -5950
rect 32750 -6070 32805 -5950
rect 32925 -6070 32970 -5950
rect 33090 -6070 33135 -5950
rect 33255 -6070 33300 -5950
rect 33420 -6070 33475 -5950
rect 33595 -6070 33640 -5950
rect 33760 -6070 33805 -5950
rect 33925 -6070 33970 -5950
rect 34090 -6070 34145 -5950
rect 34265 -6070 34310 -5950
rect 34430 -6070 34475 -5950
rect 34595 -6070 34640 -5950
rect 34760 -6070 34815 -5950
rect 34935 -6070 34980 -5950
rect 35100 -6070 35145 -5950
rect 35265 -6070 35310 -5950
rect 35430 -6070 35485 -5950
rect 35605 -6070 35650 -5950
rect 35770 -6070 35815 -5950
rect 35935 -6070 35980 -5950
rect 36100 -6070 36155 -5950
rect 36275 -6070 36285 -5950
rect 30785 -6115 36285 -6070
rect 30785 -6235 30795 -6115
rect 30915 -6235 30960 -6115
rect 31080 -6235 31125 -6115
rect 31245 -6235 31290 -6115
rect 31410 -6235 31465 -6115
rect 31585 -6235 31630 -6115
rect 31750 -6235 31795 -6115
rect 31915 -6235 31960 -6115
rect 32080 -6235 32135 -6115
rect 32255 -6235 32300 -6115
rect 32420 -6235 32465 -6115
rect 32585 -6235 32630 -6115
rect 32750 -6235 32805 -6115
rect 32925 -6235 32970 -6115
rect 33090 -6235 33135 -6115
rect 33255 -6235 33300 -6115
rect 33420 -6235 33475 -6115
rect 33595 -6235 33640 -6115
rect 33760 -6235 33805 -6115
rect 33925 -6235 33970 -6115
rect 34090 -6235 34145 -6115
rect 34265 -6235 34310 -6115
rect 34430 -6235 34475 -6115
rect 34595 -6235 34640 -6115
rect 34760 -6235 34815 -6115
rect 34935 -6235 34980 -6115
rect 35100 -6235 35145 -6115
rect 35265 -6235 35310 -6115
rect 35430 -6235 35485 -6115
rect 35605 -6235 35650 -6115
rect 35770 -6235 35815 -6115
rect 35935 -6235 35980 -6115
rect 36100 -6235 36155 -6115
rect 36275 -6235 36285 -6115
rect 30785 -6280 36285 -6235
rect 30785 -6400 30795 -6280
rect 30915 -6400 30960 -6280
rect 31080 -6400 31125 -6280
rect 31245 -6400 31290 -6280
rect 31410 -6400 31465 -6280
rect 31585 -6400 31630 -6280
rect 31750 -6400 31795 -6280
rect 31915 -6400 31960 -6280
rect 32080 -6400 32135 -6280
rect 32255 -6400 32300 -6280
rect 32420 -6400 32465 -6280
rect 32585 -6400 32630 -6280
rect 32750 -6400 32805 -6280
rect 32925 -6400 32970 -6280
rect 33090 -6400 33135 -6280
rect 33255 -6400 33300 -6280
rect 33420 -6400 33475 -6280
rect 33595 -6400 33640 -6280
rect 33760 -6400 33805 -6280
rect 33925 -6400 33970 -6280
rect 34090 -6400 34145 -6280
rect 34265 -6400 34310 -6280
rect 34430 -6400 34475 -6280
rect 34595 -6400 34640 -6280
rect 34760 -6400 34815 -6280
rect 34935 -6400 34980 -6280
rect 35100 -6400 35145 -6280
rect 35265 -6400 35310 -6280
rect 35430 -6400 35485 -6280
rect 35605 -6400 35650 -6280
rect 35770 -6400 35815 -6280
rect 35935 -6400 35980 -6280
rect 36100 -6400 36155 -6280
rect 36275 -6400 36285 -6280
rect 30785 -6455 36285 -6400
rect 30785 -6575 30795 -6455
rect 30915 -6575 30960 -6455
rect 31080 -6575 31125 -6455
rect 31245 -6575 31290 -6455
rect 31410 -6575 31465 -6455
rect 31585 -6575 31630 -6455
rect 31750 -6575 31795 -6455
rect 31915 -6575 31960 -6455
rect 32080 -6575 32135 -6455
rect 32255 -6575 32300 -6455
rect 32420 -6575 32465 -6455
rect 32585 -6575 32630 -6455
rect 32750 -6575 32805 -6455
rect 32925 -6575 32970 -6455
rect 33090 -6575 33135 -6455
rect 33255 -6575 33300 -6455
rect 33420 -6575 33475 -6455
rect 33595 -6575 33640 -6455
rect 33760 -6575 33805 -6455
rect 33925 -6575 33970 -6455
rect 34090 -6575 34145 -6455
rect 34265 -6575 34310 -6455
rect 34430 -6575 34475 -6455
rect 34595 -6575 34640 -6455
rect 34760 -6575 34815 -6455
rect 34935 -6575 34980 -6455
rect 35100 -6575 35145 -6455
rect 35265 -6575 35310 -6455
rect 35430 -6575 35485 -6455
rect 35605 -6575 35650 -6455
rect 35770 -6575 35815 -6455
rect 35935 -6575 35980 -6455
rect 36100 -6575 36155 -6455
rect 36275 -6575 36285 -6455
rect 30785 -6620 36285 -6575
rect 30785 -6740 30795 -6620
rect 30915 -6740 30960 -6620
rect 31080 -6740 31125 -6620
rect 31245 -6740 31290 -6620
rect 31410 -6740 31465 -6620
rect 31585 -6740 31630 -6620
rect 31750 -6740 31795 -6620
rect 31915 -6740 31960 -6620
rect 32080 -6740 32135 -6620
rect 32255 -6740 32300 -6620
rect 32420 -6740 32465 -6620
rect 32585 -6740 32630 -6620
rect 32750 -6740 32805 -6620
rect 32925 -6740 32970 -6620
rect 33090 -6740 33135 -6620
rect 33255 -6740 33300 -6620
rect 33420 -6740 33475 -6620
rect 33595 -6740 33640 -6620
rect 33760 -6740 33805 -6620
rect 33925 -6740 33970 -6620
rect 34090 -6740 34145 -6620
rect 34265 -6740 34310 -6620
rect 34430 -6740 34475 -6620
rect 34595 -6740 34640 -6620
rect 34760 -6740 34815 -6620
rect 34935 -6740 34980 -6620
rect 35100 -6740 35145 -6620
rect 35265 -6740 35310 -6620
rect 35430 -6740 35485 -6620
rect 35605 -6740 35650 -6620
rect 35770 -6740 35815 -6620
rect 35935 -6740 35980 -6620
rect 36100 -6740 36155 -6620
rect 36275 -6740 36285 -6620
rect 30785 -6785 36285 -6740
rect 30785 -6905 30795 -6785
rect 30915 -6905 30960 -6785
rect 31080 -6905 31125 -6785
rect 31245 -6905 31290 -6785
rect 31410 -6905 31465 -6785
rect 31585 -6905 31630 -6785
rect 31750 -6905 31795 -6785
rect 31915 -6905 31960 -6785
rect 32080 -6905 32135 -6785
rect 32255 -6905 32300 -6785
rect 32420 -6905 32465 -6785
rect 32585 -6905 32630 -6785
rect 32750 -6905 32805 -6785
rect 32925 -6905 32970 -6785
rect 33090 -6905 33135 -6785
rect 33255 -6905 33300 -6785
rect 33420 -6905 33475 -6785
rect 33595 -6905 33640 -6785
rect 33760 -6905 33805 -6785
rect 33925 -6905 33970 -6785
rect 34090 -6905 34145 -6785
rect 34265 -6905 34310 -6785
rect 34430 -6905 34475 -6785
rect 34595 -6905 34640 -6785
rect 34760 -6905 34815 -6785
rect 34935 -6905 34980 -6785
rect 35100 -6905 35145 -6785
rect 35265 -6905 35310 -6785
rect 35430 -6905 35485 -6785
rect 35605 -6905 35650 -6785
rect 35770 -6905 35815 -6785
rect 35935 -6905 35980 -6785
rect 36100 -6905 36155 -6785
rect 36275 -6905 36285 -6785
rect 30785 -6950 36285 -6905
rect 30785 -7070 30795 -6950
rect 30915 -7070 30960 -6950
rect 31080 -7070 31125 -6950
rect 31245 -7070 31290 -6950
rect 31410 -7070 31465 -6950
rect 31585 -7070 31630 -6950
rect 31750 -7070 31795 -6950
rect 31915 -7070 31960 -6950
rect 32080 -7070 32135 -6950
rect 32255 -7070 32300 -6950
rect 32420 -7070 32465 -6950
rect 32585 -7070 32630 -6950
rect 32750 -7070 32805 -6950
rect 32925 -7070 32970 -6950
rect 33090 -7070 33135 -6950
rect 33255 -7070 33300 -6950
rect 33420 -7070 33475 -6950
rect 33595 -7070 33640 -6950
rect 33760 -7070 33805 -6950
rect 33925 -7070 33970 -6950
rect 34090 -7070 34145 -6950
rect 34265 -7070 34310 -6950
rect 34430 -7070 34475 -6950
rect 34595 -7070 34640 -6950
rect 34760 -7070 34815 -6950
rect 34935 -7070 34980 -6950
rect 35100 -7070 35145 -6950
rect 35265 -7070 35310 -6950
rect 35430 -7070 35485 -6950
rect 35605 -7070 35650 -6950
rect 35770 -7070 35815 -6950
rect 35935 -7070 35980 -6950
rect 36100 -7070 36155 -6950
rect 36275 -7070 36285 -6950
rect 30785 -7125 36285 -7070
rect 30785 -7245 30795 -7125
rect 30915 -7245 30960 -7125
rect 31080 -7245 31125 -7125
rect 31245 -7245 31290 -7125
rect 31410 -7245 31465 -7125
rect 31585 -7245 31630 -7125
rect 31750 -7245 31795 -7125
rect 31915 -7245 31960 -7125
rect 32080 -7245 32135 -7125
rect 32255 -7245 32300 -7125
rect 32420 -7245 32465 -7125
rect 32585 -7245 32630 -7125
rect 32750 -7245 32805 -7125
rect 32925 -7245 32970 -7125
rect 33090 -7245 33135 -7125
rect 33255 -7245 33300 -7125
rect 33420 -7245 33475 -7125
rect 33595 -7245 33640 -7125
rect 33760 -7245 33805 -7125
rect 33925 -7245 33970 -7125
rect 34090 -7245 34145 -7125
rect 34265 -7245 34310 -7125
rect 34430 -7245 34475 -7125
rect 34595 -7245 34640 -7125
rect 34760 -7245 34815 -7125
rect 34935 -7245 34980 -7125
rect 35100 -7245 35145 -7125
rect 35265 -7245 35310 -7125
rect 35430 -7245 35485 -7125
rect 35605 -7245 35650 -7125
rect 35770 -7245 35815 -7125
rect 35935 -7245 35980 -7125
rect 36100 -7245 36155 -7125
rect 36275 -7245 36285 -7125
rect 30785 -7290 36285 -7245
rect 30785 -7410 30795 -7290
rect 30915 -7410 30960 -7290
rect 31080 -7410 31125 -7290
rect 31245 -7410 31290 -7290
rect 31410 -7410 31465 -7290
rect 31585 -7410 31630 -7290
rect 31750 -7410 31795 -7290
rect 31915 -7410 31960 -7290
rect 32080 -7410 32135 -7290
rect 32255 -7410 32300 -7290
rect 32420 -7410 32465 -7290
rect 32585 -7410 32630 -7290
rect 32750 -7410 32805 -7290
rect 32925 -7410 32970 -7290
rect 33090 -7410 33135 -7290
rect 33255 -7410 33300 -7290
rect 33420 -7410 33475 -7290
rect 33595 -7410 33640 -7290
rect 33760 -7410 33805 -7290
rect 33925 -7410 33970 -7290
rect 34090 -7410 34145 -7290
rect 34265 -7410 34310 -7290
rect 34430 -7410 34475 -7290
rect 34595 -7410 34640 -7290
rect 34760 -7410 34815 -7290
rect 34935 -7410 34980 -7290
rect 35100 -7410 35145 -7290
rect 35265 -7410 35310 -7290
rect 35430 -7410 35485 -7290
rect 35605 -7410 35650 -7290
rect 35770 -7410 35815 -7290
rect 35935 -7410 35980 -7290
rect 36100 -7410 36155 -7290
rect 36275 -7410 36285 -7290
rect 30785 -7455 36285 -7410
rect 30785 -7575 30795 -7455
rect 30915 -7575 30960 -7455
rect 31080 -7575 31125 -7455
rect 31245 -7575 31290 -7455
rect 31410 -7575 31465 -7455
rect 31585 -7575 31630 -7455
rect 31750 -7575 31795 -7455
rect 31915 -7575 31960 -7455
rect 32080 -7575 32135 -7455
rect 32255 -7575 32300 -7455
rect 32420 -7575 32465 -7455
rect 32585 -7575 32630 -7455
rect 32750 -7575 32805 -7455
rect 32925 -7575 32970 -7455
rect 33090 -7575 33135 -7455
rect 33255 -7575 33300 -7455
rect 33420 -7575 33475 -7455
rect 33595 -7575 33640 -7455
rect 33760 -7575 33805 -7455
rect 33925 -7575 33970 -7455
rect 34090 -7575 34145 -7455
rect 34265 -7575 34310 -7455
rect 34430 -7575 34475 -7455
rect 34595 -7575 34640 -7455
rect 34760 -7575 34815 -7455
rect 34935 -7575 34980 -7455
rect 35100 -7575 35145 -7455
rect 35265 -7575 35310 -7455
rect 35430 -7575 35485 -7455
rect 35605 -7575 35650 -7455
rect 35770 -7575 35815 -7455
rect 35935 -7575 35980 -7455
rect 36100 -7575 36155 -7455
rect 36275 -7575 36285 -7455
rect 30785 -7620 36285 -7575
rect 30785 -7740 30795 -7620
rect 30915 -7740 30960 -7620
rect 31080 -7740 31125 -7620
rect 31245 -7740 31290 -7620
rect 31410 -7740 31465 -7620
rect 31585 -7740 31630 -7620
rect 31750 -7740 31795 -7620
rect 31915 -7740 31960 -7620
rect 32080 -7740 32135 -7620
rect 32255 -7740 32300 -7620
rect 32420 -7740 32465 -7620
rect 32585 -7740 32630 -7620
rect 32750 -7740 32805 -7620
rect 32925 -7740 32970 -7620
rect 33090 -7740 33135 -7620
rect 33255 -7740 33300 -7620
rect 33420 -7740 33475 -7620
rect 33595 -7740 33640 -7620
rect 33760 -7740 33805 -7620
rect 33925 -7740 33970 -7620
rect 34090 -7740 34145 -7620
rect 34265 -7740 34310 -7620
rect 34430 -7740 34475 -7620
rect 34595 -7740 34640 -7620
rect 34760 -7740 34815 -7620
rect 34935 -7740 34980 -7620
rect 35100 -7740 35145 -7620
rect 35265 -7740 35310 -7620
rect 35430 -7740 35485 -7620
rect 35605 -7740 35650 -7620
rect 35770 -7740 35815 -7620
rect 35935 -7740 35980 -7620
rect 36100 -7740 36155 -7620
rect 36275 -7740 36285 -7620
rect 30785 -7795 36285 -7740
rect 30785 -7915 30795 -7795
rect 30915 -7915 30960 -7795
rect 31080 -7915 31125 -7795
rect 31245 -7915 31290 -7795
rect 31410 -7915 31465 -7795
rect 31585 -7915 31630 -7795
rect 31750 -7915 31795 -7795
rect 31915 -7915 31960 -7795
rect 32080 -7915 32135 -7795
rect 32255 -7915 32300 -7795
rect 32420 -7915 32465 -7795
rect 32585 -7915 32630 -7795
rect 32750 -7915 32805 -7795
rect 32925 -7915 32970 -7795
rect 33090 -7915 33135 -7795
rect 33255 -7915 33300 -7795
rect 33420 -7915 33475 -7795
rect 33595 -7915 33640 -7795
rect 33760 -7915 33805 -7795
rect 33925 -7915 33970 -7795
rect 34090 -7915 34145 -7795
rect 34265 -7915 34310 -7795
rect 34430 -7915 34475 -7795
rect 34595 -7915 34640 -7795
rect 34760 -7915 34815 -7795
rect 34935 -7915 34980 -7795
rect 35100 -7915 35145 -7795
rect 35265 -7915 35310 -7795
rect 35430 -7915 35485 -7795
rect 35605 -7915 35650 -7795
rect 35770 -7915 35815 -7795
rect 35935 -7915 35980 -7795
rect 36100 -7915 36155 -7795
rect 36275 -7915 36285 -7795
rect 30785 -7960 36285 -7915
rect 30785 -8080 30795 -7960
rect 30915 -8080 30960 -7960
rect 31080 -8080 31125 -7960
rect 31245 -8080 31290 -7960
rect 31410 -8080 31465 -7960
rect 31585 -8080 31630 -7960
rect 31750 -8080 31795 -7960
rect 31915 -8080 31960 -7960
rect 32080 -8080 32135 -7960
rect 32255 -8080 32300 -7960
rect 32420 -8080 32465 -7960
rect 32585 -8080 32630 -7960
rect 32750 -8080 32805 -7960
rect 32925 -8080 32970 -7960
rect 33090 -8080 33135 -7960
rect 33255 -8080 33300 -7960
rect 33420 -8080 33475 -7960
rect 33595 -8080 33640 -7960
rect 33760 -8080 33805 -7960
rect 33925 -8080 33970 -7960
rect 34090 -8080 34145 -7960
rect 34265 -8080 34310 -7960
rect 34430 -8080 34475 -7960
rect 34595 -8080 34640 -7960
rect 34760 -8080 34815 -7960
rect 34935 -8080 34980 -7960
rect 35100 -8080 35145 -7960
rect 35265 -8080 35310 -7960
rect 35430 -8080 35485 -7960
rect 35605 -8080 35650 -7960
rect 35770 -8080 35815 -7960
rect 35935 -8080 35980 -7960
rect 36100 -8080 36155 -7960
rect 36275 -8080 36285 -7960
rect 30785 -8125 36285 -8080
rect 30785 -8245 30795 -8125
rect 30915 -8245 30960 -8125
rect 31080 -8245 31125 -8125
rect 31245 -8245 31290 -8125
rect 31410 -8245 31465 -8125
rect 31585 -8245 31630 -8125
rect 31750 -8245 31795 -8125
rect 31915 -8245 31960 -8125
rect 32080 -8245 32135 -8125
rect 32255 -8245 32300 -8125
rect 32420 -8245 32465 -8125
rect 32585 -8245 32630 -8125
rect 32750 -8245 32805 -8125
rect 32925 -8245 32970 -8125
rect 33090 -8245 33135 -8125
rect 33255 -8245 33300 -8125
rect 33420 -8245 33475 -8125
rect 33595 -8245 33640 -8125
rect 33760 -8245 33805 -8125
rect 33925 -8245 33970 -8125
rect 34090 -8245 34145 -8125
rect 34265 -8245 34310 -8125
rect 34430 -8245 34475 -8125
rect 34595 -8245 34640 -8125
rect 34760 -8245 34815 -8125
rect 34935 -8245 34980 -8125
rect 35100 -8245 35145 -8125
rect 35265 -8245 35310 -8125
rect 35430 -8245 35485 -8125
rect 35605 -8245 35650 -8125
rect 35770 -8245 35815 -8125
rect 35935 -8245 35980 -8125
rect 36100 -8245 36155 -8125
rect 36275 -8245 36285 -8125
rect 30785 -8290 36285 -8245
rect 30785 -8410 30795 -8290
rect 30915 -8410 30960 -8290
rect 31080 -8410 31125 -8290
rect 31245 -8410 31290 -8290
rect 31410 -8410 31465 -8290
rect 31585 -8410 31630 -8290
rect 31750 -8410 31795 -8290
rect 31915 -8410 31960 -8290
rect 32080 -8410 32135 -8290
rect 32255 -8410 32300 -8290
rect 32420 -8410 32465 -8290
rect 32585 -8410 32630 -8290
rect 32750 -8410 32805 -8290
rect 32925 -8410 32970 -8290
rect 33090 -8410 33135 -8290
rect 33255 -8410 33300 -8290
rect 33420 -8410 33475 -8290
rect 33595 -8410 33640 -8290
rect 33760 -8410 33805 -8290
rect 33925 -8410 33970 -8290
rect 34090 -8410 34145 -8290
rect 34265 -8410 34310 -8290
rect 34430 -8410 34475 -8290
rect 34595 -8410 34640 -8290
rect 34760 -8410 34815 -8290
rect 34935 -8410 34980 -8290
rect 35100 -8410 35145 -8290
rect 35265 -8410 35310 -8290
rect 35430 -8410 35485 -8290
rect 35605 -8410 35650 -8290
rect 35770 -8410 35815 -8290
rect 35935 -8410 35980 -8290
rect 36100 -8410 36155 -8290
rect 36275 -8410 36285 -8290
rect 30785 -8465 36285 -8410
rect 30785 -8585 30795 -8465
rect 30915 -8585 30960 -8465
rect 31080 -8585 31125 -8465
rect 31245 -8585 31290 -8465
rect 31410 -8585 31465 -8465
rect 31585 -8585 31630 -8465
rect 31750 -8585 31795 -8465
rect 31915 -8585 31960 -8465
rect 32080 -8585 32135 -8465
rect 32255 -8585 32300 -8465
rect 32420 -8585 32465 -8465
rect 32585 -8585 32630 -8465
rect 32750 -8585 32805 -8465
rect 32925 -8585 32970 -8465
rect 33090 -8585 33135 -8465
rect 33255 -8585 33300 -8465
rect 33420 -8585 33475 -8465
rect 33595 -8585 33640 -8465
rect 33760 -8585 33805 -8465
rect 33925 -8585 33970 -8465
rect 34090 -8585 34145 -8465
rect 34265 -8585 34310 -8465
rect 34430 -8585 34475 -8465
rect 34595 -8585 34640 -8465
rect 34760 -8585 34815 -8465
rect 34935 -8585 34980 -8465
rect 35100 -8585 35145 -8465
rect 35265 -8585 35310 -8465
rect 35430 -8585 35485 -8465
rect 35605 -8585 35650 -8465
rect 35770 -8585 35815 -8465
rect 35935 -8585 35980 -8465
rect 36100 -8585 36155 -8465
rect 36275 -8585 36285 -8465
rect 30785 -8630 36285 -8585
rect 30785 -8750 30795 -8630
rect 30915 -8750 30960 -8630
rect 31080 -8750 31125 -8630
rect 31245 -8750 31290 -8630
rect 31410 -8750 31465 -8630
rect 31585 -8750 31630 -8630
rect 31750 -8750 31795 -8630
rect 31915 -8750 31960 -8630
rect 32080 -8750 32135 -8630
rect 32255 -8750 32300 -8630
rect 32420 -8750 32465 -8630
rect 32585 -8750 32630 -8630
rect 32750 -8750 32805 -8630
rect 32925 -8750 32970 -8630
rect 33090 -8750 33135 -8630
rect 33255 -8750 33300 -8630
rect 33420 -8750 33475 -8630
rect 33595 -8750 33640 -8630
rect 33760 -8750 33805 -8630
rect 33925 -8750 33970 -8630
rect 34090 -8750 34145 -8630
rect 34265 -8750 34310 -8630
rect 34430 -8750 34475 -8630
rect 34595 -8750 34640 -8630
rect 34760 -8750 34815 -8630
rect 34935 -8750 34980 -8630
rect 35100 -8750 35145 -8630
rect 35265 -8750 35310 -8630
rect 35430 -8750 35485 -8630
rect 35605 -8750 35650 -8630
rect 35770 -8750 35815 -8630
rect 35935 -8750 35980 -8630
rect 36100 -8750 36155 -8630
rect 36275 -8750 36285 -8630
rect 30785 -8795 36285 -8750
rect 30785 -8915 30795 -8795
rect 30915 -8915 30960 -8795
rect 31080 -8915 31125 -8795
rect 31245 -8915 31290 -8795
rect 31410 -8915 31465 -8795
rect 31585 -8915 31630 -8795
rect 31750 -8915 31795 -8795
rect 31915 -8915 31960 -8795
rect 32080 -8915 32135 -8795
rect 32255 -8915 32300 -8795
rect 32420 -8915 32465 -8795
rect 32585 -8915 32630 -8795
rect 32750 -8915 32805 -8795
rect 32925 -8915 32970 -8795
rect 33090 -8915 33135 -8795
rect 33255 -8915 33300 -8795
rect 33420 -8915 33475 -8795
rect 33595 -8915 33640 -8795
rect 33760 -8915 33805 -8795
rect 33925 -8915 33970 -8795
rect 34090 -8915 34145 -8795
rect 34265 -8915 34310 -8795
rect 34430 -8915 34475 -8795
rect 34595 -8915 34640 -8795
rect 34760 -8915 34815 -8795
rect 34935 -8915 34980 -8795
rect 35100 -8915 35145 -8795
rect 35265 -8915 35310 -8795
rect 35430 -8915 35485 -8795
rect 35605 -8915 35650 -8795
rect 35770 -8915 35815 -8795
rect 35935 -8915 35980 -8795
rect 36100 -8915 36155 -8795
rect 36275 -8915 36285 -8795
rect 30785 -8960 36285 -8915
rect 30785 -9080 30795 -8960
rect 30915 -9080 30960 -8960
rect 31080 -9080 31125 -8960
rect 31245 -9080 31290 -8960
rect 31410 -9080 31465 -8960
rect 31585 -9080 31630 -8960
rect 31750 -9080 31795 -8960
rect 31915 -9080 31960 -8960
rect 32080 -9080 32135 -8960
rect 32255 -9080 32300 -8960
rect 32420 -9080 32465 -8960
rect 32585 -9080 32630 -8960
rect 32750 -9080 32805 -8960
rect 32925 -9080 32970 -8960
rect 33090 -9080 33135 -8960
rect 33255 -9080 33300 -8960
rect 33420 -9080 33475 -8960
rect 33595 -9080 33640 -8960
rect 33760 -9080 33805 -8960
rect 33925 -9080 33970 -8960
rect 34090 -9080 34145 -8960
rect 34265 -9080 34310 -8960
rect 34430 -9080 34475 -8960
rect 34595 -9080 34640 -8960
rect 34760 -9080 34815 -8960
rect 34935 -9080 34980 -8960
rect 35100 -9080 35145 -8960
rect 35265 -9080 35310 -8960
rect 35430 -9080 35485 -8960
rect 35605 -9080 35650 -8960
rect 35770 -9080 35815 -8960
rect 35935 -9080 35980 -8960
rect 36100 -9080 36155 -8960
rect 36275 -9080 36285 -8960
rect 30785 -9135 36285 -9080
rect 30785 -9255 30795 -9135
rect 30915 -9255 30960 -9135
rect 31080 -9255 31125 -9135
rect 31245 -9255 31290 -9135
rect 31410 -9255 31465 -9135
rect 31585 -9255 31630 -9135
rect 31750 -9255 31795 -9135
rect 31915 -9255 31960 -9135
rect 32080 -9255 32135 -9135
rect 32255 -9255 32300 -9135
rect 32420 -9255 32465 -9135
rect 32585 -9255 32630 -9135
rect 32750 -9255 32805 -9135
rect 32925 -9255 32970 -9135
rect 33090 -9255 33135 -9135
rect 33255 -9255 33300 -9135
rect 33420 -9255 33475 -9135
rect 33595 -9255 33640 -9135
rect 33760 -9255 33805 -9135
rect 33925 -9255 33970 -9135
rect 34090 -9255 34145 -9135
rect 34265 -9255 34310 -9135
rect 34430 -9255 34475 -9135
rect 34595 -9255 34640 -9135
rect 34760 -9255 34815 -9135
rect 34935 -9255 34980 -9135
rect 35100 -9255 35145 -9135
rect 35265 -9255 35310 -9135
rect 35430 -9255 35485 -9135
rect 35605 -9255 35650 -9135
rect 35770 -9255 35815 -9135
rect 35935 -9255 35980 -9135
rect 36100 -9255 36155 -9135
rect 36275 -9255 36285 -9135
rect 30785 -9300 36285 -9255
rect 30785 -9420 30795 -9300
rect 30915 -9420 30960 -9300
rect 31080 -9420 31125 -9300
rect 31245 -9420 31290 -9300
rect 31410 -9420 31465 -9300
rect 31585 -9420 31630 -9300
rect 31750 -9420 31795 -9300
rect 31915 -9420 31960 -9300
rect 32080 -9420 32135 -9300
rect 32255 -9420 32300 -9300
rect 32420 -9420 32465 -9300
rect 32585 -9420 32630 -9300
rect 32750 -9420 32805 -9300
rect 32925 -9420 32970 -9300
rect 33090 -9420 33135 -9300
rect 33255 -9420 33300 -9300
rect 33420 -9420 33475 -9300
rect 33595 -9420 33640 -9300
rect 33760 -9420 33805 -9300
rect 33925 -9420 33970 -9300
rect 34090 -9420 34145 -9300
rect 34265 -9420 34310 -9300
rect 34430 -9420 34475 -9300
rect 34595 -9420 34640 -9300
rect 34760 -9420 34815 -9300
rect 34935 -9420 34980 -9300
rect 35100 -9420 35145 -9300
rect 35265 -9420 35310 -9300
rect 35430 -9420 35485 -9300
rect 35605 -9420 35650 -9300
rect 35770 -9420 35815 -9300
rect 35935 -9420 35980 -9300
rect 36100 -9420 36155 -9300
rect 36275 -9420 36285 -9300
rect 30785 -9465 36285 -9420
rect 30785 -9585 30795 -9465
rect 30915 -9585 30960 -9465
rect 31080 -9585 31125 -9465
rect 31245 -9585 31290 -9465
rect 31410 -9585 31465 -9465
rect 31585 -9585 31630 -9465
rect 31750 -9585 31795 -9465
rect 31915 -9585 31960 -9465
rect 32080 -9585 32135 -9465
rect 32255 -9585 32300 -9465
rect 32420 -9585 32465 -9465
rect 32585 -9585 32630 -9465
rect 32750 -9585 32805 -9465
rect 32925 -9585 32970 -9465
rect 33090 -9585 33135 -9465
rect 33255 -9585 33300 -9465
rect 33420 -9585 33475 -9465
rect 33595 -9585 33640 -9465
rect 33760 -9585 33805 -9465
rect 33925 -9585 33970 -9465
rect 34090 -9585 34145 -9465
rect 34265 -9585 34310 -9465
rect 34430 -9585 34475 -9465
rect 34595 -9585 34640 -9465
rect 34760 -9585 34815 -9465
rect 34935 -9585 34980 -9465
rect 35100 -9585 35145 -9465
rect 35265 -9585 35310 -9465
rect 35430 -9585 35485 -9465
rect 35605 -9585 35650 -9465
rect 35770 -9585 35815 -9465
rect 35935 -9585 35980 -9465
rect 36100 -9585 36155 -9465
rect 36275 -9585 36285 -9465
rect 30785 -9630 36285 -9585
rect 30785 -9750 30795 -9630
rect 30915 -9750 30960 -9630
rect 31080 -9750 31125 -9630
rect 31245 -9750 31290 -9630
rect 31410 -9750 31465 -9630
rect 31585 -9750 31630 -9630
rect 31750 -9750 31795 -9630
rect 31915 -9750 31960 -9630
rect 32080 -9750 32135 -9630
rect 32255 -9750 32300 -9630
rect 32420 -9750 32465 -9630
rect 32585 -9750 32630 -9630
rect 32750 -9750 32805 -9630
rect 32925 -9750 32970 -9630
rect 33090 -9750 33135 -9630
rect 33255 -9750 33300 -9630
rect 33420 -9750 33475 -9630
rect 33595 -9750 33640 -9630
rect 33760 -9750 33805 -9630
rect 33925 -9750 33970 -9630
rect 34090 -9750 34145 -9630
rect 34265 -9750 34310 -9630
rect 34430 -9750 34475 -9630
rect 34595 -9750 34640 -9630
rect 34760 -9750 34815 -9630
rect 34935 -9750 34980 -9630
rect 35100 -9750 35145 -9630
rect 35265 -9750 35310 -9630
rect 35430 -9750 35485 -9630
rect 35605 -9750 35650 -9630
rect 35770 -9750 35815 -9630
rect 35935 -9750 35980 -9630
rect 36100 -9750 36155 -9630
rect 36275 -9750 36285 -9630
rect 30785 -9760 36285 -9750
rect 36475 -4270 41975 -4260
rect 36475 -4390 36485 -4270
rect 36605 -4390 36650 -4270
rect 36770 -4390 36815 -4270
rect 36935 -4390 36980 -4270
rect 37100 -4390 37155 -4270
rect 37275 -4390 37320 -4270
rect 37440 -4390 37485 -4270
rect 37605 -4390 37650 -4270
rect 37770 -4390 37825 -4270
rect 37945 -4390 37990 -4270
rect 38110 -4390 38155 -4270
rect 38275 -4390 38320 -4270
rect 38440 -4390 38495 -4270
rect 38615 -4390 38660 -4270
rect 38780 -4390 38825 -4270
rect 38945 -4390 38990 -4270
rect 39110 -4390 39165 -4270
rect 39285 -4390 39330 -4270
rect 39450 -4390 39495 -4270
rect 39615 -4390 39660 -4270
rect 39780 -4390 39835 -4270
rect 39955 -4390 40000 -4270
rect 40120 -4390 40165 -4270
rect 40285 -4390 40330 -4270
rect 40450 -4390 40505 -4270
rect 40625 -4390 40670 -4270
rect 40790 -4390 40835 -4270
rect 40955 -4390 41000 -4270
rect 41120 -4390 41175 -4270
rect 41295 -4390 41340 -4270
rect 41460 -4390 41505 -4270
rect 41625 -4390 41670 -4270
rect 41790 -4390 41845 -4270
rect 41965 -4390 41975 -4270
rect 36475 -4445 41975 -4390
rect 36475 -4565 36485 -4445
rect 36605 -4565 36650 -4445
rect 36770 -4565 36815 -4445
rect 36935 -4565 36980 -4445
rect 37100 -4565 37155 -4445
rect 37275 -4565 37320 -4445
rect 37440 -4565 37485 -4445
rect 37605 -4565 37650 -4445
rect 37770 -4565 37825 -4445
rect 37945 -4565 37990 -4445
rect 38110 -4565 38155 -4445
rect 38275 -4565 38320 -4445
rect 38440 -4565 38495 -4445
rect 38615 -4565 38660 -4445
rect 38780 -4565 38825 -4445
rect 38945 -4565 38990 -4445
rect 39110 -4565 39165 -4445
rect 39285 -4565 39330 -4445
rect 39450 -4565 39495 -4445
rect 39615 -4565 39660 -4445
rect 39780 -4565 39835 -4445
rect 39955 -4565 40000 -4445
rect 40120 -4565 40165 -4445
rect 40285 -4565 40330 -4445
rect 40450 -4565 40505 -4445
rect 40625 -4565 40670 -4445
rect 40790 -4565 40835 -4445
rect 40955 -4565 41000 -4445
rect 41120 -4565 41175 -4445
rect 41295 -4565 41340 -4445
rect 41460 -4565 41505 -4445
rect 41625 -4565 41670 -4445
rect 41790 -4565 41845 -4445
rect 41965 -4565 41975 -4445
rect 36475 -4610 41975 -4565
rect 36475 -4730 36485 -4610
rect 36605 -4730 36650 -4610
rect 36770 -4730 36815 -4610
rect 36935 -4730 36980 -4610
rect 37100 -4730 37155 -4610
rect 37275 -4730 37320 -4610
rect 37440 -4730 37485 -4610
rect 37605 -4730 37650 -4610
rect 37770 -4730 37825 -4610
rect 37945 -4730 37990 -4610
rect 38110 -4730 38155 -4610
rect 38275 -4730 38320 -4610
rect 38440 -4730 38495 -4610
rect 38615 -4730 38660 -4610
rect 38780 -4730 38825 -4610
rect 38945 -4730 38990 -4610
rect 39110 -4730 39165 -4610
rect 39285 -4730 39330 -4610
rect 39450 -4730 39495 -4610
rect 39615 -4730 39660 -4610
rect 39780 -4730 39835 -4610
rect 39955 -4730 40000 -4610
rect 40120 -4730 40165 -4610
rect 40285 -4730 40330 -4610
rect 40450 -4730 40505 -4610
rect 40625 -4730 40670 -4610
rect 40790 -4730 40835 -4610
rect 40955 -4730 41000 -4610
rect 41120 -4730 41175 -4610
rect 41295 -4730 41340 -4610
rect 41460 -4730 41505 -4610
rect 41625 -4730 41670 -4610
rect 41790 -4730 41845 -4610
rect 41965 -4730 41975 -4610
rect 36475 -4775 41975 -4730
rect 36475 -4895 36485 -4775
rect 36605 -4895 36650 -4775
rect 36770 -4895 36815 -4775
rect 36935 -4895 36980 -4775
rect 37100 -4895 37155 -4775
rect 37275 -4895 37320 -4775
rect 37440 -4895 37485 -4775
rect 37605 -4895 37650 -4775
rect 37770 -4895 37825 -4775
rect 37945 -4895 37990 -4775
rect 38110 -4895 38155 -4775
rect 38275 -4895 38320 -4775
rect 38440 -4895 38495 -4775
rect 38615 -4895 38660 -4775
rect 38780 -4895 38825 -4775
rect 38945 -4895 38990 -4775
rect 39110 -4895 39165 -4775
rect 39285 -4895 39330 -4775
rect 39450 -4895 39495 -4775
rect 39615 -4895 39660 -4775
rect 39780 -4895 39835 -4775
rect 39955 -4895 40000 -4775
rect 40120 -4895 40165 -4775
rect 40285 -4895 40330 -4775
rect 40450 -4895 40505 -4775
rect 40625 -4895 40670 -4775
rect 40790 -4895 40835 -4775
rect 40955 -4895 41000 -4775
rect 41120 -4895 41175 -4775
rect 41295 -4895 41340 -4775
rect 41460 -4895 41505 -4775
rect 41625 -4895 41670 -4775
rect 41790 -4895 41845 -4775
rect 41965 -4895 41975 -4775
rect 36475 -4940 41975 -4895
rect 36475 -5060 36485 -4940
rect 36605 -5060 36650 -4940
rect 36770 -5060 36815 -4940
rect 36935 -5060 36980 -4940
rect 37100 -5060 37155 -4940
rect 37275 -5060 37320 -4940
rect 37440 -5060 37485 -4940
rect 37605 -5060 37650 -4940
rect 37770 -5060 37825 -4940
rect 37945 -5060 37990 -4940
rect 38110 -5060 38155 -4940
rect 38275 -5060 38320 -4940
rect 38440 -5060 38495 -4940
rect 38615 -5060 38660 -4940
rect 38780 -5060 38825 -4940
rect 38945 -5060 38990 -4940
rect 39110 -5060 39165 -4940
rect 39285 -5060 39330 -4940
rect 39450 -5060 39495 -4940
rect 39615 -5060 39660 -4940
rect 39780 -5060 39835 -4940
rect 39955 -5060 40000 -4940
rect 40120 -5060 40165 -4940
rect 40285 -5060 40330 -4940
rect 40450 -5060 40505 -4940
rect 40625 -5060 40670 -4940
rect 40790 -5060 40835 -4940
rect 40955 -5060 41000 -4940
rect 41120 -5060 41175 -4940
rect 41295 -5060 41340 -4940
rect 41460 -5060 41505 -4940
rect 41625 -5060 41670 -4940
rect 41790 -5060 41845 -4940
rect 41965 -5060 41975 -4940
rect 36475 -5115 41975 -5060
rect 36475 -5235 36485 -5115
rect 36605 -5235 36650 -5115
rect 36770 -5235 36815 -5115
rect 36935 -5235 36980 -5115
rect 37100 -5235 37155 -5115
rect 37275 -5235 37320 -5115
rect 37440 -5235 37485 -5115
rect 37605 -5235 37650 -5115
rect 37770 -5235 37825 -5115
rect 37945 -5235 37990 -5115
rect 38110 -5235 38155 -5115
rect 38275 -5235 38320 -5115
rect 38440 -5235 38495 -5115
rect 38615 -5235 38660 -5115
rect 38780 -5235 38825 -5115
rect 38945 -5235 38990 -5115
rect 39110 -5235 39165 -5115
rect 39285 -5235 39330 -5115
rect 39450 -5235 39495 -5115
rect 39615 -5235 39660 -5115
rect 39780 -5235 39835 -5115
rect 39955 -5235 40000 -5115
rect 40120 -5235 40165 -5115
rect 40285 -5235 40330 -5115
rect 40450 -5235 40505 -5115
rect 40625 -5235 40670 -5115
rect 40790 -5235 40835 -5115
rect 40955 -5235 41000 -5115
rect 41120 -5235 41175 -5115
rect 41295 -5235 41340 -5115
rect 41460 -5235 41505 -5115
rect 41625 -5235 41670 -5115
rect 41790 -5235 41845 -5115
rect 41965 -5235 41975 -5115
rect 36475 -5280 41975 -5235
rect 36475 -5400 36485 -5280
rect 36605 -5400 36650 -5280
rect 36770 -5400 36815 -5280
rect 36935 -5400 36980 -5280
rect 37100 -5400 37155 -5280
rect 37275 -5400 37320 -5280
rect 37440 -5400 37485 -5280
rect 37605 -5400 37650 -5280
rect 37770 -5400 37825 -5280
rect 37945 -5400 37990 -5280
rect 38110 -5400 38155 -5280
rect 38275 -5400 38320 -5280
rect 38440 -5400 38495 -5280
rect 38615 -5400 38660 -5280
rect 38780 -5400 38825 -5280
rect 38945 -5400 38990 -5280
rect 39110 -5400 39165 -5280
rect 39285 -5400 39330 -5280
rect 39450 -5400 39495 -5280
rect 39615 -5400 39660 -5280
rect 39780 -5400 39835 -5280
rect 39955 -5400 40000 -5280
rect 40120 -5400 40165 -5280
rect 40285 -5400 40330 -5280
rect 40450 -5400 40505 -5280
rect 40625 -5400 40670 -5280
rect 40790 -5400 40835 -5280
rect 40955 -5400 41000 -5280
rect 41120 -5400 41175 -5280
rect 41295 -5400 41340 -5280
rect 41460 -5400 41505 -5280
rect 41625 -5400 41670 -5280
rect 41790 -5400 41845 -5280
rect 41965 -5400 41975 -5280
rect 36475 -5445 41975 -5400
rect 36475 -5565 36485 -5445
rect 36605 -5565 36650 -5445
rect 36770 -5565 36815 -5445
rect 36935 -5565 36980 -5445
rect 37100 -5565 37155 -5445
rect 37275 -5565 37320 -5445
rect 37440 -5565 37485 -5445
rect 37605 -5565 37650 -5445
rect 37770 -5565 37825 -5445
rect 37945 -5565 37990 -5445
rect 38110 -5565 38155 -5445
rect 38275 -5565 38320 -5445
rect 38440 -5565 38495 -5445
rect 38615 -5565 38660 -5445
rect 38780 -5565 38825 -5445
rect 38945 -5565 38990 -5445
rect 39110 -5565 39165 -5445
rect 39285 -5565 39330 -5445
rect 39450 -5565 39495 -5445
rect 39615 -5565 39660 -5445
rect 39780 -5565 39835 -5445
rect 39955 -5565 40000 -5445
rect 40120 -5565 40165 -5445
rect 40285 -5565 40330 -5445
rect 40450 -5565 40505 -5445
rect 40625 -5565 40670 -5445
rect 40790 -5565 40835 -5445
rect 40955 -5565 41000 -5445
rect 41120 -5565 41175 -5445
rect 41295 -5565 41340 -5445
rect 41460 -5565 41505 -5445
rect 41625 -5565 41670 -5445
rect 41790 -5565 41845 -5445
rect 41965 -5565 41975 -5445
rect 36475 -5610 41975 -5565
rect 36475 -5730 36485 -5610
rect 36605 -5730 36650 -5610
rect 36770 -5730 36815 -5610
rect 36935 -5730 36980 -5610
rect 37100 -5730 37155 -5610
rect 37275 -5730 37320 -5610
rect 37440 -5730 37485 -5610
rect 37605 -5730 37650 -5610
rect 37770 -5730 37825 -5610
rect 37945 -5730 37990 -5610
rect 38110 -5730 38155 -5610
rect 38275 -5730 38320 -5610
rect 38440 -5730 38495 -5610
rect 38615 -5730 38660 -5610
rect 38780 -5730 38825 -5610
rect 38945 -5730 38990 -5610
rect 39110 -5730 39165 -5610
rect 39285 -5730 39330 -5610
rect 39450 -5730 39495 -5610
rect 39615 -5730 39660 -5610
rect 39780 -5730 39835 -5610
rect 39955 -5730 40000 -5610
rect 40120 -5730 40165 -5610
rect 40285 -5730 40330 -5610
rect 40450 -5730 40505 -5610
rect 40625 -5730 40670 -5610
rect 40790 -5730 40835 -5610
rect 40955 -5730 41000 -5610
rect 41120 -5730 41175 -5610
rect 41295 -5730 41340 -5610
rect 41460 -5730 41505 -5610
rect 41625 -5730 41670 -5610
rect 41790 -5730 41845 -5610
rect 41965 -5730 41975 -5610
rect 36475 -5785 41975 -5730
rect 36475 -5905 36485 -5785
rect 36605 -5905 36650 -5785
rect 36770 -5905 36815 -5785
rect 36935 -5905 36980 -5785
rect 37100 -5905 37155 -5785
rect 37275 -5905 37320 -5785
rect 37440 -5905 37485 -5785
rect 37605 -5905 37650 -5785
rect 37770 -5905 37825 -5785
rect 37945 -5905 37990 -5785
rect 38110 -5905 38155 -5785
rect 38275 -5905 38320 -5785
rect 38440 -5905 38495 -5785
rect 38615 -5905 38660 -5785
rect 38780 -5905 38825 -5785
rect 38945 -5905 38990 -5785
rect 39110 -5905 39165 -5785
rect 39285 -5905 39330 -5785
rect 39450 -5905 39495 -5785
rect 39615 -5905 39660 -5785
rect 39780 -5905 39835 -5785
rect 39955 -5905 40000 -5785
rect 40120 -5905 40165 -5785
rect 40285 -5905 40330 -5785
rect 40450 -5905 40505 -5785
rect 40625 -5905 40670 -5785
rect 40790 -5905 40835 -5785
rect 40955 -5905 41000 -5785
rect 41120 -5905 41175 -5785
rect 41295 -5905 41340 -5785
rect 41460 -5905 41505 -5785
rect 41625 -5905 41670 -5785
rect 41790 -5905 41845 -5785
rect 41965 -5905 41975 -5785
rect 36475 -5950 41975 -5905
rect 36475 -6070 36485 -5950
rect 36605 -6070 36650 -5950
rect 36770 -6070 36815 -5950
rect 36935 -6070 36980 -5950
rect 37100 -6070 37155 -5950
rect 37275 -6070 37320 -5950
rect 37440 -6070 37485 -5950
rect 37605 -6070 37650 -5950
rect 37770 -6070 37825 -5950
rect 37945 -6070 37990 -5950
rect 38110 -6070 38155 -5950
rect 38275 -6070 38320 -5950
rect 38440 -6070 38495 -5950
rect 38615 -6070 38660 -5950
rect 38780 -6070 38825 -5950
rect 38945 -6070 38990 -5950
rect 39110 -6070 39165 -5950
rect 39285 -6070 39330 -5950
rect 39450 -6070 39495 -5950
rect 39615 -6070 39660 -5950
rect 39780 -6070 39835 -5950
rect 39955 -6070 40000 -5950
rect 40120 -6070 40165 -5950
rect 40285 -6070 40330 -5950
rect 40450 -6070 40505 -5950
rect 40625 -6070 40670 -5950
rect 40790 -6070 40835 -5950
rect 40955 -6070 41000 -5950
rect 41120 -6070 41175 -5950
rect 41295 -6070 41340 -5950
rect 41460 -6070 41505 -5950
rect 41625 -6070 41670 -5950
rect 41790 -6070 41845 -5950
rect 41965 -6070 41975 -5950
rect 36475 -6115 41975 -6070
rect 36475 -6235 36485 -6115
rect 36605 -6235 36650 -6115
rect 36770 -6235 36815 -6115
rect 36935 -6235 36980 -6115
rect 37100 -6235 37155 -6115
rect 37275 -6235 37320 -6115
rect 37440 -6235 37485 -6115
rect 37605 -6235 37650 -6115
rect 37770 -6235 37825 -6115
rect 37945 -6235 37990 -6115
rect 38110 -6235 38155 -6115
rect 38275 -6235 38320 -6115
rect 38440 -6235 38495 -6115
rect 38615 -6235 38660 -6115
rect 38780 -6235 38825 -6115
rect 38945 -6235 38990 -6115
rect 39110 -6235 39165 -6115
rect 39285 -6235 39330 -6115
rect 39450 -6235 39495 -6115
rect 39615 -6235 39660 -6115
rect 39780 -6235 39835 -6115
rect 39955 -6235 40000 -6115
rect 40120 -6235 40165 -6115
rect 40285 -6235 40330 -6115
rect 40450 -6235 40505 -6115
rect 40625 -6235 40670 -6115
rect 40790 -6235 40835 -6115
rect 40955 -6235 41000 -6115
rect 41120 -6235 41175 -6115
rect 41295 -6235 41340 -6115
rect 41460 -6235 41505 -6115
rect 41625 -6235 41670 -6115
rect 41790 -6235 41845 -6115
rect 41965 -6235 41975 -6115
rect 36475 -6280 41975 -6235
rect 36475 -6400 36485 -6280
rect 36605 -6400 36650 -6280
rect 36770 -6400 36815 -6280
rect 36935 -6400 36980 -6280
rect 37100 -6400 37155 -6280
rect 37275 -6400 37320 -6280
rect 37440 -6400 37485 -6280
rect 37605 -6400 37650 -6280
rect 37770 -6400 37825 -6280
rect 37945 -6400 37990 -6280
rect 38110 -6400 38155 -6280
rect 38275 -6400 38320 -6280
rect 38440 -6400 38495 -6280
rect 38615 -6400 38660 -6280
rect 38780 -6400 38825 -6280
rect 38945 -6400 38990 -6280
rect 39110 -6400 39165 -6280
rect 39285 -6400 39330 -6280
rect 39450 -6400 39495 -6280
rect 39615 -6400 39660 -6280
rect 39780 -6400 39835 -6280
rect 39955 -6400 40000 -6280
rect 40120 -6400 40165 -6280
rect 40285 -6400 40330 -6280
rect 40450 -6400 40505 -6280
rect 40625 -6400 40670 -6280
rect 40790 -6400 40835 -6280
rect 40955 -6400 41000 -6280
rect 41120 -6400 41175 -6280
rect 41295 -6400 41340 -6280
rect 41460 -6400 41505 -6280
rect 41625 -6400 41670 -6280
rect 41790 -6400 41845 -6280
rect 41965 -6400 41975 -6280
rect 36475 -6455 41975 -6400
rect 36475 -6575 36485 -6455
rect 36605 -6575 36650 -6455
rect 36770 -6575 36815 -6455
rect 36935 -6575 36980 -6455
rect 37100 -6575 37155 -6455
rect 37275 -6575 37320 -6455
rect 37440 -6575 37485 -6455
rect 37605 -6575 37650 -6455
rect 37770 -6575 37825 -6455
rect 37945 -6575 37990 -6455
rect 38110 -6575 38155 -6455
rect 38275 -6575 38320 -6455
rect 38440 -6575 38495 -6455
rect 38615 -6575 38660 -6455
rect 38780 -6575 38825 -6455
rect 38945 -6575 38990 -6455
rect 39110 -6575 39165 -6455
rect 39285 -6575 39330 -6455
rect 39450 -6575 39495 -6455
rect 39615 -6575 39660 -6455
rect 39780 -6575 39835 -6455
rect 39955 -6575 40000 -6455
rect 40120 -6575 40165 -6455
rect 40285 -6575 40330 -6455
rect 40450 -6575 40505 -6455
rect 40625 -6575 40670 -6455
rect 40790 -6575 40835 -6455
rect 40955 -6575 41000 -6455
rect 41120 -6575 41175 -6455
rect 41295 -6575 41340 -6455
rect 41460 -6575 41505 -6455
rect 41625 -6575 41670 -6455
rect 41790 -6575 41845 -6455
rect 41965 -6575 41975 -6455
rect 36475 -6620 41975 -6575
rect 36475 -6740 36485 -6620
rect 36605 -6740 36650 -6620
rect 36770 -6740 36815 -6620
rect 36935 -6740 36980 -6620
rect 37100 -6740 37155 -6620
rect 37275 -6740 37320 -6620
rect 37440 -6740 37485 -6620
rect 37605 -6740 37650 -6620
rect 37770 -6740 37825 -6620
rect 37945 -6740 37990 -6620
rect 38110 -6740 38155 -6620
rect 38275 -6740 38320 -6620
rect 38440 -6740 38495 -6620
rect 38615 -6740 38660 -6620
rect 38780 -6740 38825 -6620
rect 38945 -6740 38990 -6620
rect 39110 -6740 39165 -6620
rect 39285 -6740 39330 -6620
rect 39450 -6740 39495 -6620
rect 39615 -6740 39660 -6620
rect 39780 -6740 39835 -6620
rect 39955 -6740 40000 -6620
rect 40120 -6740 40165 -6620
rect 40285 -6740 40330 -6620
rect 40450 -6740 40505 -6620
rect 40625 -6740 40670 -6620
rect 40790 -6740 40835 -6620
rect 40955 -6740 41000 -6620
rect 41120 -6740 41175 -6620
rect 41295 -6740 41340 -6620
rect 41460 -6740 41505 -6620
rect 41625 -6740 41670 -6620
rect 41790 -6740 41845 -6620
rect 41965 -6740 41975 -6620
rect 36475 -6785 41975 -6740
rect 36475 -6905 36485 -6785
rect 36605 -6905 36650 -6785
rect 36770 -6905 36815 -6785
rect 36935 -6905 36980 -6785
rect 37100 -6905 37155 -6785
rect 37275 -6905 37320 -6785
rect 37440 -6905 37485 -6785
rect 37605 -6905 37650 -6785
rect 37770 -6905 37825 -6785
rect 37945 -6905 37990 -6785
rect 38110 -6905 38155 -6785
rect 38275 -6905 38320 -6785
rect 38440 -6905 38495 -6785
rect 38615 -6905 38660 -6785
rect 38780 -6905 38825 -6785
rect 38945 -6905 38990 -6785
rect 39110 -6905 39165 -6785
rect 39285 -6905 39330 -6785
rect 39450 -6905 39495 -6785
rect 39615 -6905 39660 -6785
rect 39780 -6905 39835 -6785
rect 39955 -6905 40000 -6785
rect 40120 -6905 40165 -6785
rect 40285 -6905 40330 -6785
rect 40450 -6905 40505 -6785
rect 40625 -6905 40670 -6785
rect 40790 -6905 40835 -6785
rect 40955 -6905 41000 -6785
rect 41120 -6905 41175 -6785
rect 41295 -6905 41340 -6785
rect 41460 -6905 41505 -6785
rect 41625 -6905 41670 -6785
rect 41790 -6905 41845 -6785
rect 41965 -6905 41975 -6785
rect 36475 -6950 41975 -6905
rect 36475 -7070 36485 -6950
rect 36605 -7070 36650 -6950
rect 36770 -7070 36815 -6950
rect 36935 -7070 36980 -6950
rect 37100 -7070 37155 -6950
rect 37275 -7070 37320 -6950
rect 37440 -7070 37485 -6950
rect 37605 -7070 37650 -6950
rect 37770 -7070 37825 -6950
rect 37945 -7070 37990 -6950
rect 38110 -7070 38155 -6950
rect 38275 -7070 38320 -6950
rect 38440 -7070 38495 -6950
rect 38615 -7070 38660 -6950
rect 38780 -7070 38825 -6950
rect 38945 -7070 38990 -6950
rect 39110 -7070 39165 -6950
rect 39285 -7070 39330 -6950
rect 39450 -7070 39495 -6950
rect 39615 -7070 39660 -6950
rect 39780 -7070 39835 -6950
rect 39955 -7070 40000 -6950
rect 40120 -7070 40165 -6950
rect 40285 -7070 40330 -6950
rect 40450 -7070 40505 -6950
rect 40625 -7070 40670 -6950
rect 40790 -7070 40835 -6950
rect 40955 -7070 41000 -6950
rect 41120 -7070 41175 -6950
rect 41295 -7070 41340 -6950
rect 41460 -7070 41505 -6950
rect 41625 -7070 41670 -6950
rect 41790 -7070 41845 -6950
rect 41965 -7070 41975 -6950
rect 36475 -7125 41975 -7070
rect 36475 -7245 36485 -7125
rect 36605 -7245 36650 -7125
rect 36770 -7245 36815 -7125
rect 36935 -7245 36980 -7125
rect 37100 -7245 37155 -7125
rect 37275 -7245 37320 -7125
rect 37440 -7245 37485 -7125
rect 37605 -7245 37650 -7125
rect 37770 -7245 37825 -7125
rect 37945 -7245 37990 -7125
rect 38110 -7245 38155 -7125
rect 38275 -7245 38320 -7125
rect 38440 -7245 38495 -7125
rect 38615 -7245 38660 -7125
rect 38780 -7245 38825 -7125
rect 38945 -7245 38990 -7125
rect 39110 -7245 39165 -7125
rect 39285 -7245 39330 -7125
rect 39450 -7245 39495 -7125
rect 39615 -7245 39660 -7125
rect 39780 -7245 39835 -7125
rect 39955 -7245 40000 -7125
rect 40120 -7245 40165 -7125
rect 40285 -7245 40330 -7125
rect 40450 -7245 40505 -7125
rect 40625 -7245 40670 -7125
rect 40790 -7245 40835 -7125
rect 40955 -7245 41000 -7125
rect 41120 -7245 41175 -7125
rect 41295 -7245 41340 -7125
rect 41460 -7245 41505 -7125
rect 41625 -7245 41670 -7125
rect 41790 -7245 41845 -7125
rect 41965 -7245 41975 -7125
rect 36475 -7290 41975 -7245
rect 36475 -7410 36485 -7290
rect 36605 -7410 36650 -7290
rect 36770 -7410 36815 -7290
rect 36935 -7410 36980 -7290
rect 37100 -7410 37155 -7290
rect 37275 -7410 37320 -7290
rect 37440 -7410 37485 -7290
rect 37605 -7410 37650 -7290
rect 37770 -7410 37825 -7290
rect 37945 -7410 37990 -7290
rect 38110 -7410 38155 -7290
rect 38275 -7410 38320 -7290
rect 38440 -7410 38495 -7290
rect 38615 -7410 38660 -7290
rect 38780 -7410 38825 -7290
rect 38945 -7410 38990 -7290
rect 39110 -7410 39165 -7290
rect 39285 -7410 39330 -7290
rect 39450 -7410 39495 -7290
rect 39615 -7410 39660 -7290
rect 39780 -7410 39835 -7290
rect 39955 -7410 40000 -7290
rect 40120 -7410 40165 -7290
rect 40285 -7410 40330 -7290
rect 40450 -7410 40505 -7290
rect 40625 -7410 40670 -7290
rect 40790 -7410 40835 -7290
rect 40955 -7410 41000 -7290
rect 41120 -7410 41175 -7290
rect 41295 -7410 41340 -7290
rect 41460 -7410 41505 -7290
rect 41625 -7410 41670 -7290
rect 41790 -7410 41845 -7290
rect 41965 -7410 41975 -7290
rect 36475 -7455 41975 -7410
rect 36475 -7575 36485 -7455
rect 36605 -7575 36650 -7455
rect 36770 -7575 36815 -7455
rect 36935 -7575 36980 -7455
rect 37100 -7575 37155 -7455
rect 37275 -7575 37320 -7455
rect 37440 -7575 37485 -7455
rect 37605 -7575 37650 -7455
rect 37770 -7575 37825 -7455
rect 37945 -7575 37990 -7455
rect 38110 -7575 38155 -7455
rect 38275 -7575 38320 -7455
rect 38440 -7575 38495 -7455
rect 38615 -7575 38660 -7455
rect 38780 -7575 38825 -7455
rect 38945 -7575 38990 -7455
rect 39110 -7575 39165 -7455
rect 39285 -7575 39330 -7455
rect 39450 -7575 39495 -7455
rect 39615 -7575 39660 -7455
rect 39780 -7575 39835 -7455
rect 39955 -7575 40000 -7455
rect 40120 -7575 40165 -7455
rect 40285 -7575 40330 -7455
rect 40450 -7575 40505 -7455
rect 40625 -7575 40670 -7455
rect 40790 -7575 40835 -7455
rect 40955 -7575 41000 -7455
rect 41120 -7575 41175 -7455
rect 41295 -7575 41340 -7455
rect 41460 -7575 41505 -7455
rect 41625 -7575 41670 -7455
rect 41790 -7575 41845 -7455
rect 41965 -7575 41975 -7455
rect 36475 -7620 41975 -7575
rect 36475 -7740 36485 -7620
rect 36605 -7740 36650 -7620
rect 36770 -7740 36815 -7620
rect 36935 -7740 36980 -7620
rect 37100 -7740 37155 -7620
rect 37275 -7740 37320 -7620
rect 37440 -7740 37485 -7620
rect 37605 -7740 37650 -7620
rect 37770 -7740 37825 -7620
rect 37945 -7740 37990 -7620
rect 38110 -7740 38155 -7620
rect 38275 -7740 38320 -7620
rect 38440 -7740 38495 -7620
rect 38615 -7740 38660 -7620
rect 38780 -7740 38825 -7620
rect 38945 -7740 38990 -7620
rect 39110 -7740 39165 -7620
rect 39285 -7740 39330 -7620
rect 39450 -7740 39495 -7620
rect 39615 -7740 39660 -7620
rect 39780 -7740 39835 -7620
rect 39955 -7740 40000 -7620
rect 40120 -7740 40165 -7620
rect 40285 -7740 40330 -7620
rect 40450 -7740 40505 -7620
rect 40625 -7740 40670 -7620
rect 40790 -7740 40835 -7620
rect 40955 -7740 41000 -7620
rect 41120 -7740 41175 -7620
rect 41295 -7740 41340 -7620
rect 41460 -7740 41505 -7620
rect 41625 -7740 41670 -7620
rect 41790 -7740 41845 -7620
rect 41965 -7740 41975 -7620
rect 36475 -7795 41975 -7740
rect 36475 -7915 36485 -7795
rect 36605 -7915 36650 -7795
rect 36770 -7915 36815 -7795
rect 36935 -7915 36980 -7795
rect 37100 -7915 37155 -7795
rect 37275 -7915 37320 -7795
rect 37440 -7915 37485 -7795
rect 37605 -7915 37650 -7795
rect 37770 -7915 37825 -7795
rect 37945 -7915 37990 -7795
rect 38110 -7915 38155 -7795
rect 38275 -7915 38320 -7795
rect 38440 -7915 38495 -7795
rect 38615 -7915 38660 -7795
rect 38780 -7915 38825 -7795
rect 38945 -7915 38990 -7795
rect 39110 -7915 39165 -7795
rect 39285 -7915 39330 -7795
rect 39450 -7915 39495 -7795
rect 39615 -7915 39660 -7795
rect 39780 -7915 39835 -7795
rect 39955 -7915 40000 -7795
rect 40120 -7915 40165 -7795
rect 40285 -7915 40330 -7795
rect 40450 -7915 40505 -7795
rect 40625 -7915 40670 -7795
rect 40790 -7915 40835 -7795
rect 40955 -7915 41000 -7795
rect 41120 -7915 41175 -7795
rect 41295 -7915 41340 -7795
rect 41460 -7915 41505 -7795
rect 41625 -7915 41670 -7795
rect 41790 -7915 41845 -7795
rect 41965 -7915 41975 -7795
rect 36475 -7960 41975 -7915
rect 36475 -8080 36485 -7960
rect 36605 -8080 36650 -7960
rect 36770 -8080 36815 -7960
rect 36935 -8080 36980 -7960
rect 37100 -8080 37155 -7960
rect 37275 -8080 37320 -7960
rect 37440 -8080 37485 -7960
rect 37605 -8080 37650 -7960
rect 37770 -8080 37825 -7960
rect 37945 -8080 37990 -7960
rect 38110 -8080 38155 -7960
rect 38275 -8080 38320 -7960
rect 38440 -8080 38495 -7960
rect 38615 -8080 38660 -7960
rect 38780 -8080 38825 -7960
rect 38945 -8080 38990 -7960
rect 39110 -8080 39165 -7960
rect 39285 -8080 39330 -7960
rect 39450 -8080 39495 -7960
rect 39615 -8080 39660 -7960
rect 39780 -8080 39835 -7960
rect 39955 -8080 40000 -7960
rect 40120 -8080 40165 -7960
rect 40285 -8080 40330 -7960
rect 40450 -8080 40505 -7960
rect 40625 -8080 40670 -7960
rect 40790 -8080 40835 -7960
rect 40955 -8080 41000 -7960
rect 41120 -8080 41175 -7960
rect 41295 -8080 41340 -7960
rect 41460 -8080 41505 -7960
rect 41625 -8080 41670 -7960
rect 41790 -8080 41845 -7960
rect 41965 -8080 41975 -7960
rect 36475 -8125 41975 -8080
rect 36475 -8245 36485 -8125
rect 36605 -8245 36650 -8125
rect 36770 -8245 36815 -8125
rect 36935 -8245 36980 -8125
rect 37100 -8245 37155 -8125
rect 37275 -8245 37320 -8125
rect 37440 -8245 37485 -8125
rect 37605 -8245 37650 -8125
rect 37770 -8245 37825 -8125
rect 37945 -8245 37990 -8125
rect 38110 -8245 38155 -8125
rect 38275 -8245 38320 -8125
rect 38440 -8245 38495 -8125
rect 38615 -8245 38660 -8125
rect 38780 -8245 38825 -8125
rect 38945 -8245 38990 -8125
rect 39110 -8245 39165 -8125
rect 39285 -8245 39330 -8125
rect 39450 -8245 39495 -8125
rect 39615 -8245 39660 -8125
rect 39780 -8245 39835 -8125
rect 39955 -8245 40000 -8125
rect 40120 -8245 40165 -8125
rect 40285 -8245 40330 -8125
rect 40450 -8245 40505 -8125
rect 40625 -8245 40670 -8125
rect 40790 -8245 40835 -8125
rect 40955 -8245 41000 -8125
rect 41120 -8245 41175 -8125
rect 41295 -8245 41340 -8125
rect 41460 -8245 41505 -8125
rect 41625 -8245 41670 -8125
rect 41790 -8245 41845 -8125
rect 41965 -8245 41975 -8125
rect 36475 -8290 41975 -8245
rect 36475 -8410 36485 -8290
rect 36605 -8410 36650 -8290
rect 36770 -8410 36815 -8290
rect 36935 -8410 36980 -8290
rect 37100 -8410 37155 -8290
rect 37275 -8410 37320 -8290
rect 37440 -8410 37485 -8290
rect 37605 -8410 37650 -8290
rect 37770 -8410 37825 -8290
rect 37945 -8410 37990 -8290
rect 38110 -8410 38155 -8290
rect 38275 -8410 38320 -8290
rect 38440 -8410 38495 -8290
rect 38615 -8410 38660 -8290
rect 38780 -8410 38825 -8290
rect 38945 -8410 38990 -8290
rect 39110 -8410 39165 -8290
rect 39285 -8410 39330 -8290
rect 39450 -8410 39495 -8290
rect 39615 -8410 39660 -8290
rect 39780 -8410 39835 -8290
rect 39955 -8410 40000 -8290
rect 40120 -8410 40165 -8290
rect 40285 -8410 40330 -8290
rect 40450 -8410 40505 -8290
rect 40625 -8410 40670 -8290
rect 40790 -8410 40835 -8290
rect 40955 -8410 41000 -8290
rect 41120 -8410 41175 -8290
rect 41295 -8410 41340 -8290
rect 41460 -8410 41505 -8290
rect 41625 -8410 41670 -8290
rect 41790 -8410 41845 -8290
rect 41965 -8410 41975 -8290
rect 36475 -8465 41975 -8410
rect 36475 -8585 36485 -8465
rect 36605 -8585 36650 -8465
rect 36770 -8585 36815 -8465
rect 36935 -8585 36980 -8465
rect 37100 -8585 37155 -8465
rect 37275 -8585 37320 -8465
rect 37440 -8585 37485 -8465
rect 37605 -8585 37650 -8465
rect 37770 -8585 37825 -8465
rect 37945 -8585 37990 -8465
rect 38110 -8585 38155 -8465
rect 38275 -8585 38320 -8465
rect 38440 -8585 38495 -8465
rect 38615 -8585 38660 -8465
rect 38780 -8585 38825 -8465
rect 38945 -8585 38990 -8465
rect 39110 -8585 39165 -8465
rect 39285 -8585 39330 -8465
rect 39450 -8585 39495 -8465
rect 39615 -8585 39660 -8465
rect 39780 -8585 39835 -8465
rect 39955 -8585 40000 -8465
rect 40120 -8585 40165 -8465
rect 40285 -8585 40330 -8465
rect 40450 -8585 40505 -8465
rect 40625 -8585 40670 -8465
rect 40790 -8585 40835 -8465
rect 40955 -8585 41000 -8465
rect 41120 -8585 41175 -8465
rect 41295 -8585 41340 -8465
rect 41460 -8585 41505 -8465
rect 41625 -8585 41670 -8465
rect 41790 -8585 41845 -8465
rect 41965 -8585 41975 -8465
rect 36475 -8630 41975 -8585
rect 36475 -8750 36485 -8630
rect 36605 -8750 36650 -8630
rect 36770 -8750 36815 -8630
rect 36935 -8750 36980 -8630
rect 37100 -8750 37155 -8630
rect 37275 -8750 37320 -8630
rect 37440 -8750 37485 -8630
rect 37605 -8750 37650 -8630
rect 37770 -8750 37825 -8630
rect 37945 -8750 37990 -8630
rect 38110 -8750 38155 -8630
rect 38275 -8750 38320 -8630
rect 38440 -8750 38495 -8630
rect 38615 -8750 38660 -8630
rect 38780 -8750 38825 -8630
rect 38945 -8750 38990 -8630
rect 39110 -8750 39165 -8630
rect 39285 -8750 39330 -8630
rect 39450 -8750 39495 -8630
rect 39615 -8750 39660 -8630
rect 39780 -8750 39835 -8630
rect 39955 -8750 40000 -8630
rect 40120 -8750 40165 -8630
rect 40285 -8750 40330 -8630
rect 40450 -8750 40505 -8630
rect 40625 -8750 40670 -8630
rect 40790 -8750 40835 -8630
rect 40955 -8750 41000 -8630
rect 41120 -8750 41175 -8630
rect 41295 -8750 41340 -8630
rect 41460 -8750 41505 -8630
rect 41625 -8750 41670 -8630
rect 41790 -8750 41845 -8630
rect 41965 -8750 41975 -8630
rect 36475 -8795 41975 -8750
rect 36475 -8915 36485 -8795
rect 36605 -8915 36650 -8795
rect 36770 -8915 36815 -8795
rect 36935 -8915 36980 -8795
rect 37100 -8915 37155 -8795
rect 37275 -8915 37320 -8795
rect 37440 -8915 37485 -8795
rect 37605 -8915 37650 -8795
rect 37770 -8915 37825 -8795
rect 37945 -8915 37990 -8795
rect 38110 -8915 38155 -8795
rect 38275 -8915 38320 -8795
rect 38440 -8915 38495 -8795
rect 38615 -8915 38660 -8795
rect 38780 -8915 38825 -8795
rect 38945 -8915 38990 -8795
rect 39110 -8915 39165 -8795
rect 39285 -8915 39330 -8795
rect 39450 -8915 39495 -8795
rect 39615 -8915 39660 -8795
rect 39780 -8915 39835 -8795
rect 39955 -8915 40000 -8795
rect 40120 -8915 40165 -8795
rect 40285 -8915 40330 -8795
rect 40450 -8915 40505 -8795
rect 40625 -8915 40670 -8795
rect 40790 -8915 40835 -8795
rect 40955 -8915 41000 -8795
rect 41120 -8915 41175 -8795
rect 41295 -8915 41340 -8795
rect 41460 -8915 41505 -8795
rect 41625 -8915 41670 -8795
rect 41790 -8915 41845 -8795
rect 41965 -8915 41975 -8795
rect 36475 -8960 41975 -8915
rect 36475 -9080 36485 -8960
rect 36605 -9080 36650 -8960
rect 36770 -9080 36815 -8960
rect 36935 -9080 36980 -8960
rect 37100 -9080 37155 -8960
rect 37275 -9080 37320 -8960
rect 37440 -9080 37485 -8960
rect 37605 -9080 37650 -8960
rect 37770 -9080 37825 -8960
rect 37945 -9080 37990 -8960
rect 38110 -9080 38155 -8960
rect 38275 -9080 38320 -8960
rect 38440 -9080 38495 -8960
rect 38615 -9080 38660 -8960
rect 38780 -9080 38825 -8960
rect 38945 -9080 38990 -8960
rect 39110 -9080 39165 -8960
rect 39285 -9080 39330 -8960
rect 39450 -9080 39495 -8960
rect 39615 -9080 39660 -8960
rect 39780 -9080 39835 -8960
rect 39955 -9080 40000 -8960
rect 40120 -9080 40165 -8960
rect 40285 -9080 40330 -8960
rect 40450 -9080 40505 -8960
rect 40625 -9080 40670 -8960
rect 40790 -9080 40835 -8960
rect 40955 -9080 41000 -8960
rect 41120 -9080 41175 -8960
rect 41295 -9080 41340 -8960
rect 41460 -9080 41505 -8960
rect 41625 -9080 41670 -8960
rect 41790 -9080 41845 -8960
rect 41965 -9080 41975 -8960
rect 36475 -9135 41975 -9080
rect 36475 -9255 36485 -9135
rect 36605 -9255 36650 -9135
rect 36770 -9255 36815 -9135
rect 36935 -9255 36980 -9135
rect 37100 -9255 37155 -9135
rect 37275 -9255 37320 -9135
rect 37440 -9255 37485 -9135
rect 37605 -9255 37650 -9135
rect 37770 -9255 37825 -9135
rect 37945 -9255 37990 -9135
rect 38110 -9255 38155 -9135
rect 38275 -9255 38320 -9135
rect 38440 -9255 38495 -9135
rect 38615 -9255 38660 -9135
rect 38780 -9255 38825 -9135
rect 38945 -9255 38990 -9135
rect 39110 -9255 39165 -9135
rect 39285 -9255 39330 -9135
rect 39450 -9255 39495 -9135
rect 39615 -9255 39660 -9135
rect 39780 -9255 39835 -9135
rect 39955 -9255 40000 -9135
rect 40120 -9255 40165 -9135
rect 40285 -9255 40330 -9135
rect 40450 -9255 40505 -9135
rect 40625 -9255 40670 -9135
rect 40790 -9255 40835 -9135
rect 40955 -9255 41000 -9135
rect 41120 -9255 41175 -9135
rect 41295 -9255 41340 -9135
rect 41460 -9255 41505 -9135
rect 41625 -9255 41670 -9135
rect 41790 -9255 41845 -9135
rect 41965 -9255 41975 -9135
rect 36475 -9300 41975 -9255
rect 36475 -9420 36485 -9300
rect 36605 -9420 36650 -9300
rect 36770 -9420 36815 -9300
rect 36935 -9420 36980 -9300
rect 37100 -9420 37155 -9300
rect 37275 -9420 37320 -9300
rect 37440 -9420 37485 -9300
rect 37605 -9420 37650 -9300
rect 37770 -9420 37825 -9300
rect 37945 -9420 37990 -9300
rect 38110 -9420 38155 -9300
rect 38275 -9420 38320 -9300
rect 38440 -9420 38495 -9300
rect 38615 -9420 38660 -9300
rect 38780 -9420 38825 -9300
rect 38945 -9420 38990 -9300
rect 39110 -9420 39165 -9300
rect 39285 -9420 39330 -9300
rect 39450 -9420 39495 -9300
rect 39615 -9420 39660 -9300
rect 39780 -9420 39835 -9300
rect 39955 -9420 40000 -9300
rect 40120 -9420 40165 -9300
rect 40285 -9420 40330 -9300
rect 40450 -9420 40505 -9300
rect 40625 -9420 40670 -9300
rect 40790 -9420 40835 -9300
rect 40955 -9420 41000 -9300
rect 41120 -9420 41175 -9300
rect 41295 -9420 41340 -9300
rect 41460 -9420 41505 -9300
rect 41625 -9420 41670 -9300
rect 41790 -9420 41845 -9300
rect 41965 -9420 41975 -9300
rect 36475 -9465 41975 -9420
rect 36475 -9585 36485 -9465
rect 36605 -9585 36650 -9465
rect 36770 -9585 36815 -9465
rect 36935 -9585 36980 -9465
rect 37100 -9585 37155 -9465
rect 37275 -9585 37320 -9465
rect 37440 -9585 37485 -9465
rect 37605 -9585 37650 -9465
rect 37770 -9585 37825 -9465
rect 37945 -9585 37990 -9465
rect 38110 -9585 38155 -9465
rect 38275 -9585 38320 -9465
rect 38440 -9585 38495 -9465
rect 38615 -9585 38660 -9465
rect 38780 -9585 38825 -9465
rect 38945 -9585 38990 -9465
rect 39110 -9585 39165 -9465
rect 39285 -9585 39330 -9465
rect 39450 -9585 39495 -9465
rect 39615 -9585 39660 -9465
rect 39780 -9585 39835 -9465
rect 39955 -9585 40000 -9465
rect 40120 -9585 40165 -9465
rect 40285 -9585 40330 -9465
rect 40450 -9585 40505 -9465
rect 40625 -9585 40670 -9465
rect 40790 -9585 40835 -9465
rect 40955 -9585 41000 -9465
rect 41120 -9585 41175 -9465
rect 41295 -9585 41340 -9465
rect 41460 -9585 41505 -9465
rect 41625 -9585 41670 -9465
rect 41790 -9585 41845 -9465
rect 41965 -9585 41975 -9465
rect 36475 -9630 41975 -9585
rect 36475 -9750 36485 -9630
rect 36605 -9750 36650 -9630
rect 36770 -9750 36815 -9630
rect 36935 -9750 36980 -9630
rect 37100 -9750 37155 -9630
rect 37275 -9750 37320 -9630
rect 37440 -9750 37485 -9630
rect 37605 -9750 37650 -9630
rect 37770 -9750 37825 -9630
rect 37945 -9750 37990 -9630
rect 38110 -9750 38155 -9630
rect 38275 -9750 38320 -9630
rect 38440 -9750 38495 -9630
rect 38615 -9750 38660 -9630
rect 38780 -9750 38825 -9630
rect 38945 -9750 38990 -9630
rect 39110 -9750 39165 -9630
rect 39285 -9750 39330 -9630
rect 39450 -9750 39495 -9630
rect 39615 -9750 39660 -9630
rect 39780 -9750 39835 -9630
rect 39955 -9750 40000 -9630
rect 40120 -9750 40165 -9630
rect 40285 -9750 40330 -9630
rect 40450 -9750 40505 -9630
rect 40625 -9750 40670 -9630
rect 40790 -9750 40835 -9630
rect 40955 -9750 41000 -9630
rect 41120 -9750 41175 -9630
rect 41295 -9750 41340 -9630
rect 41460 -9750 41505 -9630
rect 41625 -9750 41670 -9630
rect 41790 -9750 41845 -9630
rect 41965 -9750 41975 -9630
rect 36475 -9760 41975 -9750
rect 42165 -4270 47665 -4260
rect 42165 -4390 42175 -4270
rect 42295 -4390 42340 -4270
rect 42460 -4390 42505 -4270
rect 42625 -4390 42670 -4270
rect 42790 -4390 42845 -4270
rect 42965 -4390 43010 -4270
rect 43130 -4390 43175 -4270
rect 43295 -4390 43340 -4270
rect 43460 -4390 43515 -4270
rect 43635 -4390 43680 -4270
rect 43800 -4390 43845 -4270
rect 43965 -4390 44010 -4270
rect 44130 -4390 44185 -4270
rect 44305 -4390 44350 -4270
rect 44470 -4390 44515 -4270
rect 44635 -4390 44680 -4270
rect 44800 -4390 44855 -4270
rect 44975 -4390 45020 -4270
rect 45140 -4390 45185 -4270
rect 45305 -4390 45350 -4270
rect 45470 -4390 45525 -4270
rect 45645 -4390 45690 -4270
rect 45810 -4390 45855 -4270
rect 45975 -4390 46020 -4270
rect 46140 -4390 46195 -4270
rect 46315 -4390 46360 -4270
rect 46480 -4390 46525 -4270
rect 46645 -4390 46690 -4270
rect 46810 -4390 46865 -4270
rect 46985 -4390 47030 -4270
rect 47150 -4390 47195 -4270
rect 47315 -4390 47360 -4270
rect 47480 -4390 47535 -4270
rect 47655 -4390 47665 -4270
rect 42165 -4445 47665 -4390
rect 42165 -4565 42175 -4445
rect 42295 -4565 42340 -4445
rect 42460 -4565 42505 -4445
rect 42625 -4565 42670 -4445
rect 42790 -4565 42845 -4445
rect 42965 -4565 43010 -4445
rect 43130 -4565 43175 -4445
rect 43295 -4565 43340 -4445
rect 43460 -4565 43515 -4445
rect 43635 -4565 43680 -4445
rect 43800 -4565 43845 -4445
rect 43965 -4565 44010 -4445
rect 44130 -4565 44185 -4445
rect 44305 -4565 44350 -4445
rect 44470 -4565 44515 -4445
rect 44635 -4565 44680 -4445
rect 44800 -4565 44855 -4445
rect 44975 -4565 45020 -4445
rect 45140 -4565 45185 -4445
rect 45305 -4565 45350 -4445
rect 45470 -4565 45525 -4445
rect 45645 -4565 45690 -4445
rect 45810 -4565 45855 -4445
rect 45975 -4565 46020 -4445
rect 46140 -4565 46195 -4445
rect 46315 -4565 46360 -4445
rect 46480 -4565 46525 -4445
rect 46645 -4565 46690 -4445
rect 46810 -4565 46865 -4445
rect 46985 -4565 47030 -4445
rect 47150 -4565 47195 -4445
rect 47315 -4565 47360 -4445
rect 47480 -4565 47535 -4445
rect 47655 -4565 47665 -4445
rect 42165 -4610 47665 -4565
rect 42165 -4730 42175 -4610
rect 42295 -4730 42340 -4610
rect 42460 -4730 42505 -4610
rect 42625 -4730 42670 -4610
rect 42790 -4730 42845 -4610
rect 42965 -4730 43010 -4610
rect 43130 -4730 43175 -4610
rect 43295 -4730 43340 -4610
rect 43460 -4730 43515 -4610
rect 43635 -4730 43680 -4610
rect 43800 -4730 43845 -4610
rect 43965 -4730 44010 -4610
rect 44130 -4730 44185 -4610
rect 44305 -4730 44350 -4610
rect 44470 -4730 44515 -4610
rect 44635 -4730 44680 -4610
rect 44800 -4730 44855 -4610
rect 44975 -4730 45020 -4610
rect 45140 -4730 45185 -4610
rect 45305 -4730 45350 -4610
rect 45470 -4730 45525 -4610
rect 45645 -4730 45690 -4610
rect 45810 -4730 45855 -4610
rect 45975 -4730 46020 -4610
rect 46140 -4730 46195 -4610
rect 46315 -4730 46360 -4610
rect 46480 -4730 46525 -4610
rect 46645 -4730 46690 -4610
rect 46810 -4730 46865 -4610
rect 46985 -4730 47030 -4610
rect 47150 -4730 47195 -4610
rect 47315 -4730 47360 -4610
rect 47480 -4730 47535 -4610
rect 47655 -4730 47665 -4610
rect 42165 -4775 47665 -4730
rect 42165 -4895 42175 -4775
rect 42295 -4895 42340 -4775
rect 42460 -4895 42505 -4775
rect 42625 -4895 42670 -4775
rect 42790 -4895 42845 -4775
rect 42965 -4895 43010 -4775
rect 43130 -4895 43175 -4775
rect 43295 -4895 43340 -4775
rect 43460 -4895 43515 -4775
rect 43635 -4895 43680 -4775
rect 43800 -4895 43845 -4775
rect 43965 -4895 44010 -4775
rect 44130 -4895 44185 -4775
rect 44305 -4895 44350 -4775
rect 44470 -4895 44515 -4775
rect 44635 -4895 44680 -4775
rect 44800 -4895 44855 -4775
rect 44975 -4895 45020 -4775
rect 45140 -4895 45185 -4775
rect 45305 -4895 45350 -4775
rect 45470 -4895 45525 -4775
rect 45645 -4895 45690 -4775
rect 45810 -4895 45855 -4775
rect 45975 -4895 46020 -4775
rect 46140 -4895 46195 -4775
rect 46315 -4895 46360 -4775
rect 46480 -4895 46525 -4775
rect 46645 -4895 46690 -4775
rect 46810 -4895 46865 -4775
rect 46985 -4895 47030 -4775
rect 47150 -4895 47195 -4775
rect 47315 -4895 47360 -4775
rect 47480 -4895 47535 -4775
rect 47655 -4895 47665 -4775
rect 42165 -4940 47665 -4895
rect 42165 -5060 42175 -4940
rect 42295 -5060 42340 -4940
rect 42460 -5060 42505 -4940
rect 42625 -5060 42670 -4940
rect 42790 -5060 42845 -4940
rect 42965 -5060 43010 -4940
rect 43130 -5060 43175 -4940
rect 43295 -5060 43340 -4940
rect 43460 -5060 43515 -4940
rect 43635 -5060 43680 -4940
rect 43800 -5060 43845 -4940
rect 43965 -5060 44010 -4940
rect 44130 -5060 44185 -4940
rect 44305 -5060 44350 -4940
rect 44470 -5060 44515 -4940
rect 44635 -5060 44680 -4940
rect 44800 -5060 44855 -4940
rect 44975 -5060 45020 -4940
rect 45140 -5060 45185 -4940
rect 45305 -5060 45350 -4940
rect 45470 -5060 45525 -4940
rect 45645 -5060 45690 -4940
rect 45810 -5060 45855 -4940
rect 45975 -5060 46020 -4940
rect 46140 -5060 46195 -4940
rect 46315 -5060 46360 -4940
rect 46480 -5060 46525 -4940
rect 46645 -5060 46690 -4940
rect 46810 -5060 46865 -4940
rect 46985 -5060 47030 -4940
rect 47150 -5060 47195 -4940
rect 47315 -5060 47360 -4940
rect 47480 -5060 47535 -4940
rect 47655 -5060 47665 -4940
rect 42165 -5115 47665 -5060
rect 42165 -5235 42175 -5115
rect 42295 -5235 42340 -5115
rect 42460 -5235 42505 -5115
rect 42625 -5235 42670 -5115
rect 42790 -5235 42845 -5115
rect 42965 -5235 43010 -5115
rect 43130 -5235 43175 -5115
rect 43295 -5235 43340 -5115
rect 43460 -5235 43515 -5115
rect 43635 -5235 43680 -5115
rect 43800 -5235 43845 -5115
rect 43965 -5235 44010 -5115
rect 44130 -5235 44185 -5115
rect 44305 -5235 44350 -5115
rect 44470 -5235 44515 -5115
rect 44635 -5235 44680 -5115
rect 44800 -5235 44855 -5115
rect 44975 -5235 45020 -5115
rect 45140 -5235 45185 -5115
rect 45305 -5235 45350 -5115
rect 45470 -5235 45525 -5115
rect 45645 -5235 45690 -5115
rect 45810 -5235 45855 -5115
rect 45975 -5235 46020 -5115
rect 46140 -5235 46195 -5115
rect 46315 -5235 46360 -5115
rect 46480 -5235 46525 -5115
rect 46645 -5235 46690 -5115
rect 46810 -5235 46865 -5115
rect 46985 -5235 47030 -5115
rect 47150 -5235 47195 -5115
rect 47315 -5235 47360 -5115
rect 47480 -5235 47535 -5115
rect 47655 -5235 47665 -5115
rect 42165 -5280 47665 -5235
rect 42165 -5400 42175 -5280
rect 42295 -5400 42340 -5280
rect 42460 -5400 42505 -5280
rect 42625 -5400 42670 -5280
rect 42790 -5400 42845 -5280
rect 42965 -5400 43010 -5280
rect 43130 -5400 43175 -5280
rect 43295 -5400 43340 -5280
rect 43460 -5400 43515 -5280
rect 43635 -5400 43680 -5280
rect 43800 -5400 43845 -5280
rect 43965 -5400 44010 -5280
rect 44130 -5400 44185 -5280
rect 44305 -5400 44350 -5280
rect 44470 -5400 44515 -5280
rect 44635 -5400 44680 -5280
rect 44800 -5400 44855 -5280
rect 44975 -5400 45020 -5280
rect 45140 -5400 45185 -5280
rect 45305 -5400 45350 -5280
rect 45470 -5400 45525 -5280
rect 45645 -5400 45690 -5280
rect 45810 -5400 45855 -5280
rect 45975 -5400 46020 -5280
rect 46140 -5400 46195 -5280
rect 46315 -5400 46360 -5280
rect 46480 -5400 46525 -5280
rect 46645 -5400 46690 -5280
rect 46810 -5400 46865 -5280
rect 46985 -5400 47030 -5280
rect 47150 -5400 47195 -5280
rect 47315 -5400 47360 -5280
rect 47480 -5400 47535 -5280
rect 47655 -5400 47665 -5280
rect 42165 -5445 47665 -5400
rect 42165 -5565 42175 -5445
rect 42295 -5565 42340 -5445
rect 42460 -5565 42505 -5445
rect 42625 -5565 42670 -5445
rect 42790 -5565 42845 -5445
rect 42965 -5565 43010 -5445
rect 43130 -5565 43175 -5445
rect 43295 -5565 43340 -5445
rect 43460 -5565 43515 -5445
rect 43635 -5565 43680 -5445
rect 43800 -5565 43845 -5445
rect 43965 -5565 44010 -5445
rect 44130 -5565 44185 -5445
rect 44305 -5565 44350 -5445
rect 44470 -5565 44515 -5445
rect 44635 -5565 44680 -5445
rect 44800 -5565 44855 -5445
rect 44975 -5565 45020 -5445
rect 45140 -5565 45185 -5445
rect 45305 -5565 45350 -5445
rect 45470 -5565 45525 -5445
rect 45645 -5565 45690 -5445
rect 45810 -5565 45855 -5445
rect 45975 -5565 46020 -5445
rect 46140 -5565 46195 -5445
rect 46315 -5565 46360 -5445
rect 46480 -5565 46525 -5445
rect 46645 -5565 46690 -5445
rect 46810 -5565 46865 -5445
rect 46985 -5565 47030 -5445
rect 47150 -5565 47195 -5445
rect 47315 -5565 47360 -5445
rect 47480 -5565 47535 -5445
rect 47655 -5565 47665 -5445
rect 42165 -5610 47665 -5565
rect 42165 -5730 42175 -5610
rect 42295 -5730 42340 -5610
rect 42460 -5730 42505 -5610
rect 42625 -5730 42670 -5610
rect 42790 -5730 42845 -5610
rect 42965 -5730 43010 -5610
rect 43130 -5730 43175 -5610
rect 43295 -5730 43340 -5610
rect 43460 -5730 43515 -5610
rect 43635 -5730 43680 -5610
rect 43800 -5730 43845 -5610
rect 43965 -5730 44010 -5610
rect 44130 -5730 44185 -5610
rect 44305 -5730 44350 -5610
rect 44470 -5730 44515 -5610
rect 44635 -5730 44680 -5610
rect 44800 -5730 44855 -5610
rect 44975 -5730 45020 -5610
rect 45140 -5730 45185 -5610
rect 45305 -5730 45350 -5610
rect 45470 -5730 45525 -5610
rect 45645 -5730 45690 -5610
rect 45810 -5730 45855 -5610
rect 45975 -5730 46020 -5610
rect 46140 -5730 46195 -5610
rect 46315 -5730 46360 -5610
rect 46480 -5730 46525 -5610
rect 46645 -5730 46690 -5610
rect 46810 -5730 46865 -5610
rect 46985 -5730 47030 -5610
rect 47150 -5730 47195 -5610
rect 47315 -5730 47360 -5610
rect 47480 -5730 47535 -5610
rect 47655 -5730 47665 -5610
rect 42165 -5785 47665 -5730
rect 42165 -5905 42175 -5785
rect 42295 -5905 42340 -5785
rect 42460 -5905 42505 -5785
rect 42625 -5905 42670 -5785
rect 42790 -5905 42845 -5785
rect 42965 -5905 43010 -5785
rect 43130 -5905 43175 -5785
rect 43295 -5905 43340 -5785
rect 43460 -5905 43515 -5785
rect 43635 -5905 43680 -5785
rect 43800 -5905 43845 -5785
rect 43965 -5905 44010 -5785
rect 44130 -5905 44185 -5785
rect 44305 -5905 44350 -5785
rect 44470 -5905 44515 -5785
rect 44635 -5905 44680 -5785
rect 44800 -5905 44855 -5785
rect 44975 -5905 45020 -5785
rect 45140 -5905 45185 -5785
rect 45305 -5905 45350 -5785
rect 45470 -5905 45525 -5785
rect 45645 -5905 45690 -5785
rect 45810 -5905 45855 -5785
rect 45975 -5905 46020 -5785
rect 46140 -5905 46195 -5785
rect 46315 -5905 46360 -5785
rect 46480 -5905 46525 -5785
rect 46645 -5905 46690 -5785
rect 46810 -5905 46865 -5785
rect 46985 -5905 47030 -5785
rect 47150 -5905 47195 -5785
rect 47315 -5905 47360 -5785
rect 47480 -5905 47535 -5785
rect 47655 -5905 47665 -5785
rect 42165 -5950 47665 -5905
rect 42165 -6070 42175 -5950
rect 42295 -6070 42340 -5950
rect 42460 -6070 42505 -5950
rect 42625 -6070 42670 -5950
rect 42790 -6070 42845 -5950
rect 42965 -6070 43010 -5950
rect 43130 -6070 43175 -5950
rect 43295 -6070 43340 -5950
rect 43460 -6070 43515 -5950
rect 43635 -6070 43680 -5950
rect 43800 -6070 43845 -5950
rect 43965 -6070 44010 -5950
rect 44130 -6070 44185 -5950
rect 44305 -6070 44350 -5950
rect 44470 -6070 44515 -5950
rect 44635 -6070 44680 -5950
rect 44800 -6070 44855 -5950
rect 44975 -6070 45020 -5950
rect 45140 -6070 45185 -5950
rect 45305 -6070 45350 -5950
rect 45470 -6070 45525 -5950
rect 45645 -6070 45690 -5950
rect 45810 -6070 45855 -5950
rect 45975 -6070 46020 -5950
rect 46140 -6070 46195 -5950
rect 46315 -6070 46360 -5950
rect 46480 -6070 46525 -5950
rect 46645 -6070 46690 -5950
rect 46810 -6070 46865 -5950
rect 46985 -6070 47030 -5950
rect 47150 -6070 47195 -5950
rect 47315 -6070 47360 -5950
rect 47480 -6070 47535 -5950
rect 47655 -6070 47665 -5950
rect 42165 -6115 47665 -6070
rect 42165 -6235 42175 -6115
rect 42295 -6235 42340 -6115
rect 42460 -6235 42505 -6115
rect 42625 -6235 42670 -6115
rect 42790 -6235 42845 -6115
rect 42965 -6235 43010 -6115
rect 43130 -6235 43175 -6115
rect 43295 -6235 43340 -6115
rect 43460 -6235 43515 -6115
rect 43635 -6235 43680 -6115
rect 43800 -6235 43845 -6115
rect 43965 -6235 44010 -6115
rect 44130 -6235 44185 -6115
rect 44305 -6235 44350 -6115
rect 44470 -6235 44515 -6115
rect 44635 -6235 44680 -6115
rect 44800 -6235 44855 -6115
rect 44975 -6235 45020 -6115
rect 45140 -6235 45185 -6115
rect 45305 -6235 45350 -6115
rect 45470 -6235 45525 -6115
rect 45645 -6235 45690 -6115
rect 45810 -6235 45855 -6115
rect 45975 -6235 46020 -6115
rect 46140 -6235 46195 -6115
rect 46315 -6235 46360 -6115
rect 46480 -6235 46525 -6115
rect 46645 -6235 46690 -6115
rect 46810 -6235 46865 -6115
rect 46985 -6235 47030 -6115
rect 47150 -6235 47195 -6115
rect 47315 -6235 47360 -6115
rect 47480 -6235 47535 -6115
rect 47655 -6235 47665 -6115
rect 42165 -6280 47665 -6235
rect 42165 -6400 42175 -6280
rect 42295 -6400 42340 -6280
rect 42460 -6400 42505 -6280
rect 42625 -6400 42670 -6280
rect 42790 -6400 42845 -6280
rect 42965 -6400 43010 -6280
rect 43130 -6400 43175 -6280
rect 43295 -6400 43340 -6280
rect 43460 -6400 43515 -6280
rect 43635 -6400 43680 -6280
rect 43800 -6400 43845 -6280
rect 43965 -6400 44010 -6280
rect 44130 -6400 44185 -6280
rect 44305 -6400 44350 -6280
rect 44470 -6400 44515 -6280
rect 44635 -6400 44680 -6280
rect 44800 -6400 44855 -6280
rect 44975 -6400 45020 -6280
rect 45140 -6400 45185 -6280
rect 45305 -6400 45350 -6280
rect 45470 -6400 45525 -6280
rect 45645 -6400 45690 -6280
rect 45810 -6400 45855 -6280
rect 45975 -6400 46020 -6280
rect 46140 -6400 46195 -6280
rect 46315 -6400 46360 -6280
rect 46480 -6400 46525 -6280
rect 46645 -6400 46690 -6280
rect 46810 -6400 46865 -6280
rect 46985 -6400 47030 -6280
rect 47150 -6400 47195 -6280
rect 47315 -6400 47360 -6280
rect 47480 -6400 47535 -6280
rect 47655 -6400 47665 -6280
rect 42165 -6455 47665 -6400
rect 42165 -6575 42175 -6455
rect 42295 -6575 42340 -6455
rect 42460 -6575 42505 -6455
rect 42625 -6575 42670 -6455
rect 42790 -6575 42845 -6455
rect 42965 -6575 43010 -6455
rect 43130 -6575 43175 -6455
rect 43295 -6575 43340 -6455
rect 43460 -6575 43515 -6455
rect 43635 -6575 43680 -6455
rect 43800 -6575 43845 -6455
rect 43965 -6575 44010 -6455
rect 44130 -6575 44185 -6455
rect 44305 -6575 44350 -6455
rect 44470 -6575 44515 -6455
rect 44635 -6575 44680 -6455
rect 44800 -6575 44855 -6455
rect 44975 -6575 45020 -6455
rect 45140 -6575 45185 -6455
rect 45305 -6575 45350 -6455
rect 45470 -6575 45525 -6455
rect 45645 -6575 45690 -6455
rect 45810 -6575 45855 -6455
rect 45975 -6575 46020 -6455
rect 46140 -6575 46195 -6455
rect 46315 -6575 46360 -6455
rect 46480 -6575 46525 -6455
rect 46645 -6575 46690 -6455
rect 46810 -6575 46865 -6455
rect 46985 -6575 47030 -6455
rect 47150 -6575 47195 -6455
rect 47315 -6575 47360 -6455
rect 47480 -6575 47535 -6455
rect 47655 -6575 47665 -6455
rect 42165 -6620 47665 -6575
rect 42165 -6740 42175 -6620
rect 42295 -6740 42340 -6620
rect 42460 -6740 42505 -6620
rect 42625 -6740 42670 -6620
rect 42790 -6740 42845 -6620
rect 42965 -6740 43010 -6620
rect 43130 -6740 43175 -6620
rect 43295 -6740 43340 -6620
rect 43460 -6740 43515 -6620
rect 43635 -6740 43680 -6620
rect 43800 -6740 43845 -6620
rect 43965 -6740 44010 -6620
rect 44130 -6740 44185 -6620
rect 44305 -6740 44350 -6620
rect 44470 -6740 44515 -6620
rect 44635 -6740 44680 -6620
rect 44800 -6740 44855 -6620
rect 44975 -6740 45020 -6620
rect 45140 -6740 45185 -6620
rect 45305 -6740 45350 -6620
rect 45470 -6740 45525 -6620
rect 45645 -6740 45690 -6620
rect 45810 -6740 45855 -6620
rect 45975 -6740 46020 -6620
rect 46140 -6740 46195 -6620
rect 46315 -6740 46360 -6620
rect 46480 -6740 46525 -6620
rect 46645 -6740 46690 -6620
rect 46810 -6740 46865 -6620
rect 46985 -6740 47030 -6620
rect 47150 -6740 47195 -6620
rect 47315 -6740 47360 -6620
rect 47480 -6740 47535 -6620
rect 47655 -6740 47665 -6620
rect 42165 -6785 47665 -6740
rect 42165 -6905 42175 -6785
rect 42295 -6905 42340 -6785
rect 42460 -6905 42505 -6785
rect 42625 -6905 42670 -6785
rect 42790 -6905 42845 -6785
rect 42965 -6905 43010 -6785
rect 43130 -6905 43175 -6785
rect 43295 -6905 43340 -6785
rect 43460 -6905 43515 -6785
rect 43635 -6905 43680 -6785
rect 43800 -6905 43845 -6785
rect 43965 -6905 44010 -6785
rect 44130 -6905 44185 -6785
rect 44305 -6905 44350 -6785
rect 44470 -6905 44515 -6785
rect 44635 -6905 44680 -6785
rect 44800 -6905 44855 -6785
rect 44975 -6905 45020 -6785
rect 45140 -6905 45185 -6785
rect 45305 -6905 45350 -6785
rect 45470 -6905 45525 -6785
rect 45645 -6905 45690 -6785
rect 45810 -6905 45855 -6785
rect 45975 -6905 46020 -6785
rect 46140 -6905 46195 -6785
rect 46315 -6905 46360 -6785
rect 46480 -6905 46525 -6785
rect 46645 -6905 46690 -6785
rect 46810 -6905 46865 -6785
rect 46985 -6905 47030 -6785
rect 47150 -6905 47195 -6785
rect 47315 -6905 47360 -6785
rect 47480 -6905 47535 -6785
rect 47655 -6905 47665 -6785
rect 42165 -6950 47665 -6905
rect 42165 -7070 42175 -6950
rect 42295 -7070 42340 -6950
rect 42460 -7070 42505 -6950
rect 42625 -7070 42670 -6950
rect 42790 -7070 42845 -6950
rect 42965 -7070 43010 -6950
rect 43130 -7070 43175 -6950
rect 43295 -7070 43340 -6950
rect 43460 -7070 43515 -6950
rect 43635 -7070 43680 -6950
rect 43800 -7070 43845 -6950
rect 43965 -7070 44010 -6950
rect 44130 -7070 44185 -6950
rect 44305 -7070 44350 -6950
rect 44470 -7070 44515 -6950
rect 44635 -7070 44680 -6950
rect 44800 -7070 44855 -6950
rect 44975 -7070 45020 -6950
rect 45140 -7070 45185 -6950
rect 45305 -7070 45350 -6950
rect 45470 -7070 45525 -6950
rect 45645 -7070 45690 -6950
rect 45810 -7070 45855 -6950
rect 45975 -7070 46020 -6950
rect 46140 -7070 46195 -6950
rect 46315 -7070 46360 -6950
rect 46480 -7070 46525 -6950
rect 46645 -7070 46690 -6950
rect 46810 -7070 46865 -6950
rect 46985 -7070 47030 -6950
rect 47150 -7070 47195 -6950
rect 47315 -7070 47360 -6950
rect 47480 -7070 47535 -6950
rect 47655 -7070 47665 -6950
rect 42165 -7125 47665 -7070
rect 42165 -7245 42175 -7125
rect 42295 -7245 42340 -7125
rect 42460 -7245 42505 -7125
rect 42625 -7245 42670 -7125
rect 42790 -7245 42845 -7125
rect 42965 -7245 43010 -7125
rect 43130 -7245 43175 -7125
rect 43295 -7245 43340 -7125
rect 43460 -7245 43515 -7125
rect 43635 -7245 43680 -7125
rect 43800 -7245 43845 -7125
rect 43965 -7245 44010 -7125
rect 44130 -7245 44185 -7125
rect 44305 -7245 44350 -7125
rect 44470 -7245 44515 -7125
rect 44635 -7245 44680 -7125
rect 44800 -7245 44855 -7125
rect 44975 -7245 45020 -7125
rect 45140 -7245 45185 -7125
rect 45305 -7245 45350 -7125
rect 45470 -7245 45525 -7125
rect 45645 -7245 45690 -7125
rect 45810 -7245 45855 -7125
rect 45975 -7245 46020 -7125
rect 46140 -7245 46195 -7125
rect 46315 -7245 46360 -7125
rect 46480 -7245 46525 -7125
rect 46645 -7245 46690 -7125
rect 46810 -7245 46865 -7125
rect 46985 -7245 47030 -7125
rect 47150 -7245 47195 -7125
rect 47315 -7245 47360 -7125
rect 47480 -7245 47535 -7125
rect 47655 -7245 47665 -7125
rect 42165 -7290 47665 -7245
rect 42165 -7410 42175 -7290
rect 42295 -7410 42340 -7290
rect 42460 -7410 42505 -7290
rect 42625 -7410 42670 -7290
rect 42790 -7410 42845 -7290
rect 42965 -7410 43010 -7290
rect 43130 -7410 43175 -7290
rect 43295 -7410 43340 -7290
rect 43460 -7410 43515 -7290
rect 43635 -7410 43680 -7290
rect 43800 -7410 43845 -7290
rect 43965 -7410 44010 -7290
rect 44130 -7410 44185 -7290
rect 44305 -7410 44350 -7290
rect 44470 -7410 44515 -7290
rect 44635 -7410 44680 -7290
rect 44800 -7410 44855 -7290
rect 44975 -7410 45020 -7290
rect 45140 -7410 45185 -7290
rect 45305 -7410 45350 -7290
rect 45470 -7410 45525 -7290
rect 45645 -7410 45690 -7290
rect 45810 -7410 45855 -7290
rect 45975 -7410 46020 -7290
rect 46140 -7410 46195 -7290
rect 46315 -7410 46360 -7290
rect 46480 -7410 46525 -7290
rect 46645 -7410 46690 -7290
rect 46810 -7410 46865 -7290
rect 46985 -7410 47030 -7290
rect 47150 -7410 47195 -7290
rect 47315 -7410 47360 -7290
rect 47480 -7410 47535 -7290
rect 47655 -7410 47665 -7290
rect 42165 -7455 47665 -7410
rect 42165 -7575 42175 -7455
rect 42295 -7575 42340 -7455
rect 42460 -7575 42505 -7455
rect 42625 -7575 42670 -7455
rect 42790 -7575 42845 -7455
rect 42965 -7575 43010 -7455
rect 43130 -7575 43175 -7455
rect 43295 -7575 43340 -7455
rect 43460 -7575 43515 -7455
rect 43635 -7575 43680 -7455
rect 43800 -7575 43845 -7455
rect 43965 -7575 44010 -7455
rect 44130 -7575 44185 -7455
rect 44305 -7575 44350 -7455
rect 44470 -7575 44515 -7455
rect 44635 -7575 44680 -7455
rect 44800 -7575 44855 -7455
rect 44975 -7575 45020 -7455
rect 45140 -7575 45185 -7455
rect 45305 -7575 45350 -7455
rect 45470 -7575 45525 -7455
rect 45645 -7575 45690 -7455
rect 45810 -7575 45855 -7455
rect 45975 -7575 46020 -7455
rect 46140 -7575 46195 -7455
rect 46315 -7575 46360 -7455
rect 46480 -7575 46525 -7455
rect 46645 -7575 46690 -7455
rect 46810 -7575 46865 -7455
rect 46985 -7575 47030 -7455
rect 47150 -7575 47195 -7455
rect 47315 -7575 47360 -7455
rect 47480 -7575 47535 -7455
rect 47655 -7575 47665 -7455
rect 42165 -7620 47665 -7575
rect 42165 -7740 42175 -7620
rect 42295 -7740 42340 -7620
rect 42460 -7740 42505 -7620
rect 42625 -7740 42670 -7620
rect 42790 -7740 42845 -7620
rect 42965 -7740 43010 -7620
rect 43130 -7740 43175 -7620
rect 43295 -7740 43340 -7620
rect 43460 -7740 43515 -7620
rect 43635 -7740 43680 -7620
rect 43800 -7740 43845 -7620
rect 43965 -7740 44010 -7620
rect 44130 -7740 44185 -7620
rect 44305 -7740 44350 -7620
rect 44470 -7740 44515 -7620
rect 44635 -7740 44680 -7620
rect 44800 -7740 44855 -7620
rect 44975 -7740 45020 -7620
rect 45140 -7740 45185 -7620
rect 45305 -7740 45350 -7620
rect 45470 -7740 45525 -7620
rect 45645 -7740 45690 -7620
rect 45810 -7740 45855 -7620
rect 45975 -7740 46020 -7620
rect 46140 -7740 46195 -7620
rect 46315 -7740 46360 -7620
rect 46480 -7740 46525 -7620
rect 46645 -7740 46690 -7620
rect 46810 -7740 46865 -7620
rect 46985 -7740 47030 -7620
rect 47150 -7740 47195 -7620
rect 47315 -7740 47360 -7620
rect 47480 -7740 47535 -7620
rect 47655 -7740 47665 -7620
rect 42165 -7795 47665 -7740
rect 42165 -7915 42175 -7795
rect 42295 -7915 42340 -7795
rect 42460 -7915 42505 -7795
rect 42625 -7915 42670 -7795
rect 42790 -7915 42845 -7795
rect 42965 -7915 43010 -7795
rect 43130 -7915 43175 -7795
rect 43295 -7915 43340 -7795
rect 43460 -7915 43515 -7795
rect 43635 -7915 43680 -7795
rect 43800 -7915 43845 -7795
rect 43965 -7915 44010 -7795
rect 44130 -7915 44185 -7795
rect 44305 -7915 44350 -7795
rect 44470 -7915 44515 -7795
rect 44635 -7915 44680 -7795
rect 44800 -7915 44855 -7795
rect 44975 -7915 45020 -7795
rect 45140 -7915 45185 -7795
rect 45305 -7915 45350 -7795
rect 45470 -7915 45525 -7795
rect 45645 -7915 45690 -7795
rect 45810 -7915 45855 -7795
rect 45975 -7915 46020 -7795
rect 46140 -7915 46195 -7795
rect 46315 -7915 46360 -7795
rect 46480 -7915 46525 -7795
rect 46645 -7915 46690 -7795
rect 46810 -7915 46865 -7795
rect 46985 -7915 47030 -7795
rect 47150 -7915 47195 -7795
rect 47315 -7915 47360 -7795
rect 47480 -7915 47535 -7795
rect 47655 -7915 47665 -7795
rect 42165 -7960 47665 -7915
rect 42165 -8080 42175 -7960
rect 42295 -8080 42340 -7960
rect 42460 -8080 42505 -7960
rect 42625 -8080 42670 -7960
rect 42790 -8080 42845 -7960
rect 42965 -8080 43010 -7960
rect 43130 -8080 43175 -7960
rect 43295 -8080 43340 -7960
rect 43460 -8080 43515 -7960
rect 43635 -8080 43680 -7960
rect 43800 -8080 43845 -7960
rect 43965 -8080 44010 -7960
rect 44130 -8080 44185 -7960
rect 44305 -8080 44350 -7960
rect 44470 -8080 44515 -7960
rect 44635 -8080 44680 -7960
rect 44800 -8080 44855 -7960
rect 44975 -8080 45020 -7960
rect 45140 -8080 45185 -7960
rect 45305 -8080 45350 -7960
rect 45470 -8080 45525 -7960
rect 45645 -8080 45690 -7960
rect 45810 -8080 45855 -7960
rect 45975 -8080 46020 -7960
rect 46140 -8080 46195 -7960
rect 46315 -8080 46360 -7960
rect 46480 -8080 46525 -7960
rect 46645 -8080 46690 -7960
rect 46810 -8080 46865 -7960
rect 46985 -8080 47030 -7960
rect 47150 -8080 47195 -7960
rect 47315 -8080 47360 -7960
rect 47480 -8080 47535 -7960
rect 47655 -8080 47665 -7960
rect 42165 -8125 47665 -8080
rect 42165 -8245 42175 -8125
rect 42295 -8245 42340 -8125
rect 42460 -8245 42505 -8125
rect 42625 -8245 42670 -8125
rect 42790 -8245 42845 -8125
rect 42965 -8245 43010 -8125
rect 43130 -8245 43175 -8125
rect 43295 -8245 43340 -8125
rect 43460 -8245 43515 -8125
rect 43635 -8245 43680 -8125
rect 43800 -8245 43845 -8125
rect 43965 -8245 44010 -8125
rect 44130 -8245 44185 -8125
rect 44305 -8245 44350 -8125
rect 44470 -8245 44515 -8125
rect 44635 -8245 44680 -8125
rect 44800 -8245 44855 -8125
rect 44975 -8245 45020 -8125
rect 45140 -8245 45185 -8125
rect 45305 -8245 45350 -8125
rect 45470 -8245 45525 -8125
rect 45645 -8245 45690 -8125
rect 45810 -8245 45855 -8125
rect 45975 -8245 46020 -8125
rect 46140 -8245 46195 -8125
rect 46315 -8245 46360 -8125
rect 46480 -8245 46525 -8125
rect 46645 -8245 46690 -8125
rect 46810 -8245 46865 -8125
rect 46985 -8245 47030 -8125
rect 47150 -8245 47195 -8125
rect 47315 -8245 47360 -8125
rect 47480 -8245 47535 -8125
rect 47655 -8245 47665 -8125
rect 42165 -8290 47665 -8245
rect 42165 -8410 42175 -8290
rect 42295 -8410 42340 -8290
rect 42460 -8410 42505 -8290
rect 42625 -8410 42670 -8290
rect 42790 -8410 42845 -8290
rect 42965 -8410 43010 -8290
rect 43130 -8410 43175 -8290
rect 43295 -8410 43340 -8290
rect 43460 -8410 43515 -8290
rect 43635 -8410 43680 -8290
rect 43800 -8410 43845 -8290
rect 43965 -8410 44010 -8290
rect 44130 -8410 44185 -8290
rect 44305 -8410 44350 -8290
rect 44470 -8410 44515 -8290
rect 44635 -8410 44680 -8290
rect 44800 -8410 44855 -8290
rect 44975 -8410 45020 -8290
rect 45140 -8410 45185 -8290
rect 45305 -8410 45350 -8290
rect 45470 -8410 45525 -8290
rect 45645 -8410 45690 -8290
rect 45810 -8410 45855 -8290
rect 45975 -8410 46020 -8290
rect 46140 -8410 46195 -8290
rect 46315 -8410 46360 -8290
rect 46480 -8410 46525 -8290
rect 46645 -8410 46690 -8290
rect 46810 -8410 46865 -8290
rect 46985 -8410 47030 -8290
rect 47150 -8410 47195 -8290
rect 47315 -8410 47360 -8290
rect 47480 -8410 47535 -8290
rect 47655 -8410 47665 -8290
rect 42165 -8465 47665 -8410
rect 42165 -8585 42175 -8465
rect 42295 -8585 42340 -8465
rect 42460 -8585 42505 -8465
rect 42625 -8585 42670 -8465
rect 42790 -8585 42845 -8465
rect 42965 -8585 43010 -8465
rect 43130 -8585 43175 -8465
rect 43295 -8585 43340 -8465
rect 43460 -8585 43515 -8465
rect 43635 -8585 43680 -8465
rect 43800 -8585 43845 -8465
rect 43965 -8585 44010 -8465
rect 44130 -8585 44185 -8465
rect 44305 -8585 44350 -8465
rect 44470 -8585 44515 -8465
rect 44635 -8585 44680 -8465
rect 44800 -8585 44855 -8465
rect 44975 -8585 45020 -8465
rect 45140 -8585 45185 -8465
rect 45305 -8585 45350 -8465
rect 45470 -8585 45525 -8465
rect 45645 -8585 45690 -8465
rect 45810 -8585 45855 -8465
rect 45975 -8585 46020 -8465
rect 46140 -8585 46195 -8465
rect 46315 -8585 46360 -8465
rect 46480 -8585 46525 -8465
rect 46645 -8585 46690 -8465
rect 46810 -8585 46865 -8465
rect 46985 -8585 47030 -8465
rect 47150 -8585 47195 -8465
rect 47315 -8585 47360 -8465
rect 47480 -8585 47535 -8465
rect 47655 -8585 47665 -8465
rect 42165 -8630 47665 -8585
rect 42165 -8750 42175 -8630
rect 42295 -8750 42340 -8630
rect 42460 -8750 42505 -8630
rect 42625 -8750 42670 -8630
rect 42790 -8750 42845 -8630
rect 42965 -8750 43010 -8630
rect 43130 -8750 43175 -8630
rect 43295 -8750 43340 -8630
rect 43460 -8750 43515 -8630
rect 43635 -8750 43680 -8630
rect 43800 -8750 43845 -8630
rect 43965 -8750 44010 -8630
rect 44130 -8750 44185 -8630
rect 44305 -8750 44350 -8630
rect 44470 -8750 44515 -8630
rect 44635 -8750 44680 -8630
rect 44800 -8750 44855 -8630
rect 44975 -8750 45020 -8630
rect 45140 -8750 45185 -8630
rect 45305 -8750 45350 -8630
rect 45470 -8750 45525 -8630
rect 45645 -8750 45690 -8630
rect 45810 -8750 45855 -8630
rect 45975 -8750 46020 -8630
rect 46140 -8750 46195 -8630
rect 46315 -8750 46360 -8630
rect 46480 -8750 46525 -8630
rect 46645 -8750 46690 -8630
rect 46810 -8750 46865 -8630
rect 46985 -8750 47030 -8630
rect 47150 -8750 47195 -8630
rect 47315 -8750 47360 -8630
rect 47480 -8750 47535 -8630
rect 47655 -8750 47665 -8630
rect 42165 -8795 47665 -8750
rect 42165 -8915 42175 -8795
rect 42295 -8915 42340 -8795
rect 42460 -8915 42505 -8795
rect 42625 -8915 42670 -8795
rect 42790 -8915 42845 -8795
rect 42965 -8915 43010 -8795
rect 43130 -8915 43175 -8795
rect 43295 -8915 43340 -8795
rect 43460 -8915 43515 -8795
rect 43635 -8915 43680 -8795
rect 43800 -8915 43845 -8795
rect 43965 -8915 44010 -8795
rect 44130 -8915 44185 -8795
rect 44305 -8915 44350 -8795
rect 44470 -8915 44515 -8795
rect 44635 -8915 44680 -8795
rect 44800 -8915 44855 -8795
rect 44975 -8915 45020 -8795
rect 45140 -8915 45185 -8795
rect 45305 -8915 45350 -8795
rect 45470 -8915 45525 -8795
rect 45645 -8915 45690 -8795
rect 45810 -8915 45855 -8795
rect 45975 -8915 46020 -8795
rect 46140 -8915 46195 -8795
rect 46315 -8915 46360 -8795
rect 46480 -8915 46525 -8795
rect 46645 -8915 46690 -8795
rect 46810 -8915 46865 -8795
rect 46985 -8915 47030 -8795
rect 47150 -8915 47195 -8795
rect 47315 -8915 47360 -8795
rect 47480 -8915 47535 -8795
rect 47655 -8915 47665 -8795
rect 42165 -8960 47665 -8915
rect 42165 -9080 42175 -8960
rect 42295 -9080 42340 -8960
rect 42460 -9080 42505 -8960
rect 42625 -9080 42670 -8960
rect 42790 -9080 42845 -8960
rect 42965 -9080 43010 -8960
rect 43130 -9080 43175 -8960
rect 43295 -9080 43340 -8960
rect 43460 -9080 43515 -8960
rect 43635 -9080 43680 -8960
rect 43800 -9080 43845 -8960
rect 43965 -9080 44010 -8960
rect 44130 -9080 44185 -8960
rect 44305 -9080 44350 -8960
rect 44470 -9080 44515 -8960
rect 44635 -9080 44680 -8960
rect 44800 -9080 44855 -8960
rect 44975 -9080 45020 -8960
rect 45140 -9080 45185 -8960
rect 45305 -9080 45350 -8960
rect 45470 -9080 45525 -8960
rect 45645 -9080 45690 -8960
rect 45810 -9080 45855 -8960
rect 45975 -9080 46020 -8960
rect 46140 -9080 46195 -8960
rect 46315 -9080 46360 -8960
rect 46480 -9080 46525 -8960
rect 46645 -9080 46690 -8960
rect 46810 -9080 46865 -8960
rect 46985 -9080 47030 -8960
rect 47150 -9080 47195 -8960
rect 47315 -9080 47360 -8960
rect 47480 -9080 47535 -8960
rect 47655 -9080 47665 -8960
rect 42165 -9135 47665 -9080
rect 42165 -9255 42175 -9135
rect 42295 -9255 42340 -9135
rect 42460 -9255 42505 -9135
rect 42625 -9255 42670 -9135
rect 42790 -9255 42845 -9135
rect 42965 -9255 43010 -9135
rect 43130 -9255 43175 -9135
rect 43295 -9255 43340 -9135
rect 43460 -9255 43515 -9135
rect 43635 -9255 43680 -9135
rect 43800 -9255 43845 -9135
rect 43965 -9255 44010 -9135
rect 44130 -9255 44185 -9135
rect 44305 -9255 44350 -9135
rect 44470 -9255 44515 -9135
rect 44635 -9255 44680 -9135
rect 44800 -9255 44855 -9135
rect 44975 -9255 45020 -9135
rect 45140 -9255 45185 -9135
rect 45305 -9255 45350 -9135
rect 45470 -9255 45525 -9135
rect 45645 -9255 45690 -9135
rect 45810 -9255 45855 -9135
rect 45975 -9255 46020 -9135
rect 46140 -9255 46195 -9135
rect 46315 -9255 46360 -9135
rect 46480 -9255 46525 -9135
rect 46645 -9255 46690 -9135
rect 46810 -9255 46865 -9135
rect 46985 -9255 47030 -9135
rect 47150 -9255 47195 -9135
rect 47315 -9255 47360 -9135
rect 47480 -9255 47535 -9135
rect 47655 -9255 47665 -9135
rect 42165 -9300 47665 -9255
rect 42165 -9420 42175 -9300
rect 42295 -9420 42340 -9300
rect 42460 -9420 42505 -9300
rect 42625 -9420 42670 -9300
rect 42790 -9420 42845 -9300
rect 42965 -9420 43010 -9300
rect 43130 -9420 43175 -9300
rect 43295 -9420 43340 -9300
rect 43460 -9420 43515 -9300
rect 43635 -9420 43680 -9300
rect 43800 -9420 43845 -9300
rect 43965 -9420 44010 -9300
rect 44130 -9420 44185 -9300
rect 44305 -9420 44350 -9300
rect 44470 -9420 44515 -9300
rect 44635 -9420 44680 -9300
rect 44800 -9420 44855 -9300
rect 44975 -9420 45020 -9300
rect 45140 -9420 45185 -9300
rect 45305 -9420 45350 -9300
rect 45470 -9420 45525 -9300
rect 45645 -9420 45690 -9300
rect 45810 -9420 45855 -9300
rect 45975 -9420 46020 -9300
rect 46140 -9420 46195 -9300
rect 46315 -9420 46360 -9300
rect 46480 -9420 46525 -9300
rect 46645 -9420 46690 -9300
rect 46810 -9420 46865 -9300
rect 46985 -9420 47030 -9300
rect 47150 -9420 47195 -9300
rect 47315 -9420 47360 -9300
rect 47480 -9420 47535 -9300
rect 47655 -9420 47665 -9300
rect 42165 -9465 47665 -9420
rect 42165 -9585 42175 -9465
rect 42295 -9585 42340 -9465
rect 42460 -9585 42505 -9465
rect 42625 -9585 42670 -9465
rect 42790 -9585 42845 -9465
rect 42965 -9585 43010 -9465
rect 43130 -9585 43175 -9465
rect 43295 -9585 43340 -9465
rect 43460 -9585 43515 -9465
rect 43635 -9585 43680 -9465
rect 43800 -9585 43845 -9465
rect 43965 -9585 44010 -9465
rect 44130 -9585 44185 -9465
rect 44305 -9585 44350 -9465
rect 44470 -9585 44515 -9465
rect 44635 -9585 44680 -9465
rect 44800 -9585 44855 -9465
rect 44975 -9585 45020 -9465
rect 45140 -9585 45185 -9465
rect 45305 -9585 45350 -9465
rect 45470 -9585 45525 -9465
rect 45645 -9585 45690 -9465
rect 45810 -9585 45855 -9465
rect 45975 -9585 46020 -9465
rect 46140 -9585 46195 -9465
rect 46315 -9585 46360 -9465
rect 46480 -9585 46525 -9465
rect 46645 -9585 46690 -9465
rect 46810 -9585 46865 -9465
rect 46985 -9585 47030 -9465
rect 47150 -9585 47195 -9465
rect 47315 -9585 47360 -9465
rect 47480 -9585 47535 -9465
rect 47655 -9585 47665 -9465
rect 42165 -9630 47665 -9585
rect 42165 -9750 42175 -9630
rect 42295 -9750 42340 -9630
rect 42460 -9750 42505 -9630
rect 42625 -9750 42670 -9630
rect 42790 -9750 42845 -9630
rect 42965 -9750 43010 -9630
rect 43130 -9750 43175 -9630
rect 43295 -9750 43340 -9630
rect 43460 -9750 43515 -9630
rect 43635 -9750 43680 -9630
rect 43800 -9750 43845 -9630
rect 43965 -9750 44010 -9630
rect 44130 -9750 44185 -9630
rect 44305 -9750 44350 -9630
rect 44470 -9750 44515 -9630
rect 44635 -9750 44680 -9630
rect 44800 -9750 44855 -9630
rect 44975 -9750 45020 -9630
rect 45140 -9750 45185 -9630
rect 45305 -9750 45350 -9630
rect 45470 -9750 45525 -9630
rect 45645 -9750 45690 -9630
rect 45810 -9750 45855 -9630
rect 45975 -9750 46020 -9630
rect 46140 -9750 46195 -9630
rect 46315 -9750 46360 -9630
rect 46480 -9750 46525 -9630
rect 46645 -9750 46690 -9630
rect 46810 -9750 46865 -9630
rect 46985 -9750 47030 -9630
rect 47150 -9750 47195 -9630
rect 47315 -9750 47360 -9630
rect 47480 -9750 47535 -9630
rect 47655 -9750 47665 -9630
rect 42165 -9760 47665 -9750
rect 47855 -4270 53355 -4260
rect 47855 -4390 47865 -4270
rect 47985 -4390 48030 -4270
rect 48150 -4390 48195 -4270
rect 48315 -4390 48360 -4270
rect 48480 -4390 48535 -4270
rect 48655 -4390 48700 -4270
rect 48820 -4390 48865 -4270
rect 48985 -4390 49030 -4270
rect 49150 -4390 49205 -4270
rect 49325 -4390 49370 -4270
rect 49490 -4390 49535 -4270
rect 49655 -4390 49700 -4270
rect 49820 -4390 49875 -4270
rect 49995 -4390 50040 -4270
rect 50160 -4390 50205 -4270
rect 50325 -4390 50370 -4270
rect 50490 -4390 50545 -4270
rect 50665 -4390 50710 -4270
rect 50830 -4390 50875 -4270
rect 50995 -4390 51040 -4270
rect 51160 -4390 51215 -4270
rect 51335 -4390 51380 -4270
rect 51500 -4390 51545 -4270
rect 51665 -4390 51710 -4270
rect 51830 -4390 51885 -4270
rect 52005 -4390 52050 -4270
rect 52170 -4390 52215 -4270
rect 52335 -4390 52380 -4270
rect 52500 -4390 52555 -4270
rect 52675 -4390 52720 -4270
rect 52840 -4390 52885 -4270
rect 53005 -4390 53050 -4270
rect 53170 -4390 53225 -4270
rect 53345 -4390 53355 -4270
rect 47855 -4445 53355 -4390
rect 47855 -4565 47865 -4445
rect 47985 -4565 48030 -4445
rect 48150 -4565 48195 -4445
rect 48315 -4565 48360 -4445
rect 48480 -4565 48535 -4445
rect 48655 -4565 48700 -4445
rect 48820 -4565 48865 -4445
rect 48985 -4565 49030 -4445
rect 49150 -4565 49205 -4445
rect 49325 -4565 49370 -4445
rect 49490 -4565 49535 -4445
rect 49655 -4565 49700 -4445
rect 49820 -4565 49875 -4445
rect 49995 -4565 50040 -4445
rect 50160 -4565 50205 -4445
rect 50325 -4565 50370 -4445
rect 50490 -4565 50545 -4445
rect 50665 -4565 50710 -4445
rect 50830 -4565 50875 -4445
rect 50995 -4565 51040 -4445
rect 51160 -4565 51215 -4445
rect 51335 -4565 51380 -4445
rect 51500 -4565 51545 -4445
rect 51665 -4565 51710 -4445
rect 51830 -4565 51885 -4445
rect 52005 -4565 52050 -4445
rect 52170 -4565 52215 -4445
rect 52335 -4565 52380 -4445
rect 52500 -4565 52555 -4445
rect 52675 -4565 52720 -4445
rect 52840 -4565 52885 -4445
rect 53005 -4565 53050 -4445
rect 53170 -4565 53225 -4445
rect 53345 -4565 53355 -4445
rect 47855 -4610 53355 -4565
rect 47855 -4730 47865 -4610
rect 47985 -4730 48030 -4610
rect 48150 -4730 48195 -4610
rect 48315 -4730 48360 -4610
rect 48480 -4730 48535 -4610
rect 48655 -4730 48700 -4610
rect 48820 -4730 48865 -4610
rect 48985 -4730 49030 -4610
rect 49150 -4730 49205 -4610
rect 49325 -4730 49370 -4610
rect 49490 -4730 49535 -4610
rect 49655 -4730 49700 -4610
rect 49820 -4730 49875 -4610
rect 49995 -4730 50040 -4610
rect 50160 -4730 50205 -4610
rect 50325 -4730 50370 -4610
rect 50490 -4730 50545 -4610
rect 50665 -4730 50710 -4610
rect 50830 -4730 50875 -4610
rect 50995 -4730 51040 -4610
rect 51160 -4730 51215 -4610
rect 51335 -4730 51380 -4610
rect 51500 -4730 51545 -4610
rect 51665 -4730 51710 -4610
rect 51830 -4730 51885 -4610
rect 52005 -4730 52050 -4610
rect 52170 -4730 52215 -4610
rect 52335 -4730 52380 -4610
rect 52500 -4730 52555 -4610
rect 52675 -4730 52720 -4610
rect 52840 -4730 52885 -4610
rect 53005 -4730 53050 -4610
rect 53170 -4730 53225 -4610
rect 53345 -4730 53355 -4610
rect 47855 -4775 53355 -4730
rect 47855 -4895 47865 -4775
rect 47985 -4895 48030 -4775
rect 48150 -4895 48195 -4775
rect 48315 -4895 48360 -4775
rect 48480 -4895 48535 -4775
rect 48655 -4895 48700 -4775
rect 48820 -4895 48865 -4775
rect 48985 -4895 49030 -4775
rect 49150 -4895 49205 -4775
rect 49325 -4895 49370 -4775
rect 49490 -4895 49535 -4775
rect 49655 -4895 49700 -4775
rect 49820 -4895 49875 -4775
rect 49995 -4895 50040 -4775
rect 50160 -4895 50205 -4775
rect 50325 -4895 50370 -4775
rect 50490 -4895 50545 -4775
rect 50665 -4895 50710 -4775
rect 50830 -4895 50875 -4775
rect 50995 -4895 51040 -4775
rect 51160 -4895 51215 -4775
rect 51335 -4895 51380 -4775
rect 51500 -4895 51545 -4775
rect 51665 -4895 51710 -4775
rect 51830 -4895 51885 -4775
rect 52005 -4895 52050 -4775
rect 52170 -4895 52215 -4775
rect 52335 -4895 52380 -4775
rect 52500 -4895 52555 -4775
rect 52675 -4895 52720 -4775
rect 52840 -4895 52885 -4775
rect 53005 -4895 53050 -4775
rect 53170 -4895 53225 -4775
rect 53345 -4895 53355 -4775
rect 47855 -4940 53355 -4895
rect 47855 -5060 47865 -4940
rect 47985 -5060 48030 -4940
rect 48150 -5060 48195 -4940
rect 48315 -5060 48360 -4940
rect 48480 -5060 48535 -4940
rect 48655 -5060 48700 -4940
rect 48820 -5060 48865 -4940
rect 48985 -5060 49030 -4940
rect 49150 -5060 49205 -4940
rect 49325 -5060 49370 -4940
rect 49490 -5060 49535 -4940
rect 49655 -5060 49700 -4940
rect 49820 -5060 49875 -4940
rect 49995 -5060 50040 -4940
rect 50160 -5060 50205 -4940
rect 50325 -5060 50370 -4940
rect 50490 -5060 50545 -4940
rect 50665 -5060 50710 -4940
rect 50830 -5060 50875 -4940
rect 50995 -5060 51040 -4940
rect 51160 -5060 51215 -4940
rect 51335 -5060 51380 -4940
rect 51500 -5060 51545 -4940
rect 51665 -5060 51710 -4940
rect 51830 -5060 51885 -4940
rect 52005 -5060 52050 -4940
rect 52170 -5060 52215 -4940
rect 52335 -5060 52380 -4940
rect 52500 -5060 52555 -4940
rect 52675 -5060 52720 -4940
rect 52840 -5060 52885 -4940
rect 53005 -5060 53050 -4940
rect 53170 -5060 53225 -4940
rect 53345 -5060 53355 -4940
rect 47855 -5115 53355 -5060
rect 47855 -5235 47865 -5115
rect 47985 -5235 48030 -5115
rect 48150 -5235 48195 -5115
rect 48315 -5235 48360 -5115
rect 48480 -5235 48535 -5115
rect 48655 -5235 48700 -5115
rect 48820 -5235 48865 -5115
rect 48985 -5235 49030 -5115
rect 49150 -5235 49205 -5115
rect 49325 -5235 49370 -5115
rect 49490 -5235 49535 -5115
rect 49655 -5235 49700 -5115
rect 49820 -5235 49875 -5115
rect 49995 -5235 50040 -5115
rect 50160 -5235 50205 -5115
rect 50325 -5235 50370 -5115
rect 50490 -5235 50545 -5115
rect 50665 -5235 50710 -5115
rect 50830 -5235 50875 -5115
rect 50995 -5235 51040 -5115
rect 51160 -5235 51215 -5115
rect 51335 -5235 51380 -5115
rect 51500 -5235 51545 -5115
rect 51665 -5235 51710 -5115
rect 51830 -5235 51885 -5115
rect 52005 -5235 52050 -5115
rect 52170 -5235 52215 -5115
rect 52335 -5235 52380 -5115
rect 52500 -5235 52555 -5115
rect 52675 -5235 52720 -5115
rect 52840 -5235 52885 -5115
rect 53005 -5235 53050 -5115
rect 53170 -5235 53225 -5115
rect 53345 -5235 53355 -5115
rect 47855 -5280 53355 -5235
rect 47855 -5400 47865 -5280
rect 47985 -5400 48030 -5280
rect 48150 -5400 48195 -5280
rect 48315 -5400 48360 -5280
rect 48480 -5400 48535 -5280
rect 48655 -5400 48700 -5280
rect 48820 -5400 48865 -5280
rect 48985 -5400 49030 -5280
rect 49150 -5400 49205 -5280
rect 49325 -5400 49370 -5280
rect 49490 -5400 49535 -5280
rect 49655 -5400 49700 -5280
rect 49820 -5400 49875 -5280
rect 49995 -5400 50040 -5280
rect 50160 -5400 50205 -5280
rect 50325 -5400 50370 -5280
rect 50490 -5400 50545 -5280
rect 50665 -5400 50710 -5280
rect 50830 -5400 50875 -5280
rect 50995 -5400 51040 -5280
rect 51160 -5400 51215 -5280
rect 51335 -5400 51380 -5280
rect 51500 -5400 51545 -5280
rect 51665 -5400 51710 -5280
rect 51830 -5400 51885 -5280
rect 52005 -5400 52050 -5280
rect 52170 -5400 52215 -5280
rect 52335 -5400 52380 -5280
rect 52500 -5400 52555 -5280
rect 52675 -5400 52720 -5280
rect 52840 -5400 52885 -5280
rect 53005 -5400 53050 -5280
rect 53170 -5400 53225 -5280
rect 53345 -5400 53355 -5280
rect 47855 -5445 53355 -5400
rect 47855 -5565 47865 -5445
rect 47985 -5565 48030 -5445
rect 48150 -5565 48195 -5445
rect 48315 -5565 48360 -5445
rect 48480 -5565 48535 -5445
rect 48655 -5565 48700 -5445
rect 48820 -5565 48865 -5445
rect 48985 -5565 49030 -5445
rect 49150 -5565 49205 -5445
rect 49325 -5565 49370 -5445
rect 49490 -5565 49535 -5445
rect 49655 -5565 49700 -5445
rect 49820 -5565 49875 -5445
rect 49995 -5565 50040 -5445
rect 50160 -5565 50205 -5445
rect 50325 -5565 50370 -5445
rect 50490 -5565 50545 -5445
rect 50665 -5565 50710 -5445
rect 50830 -5565 50875 -5445
rect 50995 -5565 51040 -5445
rect 51160 -5565 51215 -5445
rect 51335 -5565 51380 -5445
rect 51500 -5565 51545 -5445
rect 51665 -5565 51710 -5445
rect 51830 -5565 51885 -5445
rect 52005 -5565 52050 -5445
rect 52170 -5565 52215 -5445
rect 52335 -5565 52380 -5445
rect 52500 -5565 52555 -5445
rect 52675 -5565 52720 -5445
rect 52840 -5565 52885 -5445
rect 53005 -5565 53050 -5445
rect 53170 -5565 53225 -5445
rect 53345 -5565 53355 -5445
rect 47855 -5610 53355 -5565
rect 47855 -5730 47865 -5610
rect 47985 -5730 48030 -5610
rect 48150 -5730 48195 -5610
rect 48315 -5730 48360 -5610
rect 48480 -5730 48535 -5610
rect 48655 -5730 48700 -5610
rect 48820 -5730 48865 -5610
rect 48985 -5730 49030 -5610
rect 49150 -5730 49205 -5610
rect 49325 -5730 49370 -5610
rect 49490 -5730 49535 -5610
rect 49655 -5730 49700 -5610
rect 49820 -5730 49875 -5610
rect 49995 -5730 50040 -5610
rect 50160 -5730 50205 -5610
rect 50325 -5730 50370 -5610
rect 50490 -5730 50545 -5610
rect 50665 -5730 50710 -5610
rect 50830 -5730 50875 -5610
rect 50995 -5730 51040 -5610
rect 51160 -5730 51215 -5610
rect 51335 -5730 51380 -5610
rect 51500 -5730 51545 -5610
rect 51665 -5730 51710 -5610
rect 51830 -5730 51885 -5610
rect 52005 -5730 52050 -5610
rect 52170 -5730 52215 -5610
rect 52335 -5730 52380 -5610
rect 52500 -5730 52555 -5610
rect 52675 -5730 52720 -5610
rect 52840 -5730 52885 -5610
rect 53005 -5730 53050 -5610
rect 53170 -5730 53225 -5610
rect 53345 -5730 53355 -5610
rect 47855 -5785 53355 -5730
rect 47855 -5905 47865 -5785
rect 47985 -5905 48030 -5785
rect 48150 -5905 48195 -5785
rect 48315 -5905 48360 -5785
rect 48480 -5905 48535 -5785
rect 48655 -5905 48700 -5785
rect 48820 -5905 48865 -5785
rect 48985 -5905 49030 -5785
rect 49150 -5905 49205 -5785
rect 49325 -5905 49370 -5785
rect 49490 -5905 49535 -5785
rect 49655 -5905 49700 -5785
rect 49820 -5905 49875 -5785
rect 49995 -5905 50040 -5785
rect 50160 -5905 50205 -5785
rect 50325 -5905 50370 -5785
rect 50490 -5905 50545 -5785
rect 50665 -5905 50710 -5785
rect 50830 -5905 50875 -5785
rect 50995 -5905 51040 -5785
rect 51160 -5905 51215 -5785
rect 51335 -5905 51380 -5785
rect 51500 -5905 51545 -5785
rect 51665 -5905 51710 -5785
rect 51830 -5905 51885 -5785
rect 52005 -5905 52050 -5785
rect 52170 -5905 52215 -5785
rect 52335 -5905 52380 -5785
rect 52500 -5905 52555 -5785
rect 52675 -5905 52720 -5785
rect 52840 -5905 52885 -5785
rect 53005 -5905 53050 -5785
rect 53170 -5905 53225 -5785
rect 53345 -5905 53355 -5785
rect 47855 -5950 53355 -5905
rect 47855 -6070 47865 -5950
rect 47985 -6070 48030 -5950
rect 48150 -6070 48195 -5950
rect 48315 -6070 48360 -5950
rect 48480 -6070 48535 -5950
rect 48655 -6070 48700 -5950
rect 48820 -6070 48865 -5950
rect 48985 -6070 49030 -5950
rect 49150 -6070 49205 -5950
rect 49325 -6070 49370 -5950
rect 49490 -6070 49535 -5950
rect 49655 -6070 49700 -5950
rect 49820 -6070 49875 -5950
rect 49995 -6070 50040 -5950
rect 50160 -6070 50205 -5950
rect 50325 -6070 50370 -5950
rect 50490 -6070 50545 -5950
rect 50665 -6070 50710 -5950
rect 50830 -6070 50875 -5950
rect 50995 -6070 51040 -5950
rect 51160 -6070 51215 -5950
rect 51335 -6070 51380 -5950
rect 51500 -6070 51545 -5950
rect 51665 -6070 51710 -5950
rect 51830 -6070 51885 -5950
rect 52005 -6070 52050 -5950
rect 52170 -6070 52215 -5950
rect 52335 -6070 52380 -5950
rect 52500 -6070 52555 -5950
rect 52675 -6070 52720 -5950
rect 52840 -6070 52885 -5950
rect 53005 -6070 53050 -5950
rect 53170 -6070 53225 -5950
rect 53345 -6070 53355 -5950
rect 47855 -6115 53355 -6070
rect 47855 -6235 47865 -6115
rect 47985 -6235 48030 -6115
rect 48150 -6235 48195 -6115
rect 48315 -6235 48360 -6115
rect 48480 -6235 48535 -6115
rect 48655 -6235 48700 -6115
rect 48820 -6235 48865 -6115
rect 48985 -6235 49030 -6115
rect 49150 -6235 49205 -6115
rect 49325 -6235 49370 -6115
rect 49490 -6235 49535 -6115
rect 49655 -6235 49700 -6115
rect 49820 -6235 49875 -6115
rect 49995 -6235 50040 -6115
rect 50160 -6235 50205 -6115
rect 50325 -6235 50370 -6115
rect 50490 -6235 50545 -6115
rect 50665 -6235 50710 -6115
rect 50830 -6235 50875 -6115
rect 50995 -6235 51040 -6115
rect 51160 -6235 51215 -6115
rect 51335 -6235 51380 -6115
rect 51500 -6235 51545 -6115
rect 51665 -6235 51710 -6115
rect 51830 -6235 51885 -6115
rect 52005 -6235 52050 -6115
rect 52170 -6235 52215 -6115
rect 52335 -6235 52380 -6115
rect 52500 -6235 52555 -6115
rect 52675 -6235 52720 -6115
rect 52840 -6235 52885 -6115
rect 53005 -6235 53050 -6115
rect 53170 -6235 53225 -6115
rect 53345 -6235 53355 -6115
rect 47855 -6280 53355 -6235
rect 47855 -6400 47865 -6280
rect 47985 -6400 48030 -6280
rect 48150 -6400 48195 -6280
rect 48315 -6400 48360 -6280
rect 48480 -6400 48535 -6280
rect 48655 -6400 48700 -6280
rect 48820 -6400 48865 -6280
rect 48985 -6400 49030 -6280
rect 49150 -6400 49205 -6280
rect 49325 -6400 49370 -6280
rect 49490 -6400 49535 -6280
rect 49655 -6400 49700 -6280
rect 49820 -6400 49875 -6280
rect 49995 -6400 50040 -6280
rect 50160 -6400 50205 -6280
rect 50325 -6400 50370 -6280
rect 50490 -6400 50545 -6280
rect 50665 -6400 50710 -6280
rect 50830 -6400 50875 -6280
rect 50995 -6400 51040 -6280
rect 51160 -6400 51215 -6280
rect 51335 -6400 51380 -6280
rect 51500 -6400 51545 -6280
rect 51665 -6400 51710 -6280
rect 51830 -6400 51885 -6280
rect 52005 -6400 52050 -6280
rect 52170 -6400 52215 -6280
rect 52335 -6400 52380 -6280
rect 52500 -6400 52555 -6280
rect 52675 -6400 52720 -6280
rect 52840 -6400 52885 -6280
rect 53005 -6400 53050 -6280
rect 53170 -6400 53225 -6280
rect 53345 -6400 53355 -6280
rect 47855 -6455 53355 -6400
rect 47855 -6575 47865 -6455
rect 47985 -6575 48030 -6455
rect 48150 -6575 48195 -6455
rect 48315 -6575 48360 -6455
rect 48480 -6575 48535 -6455
rect 48655 -6575 48700 -6455
rect 48820 -6575 48865 -6455
rect 48985 -6575 49030 -6455
rect 49150 -6575 49205 -6455
rect 49325 -6575 49370 -6455
rect 49490 -6575 49535 -6455
rect 49655 -6575 49700 -6455
rect 49820 -6575 49875 -6455
rect 49995 -6575 50040 -6455
rect 50160 -6575 50205 -6455
rect 50325 -6575 50370 -6455
rect 50490 -6575 50545 -6455
rect 50665 -6575 50710 -6455
rect 50830 -6575 50875 -6455
rect 50995 -6575 51040 -6455
rect 51160 -6575 51215 -6455
rect 51335 -6575 51380 -6455
rect 51500 -6575 51545 -6455
rect 51665 -6575 51710 -6455
rect 51830 -6575 51885 -6455
rect 52005 -6575 52050 -6455
rect 52170 -6575 52215 -6455
rect 52335 -6575 52380 -6455
rect 52500 -6575 52555 -6455
rect 52675 -6575 52720 -6455
rect 52840 -6575 52885 -6455
rect 53005 -6575 53050 -6455
rect 53170 -6575 53225 -6455
rect 53345 -6575 53355 -6455
rect 47855 -6620 53355 -6575
rect 47855 -6740 47865 -6620
rect 47985 -6740 48030 -6620
rect 48150 -6740 48195 -6620
rect 48315 -6740 48360 -6620
rect 48480 -6740 48535 -6620
rect 48655 -6740 48700 -6620
rect 48820 -6740 48865 -6620
rect 48985 -6740 49030 -6620
rect 49150 -6740 49205 -6620
rect 49325 -6740 49370 -6620
rect 49490 -6740 49535 -6620
rect 49655 -6740 49700 -6620
rect 49820 -6740 49875 -6620
rect 49995 -6740 50040 -6620
rect 50160 -6740 50205 -6620
rect 50325 -6740 50370 -6620
rect 50490 -6740 50545 -6620
rect 50665 -6740 50710 -6620
rect 50830 -6740 50875 -6620
rect 50995 -6740 51040 -6620
rect 51160 -6740 51215 -6620
rect 51335 -6740 51380 -6620
rect 51500 -6740 51545 -6620
rect 51665 -6740 51710 -6620
rect 51830 -6740 51885 -6620
rect 52005 -6740 52050 -6620
rect 52170 -6740 52215 -6620
rect 52335 -6740 52380 -6620
rect 52500 -6740 52555 -6620
rect 52675 -6740 52720 -6620
rect 52840 -6740 52885 -6620
rect 53005 -6740 53050 -6620
rect 53170 -6740 53225 -6620
rect 53345 -6740 53355 -6620
rect 47855 -6785 53355 -6740
rect 47855 -6905 47865 -6785
rect 47985 -6905 48030 -6785
rect 48150 -6905 48195 -6785
rect 48315 -6905 48360 -6785
rect 48480 -6905 48535 -6785
rect 48655 -6905 48700 -6785
rect 48820 -6905 48865 -6785
rect 48985 -6905 49030 -6785
rect 49150 -6905 49205 -6785
rect 49325 -6905 49370 -6785
rect 49490 -6905 49535 -6785
rect 49655 -6905 49700 -6785
rect 49820 -6905 49875 -6785
rect 49995 -6905 50040 -6785
rect 50160 -6905 50205 -6785
rect 50325 -6905 50370 -6785
rect 50490 -6905 50545 -6785
rect 50665 -6905 50710 -6785
rect 50830 -6905 50875 -6785
rect 50995 -6905 51040 -6785
rect 51160 -6905 51215 -6785
rect 51335 -6905 51380 -6785
rect 51500 -6905 51545 -6785
rect 51665 -6905 51710 -6785
rect 51830 -6905 51885 -6785
rect 52005 -6905 52050 -6785
rect 52170 -6905 52215 -6785
rect 52335 -6905 52380 -6785
rect 52500 -6905 52555 -6785
rect 52675 -6905 52720 -6785
rect 52840 -6905 52885 -6785
rect 53005 -6905 53050 -6785
rect 53170 -6905 53225 -6785
rect 53345 -6905 53355 -6785
rect 47855 -6950 53355 -6905
rect 47855 -7070 47865 -6950
rect 47985 -7070 48030 -6950
rect 48150 -7070 48195 -6950
rect 48315 -7070 48360 -6950
rect 48480 -7070 48535 -6950
rect 48655 -7070 48700 -6950
rect 48820 -7070 48865 -6950
rect 48985 -7070 49030 -6950
rect 49150 -7070 49205 -6950
rect 49325 -7070 49370 -6950
rect 49490 -7070 49535 -6950
rect 49655 -7070 49700 -6950
rect 49820 -7070 49875 -6950
rect 49995 -7070 50040 -6950
rect 50160 -7070 50205 -6950
rect 50325 -7070 50370 -6950
rect 50490 -7070 50545 -6950
rect 50665 -7070 50710 -6950
rect 50830 -7070 50875 -6950
rect 50995 -7070 51040 -6950
rect 51160 -7070 51215 -6950
rect 51335 -7070 51380 -6950
rect 51500 -7070 51545 -6950
rect 51665 -7070 51710 -6950
rect 51830 -7070 51885 -6950
rect 52005 -7070 52050 -6950
rect 52170 -7070 52215 -6950
rect 52335 -7070 52380 -6950
rect 52500 -7070 52555 -6950
rect 52675 -7070 52720 -6950
rect 52840 -7070 52885 -6950
rect 53005 -7070 53050 -6950
rect 53170 -7070 53225 -6950
rect 53345 -7070 53355 -6950
rect 47855 -7125 53355 -7070
rect 47855 -7245 47865 -7125
rect 47985 -7245 48030 -7125
rect 48150 -7245 48195 -7125
rect 48315 -7245 48360 -7125
rect 48480 -7245 48535 -7125
rect 48655 -7245 48700 -7125
rect 48820 -7245 48865 -7125
rect 48985 -7245 49030 -7125
rect 49150 -7245 49205 -7125
rect 49325 -7245 49370 -7125
rect 49490 -7245 49535 -7125
rect 49655 -7245 49700 -7125
rect 49820 -7245 49875 -7125
rect 49995 -7245 50040 -7125
rect 50160 -7245 50205 -7125
rect 50325 -7245 50370 -7125
rect 50490 -7245 50545 -7125
rect 50665 -7245 50710 -7125
rect 50830 -7245 50875 -7125
rect 50995 -7245 51040 -7125
rect 51160 -7245 51215 -7125
rect 51335 -7245 51380 -7125
rect 51500 -7245 51545 -7125
rect 51665 -7245 51710 -7125
rect 51830 -7245 51885 -7125
rect 52005 -7245 52050 -7125
rect 52170 -7245 52215 -7125
rect 52335 -7245 52380 -7125
rect 52500 -7245 52555 -7125
rect 52675 -7245 52720 -7125
rect 52840 -7245 52885 -7125
rect 53005 -7245 53050 -7125
rect 53170 -7245 53225 -7125
rect 53345 -7245 53355 -7125
rect 47855 -7290 53355 -7245
rect 47855 -7410 47865 -7290
rect 47985 -7410 48030 -7290
rect 48150 -7410 48195 -7290
rect 48315 -7410 48360 -7290
rect 48480 -7410 48535 -7290
rect 48655 -7410 48700 -7290
rect 48820 -7410 48865 -7290
rect 48985 -7410 49030 -7290
rect 49150 -7410 49205 -7290
rect 49325 -7410 49370 -7290
rect 49490 -7410 49535 -7290
rect 49655 -7410 49700 -7290
rect 49820 -7410 49875 -7290
rect 49995 -7410 50040 -7290
rect 50160 -7410 50205 -7290
rect 50325 -7410 50370 -7290
rect 50490 -7410 50545 -7290
rect 50665 -7410 50710 -7290
rect 50830 -7410 50875 -7290
rect 50995 -7410 51040 -7290
rect 51160 -7410 51215 -7290
rect 51335 -7410 51380 -7290
rect 51500 -7410 51545 -7290
rect 51665 -7410 51710 -7290
rect 51830 -7410 51885 -7290
rect 52005 -7410 52050 -7290
rect 52170 -7410 52215 -7290
rect 52335 -7410 52380 -7290
rect 52500 -7410 52555 -7290
rect 52675 -7410 52720 -7290
rect 52840 -7410 52885 -7290
rect 53005 -7410 53050 -7290
rect 53170 -7410 53225 -7290
rect 53345 -7410 53355 -7290
rect 47855 -7455 53355 -7410
rect 47855 -7575 47865 -7455
rect 47985 -7575 48030 -7455
rect 48150 -7575 48195 -7455
rect 48315 -7575 48360 -7455
rect 48480 -7575 48535 -7455
rect 48655 -7575 48700 -7455
rect 48820 -7575 48865 -7455
rect 48985 -7575 49030 -7455
rect 49150 -7575 49205 -7455
rect 49325 -7575 49370 -7455
rect 49490 -7575 49535 -7455
rect 49655 -7575 49700 -7455
rect 49820 -7575 49875 -7455
rect 49995 -7575 50040 -7455
rect 50160 -7575 50205 -7455
rect 50325 -7575 50370 -7455
rect 50490 -7575 50545 -7455
rect 50665 -7575 50710 -7455
rect 50830 -7575 50875 -7455
rect 50995 -7575 51040 -7455
rect 51160 -7575 51215 -7455
rect 51335 -7575 51380 -7455
rect 51500 -7575 51545 -7455
rect 51665 -7575 51710 -7455
rect 51830 -7575 51885 -7455
rect 52005 -7575 52050 -7455
rect 52170 -7575 52215 -7455
rect 52335 -7575 52380 -7455
rect 52500 -7575 52555 -7455
rect 52675 -7575 52720 -7455
rect 52840 -7575 52885 -7455
rect 53005 -7575 53050 -7455
rect 53170 -7575 53225 -7455
rect 53345 -7575 53355 -7455
rect 47855 -7620 53355 -7575
rect 47855 -7740 47865 -7620
rect 47985 -7740 48030 -7620
rect 48150 -7740 48195 -7620
rect 48315 -7740 48360 -7620
rect 48480 -7740 48535 -7620
rect 48655 -7740 48700 -7620
rect 48820 -7740 48865 -7620
rect 48985 -7740 49030 -7620
rect 49150 -7740 49205 -7620
rect 49325 -7740 49370 -7620
rect 49490 -7740 49535 -7620
rect 49655 -7740 49700 -7620
rect 49820 -7740 49875 -7620
rect 49995 -7740 50040 -7620
rect 50160 -7740 50205 -7620
rect 50325 -7740 50370 -7620
rect 50490 -7740 50545 -7620
rect 50665 -7740 50710 -7620
rect 50830 -7740 50875 -7620
rect 50995 -7740 51040 -7620
rect 51160 -7740 51215 -7620
rect 51335 -7740 51380 -7620
rect 51500 -7740 51545 -7620
rect 51665 -7740 51710 -7620
rect 51830 -7740 51885 -7620
rect 52005 -7740 52050 -7620
rect 52170 -7740 52215 -7620
rect 52335 -7740 52380 -7620
rect 52500 -7740 52555 -7620
rect 52675 -7740 52720 -7620
rect 52840 -7740 52885 -7620
rect 53005 -7740 53050 -7620
rect 53170 -7740 53225 -7620
rect 53345 -7740 53355 -7620
rect 47855 -7795 53355 -7740
rect 47855 -7915 47865 -7795
rect 47985 -7915 48030 -7795
rect 48150 -7915 48195 -7795
rect 48315 -7915 48360 -7795
rect 48480 -7915 48535 -7795
rect 48655 -7915 48700 -7795
rect 48820 -7915 48865 -7795
rect 48985 -7915 49030 -7795
rect 49150 -7915 49205 -7795
rect 49325 -7915 49370 -7795
rect 49490 -7915 49535 -7795
rect 49655 -7915 49700 -7795
rect 49820 -7915 49875 -7795
rect 49995 -7915 50040 -7795
rect 50160 -7915 50205 -7795
rect 50325 -7915 50370 -7795
rect 50490 -7915 50545 -7795
rect 50665 -7915 50710 -7795
rect 50830 -7915 50875 -7795
rect 50995 -7915 51040 -7795
rect 51160 -7915 51215 -7795
rect 51335 -7915 51380 -7795
rect 51500 -7915 51545 -7795
rect 51665 -7915 51710 -7795
rect 51830 -7915 51885 -7795
rect 52005 -7915 52050 -7795
rect 52170 -7915 52215 -7795
rect 52335 -7915 52380 -7795
rect 52500 -7915 52555 -7795
rect 52675 -7915 52720 -7795
rect 52840 -7915 52885 -7795
rect 53005 -7915 53050 -7795
rect 53170 -7915 53225 -7795
rect 53345 -7915 53355 -7795
rect 47855 -7960 53355 -7915
rect 47855 -8080 47865 -7960
rect 47985 -8080 48030 -7960
rect 48150 -8080 48195 -7960
rect 48315 -8080 48360 -7960
rect 48480 -8080 48535 -7960
rect 48655 -8080 48700 -7960
rect 48820 -8080 48865 -7960
rect 48985 -8080 49030 -7960
rect 49150 -8080 49205 -7960
rect 49325 -8080 49370 -7960
rect 49490 -8080 49535 -7960
rect 49655 -8080 49700 -7960
rect 49820 -8080 49875 -7960
rect 49995 -8080 50040 -7960
rect 50160 -8080 50205 -7960
rect 50325 -8080 50370 -7960
rect 50490 -8080 50545 -7960
rect 50665 -8080 50710 -7960
rect 50830 -8080 50875 -7960
rect 50995 -8080 51040 -7960
rect 51160 -8080 51215 -7960
rect 51335 -8080 51380 -7960
rect 51500 -8080 51545 -7960
rect 51665 -8080 51710 -7960
rect 51830 -8080 51885 -7960
rect 52005 -8080 52050 -7960
rect 52170 -8080 52215 -7960
rect 52335 -8080 52380 -7960
rect 52500 -8080 52555 -7960
rect 52675 -8080 52720 -7960
rect 52840 -8080 52885 -7960
rect 53005 -8080 53050 -7960
rect 53170 -8080 53225 -7960
rect 53345 -8080 53355 -7960
rect 47855 -8125 53355 -8080
rect 47855 -8245 47865 -8125
rect 47985 -8245 48030 -8125
rect 48150 -8245 48195 -8125
rect 48315 -8245 48360 -8125
rect 48480 -8245 48535 -8125
rect 48655 -8245 48700 -8125
rect 48820 -8245 48865 -8125
rect 48985 -8245 49030 -8125
rect 49150 -8245 49205 -8125
rect 49325 -8245 49370 -8125
rect 49490 -8245 49535 -8125
rect 49655 -8245 49700 -8125
rect 49820 -8245 49875 -8125
rect 49995 -8245 50040 -8125
rect 50160 -8245 50205 -8125
rect 50325 -8245 50370 -8125
rect 50490 -8245 50545 -8125
rect 50665 -8245 50710 -8125
rect 50830 -8245 50875 -8125
rect 50995 -8245 51040 -8125
rect 51160 -8245 51215 -8125
rect 51335 -8245 51380 -8125
rect 51500 -8245 51545 -8125
rect 51665 -8245 51710 -8125
rect 51830 -8245 51885 -8125
rect 52005 -8245 52050 -8125
rect 52170 -8245 52215 -8125
rect 52335 -8245 52380 -8125
rect 52500 -8245 52555 -8125
rect 52675 -8245 52720 -8125
rect 52840 -8245 52885 -8125
rect 53005 -8245 53050 -8125
rect 53170 -8245 53225 -8125
rect 53345 -8245 53355 -8125
rect 47855 -8290 53355 -8245
rect 47855 -8410 47865 -8290
rect 47985 -8410 48030 -8290
rect 48150 -8410 48195 -8290
rect 48315 -8410 48360 -8290
rect 48480 -8410 48535 -8290
rect 48655 -8410 48700 -8290
rect 48820 -8410 48865 -8290
rect 48985 -8410 49030 -8290
rect 49150 -8410 49205 -8290
rect 49325 -8410 49370 -8290
rect 49490 -8410 49535 -8290
rect 49655 -8410 49700 -8290
rect 49820 -8410 49875 -8290
rect 49995 -8410 50040 -8290
rect 50160 -8410 50205 -8290
rect 50325 -8410 50370 -8290
rect 50490 -8410 50545 -8290
rect 50665 -8410 50710 -8290
rect 50830 -8410 50875 -8290
rect 50995 -8410 51040 -8290
rect 51160 -8410 51215 -8290
rect 51335 -8410 51380 -8290
rect 51500 -8410 51545 -8290
rect 51665 -8410 51710 -8290
rect 51830 -8410 51885 -8290
rect 52005 -8410 52050 -8290
rect 52170 -8410 52215 -8290
rect 52335 -8410 52380 -8290
rect 52500 -8410 52555 -8290
rect 52675 -8410 52720 -8290
rect 52840 -8410 52885 -8290
rect 53005 -8410 53050 -8290
rect 53170 -8410 53225 -8290
rect 53345 -8410 53355 -8290
rect 47855 -8465 53355 -8410
rect 47855 -8585 47865 -8465
rect 47985 -8585 48030 -8465
rect 48150 -8585 48195 -8465
rect 48315 -8585 48360 -8465
rect 48480 -8585 48535 -8465
rect 48655 -8585 48700 -8465
rect 48820 -8585 48865 -8465
rect 48985 -8585 49030 -8465
rect 49150 -8585 49205 -8465
rect 49325 -8585 49370 -8465
rect 49490 -8585 49535 -8465
rect 49655 -8585 49700 -8465
rect 49820 -8585 49875 -8465
rect 49995 -8585 50040 -8465
rect 50160 -8585 50205 -8465
rect 50325 -8585 50370 -8465
rect 50490 -8585 50545 -8465
rect 50665 -8585 50710 -8465
rect 50830 -8585 50875 -8465
rect 50995 -8585 51040 -8465
rect 51160 -8585 51215 -8465
rect 51335 -8585 51380 -8465
rect 51500 -8585 51545 -8465
rect 51665 -8585 51710 -8465
rect 51830 -8585 51885 -8465
rect 52005 -8585 52050 -8465
rect 52170 -8585 52215 -8465
rect 52335 -8585 52380 -8465
rect 52500 -8585 52555 -8465
rect 52675 -8585 52720 -8465
rect 52840 -8585 52885 -8465
rect 53005 -8585 53050 -8465
rect 53170 -8585 53225 -8465
rect 53345 -8585 53355 -8465
rect 47855 -8630 53355 -8585
rect 47855 -8750 47865 -8630
rect 47985 -8750 48030 -8630
rect 48150 -8750 48195 -8630
rect 48315 -8750 48360 -8630
rect 48480 -8750 48535 -8630
rect 48655 -8750 48700 -8630
rect 48820 -8750 48865 -8630
rect 48985 -8750 49030 -8630
rect 49150 -8750 49205 -8630
rect 49325 -8750 49370 -8630
rect 49490 -8750 49535 -8630
rect 49655 -8750 49700 -8630
rect 49820 -8750 49875 -8630
rect 49995 -8750 50040 -8630
rect 50160 -8750 50205 -8630
rect 50325 -8750 50370 -8630
rect 50490 -8750 50545 -8630
rect 50665 -8750 50710 -8630
rect 50830 -8750 50875 -8630
rect 50995 -8750 51040 -8630
rect 51160 -8750 51215 -8630
rect 51335 -8750 51380 -8630
rect 51500 -8750 51545 -8630
rect 51665 -8750 51710 -8630
rect 51830 -8750 51885 -8630
rect 52005 -8750 52050 -8630
rect 52170 -8750 52215 -8630
rect 52335 -8750 52380 -8630
rect 52500 -8750 52555 -8630
rect 52675 -8750 52720 -8630
rect 52840 -8750 52885 -8630
rect 53005 -8750 53050 -8630
rect 53170 -8750 53225 -8630
rect 53345 -8750 53355 -8630
rect 47855 -8795 53355 -8750
rect 47855 -8915 47865 -8795
rect 47985 -8915 48030 -8795
rect 48150 -8915 48195 -8795
rect 48315 -8915 48360 -8795
rect 48480 -8915 48535 -8795
rect 48655 -8915 48700 -8795
rect 48820 -8915 48865 -8795
rect 48985 -8915 49030 -8795
rect 49150 -8915 49205 -8795
rect 49325 -8915 49370 -8795
rect 49490 -8915 49535 -8795
rect 49655 -8915 49700 -8795
rect 49820 -8915 49875 -8795
rect 49995 -8915 50040 -8795
rect 50160 -8915 50205 -8795
rect 50325 -8915 50370 -8795
rect 50490 -8915 50545 -8795
rect 50665 -8915 50710 -8795
rect 50830 -8915 50875 -8795
rect 50995 -8915 51040 -8795
rect 51160 -8915 51215 -8795
rect 51335 -8915 51380 -8795
rect 51500 -8915 51545 -8795
rect 51665 -8915 51710 -8795
rect 51830 -8915 51885 -8795
rect 52005 -8915 52050 -8795
rect 52170 -8915 52215 -8795
rect 52335 -8915 52380 -8795
rect 52500 -8915 52555 -8795
rect 52675 -8915 52720 -8795
rect 52840 -8915 52885 -8795
rect 53005 -8915 53050 -8795
rect 53170 -8915 53225 -8795
rect 53345 -8915 53355 -8795
rect 47855 -8960 53355 -8915
rect 47855 -9080 47865 -8960
rect 47985 -9080 48030 -8960
rect 48150 -9080 48195 -8960
rect 48315 -9080 48360 -8960
rect 48480 -9080 48535 -8960
rect 48655 -9080 48700 -8960
rect 48820 -9080 48865 -8960
rect 48985 -9080 49030 -8960
rect 49150 -9080 49205 -8960
rect 49325 -9080 49370 -8960
rect 49490 -9080 49535 -8960
rect 49655 -9080 49700 -8960
rect 49820 -9080 49875 -8960
rect 49995 -9080 50040 -8960
rect 50160 -9080 50205 -8960
rect 50325 -9080 50370 -8960
rect 50490 -9080 50545 -8960
rect 50665 -9080 50710 -8960
rect 50830 -9080 50875 -8960
rect 50995 -9080 51040 -8960
rect 51160 -9080 51215 -8960
rect 51335 -9080 51380 -8960
rect 51500 -9080 51545 -8960
rect 51665 -9080 51710 -8960
rect 51830 -9080 51885 -8960
rect 52005 -9080 52050 -8960
rect 52170 -9080 52215 -8960
rect 52335 -9080 52380 -8960
rect 52500 -9080 52555 -8960
rect 52675 -9080 52720 -8960
rect 52840 -9080 52885 -8960
rect 53005 -9080 53050 -8960
rect 53170 -9080 53225 -8960
rect 53345 -9080 53355 -8960
rect 47855 -9135 53355 -9080
rect 47855 -9255 47865 -9135
rect 47985 -9255 48030 -9135
rect 48150 -9255 48195 -9135
rect 48315 -9255 48360 -9135
rect 48480 -9255 48535 -9135
rect 48655 -9255 48700 -9135
rect 48820 -9255 48865 -9135
rect 48985 -9255 49030 -9135
rect 49150 -9255 49205 -9135
rect 49325 -9255 49370 -9135
rect 49490 -9255 49535 -9135
rect 49655 -9255 49700 -9135
rect 49820 -9255 49875 -9135
rect 49995 -9255 50040 -9135
rect 50160 -9255 50205 -9135
rect 50325 -9255 50370 -9135
rect 50490 -9255 50545 -9135
rect 50665 -9255 50710 -9135
rect 50830 -9255 50875 -9135
rect 50995 -9255 51040 -9135
rect 51160 -9255 51215 -9135
rect 51335 -9255 51380 -9135
rect 51500 -9255 51545 -9135
rect 51665 -9255 51710 -9135
rect 51830 -9255 51885 -9135
rect 52005 -9255 52050 -9135
rect 52170 -9255 52215 -9135
rect 52335 -9255 52380 -9135
rect 52500 -9255 52555 -9135
rect 52675 -9255 52720 -9135
rect 52840 -9255 52885 -9135
rect 53005 -9255 53050 -9135
rect 53170 -9255 53225 -9135
rect 53345 -9255 53355 -9135
rect 47855 -9300 53355 -9255
rect 47855 -9420 47865 -9300
rect 47985 -9420 48030 -9300
rect 48150 -9420 48195 -9300
rect 48315 -9420 48360 -9300
rect 48480 -9420 48535 -9300
rect 48655 -9420 48700 -9300
rect 48820 -9420 48865 -9300
rect 48985 -9420 49030 -9300
rect 49150 -9420 49205 -9300
rect 49325 -9420 49370 -9300
rect 49490 -9420 49535 -9300
rect 49655 -9420 49700 -9300
rect 49820 -9420 49875 -9300
rect 49995 -9420 50040 -9300
rect 50160 -9420 50205 -9300
rect 50325 -9420 50370 -9300
rect 50490 -9420 50545 -9300
rect 50665 -9420 50710 -9300
rect 50830 -9420 50875 -9300
rect 50995 -9420 51040 -9300
rect 51160 -9420 51215 -9300
rect 51335 -9420 51380 -9300
rect 51500 -9420 51545 -9300
rect 51665 -9420 51710 -9300
rect 51830 -9420 51885 -9300
rect 52005 -9420 52050 -9300
rect 52170 -9420 52215 -9300
rect 52335 -9420 52380 -9300
rect 52500 -9420 52555 -9300
rect 52675 -9420 52720 -9300
rect 52840 -9420 52885 -9300
rect 53005 -9420 53050 -9300
rect 53170 -9420 53225 -9300
rect 53345 -9420 53355 -9300
rect 47855 -9465 53355 -9420
rect 47855 -9585 47865 -9465
rect 47985 -9585 48030 -9465
rect 48150 -9585 48195 -9465
rect 48315 -9585 48360 -9465
rect 48480 -9585 48535 -9465
rect 48655 -9585 48700 -9465
rect 48820 -9585 48865 -9465
rect 48985 -9585 49030 -9465
rect 49150 -9585 49205 -9465
rect 49325 -9585 49370 -9465
rect 49490 -9585 49535 -9465
rect 49655 -9585 49700 -9465
rect 49820 -9585 49875 -9465
rect 49995 -9585 50040 -9465
rect 50160 -9585 50205 -9465
rect 50325 -9585 50370 -9465
rect 50490 -9585 50545 -9465
rect 50665 -9585 50710 -9465
rect 50830 -9585 50875 -9465
rect 50995 -9585 51040 -9465
rect 51160 -9585 51215 -9465
rect 51335 -9585 51380 -9465
rect 51500 -9585 51545 -9465
rect 51665 -9585 51710 -9465
rect 51830 -9585 51885 -9465
rect 52005 -9585 52050 -9465
rect 52170 -9585 52215 -9465
rect 52335 -9585 52380 -9465
rect 52500 -9585 52555 -9465
rect 52675 -9585 52720 -9465
rect 52840 -9585 52885 -9465
rect 53005 -9585 53050 -9465
rect 53170 -9585 53225 -9465
rect 53345 -9585 53355 -9465
rect 47855 -9630 53355 -9585
rect 47855 -9750 47865 -9630
rect 47985 -9750 48030 -9630
rect 48150 -9750 48195 -9630
rect 48315 -9750 48360 -9630
rect 48480 -9750 48535 -9630
rect 48655 -9750 48700 -9630
rect 48820 -9750 48865 -9630
rect 48985 -9750 49030 -9630
rect 49150 -9750 49205 -9630
rect 49325 -9750 49370 -9630
rect 49490 -9750 49535 -9630
rect 49655 -9750 49700 -9630
rect 49820 -9750 49875 -9630
rect 49995 -9750 50040 -9630
rect 50160 -9750 50205 -9630
rect 50325 -9750 50370 -9630
rect 50490 -9750 50545 -9630
rect 50665 -9750 50710 -9630
rect 50830 -9750 50875 -9630
rect 50995 -9750 51040 -9630
rect 51160 -9750 51215 -9630
rect 51335 -9750 51380 -9630
rect 51500 -9750 51545 -9630
rect 51665 -9750 51710 -9630
rect 51830 -9750 51885 -9630
rect 52005 -9750 52050 -9630
rect 52170 -9750 52215 -9630
rect 52335 -9750 52380 -9630
rect 52500 -9750 52555 -9630
rect 52675 -9750 52720 -9630
rect 52840 -9750 52885 -9630
rect 53005 -9750 53050 -9630
rect 53170 -9750 53225 -9630
rect 53345 -9750 53355 -9630
rect 47855 -9760 53355 -9750
rect 30785 -10050 36285 -10040
rect 30785 -10170 30795 -10050
rect 30915 -10170 30970 -10050
rect 31090 -10170 31135 -10050
rect 31255 -10170 31300 -10050
rect 31420 -10170 31465 -10050
rect 31585 -10170 31640 -10050
rect 31760 -10170 31805 -10050
rect 31925 -10170 31970 -10050
rect 32090 -10170 32135 -10050
rect 32255 -10170 32310 -10050
rect 32430 -10170 32475 -10050
rect 32595 -10170 32640 -10050
rect 32760 -10170 32805 -10050
rect 32925 -10170 32980 -10050
rect 33100 -10170 33145 -10050
rect 33265 -10170 33310 -10050
rect 33430 -10170 33475 -10050
rect 33595 -10170 33650 -10050
rect 33770 -10170 33815 -10050
rect 33935 -10170 33980 -10050
rect 34100 -10170 34145 -10050
rect 34265 -10170 34320 -10050
rect 34440 -10170 34485 -10050
rect 34605 -10170 34650 -10050
rect 34770 -10170 34815 -10050
rect 34935 -10170 34990 -10050
rect 35110 -10170 35155 -10050
rect 35275 -10170 35320 -10050
rect 35440 -10170 35485 -10050
rect 35605 -10170 35660 -10050
rect 35780 -10170 35825 -10050
rect 35945 -10170 35990 -10050
rect 36110 -10170 36155 -10050
rect 36275 -10170 36285 -10050
rect 30785 -10215 36285 -10170
rect 30785 -10335 30795 -10215
rect 30915 -10335 30970 -10215
rect 31090 -10335 31135 -10215
rect 31255 -10335 31300 -10215
rect 31420 -10335 31465 -10215
rect 31585 -10335 31640 -10215
rect 31760 -10335 31805 -10215
rect 31925 -10335 31970 -10215
rect 32090 -10335 32135 -10215
rect 32255 -10335 32310 -10215
rect 32430 -10335 32475 -10215
rect 32595 -10335 32640 -10215
rect 32760 -10335 32805 -10215
rect 32925 -10335 32980 -10215
rect 33100 -10335 33145 -10215
rect 33265 -10335 33310 -10215
rect 33430 -10335 33475 -10215
rect 33595 -10335 33650 -10215
rect 33770 -10335 33815 -10215
rect 33935 -10335 33980 -10215
rect 34100 -10335 34145 -10215
rect 34265 -10335 34320 -10215
rect 34440 -10335 34485 -10215
rect 34605 -10335 34650 -10215
rect 34770 -10335 34815 -10215
rect 34935 -10335 34990 -10215
rect 35110 -10335 35155 -10215
rect 35275 -10335 35320 -10215
rect 35440 -10335 35485 -10215
rect 35605 -10335 35660 -10215
rect 35780 -10335 35825 -10215
rect 35945 -10335 35990 -10215
rect 36110 -10335 36155 -10215
rect 36275 -10335 36285 -10215
rect 30785 -10380 36285 -10335
rect 30785 -10500 30795 -10380
rect 30915 -10500 30970 -10380
rect 31090 -10500 31135 -10380
rect 31255 -10500 31300 -10380
rect 31420 -10500 31465 -10380
rect 31585 -10500 31640 -10380
rect 31760 -10500 31805 -10380
rect 31925 -10500 31970 -10380
rect 32090 -10500 32135 -10380
rect 32255 -10500 32310 -10380
rect 32430 -10500 32475 -10380
rect 32595 -10500 32640 -10380
rect 32760 -10500 32805 -10380
rect 32925 -10500 32980 -10380
rect 33100 -10500 33145 -10380
rect 33265 -10500 33310 -10380
rect 33430 -10500 33475 -10380
rect 33595 -10500 33650 -10380
rect 33770 -10500 33815 -10380
rect 33935 -10500 33980 -10380
rect 34100 -10500 34145 -10380
rect 34265 -10500 34320 -10380
rect 34440 -10500 34485 -10380
rect 34605 -10500 34650 -10380
rect 34770 -10500 34815 -10380
rect 34935 -10500 34990 -10380
rect 35110 -10500 35155 -10380
rect 35275 -10500 35320 -10380
rect 35440 -10500 35485 -10380
rect 35605 -10500 35660 -10380
rect 35780 -10500 35825 -10380
rect 35945 -10500 35990 -10380
rect 36110 -10500 36155 -10380
rect 36275 -10500 36285 -10380
rect 30785 -10545 36285 -10500
rect 30785 -10665 30795 -10545
rect 30915 -10665 30970 -10545
rect 31090 -10665 31135 -10545
rect 31255 -10665 31300 -10545
rect 31420 -10665 31465 -10545
rect 31585 -10665 31640 -10545
rect 31760 -10665 31805 -10545
rect 31925 -10665 31970 -10545
rect 32090 -10665 32135 -10545
rect 32255 -10665 32310 -10545
rect 32430 -10665 32475 -10545
rect 32595 -10665 32640 -10545
rect 32760 -10665 32805 -10545
rect 32925 -10665 32980 -10545
rect 33100 -10665 33145 -10545
rect 33265 -10665 33310 -10545
rect 33430 -10665 33475 -10545
rect 33595 -10665 33650 -10545
rect 33770 -10665 33815 -10545
rect 33935 -10665 33980 -10545
rect 34100 -10665 34145 -10545
rect 34265 -10665 34320 -10545
rect 34440 -10665 34485 -10545
rect 34605 -10665 34650 -10545
rect 34770 -10665 34815 -10545
rect 34935 -10665 34990 -10545
rect 35110 -10665 35155 -10545
rect 35275 -10665 35320 -10545
rect 35440 -10665 35485 -10545
rect 35605 -10665 35660 -10545
rect 35780 -10665 35825 -10545
rect 35945 -10665 35990 -10545
rect 36110 -10665 36155 -10545
rect 36275 -10665 36285 -10545
rect 30785 -10720 36285 -10665
rect 30785 -10840 30795 -10720
rect 30915 -10840 30970 -10720
rect 31090 -10840 31135 -10720
rect 31255 -10840 31300 -10720
rect 31420 -10840 31465 -10720
rect 31585 -10840 31640 -10720
rect 31760 -10840 31805 -10720
rect 31925 -10840 31970 -10720
rect 32090 -10840 32135 -10720
rect 32255 -10840 32310 -10720
rect 32430 -10840 32475 -10720
rect 32595 -10840 32640 -10720
rect 32760 -10840 32805 -10720
rect 32925 -10840 32980 -10720
rect 33100 -10840 33145 -10720
rect 33265 -10840 33310 -10720
rect 33430 -10840 33475 -10720
rect 33595 -10840 33650 -10720
rect 33770 -10840 33815 -10720
rect 33935 -10840 33980 -10720
rect 34100 -10840 34145 -10720
rect 34265 -10840 34320 -10720
rect 34440 -10840 34485 -10720
rect 34605 -10840 34650 -10720
rect 34770 -10840 34815 -10720
rect 34935 -10840 34990 -10720
rect 35110 -10840 35155 -10720
rect 35275 -10840 35320 -10720
rect 35440 -10840 35485 -10720
rect 35605 -10840 35660 -10720
rect 35780 -10840 35825 -10720
rect 35945 -10840 35990 -10720
rect 36110 -10840 36155 -10720
rect 36275 -10840 36285 -10720
rect 30785 -10885 36285 -10840
rect 30785 -11005 30795 -10885
rect 30915 -11005 30970 -10885
rect 31090 -11005 31135 -10885
rect 31255 -11005 31300 -10885
rect 31420 -11005 31465 -10885
rect 31585 -11005 31640 -10885
rect 31760 -11005 31805 -10885
rect 31925 -11005 31970 -10885
rect 32090 -11005 32135 -10885
rect 32255 -11005 32310 -10885
rect 32430 -11005 32475 -10885
rect 32595 -11005 32640 -10885
rect 32760 -11005 32805 -10885
rect 32925 -11005 32980 -10885
rect 33100 -11005 33145 -10885
rect 33265 -11005 33310 -10885
rect 33430 -11005 33475 -10885
rect 33595 -11005 33650 -10885
rect 33770 -11005 33815 -10885
rect 33935 -11005 33980 -10885
rect 34100 -11005 34145 -10885
rect 34265 -11005 34320 -10885
rect 34440 -11005 34485 -10885
rect 34605 -11005 34650 -10885
rect 34770 -11005 34815 -10885
rect 34935 -11005 34990 -10885
rect 35110 -11005 35155 -10885
rect 35275 -11005 35320 -10885
rect 35440 -11005 35485 -10885
rect 35605 -11005 35660 -10885
rect 35780 -11005 35825 -10885
rect 35945 -11005 35990 -10885
rect 36110 -11005 36155 -10885
rect 36275 -11005 36285 -10885
rect 30785 -11050 36285 -11005
rect 30785 -11170 30795 -11050
rect 30915 -11170 30970 -11050
rect 31090 -11170 31135 -11050
rect 31255 -11170 31300 -11050
rect 31420 -11170 31465 -11050
rect 31585 -11170 31640 -11050
rect 31760 -11170 31805 -11050
rect 31925 -11170 31970 -11050
rect 32090 -11170 32135 -11050
rect 32255 -11170 32310 -11050
rect 32430 -11170 32475 -11050
rect 32595 -11170 32640 -11050
rect 32760 -11170 32805 -11050
rect 32925 -11170 32980 -11050
rect 33100 -11170 33145 -11050
rect 33265 -11170 33310 -11050
rect 33430 -11170 33475 -11050
rect 33595 -11170 33650 -11050
rect 33770 -11170 33815 -11050
rect 33935 -11170 33980 -11050
rect 34100 -11170 34145 -11050
rect 34265 -11170 34320 -11050
rect 34440 -11170 34485 -11050
rect 34605 -11170 34650 -11050
rect 34770 -11170 34815 -11050
rect 34935 -11170 34990 -11050
rect 35110 -11170 35155 -11050
rect 35275 -11170 35320 -11050
rect 35440 -11170 35485 -11050
rect 35605 -11170 35660 -11050
rect 35780 -11170 35825 -11050
rect 35945 -11170 35990 -11050
rect 36110 -11170 36155 -11050
rect 36275 -11170 36285 -11050
rect 30785 -11215 36285 -11170
rect 30785 -11335 30795 -11215
rect 30915 -11335 30970 -11215
rect 31090 -11335 31135 -11215
rect 31255 -11335 31300 -11215
rect 31420 -11335 31465 -11215
rect 31585 -11335 31640 -11215
rect 31760 -11335 31805 -11215
rect 31925 -11335 31970 -11215
rect 32090 -11335 32135 -11215
rect 32255 -11335 32310 -11215
rect 32430 -11335 32475 -11215
rect 32595 -11335 32640 -11215
rect 32760 -11335 32805 -11215
rect 32925 -11335 32980 -11215
rect 33100 -11335 33145 -11215
rect 33265 -11335 33310 -11215
rect 33430 -11335 33475 -11215
rect 33595 -11335 33650 -11215
rect 33770 -11335 33815 -11215
rect 33935 -11335 33980 -11215
rect 34100 -11335 34145 -11215
rect 34265 -11335 34320 -11215
rect 34440 -11335 34485 -11215
rect 34605 -11335 34650 -11215
rect 34770 -11335 34815 -11215
rect 34935 -11335 34990 -11215
rect 35110 -11335 35155 -11215
rect 35275 -11335 35320 -11215
rect 35440 -11335 35485 -11215
rect 35605 -11335 35660 -11215
rect 35780 -11335 35825 -11215
rect 35945 -11335 35990 -11215
rect 36110 -11335 36155 -11215
rect 36275 -11335 36285 -11215
rect 30785 -11390 36285 -11335
rect 30785 -11510 30795 -11390
rect 30915 -11510 30970 -11390
rect 31090 -11510 31135 -11390
rect 31255 -11510 31300 -11390
rect 31420 -11510 31465 -11390
rect 31585 -11510 31640 -11390
rect 31760 -11510 31805 -11390
rect 31925 -11510 31970 -11390
rect 32090 -11510 32135 -11390
rect 32255 -11510 32310 -11390
rect 32430 -11510 32475 -11390
rect 32595 -11510 32640 -11390
rect 32760 -11510 32805 -11390
rect 32925 -11510 32980 -11390
rect 33100 -11510 33145 -11390
rect 33265 -11510 33310 -11390
rect 33430 -11510 33475 -11390
rect 33595 -11510 33650 -11390
rect 33770 -11510 33815 -11390
rect 33935 -11510 33980 -11390
rect 34100 -11510 34145 -11390
rect 34265 -11510 34320 -11390
rect 34440 -11510 34485 -11390
rect 34605 -11510 34650 -11390
rect 34770 -11510 34815 -11390
rect 34935 -11510 34990 -11390
rect 35110 -11510 35155 -11390
rect 35275 -11510 35320 -11390
rect 35440 -11510 35485 -11390
rect 35605 -11510 35660 -11390
rect 35780 -11510 35825 -11390
rect 35945 -11510 35990 -11390
rect 36110 -11510 36155 -11390
rect 36275 -11510 36285 -11390
rect 30785 -11555 36285 -11510
rect 30785 -11675 30795 -11555
rect 30915 -11675 30970 -11555
rect 31090 -11675 31135 -11555
rect 31255 -11675 31300 -11555
rect 31420 -11675 31465 -11555
rect 31585 -11675 31640 -11555
rect 31760 -11675 31805 -11555
rect 31925 -11675 31970 -11555
rect 32090 -11675 32135 -11555
rect 32255 -11675 32310 -11555
rect 32430 -11675 32475 -11555
rect 32595 -11675 32640 -11555
rect 32760 -11675 32805 -11555
rect 32925 -11675 32980 -11555
rect 33100 -11675 33145 -11555
rect 33265 -11675 33310 -11555
rect 33430 -11675 33475 -11555
rect 33595 -11675 33650 -11555
rect 33770 -11675 33815 -11555
rect 33935 -11675 33980 -11555
rect 34100 -11675 34145 -11555
rect 34265 -11675 34320 -11555
rect 34440 -11675 34485 -11555
rect 34605 -11675 34650 -11555
rect 34770 -11675 34815 -11555
rect 34935 -11675 34990 -11555
rect 35110 -11675 35155 -11555
rect 35275 -11675 35320 -11555
rect 35440 -11675 35485 -11555
rect 35605 -11675 35660 -11555
rect 35780 -11675 35825 -11555
rect 35945 -11675 35990 -11555
rect 36110 -11675 36155 -11555
rect 36275 -11675 36285 -11555
rect 30785 -11720 36285 -11675
rect 30785 -11840 30795 -11720
rect 30915 -11840 30970 -11720
rect 31090 -11840 31135 -11720
rect 31255 -11840 31300 -11720
rect 31420 -11840 31465 -11720
rect 31585 -11840 31640 -11720
rect 31760 -11840 31805 -11720
rect 31925 -11840 31970 -11720
rect 32090 -11840 32135 -11720
rect 32255 -11840 32310 -11720
rect 32430 -11840 32475 -11720
rect 32595 -11840 32640 -11720
rect 32760 -11840 32805 -11720
rect 32925 -11840 32980 -11720
rect 33100 -11840 33145 -11720
rect 33265 -11840 33310 -11720
rect 33430 -11840 33475 -11720
rect 33595 -11840 33650 -11720
rect 33770 -11840 33815 -11720
rect 33935 -11840 33980 -11720
rect 34100 -11840 34145 -11720
rect 34265 -11840 34320 -11720
rect 34440 -11840 34485 -11720
rect 34605 -11840 34650 -11720
rect 34770 -11840 34815 -11720
rect 34935 -11840 34990 -11720
rect 35110 -11840 35155 -11720
rect 35275 -11840 35320 -11720
rect 35440 -11840 35485 -11720
rect 35605 -11840 35660 -11720
rect 35780 -11840 35825 -11720
rect 35945 -11840 35990 -11720
rect 36110 -11840 36155 -11720
rect 36275 -11840 36285 -11720
rect 30785 -11885 36285 -11840
rect 30785 -12005 30795 -11885
rect 30915 -12005 30970 -11885
rect 31090 -12005 31135 -11885
rect 31255 -12005 31300 -11885
rect 31420 -12005 31465 -11885
rect 31585 -12005 31640 -11885
rect 31760 -12005 31805 -11885
rect 31925 -12005 31970 -11885
rect 32090 -12005 32135 -11885
rect 32255 -12005 32310 -11885
rect 32430 -12005 32475 -11885
rect 32595 -12005 32640 -11885
rect 32760 -12005 32805 -11885
rect 32925 -12005 32980 -11885
rect 33100 -12005 33145 -11885
rect 33265 -12005 33310 -11885
rect 33430 -12005 33475 -11885
rect 33595 -12005 33650 -11885
rect 33770 -12005 33815 -11885
rect 33935 -12005 33980 -11885
rect 34100 -12005 34145 -11885
rect 34265 -12005 34320 -11885
rect 34440 -12005 34485 -11885
rect 34605 -12005 34650 -11885
rect 34770 -12005 34815 -11885
rect 34935 -12005 34990 -11885
rect 35110 -12005 35155 -11885
rect 35275 -12005 35320 -11885
rect 35440 -12005 35485 -11885
rect 35605 -12005 35660 -11885
rect 35780 -12005 35825 -11885
rect 35945 -12005 35990 -11885
rect 36110 -12005 36155 -11885
rect 36275 -12005 36285 -11885
rect 30785 -12060 36285 -12005
rect 30785 -12180 30795 -12060
rect 30915 -12180 30970 -12060
rect 31090 -12180 31135 -12060
rect 31255 -12180 31300 -12060
rect 31420 -12180 31465 -12060
rect 31585 -12180 31640 -12060
rect 31760 -12180 31805 -12060
rect 31925 -12180 31970 -12060
rect 32090 -12180 32135 -12060
rect 32255 -12180 32310 -12060
rect 32430 -12180 32475 -12060
rect 32595 -12180 32640 -12060
rect 32760 -12180 32805 -12060
rect 32925 -12180 32980 -12060
rect 33100 -12180 33145 -12060
rect 33265 -12180 33310 -12060
rect 33430 -12180 33475 -12060
rect 33595 -12180 33650 -12060
rect 33770 -12180 33815 -12060
rect 33935 -12180 33980 -12060
rect 34100 -12180 34145 -12060
rect 34265 -12180 34320 -12060
rect 34440 -12180 34485 -12060
rect 34605 -12180 34650 -12060
rect 34770 -12180 34815 -12060
rect 34935 -12180 34990 -12060
rect 35110 -12180 35155 -12060
rect 35275 -12180 35320 -12060
rect 35440 -12180 35485 -12060
rect 35605 -12180 35660 -12060
rect 35780 -12180 35825 -12060
rect 35945 -12180 35990 -12060
rect 36110 -12180 36155 -12060
rect 36275 -12180 36285 -12060
rect 30785 -12225 36285 -12180
rect 30785 -12345 30795 -12225
rect 30915 -12345 30970 -12225
rect 31090 -12345 31135 -12225
rect 31255 -12345 31300 -12225
rect 31420 -12345 31465 -12225
rect 31585 -12345 31640 -12225
rect 31760 -12345 31805 -12225
rect 31925 -12345 31970 -12225
rect 32090 -12345 32135 -12225
rect 32255 -12345 32310 -12225
rect 32430 -12345 32475 -12225
rect 32595 -12345 32640 -12225
rect 32760 -12345 32805 -12225
rect 32925 -12345 32980 -12225
rect 33100 -12345 33145 -12225
rect 33265 -12345 33310 -12225
rect 33430 -12345 33475 -12225
rect 33595 -12345 33650 -12225
rect 33770 -12345 33815 -12225
rect 33935 -12345 33980 -12225
rect 34100 -12345 34145 -12225
rect 34265 -12345 34320 -12225
rect 34440 -12345 34485 -12225
rect 34605 -12345 34650 -12225
rect 34770 -12345 34815 -12225
rect 34935 -12345 34990 -12225
rect 35110 -12345 35155 -12225
rect 35275 -12345 35320 -12225
rect 35440 -12345 35485 -12225
rect 35605 -12345 35660 -12225
rect 35780 -12345 35825 -12225
rect 35945 -12345 35990 -12225
rect 36110 -12345 36155 -12225
rect 36275 -12345 36285 -12225
rect 30785 -12390 36285 -12345
rect 30785 -12510 30795 -12390
rect 30915 -12510 30970 -12390
rect 31090 -12510 31135 -12390
rect 31255 -12510 31300 -12390
rect 31420 -12510 31465 -12390
rect 31585 -12510 31640 -12390
rect 31760 -12510 31805 -12390
rect 31925 -12510 31970 -12390
rect 32090 -12510 32135 -12390
rect 32255 -12510 32310 -12390
rect 32430 -12510 32475 -12390
rect 32595 -12510 32640 -12390
rect 32760 -12510 32805 -12390
rect 32925 -12510 32980 -12390
rect 33100 -12510 33145 -12390
rect 33265 -12510 33310 -12390
rect 33430 -12510 33475 -12390
rect 33595 -12510 33650 -12390
rect 33770 -12510 33815 -12390
rect 33935 -12510 33980 -12390
rect 34100 -12510 34145 -12390
rect 34265 -12510 34320 -12390
rect 34440 -12510 34485 -12390
rect 34605 -12510 34650 -12390
rect 34770 -12510 34815 -12390
rect 34935 -12510 34990 -12390
rect 35110 -12510 35155 -12390
rect 35275 -12510 35320 -12390
rect 35440 -12510 35485 -12390
rect 35605 -12510 35660 -12390
rect 35780 -12510 35825 -12390
rect 35945 -12510 35990 -12390
rect 36110 -12510 36155 -12390
rect 36275 -12510 36285 -12390
rect 30785 -12555 36285 -12510
rect 30785 -12675 30795 -12555
rect 30915 -12675 30970 -12555
rect 31090 -12675 31135 -12555
rect 31255 -12675 31300 -12555
rect 31420 -12675 31465 -12555
rect 31585 -12675 31640 -12555
rect 31760 -12675 31805 -12555
rect 31925 -12675 31970 -12555
rect 32090 -12675 32135 -12555
rect 32255 -12675 32310 -12555
rect 32430 -12675 32475 -12555
rect 32595 -12675 32640 -12555
rect 32760 -12675 32805 -12555
rect 32925 -12675 32980 -12555
rect 33100 -12675 33145 -12555
rect 33265 -12675 33310 -12555
rect 33430 -12675 33475 -12555
rect 33595 -12675 33650 -12555
rect 33770 -12675 33815 -12555
rect 33935 -12675 33980 -12555
rect 34100 -12675 34145 -12555
rect 34265 -12675 34320 -12555
rect 34440 -12675 34485 -12555
rect 34605 -12675 34650 -12555
rect 34770 -12675 34815 -12555
rect 34935 -12675 34990 -12555
rect 35110 -12675 35155 -12555
rect 35275 -12675 35320 -12555
rect 35440 -12675 35485 -12555
rect 35605 -12675 35660 -12555
rect 35780 -12675 35825 -12555
rect 35945 -12675 35990 -12555
rect 36110 -12675 36155 -12555
rect 36275 -12675 36285 -12555
rect 30785 -12730 36285 -12675
rect 30785 -12850 30795 -12730
rect 30915 -12850 30970 -12730
rect 31090 -12850 31135 -12730
rect 31255 -12850 31300 -12730
rect 31420 -12850 31465 -12730
rect 31585 -12850 31640 -12730
rect 31760 -12850 31805 -12730
rect 31925 -12850 31970 -12730
rect 32090 -12850 32135 -12730
rect 32255 -12850 32310 -12730
rect 32430 -12850 32475 -12730
rect 32595 -12850 32640 -12730
rect 32760 -12850 32805 -12730
rect 32925 -12850 32980 -12730
rect 33100 -12850 33145 -12730
rect 33265 -12850 33310 -12730
rect 33430 -12850 33475 -12730
rect 33595 -12850 33650 -12730
rect 33770 -12850 33815 -12730
rect 33935 -12850 33980 -12730
rect 34100 -12850 34145 -12730
rect 34265 -12850 34320 -12730
rect 34440 -12850 34485 -12730
rect 34605 -12850 34650 -12730
rect 34770 -12850 34815 -12730
rect 34935 -12850 34990 -12730
rect 35110 -12850 35155 -12730
rect 35275 -12850 35320 -12730
rect 35440 -12850 35485 -12730
rect 35605 -12850 35660 -12730
rect 35780 -12850 35825 -12730
rect 35945 -12850 35990 -12730
rect 36110 -12850 36155 -12730
rect 36275 -12850 36285 -12730
rect 30785 -12895 36285 -12850
rect 30785 -13015 30795 -12895
rect 30915 -13015 30970 -12895
rect 31090 -13015 31135 -12895
rect 31255 -13015 31300 -12895
rect 31420 -13015 31465 -12895
rect 31585 -13015 31640 -12895
rect 31760 -13015 31805 -12895
rect 31925 -13015 31970 -12895
rect 32090 -13015 32135 -12895
rect 32255 -13015 32310 -12895
rect 32430 -13015 32475 -12895
rect 32595 -13015 32640 -12895
rect 32760 -13015 32805 -12895
rect 32925 -13015 32980 -12895
rect 33100 -13015 33145 -12895
rect 33265 -13015 33310 -12895
rect 33430 -13015 33475 -12895
rect 33595 -13015 33650 -12895
rect 33770 -13015 33815 -12895
rect 33935 -13015 33980 -12895
rect 34100 -13015 34145 -12895
rect 34265 -13015 34320 -12895
rect 34440 -13015 34485 -12895
rect 34605 -13015 34650 -12895
rect 34770 -13015 34815 -12895
rect 34935 -13015 34990 -12895
rect 35110 -13015 35155 -12895
rect 35275 -13015 35320 -12895
rect 35440 -13015 35485 -12895
rect 35605 -13015 35660 -12895
rect 35780 -13015 35825 -12895
rect 35945 -13015 35990 -12895
rect 36110 -13015 36155 -12895
rect 36275 -13015 36285 -12895
rect 30785 -13060 36285 -13015
rect 30785 -13180 30795 -13060
rect 30915 -13180 30970 -13060
rect 31090 -13180 31135 -13060
rect 31255 -13180 31300 -13060
rect 31420 -13180 31465 -13060
rect 31585 -13180 31640 -13060
rect 31760 -13180 31805 -13060
rect 31925 -13180 31970 -13060
rect 32090 -13180 32135 -13060
rect 32255 -13180 32310 -13060
rect 32430 -13180 32475 -13060
rect 32595 -13180 32640 -13060
rect 32760 -13180 32805 -13060
rect 32925 -13180 32980 -13060
rect 33100 -13180 33145 -13060
rect 33265 -13180 33310 -13060
rect 33430 -13180 33475 -13060
rect 33595 -13180 33650 -13060
rect 33770 -13180 33815 -13060
rect 33935 -13180 33980 -13060
rect 34100 -13180 34145 -13060
rect 34265 -13180 34320 -13060
rect 34440 -13180 34485 -13060
rect 34605 -13180 34650 -13060
rect 34770 -13180 34815 -13060
rect 34935 -13180 34990 -13060
rect 35110 -13180 35155 -13060
rect 35275 -13180 35320 -13060
rect 35440 -13180 35485 -13060
rect 35605 -13180 35660 -13060
rect 35780 -13180 35825 -13060
rect 35945 -13180 35990 -13060
rect 36110 -13180 36155 -13060
rect 36275 -13180 36285 -13060
rect 30785 -13225 36285 -13180
rect 30785 -13345 30795 -13225
rect 30915 -13345 30970 -13225
rect 31090 -13345 31135 -13225
rect 31255 -13345 31300 -13225
rect 31420 -13345 31465 -13225
rect 31585 -13345 31640 -13225
rect 31760 -13345 31805 -13225
rect 31925 -13345 31970 -13225
rect 32090 -13345 32135 -13225
rect 32255 -13345 32310 -13225
rect 32430 -13345 32475 -13225
rect 32595 -13345 32640 -13225
rect 32760 -13345 32805 -13225
rect 32925 -13345 32980 -13225
rect 33100 -13345 33145 -13225
rect 33265 -13345 33310 -13225
rect 33430 -13345 33475 -13225
rect 33595 -13345 33650 -13225
rect 33770 -13345 33815 -13225
rect 33935 -13345 33980 -13225
rect 34100 -13345 34145 -13225
rect 34265 -13345 34320 -13225
rect 34440 -13345 34485 -13225
rect 34605 -13345 34650 -13225
rect 34770 -13345 34815 -13225
rect 34935 -13345 34990 -13225
rect 35110 -13345 35155 -13225
rect 35275 -13345 35320 -13225
rect 35440 -13345 35485 -13225
rect 35605 -13345 35660 -13225
rect 35780 -13345 35825 -13225
rect 35945 -13345 35990 -13225
rect 36110 -13345 36155 -13225
rect 36275 -13345 36285 -13225
rect 30785 -13400 36285 -13345
rect 30785 -13520 30795 -13400
rect 30915 -13520 30970 -13400
rect 31090 -13520 31135 -13400
rect 31255 -13520 31300 -13400
rect 31420 -13520 31465 -13400
rect 31585 -13520 31640 -13400
rect 31760 -13520 31805 -13400
rect 31925 -13520 31970 -13400
rect 32090 -13520 32135 -13400
rect 32255 -13520 32310 -13400
rect 32430 -13520 32475 -13400
rect 32595 -13520 32640 -13400
rect 32760 -13520 32805 -13400
rect 32925 -13520 32980 -13400
rect 33100 -13520 33145 -13400
rect 33265 -13520 33310 -13400
rect 33430 -13520 33475 -13400
rect 33595 -13520 33650 -13400
rect 33770 -13520 33815 -13400
rect 33935 -13520 33980 -13400
rect 34100 -13520 34145 -13400
rect 34265 -13520 34320 -13400
rect 34440 -13520 34485 -13400
rect 34605 -13520 34650 -13400
rect 34770 -13520 34815 -13400
rect 34935 -13520 34990 -13400
rect 35110 -13520 35155 -13400
rect 35275 -13520 35320 -13400
rect 35440 -13520 35485 -13400
rect 35605 -13520 35660 -13400
rect 35780 -13520 35825 -13400
rect 35945 -13520 35990 -13400
rect 36110 -13520 36155 -13400
rect 36275 -13520 36285 -13400
rect 30785 -13565 36285 -13520
rect 30785 -13685 30795 -13565
rect 30915 -13685 30970 -13565
rect 31090 -13685 31135 -13565
rect 31255 -13685 31300 -13565
rect 31420 -13685 31465 -13565
rect 31585 -13685 31640 -13565
rect 31760 -13685 31805 -13565
rect 31925 -13685 31970 -13565
rect 32090 -13685 32135 -13565
rect 32255 -13685 32310 -13565
rect 32430 -13685 32475 -13565
rect 32595 -13685 32640 -13565
rect 32760 -13685 32805 -13565
rect 32925 -13685 32980 -13565
rect 33100 -13685 33145 -13565
rect 33265 -13685 33310 -13565
rect 33430 -13685 33475 -13565
rect 33595 -13685 33650 -13565
rect 33770 -13685 33815 -13565
rect 33935 -13685 33980 -13565
rect 34100 -13685 34145 -13565
rect 34265 -13685 34320 -13565
rect 34440 -13685 34485 -13565
rect 34605 -13685 34650 -13565
rect 34770 -13685 34815 -13565
rect 34935 -13685 34990 -13565
rect 35110 -13685 35155 -13565
rect 35275 -13685 35320 -13565
rect 35440 -13685 35485 -13565
rect 35605 -13685 35660 -13565
rect 35780 -13685 35825 -13565
rect 35945 -13685 35990 -13565
rect 36110 -13685 36155 -13565
rect 36275 -13685 36285 -13565
rect 30785 -13730 36285 -13685
rect 30785 -13850 30795 -13730
rect 30915 -13850 30970 -13730
rect 31090 -13850 31135 -13730
rect 31255 -13850 31300 -13730
rect 31420 -13850 31465 -13730
rect 31585 -13850 31640 -13730
rect 31760 -13850 31805 -13730
rect 31925 -13850 31970 -13730
rect 32090 -13850 32135 -13730
rect 32255 -13850 32310 -13730
rect 32430 -13850 32475 -13730
rect 32595 -13850 32640 -13730
rect 32760 -13850 32805 -13730
rect 32925 -13850 32980 -13730
rect 33100 -13850 33145 -13730
rect 33265 -13850 33310 -13730
rect 33430 -13850 33475 -13730
rect 33595 -13850 33650 -13730
rect 33770 -13850 33815 -13730
rect 33935 -13850 33980 -13730
rect 34100 -13850 34145 -13730
rect 34265 -13850 34320 -13730
rect 34440 -13850 34485 -13730
rect 34605 -13850 34650 -13730
rect 34770 -13850 34815 -13730
rect 34935 -13850 34990 -13730
rect 35110 -13850 35155 -13730
rect 35275 -13850 35320 -13730
rect 35440 -13850 35485 -13730
rect 35605 -13850 35660 -13730
rect 35780 -13850 35825 -13730
rect 35945 -13850 35990 -13730
rect 36110 -13850 36155 -13730
rect 36275 -13850 36285 -13730
rect 30785 -13895 36285 -13850
rect 30785 -14015 30795 -13895
rect 30915 -14015 30970 -13895
rect 31090 -14015 31135 -13895
rect 31255 -14015 31300 -13895
rect 31420 -14015 31465 -13895
rect 31585 -14015 31640 -13895
rect 31760 -14015 31805 -13895
rect 31925 -14015 31970 -13895
rect 32090 -14015 32135 -13895
rect 32255 -14015 32310 -13895
rect 32430 -14015 32475 -13895
rect 32595 -14015 32640 -13895
rect 32760 -14015 32805 -13895
rect 32925 -14015 32980 -13895
rect 33100 -14015 33145 -13895
rect 33265 -14015 33310 -13895
rect 33430 -14015 33475 -13895
rect 33595 -14015 33650 -13895
rect 33770 -14015 33815 -13895
rect 33935 -14015 33980 -13895
rect 34100 -14015 34145 -13895
rect 34265 -14015 34320 -13895
rect 34440 -14015 34485 -13895
rect 34605 -14015 34650 -13895
rect 34770 -14015 34815 -13895
rect 34935 -14015 34990 -13895
rect 35110 -14015 35155 -13895
rect 35275 -14015 35320 -13895
rect 35440 -14015 35485 -13895
rect 35605 -14015 35660 -13895
rect 35780 -14015 35825 -13895
rect 35945 -14015 35990 -13895
rect 36110 -14015 36155 -13895
rect 36275 -14015 36285 -13895
rect 30785 -14070 36285 -14015
rect 30785 -14190 30795 -14070
rect 30915 -14190 30970 -14070
rect 31090 -14190 31135 -14070
rect 31255 -14190 31300 -14070
rect 31420 -14190 31465 -14070
rect 31585 -14190 31640 -14070
rect 31760 -14190 31805 -14070
rect 31925 -14190 31970 -14070
rect 32090 -14190 32135 -14070
rect 32255 -14190 32310 -14070
rect 32430 -14190 32475 -14070
rect 32595 -14190 32640 -14070
rect 32760 -14190 32805 -14070
rect 32925 -14190 32980 -14070
rect 33100 -14190 33145 -14070
rect 33265 -14190 33310 -14070
rect 33430 -14190 33475 -14070
rect 33595 -14190 33650 -14070
rect 33770 -14190 33815 -14070
rect 33935 -14190 33980 -14070
rect 34100 -14190 34145 -14070
rect 34265 -14190 34320 -14070
rect 34440 -14190 34485 -14070
rect 34605 -14190 34650 -14070
rect 34770 -14190 34815 -14070
rect 34935 -14190 34990 -14070
rect 35110 -14190 35155 -14070
rect 35275 -14190 35320 -14070
rect 35440 -14190 35485 -14070
rect 35605 -14190 35660 -14070
rect 35780 -14190 35825 -14070
rect 35945 -14190 35990 -14070
rect 36110 -14190 36155 -14070
rect 36275 -14190 36285 -14070
rect 30785 -14235 36285 -14190
rect 30785 -14355 30795 -14235
rect 30915 -14355 30970 -14235
rect 31090 -14355 31135 -14235
rect 31255 -14355 31300 -14235
rect 31420 -14355 31465 -14235
rect 31585 -14355 31640 -14235
rect 31760 -14355 31805 -14235
rect 31925 -14355 31970 -14235
rect 32090 -14355 32135 -14235
rect 32255 -14355 32310 -14235
rect 32430 -14355 32475 -14235
rect 32595 -14355 32640 -14235
rect 32760 -14355 32805 -14235
rect 32925 -14355 32980 -14235
rect 33100 -14355 33145 -14235
rect 33265 -14355 33310 -14235
rect 33430 -14355 33475 -14235
rect 33595 -14355 33650 -14235
rect 33770 -14355 33815 -14235
rect 33935 -14355 33980 -14235
rect 34100 -14355 34145 -14235
rect 34265 -14355 34320 -14235
rect 34440 -14355 34485 -14235
rect 34605 -14355 34650 -14235
rect 34770 -14355 34815 -14235
rect 34935 -14355 34990 -14235
rect 35110 -14355 35155 -14235
rect 35275 -14355 35320 -14235
rect 35440 -14355 35485 -14235
rect 35605 -14355 35660 -14235
rect 35780 -14355 35825 -14235
rect 35945 -14355 35990 -14235
rect 36110 -14355 36155 -14235
rect 36275 -14355 36285 -14235
rect 30785 -14400 36285 -14355
rect 30785 -14520 30795 -14400
rect 30915 -14520 30970 -14400
rect 31090 -14520 31135 -14400
rect 31255 -14520 31300 -14400
rect 31420 -14520 31465 -14400
rect 31585 -14520 31640 -14400
rect 31760 -14520 31805 -14400
rect 31925 -14520 31970 -14400
rect 32090 -14520 32135 -14400
rect 32255 -14520 32310 -14400
rect 32430 -14520 32475 -14400
rect 32595 -14520 32640 -14400
rect 32760 -14520 32805 -14400
rect 32925 -14520 32980 -14400
rect 33100 -14520 33145 -14400
rect 33265 -14520 33310 -14400
rect 33430 -14520 33475 -14400
rect 33595 -14520 33650 -14400
rect 33770 -14520 33815 -14400
rect 33935 -14520 33980 -14400
rect 34100 -14520 34145 -14400
rect 34265 -14520 34320 -14400
rect 34440 -14520 34485 -14400
rect 34605 -14520 34650 -14400
rect 34770 -14520 34815 -14400
rect 34935 -14520 34990 -14400
rect 35110 -14520 35155 -14400
rect 35275 -14520 35320 -14400
rect 35440 -14520 35485 -14400
rect 35605 -14520 35660 -14400
rect 35780 -14520 35825 -14400
rect 35945 -14520 35990 -14400
rect 36110 -14520 36155 -14400
rect 36275 -14520 36285 -14400
rect 30785 -14565 36285 -14520
rect 30785 -14685 30795 -14565
rect 30915 -14685 30970 -14565
rect 31090 -14685 31135 -14565
rect 31255 -14685 31300 -14565
rect 31420 -14685 31465 -14565
rect 31585 -14685 31640 -14565
rect 31760 -14685 31805 -14565
rect 31925 -14685 31970 -14565
rect 32090 -14685 32135 -14565
rect 32255 -14685 32310 -14565
rect 32430 -14685 32475 -14565
rect 32595 -14685 32640 -14565
rect 32760 -14685 32805 -14565
rect 32925 -14685 32980 -14565
rect 33100 -14685 33145 -14565
rect 33265 -14685 33310 -14565
rect 33430 -14685 33475 -14565
rect 33595 -14685 33650 -14565
rect 33770 -14685 33815 -14565
rect 33935 -14685 33980 -14565
rect 34100 -14685 34145 -14565
rect 34265 -14685 34320 -14565
rect 34440 -14685 34485 -14565
rect 34605 -14685 34650 -14565
rect 34770 -14685 34815 -14565
rect 34935 -14685 34990 -14565
rect 35110 -14685 35155 -14565
rect 35275 -14685 35320 -14565
rect 35440 -14685 35485 -14565
rect 35605 -14685 35660 -14565
rect 35780 -14685 35825 -14565
rect 35945 -14685 35990 -14565
rect 36110 -14685 36155 -14565
rect 36275 -14685 36285 -14565
rect 30785 -14740 36285 -14685
rect 30785 -14860 30795 -14740
rect 30915 -14860 30970 -14740
rect 31090 -14860 31135 -14740
rect 31255 -14860 31300 -14740
rect 31420 -14860 31465 -14740
rect 31585 -14860 31640 -14740
rect 31760 -14860 31805 -14740
rect 31925 -14860 31970 -14740
rect 32090 -14860 32135 -14740
rect 32255 -14860 32310 -14740
rect 32430 -14860 32475 -14740
rect 32595 -14860 32640 -14740
rect 32760 -14860 32805 -14740
rect 32925 -14860 32980 -14740
rect 33100 -14860 33145 -14740
rect 33265 -14860 33310 -14740
rect 33430 -14860 33475 -14740
rect 33595 -14860 33650 -14740
rect 33770 -14860 33815 -14740
rect 33935 -14860 33980 -14740
rect 34100 -14860 34145 -14740
rect 34265 -14860 34320 -14740
rect 34440 -14860 34485 -14740
rect 34605 -14860 34650 -14740
rect 34770 -14860 34815 -14740
rect 34935 -14860 34990 -14740
rect 35110 -14860 35155 -14740
rect 35275 -14860 35320 -14740
rect 35440 -14860 35485 -14740
rect 35605 -14860 35660 -14740
rect 35780 -14860 35825 -14740
rect 35945 -14860 35990 -14740
rect 36110 -14860 36155 -14740
rect 36275 -14860 36285 -14740
rect 30785 -14905 36285 -14860
rect 30785 -15025 30795 -14905
rect 30915 -15025 30970 -14905
rect 31090 -15025 31135 -14905
rect 31255 -15025 31300 -14905
rect 31420 -15025 31465 -14905
rect 31585 -15025 31640 -14905
rect 31760 -15025 31805 -14905
rect 31925 -15025 31970 -14905
rect 32090 -15025 32135 -14905
rect 32255 -15025 32310 -14905
rect 32430 -15025 32475 -14905
rect 32595 -15025 32640 -14905
rect 32760 -15025 32805 -14905
rect 32925 -15025 32980 -14905
rect 33100 -15025 33145 -14905
rect 33265 -15025 33310 -14905
rect 33430 -15025 33475 -14905
rect 33595 -15025 33650 -14905
rect 33770 -15025 33815 -14905
rect 33935 -15025 33980 -14905
rect 34100 -15025 34145 -14905
rect 34265 -15025 34320 -14905
rect 34440 -15025 34485 -14905
rect 34605 -15025 34650 -14905
rect 34770 -15025 34815 -14905
rect 34935 -15025 34990 -14905
rect 35110 -15025 35155 -14905
rect 35275 -15025 35320 -14905
rect 35440 -15025 35485 -14905
rect 35605 -15025 35660 -14905
rect 35780 -15025 35825 -14905
rect 35945 -15025 35990 -14905
rect 36110 -15025 36155 -14905
rect 36275 -15025 36285 -14905
rect 30785 -15070 36285 -15025
rect 30785 -15190 30795 -15070
rect 30915 -15190 30970 -15070
rect 31090 -15190 31135 -15070
rect 31255 -15190 31300 -15070
rect 31420 -15190 31465 -15070
rect 31585 -15190 31640 -15070
rect 31760 -15190 31805 -15070
rect 31925 -15190 31970 -15070
rect 32090 -15190 32135 -15070
rect 32255 -15190 32310 -15070
rect 32430 -15190 32475 -15070
rect 32595 -15190 32640 -15070
rect 32760 -15190 32805 -15070
rect 32925 -15190 32980 -15070
rect 33100 -15190 33145 -15070
rect 33265 -15190 33310 -15070
rect 33430 -15190 33475 -15070
rect 33595 -15190 33650 -15070
rect 33770 -15190 33815 -15070
rect 33935 -15190 33980 -15070
rect 34100 -15190 34145 -15070
rect 34265 -15190 34320 -15070
rect 34440 -15190 34485 -15070
rect 34605 -15190 34650 -15070
rect 34770 -15190 34815 -15070
rect 34935 -15190 34990 -15070
rect 35110 -15190 35155 -15070
rect 35275 -15190 35320 -15070
rect 35440 -15190 35485 -15070
rect 35605 -15190 35660 -15070
rect 35780 -15190 35825 -15070
rect 35945 -15190 35990 -15070
rect 36110 -15190 36155 -15070
rect 36275 -15190 36285 -15070
rect 30785 -15235 36285 -15190
rect 30785 -15355 30795 -15235
rect 30915 -15355 30970 -15235
rect 31090 -15355 31135 -15235
rect 31255 -15355 31300 -15235
rect 31420 -15355 31465 -15235
rect 31585 -15355 31640 -15235
rect 31760 -15355 31805 -15235
rect 31925 -15355 31970 -15235
rect 32090 -15355 32135 -15235
rect 32255 -15355 32310 -15235
rect 32430 -15355 32475 -15235
rect 32595 -15355 32640 -15235
rect 32760 -15355 32805 -15235
rect 32925 -15355 32980 -15235
rect 33100 -15355 33145 -15235
rect 33265 -15355 33310 -15235
rect 33430 -15355 33475 -15235
rect 33595 -15355 33650 -15235
rect 33770 -15355 33815 -15235
rect 33935 -15355 33980 -15235
rect 34100 -15355 34145 -15235
rect 34265 -15355 34320 -15235
rect 34440 -15355 34485 -15235
rect 34605 -15355 34650 -15235
rect 34770 -15355 34815 -15235
rect 34935 -15355 34990 -15235
rect 35110 -15355 35155 -15235
rect 35275 -15355 35320 -15235
rect 35440 -15355 35485 -15235
rect 35605 -15355 35660 -15235
rect 35780 -15355 35825 -15235
rect 35945 -15355 35990 -15235
rect 36110 -15355 36155 -15235
rect 36275 -15355 36285 -15235
rect 30785 -15410 36285 -15355
rect 30785 -15530 30795 -15410
rect 30915 -15530 30970 -15410
rect 31090 -15530 31135 -15410
rect 31255 -15530 31300 -15410
rect 31420 -15530 31465 -15410
rect 31585 -15530 31640 -15410
rect 31760 -15530 31805 -15410
rect 31925 -15530 31970 -15410
rect 32090 -15530 32135 -15410
rect 32255 -15530 32310 -15410
rect 32430 -15530 32475 -15410
rect 32595 -15530 32640 -15410
rect 32760 -15530 32805 -15410
rect 32925 -15530 32980 -15410
rect 33100 -15530 33145 -15410
rect 33265 -15530 33310 -15410
rect 33430 -15530 33475 -15410
rect 33595 -15530 33650 -15410
rect 33770 -15530 33815 -15410
rect 33935 -15530 33980 -15410
rect 34100 -15530 34145 -15410
rect 34265 -15530 34320 -15410
rect 34440 -15530 34485 -15410
rect 34605 -15530 34650 -15410
rect 34770 -15530 34815 -15410
rect 34935 -15530 34990 -15410
rect 35110 -15530 35155 -15410
rect 35275 -15530 35320 -15410
rect 35440 -15530 35485 -15410
rect 35605 -15530 35660 -15410
rect 35780 -15530 35825 -15410
rect 35945 -15530 35990 -15410
rect 36110 -15530 36155 -15410
rect 36275 -15530 36285 -15410
rect 30785 -15540 36285 -15530
rect 36475 -10050 41975 -10040
rect 36475 -10170 36485 -10050
rect 36605 -10170 36660 -10050
rect 36780 -10170 36825 -10050
rect 36945 -10170 36990 -10050
rect 37110 -10170 37155 -10050
rect 37275 -10170 37330 -10050
rect 37450 -10170 37495 -10050
rect 37615 -10170 37660 -10050
rect 37780 -10170 37825 -10050
rect 37945 -10170 38000 -10050
rect 38120 -10170 38165 -10050
rect 38285 -10170 38330 -10050
rect 38450 -10170 38495 -10050
rect 38615 -10170 38670 -10050
rect 38790 -10170 38835 -10050
rect 38955 -10170 39000 -10050
rect 39120 -10170 39165 -10050
rect 39285 -10170 39340 -10050
rect 39460 -10170 39505 -10050
rect 39625 -10170 39670 -10050
rect 39790 -10170 39835 -10050
rect 39955 -10170 40010 -10050
rect 40130 -10170 40175 -10050
rect 40295 -10170 40340 -10050
rect 40460 -10170 40505 -10050
rect 40625 -10170 40680 -10050
rect 40800 -10170 40845 -10050
rect 40965 -10170 41010 -10050
rect 41130 -10170 41175 -10050
rect 41295 -10170 41350 -10050
rect 41470 -10170 41515 -10050
rect 41635 -10170 41680 -10050
rect 41800 -10170 41845 -10050
rect 41965 -10170 41975 -10050
rect 36475 -10215 41975 -10170
rect 36475 -10335 36485 -10215
rect 36605 -10335 36660 -10215
rect 36780 -10335 36825 -10215
rect 36945 -10335 36990 -10215
rect 37110 -10335 37155 -10215
rect 37275 -10335 37330 -10215
rect 37450 -10335 37495 -10215
rect 37615 -10335 37660 -10215
rect 37780 -10335 37825 -10215
rect 37945 -10335 38000 -10215
rect 38120 -10335 38165 -10215
rect 38285 -10335 38330 -10215
rect 38450 -10335 38495 -10215
rect 38615 -10335 38670 -10215
rect 38790 -10335 38835 -10215
rect 38955 -10335 39000 -10215
rect 39120 -10335 39165 -10215
rect 39285 -10335 39340 -10215
rect 39460 -10335 39505 -10215
rect 39625 -10335 39670 -10215
rect 39790 -10335 39835 -10215
rect 39955 -10335 40010 -10215
rect 40130 -10335 40175 -10215
rect 40295 -10335 40340 -10215
rect 40460 -10335 40505 -10215
rect 40625 -10335 40680 -10215
rect 40800 -10335 40845 -10215
rect 40965 -10335 41010 -10215
rect 41130 -10335 41175 -10215
rect 41295 -10335 41350 -10215
rect 41470 -10335 41515 -10215
rect 41635 -10335 41680 -10215
rect 41800 -10335 41845 -10215
rect 41965 -10335 41975 -10215
rect 36475 -10380 41975 -10335
rect 36475 -10500 36485 -10380
rect 36605 -10500 36660 -10380
rect 36780 -10500 36825 -10380
rect 36945 -10500 36990 -10380
rect 37110 -10500 37155 -10380
rect 37275 -10500 37330 -10380
rect 37450 -10500 37495 -10380
rect 37615 -10500 37660 -10380
rect 37780 -10500 37825 -10380
rect 37945 -10500 38000 -10380
rect 38120 -10500 38165 -10380
rect 38285 -10500 38330 -10380
rect 38450 -10500 38495 -10380
rect 38615 -10500 38670 -10380
rect 38790 -10500 38835 -10380
rect 38955 -10500 39000 -10380
rect 39120 -10500 39165 -10380
rect 39285 -10500 39340 -10380
rect 39460 -10500 39505 -10380
rect 39625 -10500 39670 -10380
rect 39790 -10500 39835 -10380
rect 39955 -10500 40010 -10380
rect 40130 -10500 40175 -10380
rect 40295 -10500 40340 -10380
rect 40460 -10500 40505 -10380
rect 40625 -10500 40680 -10380
rect 40800 -10500 40845 -10380
rect 40965 -10500 41010 -10380
rect 41130 -10500 41175 -10380
rect 41295 -10500 41350 -10380
rect 41470 -10500 41515 -10380
rect 41635 -10500 41680 -10380
rect 41800 -10500 41845 -10380
rect 41965 -10500 41975 -10380
rect 36475 -10545 41975 -10500
rect 36475 -10665 36485 -10545
rect 36605 -10665 36660 -10545
rect 36780 -10665 36825 -10545
rect 36945 -10665 36990 -10545
rect 37110 -10665 37155 -10545
rect 37275 -10665 37330 -10545
rect 37450 -10665 37495 -10545
rect 37615 -10665 37660 -10545
rect 37780 -10665 37825 -10545
rect 37945 -10665 38000 -10545
rect 38120 -10665 38165 -10545
rect 38285 -10665 38330 -10545
rect 38450 -10665 38495 -10545
rect 38615 -10665 38670 -10545
rect 38790 -10665 38835 -10545
rect 38955 -10665 39000 -10545
rect 39120 -10665 39165 -10545
rect 39285 -10665 39340 -10545
rect 39460 -10665 39505 -10545
rect 39625 -10665 39670 -10545
rect 39790 -10665 39835 -10545
rect 39955 -10665 40010 -10545
rect 40130 -10665 40175 -10545
rect 40295 -10665 40340 -10545
rect 40460 -10665 40505 -10545
rect 40625 -10665 40680 -10545
rect 40800 -10665 40845 -10545
rect 40965 -10665 41010 -10545
rect 41130 -10665 41175 -10545
rect 41295 -10665 41350 -10545
rect 41470 -10665 41515 -10545
rect 41635 -10665 41680 -10545
rect 41800 -10665 41845 -10545
rect 41965 -10665 41975 -10545
rect 36475 -10720 41975 -10665
rect 36475 -10840 36485 -10720
rect 36605 -10840 36660 -10720
rect 36780 -10840 36825 -10720
rect 36945 -10840 36990 -10720
rect 37110 -10840 37155 -10720
rect 37275 -10840 37330 -10720
rect 37450 -10840 37495 -10720
rect 37615 -10840 37660 -10720
rect 37780 -10840 37825 -10720
rect 37945 -10840 38000 -10720
rect 38120 -10840 38165 -10720
rect 38285 -10840 38330 -10720
rect 38450 -10840 38495 -10720
rect 38615 -10840 38670 -10720
rect 38790 -10840 38835 -10720
rect 38955 -10840 39000 -10720
rect 39120 -10840 39165 -10720
rect 39285 -10840 39340 -10720
rect 39460 -10840 39505 -10720
rect 39625 -10840 39670 -10720
rect 39790 -10840 39835 -10720
rect 39955 -10840 40010 -10720
rect 40130 -10840 40175 -10720
rect 40295 -10840 40340 -10720
rect 40460 -10840 40505 -10720
rect 40625 -10840 40680 -10720
rect 40800 -10840 40845 -10720
rect 40965 -10840 41010 -10720
rect 41130 -10840 41175 -10720
rect 41295 -10840 41350 -10720
rect 41470 -10840 41515 -10720
rect 41635 -10840 41680 -10720
rect 41800 -10840 41845 -10720
rect 41965 -10840 41975 -10720
rect 36475 -10885 41975 -10840
rect 36475 -11005 36485 -10885
rect 36605 -11005 36660 -10885
rect 36780 -11005 36825 -10885
rect 36945 -11005 36990 -10885
rect 37110 -11005 37155 -10885
rect 37275 -11005 37330 -10885
rect 37450 -11005 37495 -10885
rect 37615 -11005 37660 -10885
rect 37780 -11005 37825 -10885
rect 37945 -11005 38000 -10885
rect 38120 -11005 38165 -10885
rect 38285 -11005 38330 -10885
rect 38450 -11005 38495 -10885
rect 38615 -11005 38670 -10885
rect 38790 -11005 38835 -10885
rect 38955 -11005 39000 -10885
rect 39120 -11005 39165 -10885
rect 39285 -11005 39340 -10885
rect 39460 -11005 39505 -10885
rect 39625 -11005 39670 -10885
rect 39790 -11005 39835 -10885
rect 39955 -11005 40010 -10885
rect 40130 -11005 40175 -10885
rect 40295 -11005 40340 -10885
rect 40460 -11005 40505 -10885
rect 40625 -11005 40680 -10885
rect 40800 -11005 40845 -10885
rect 40965 -11005 41010 -10885
rect 41130 -11005 41175 -10885
rect 41295 -11005 41350 -10885
rect 41470 -11005 41515 -10885
rect 41635 -11005 41680 -10885
rect 41800 -11005 41845 -10885
rect 41965 -11005 41975 -10885
rect 36475 -11050 41975 -11005
rect 36475 -11170 36485 -11050
rect 36605 -11170 36660 -11050
rect 36780 -11170 36825 -11050
rect 36945 -11170 36990 -11050
rect 37110 -11170 37155 -11050
rect 37275 -11170 37330 -11050
rect 37450 -11170 37495 -11050
rect 37615 -11170 37660 -11050
rect 37780 -11170 37825 -11050
rect 37945 -11170 38000 -11050
rect 38120 -11170 38165 -11050
rect 38285 -11170 38330 -11050
rect 38450 -11170 38495 -11050
rect 38615 -11170 38670 -11050
rect 38790 -11170 38835 -11050
rect 38955 -11170 39000 -11050
rect 39120 -11170 39165 -11050
rect 39285 -11170 39340 -11050
rect 39460 -11170 39505 -11050
rect 39625 -11170 39670 -11050
rect 39790 -11170 39835 -11050
rect 39955 -11170 40010 -11050
rect 40130 -11170 40175 -11050
rect 40295 -11170 40340 -11050
rect 40460 -11170 40505 -11050
rect 40625 -11170 40680 -11050
rect 40800 -11170 40845 -11050
rect 40965 -11170 41010 -11050
rect 41130 -11170 41175 -11050
rect 41295 -11170 41350 -11050
rect 41470 -11170 41515 -11050
rect 41635 -11170 41680 -11050
rect 41800 -11170 41845 -11050
rect 41965 -11170 41975 -11050
rect 36475 -11215 41975 -11170
rect 36475 -11335 36485 -11215
rect 36605 -11335 36660 -11215
rect 36780 -11335 36825 -11215
rect 36945 -11335 36990 -11215
rect 37110 -11335 37155 -11215
rect 37275 -11335 37330 -11215
rect 37450 -11335 37495 -11215
rect 37615 -11335 37660 -11215
rect 37780 -11335 37825 -11215
rect 37945 -11335 38000 -11215
rect 38120 -11335 38165 -11215
rect 38285 -11335 38330 -11215
rect 38450 -11335 38495 -11215
rect 38615 -11335 38670 -11215
rect 38790 -11335 38835 -11215
rect 38955 -11335 39000 -11215
rect 39120 -11335 39165 -11215
rect 39285 -11335 39340 -11215
rect 39460 -11335 39505 -11215
rect 39625 -11335 39670 -11215
rect 39790 -11335 39835 -11215
rect 39955 -11335 40010 -11215
rect 40130 -11335 40175 -11215
rect 40295 -11335 40340 -11215
rect 40460 -11335 40505 -11215
rect 40625 -11335 40680 -11215
rect 40800 -11335 40845 -11215
rect 40965 -11335 41010 -11215
rect 41130 -11335 41175 -11215
rect 41295 -11335 41350 -11215
rect 41470 -11335 41515 -11215
rect 41635 -11335 41680 -11215
rect 41800 -11335 41845 -11215
rect 41965 -11335 41975 -11215
rect 36475 -11390 41975 -11335
rect 36475 -11510 36485 -11390
rect 36605 -11510 36660 -11390
rect 36780 -11510 36825 -11390
rect 36945 -11510 36990 -11390
rect 37110 -11510 37155 -11390
rect 37275 -11510 37330 -11390
rect 37450 -11510 37495 -11390
rect 37615 -11510 37660 -11390
rect 37780 -11510 37825 -11390
rect 37945 -11510 38000 -11390
rect 38120 -11510 38165 -11390
rect 38285 -11510 38330 -11390
rect 38450 -11510 38495 -11390
rect 38615 -11510 38670 -11390
rect 38790 -11510 38835 -11390
rect 38955 -11510 39000 -11390
rect 39120 -11510 39165 -11390
rect 39285 -11510 39340 -11390
rect 39460 -11510 39505 -11390
rect 39625 -11510 39670 -11390
rect 39790 -11510 39835 -11390
rect 39955 -11510 40010 -11390
rect 40130 -11510 40175 -11390
rect 40295 -11510 40340 -11390
rect 40460 -11510 40505 -11390
rect 40625 -11510 40680 -11390
rect 40800 -11510 40845 -11390
rect 40965 -11510 41010 -11390
rect 41130 -11510 41175 -11390
rect 41295 -11510 41350 -11390
rect 41470 -11510 41515 -11390
rect 41635 -11510 41680 -11390
rect 41800 -11510 41845 -11390
rect 41965 -11510 41975 -11390
rect 36475 -11555 41975 -11510
rect 36475 -11675 36485 -11555
rect 36605 -11675 36660 -11555
rect 36780 -11675 36825 -11555
rect 36945 -11675 36990 -11555
rect 37110 -11675 37155 -11555
rect 37275 -11675 37330 -11555
rect 37450 -11675 37495 -11555
rect 37615 -11675 37660 -11555
rect 37780 -11675 37825 -11555
rect 37945 -11675 38000 -11555
rect 38120 -11675 38165 -11555
rect 38285 -11675 38330 -11555
rect 38450 -11675 38495 -11555
rect 38615 -11675 38670 -11555
rect 38790 -11675 38835 -11555
rect 38955 -11675 39000 -11555
rect 39120 -11675 39165 -11555
rect 39285 -11675 39340 -11555
rect 39460 -11675 39505 -11555
rect 39625 -11675 39670 -11555
rect 39790 -11675 39835 -11555
rect 39955 -11675 40010 -11555
rect 40130 -11675 40175 -11555
rect 40295 -11675 40340 -11555
rect 40460 -11675 40505 -11555
rect 40625 -11675 40680 -11555
rect 40800 -11675 40845 -11555
rect 40965 -11675 41010 -11555
rect 41130 -11675 41175 -11555
rect 41295 -11675 41350 -11555
rect 41470 -11675 41515 -11555
rect 41635 -11675 41680 -11555
rect 41800 -11675 41845 -11555
rect 41965 -11675 41975 -11555
rect 36475 -11720 41975 -11675
rect 36475 -11840 36485 -11720
rect 36605 -11840 36660 -11720
rect 36780 -11840 36825 -11720
rect 36945 -11840 36990 -11720
rect 37110 -11840 37155 -11720
rect 37275 -11840 37330 -11720
rect 37450 -11840 37495 -11720
rect 37615 -11840 37660 -11720
rect 37780 -11840 37825 -11720
rect 37945 -11840 38000 -11720
rect 38120 -11840 38165 -11720
rect 38285 -11840 38330 -11720
rect 38450 -11840 38495 -11720
rect 38615 -11840 38670 -11720
rect 38790 -11840 38835 -11720
rect 38955 -11840 39000 -11720
rect 39120 -11840 39165 -11720
rect 39285 -11840 39340 -11720
rect 39460 -11840 39505 -11720
rect 39625 -11840 39670 -11720
rect 39790 -11840 39835 -11720
rect 39955 -11840 40010 -11720
rect 40130 -11840 40175 -11720
rect 40295 -11840 40340 -11720
rect 40460 -11840 40505 -11720
rect 40625 -11840 40680 -11720
rect 40800 -11840 40845 -11720
rect 40965 -11840 41010 -11720
rect 41130 -11840 41175 -11720
rect 41295 -11840 41350 -11720
rect 41470 -11840 41515 -11720
rect 41635 -11840 41680 -11720
rect 41800 -11840 41845 -11720
rect 41965 -11840 41975 -11720
rect 36475 -11885 41975 -11840
rect 36475 -12005 36485 -11885
rect 36605 -12005 36660 -11885
rect 36780 -12005 36825 -11885
rect 36945 -12005 36990 -11885
rect 37110 -12005 37155 -11885
rect 37275 -12005 37330 -11885
rect 37450 -12005 37495 -11885
rect 37615 -12005 37660 -11885
rect 37780 -12005 37825 -11885
rect 37945 -12005 38000 -11885
rect 38120 -12005 38165 -11885
rect 38285 -12005 38330 -11885
rect 38450 -12005 38495 -11885
rect 38615 -12005 38670 -11885
rect 38790 -12005 38835 -11885
rect 38955 -12005 39000 -11885
rect 39120 -12005 39165 -11885
rect 39285 -12005 39340 -11885
rect 39460 -12005 39505 -11885
rect 39625 -12005 39670 -11885
rect 39790 -12005 39835 -11885
rect 39955 -12005 40010 -11885
rect 40130 -12005 40175 -11885
rect 40295 -12005 40340 -11885
rect 40460 -12005 40505 -11885
rect 40625 -12005 40680 -11885
rect 40800 -12005 40845 -11885
rect 40965 -12005 41010 -11885
rect 41130 -12005 41175 -11885
rect 41295 -12005 41350 -11885
rect 41470 -12005 41515 -11885
rect 41635 -12005 41680 -11885
rect 41800 -12005 41845 -11885
rect 41965 -12005 41975 -11885
rect 36475 -12060 41975 -12005
rect 36475 -12180 36485 -12060
rect 36605 -12180 36660 -12060
rect 36780 -12180 36825 -12060
rect 36945 -12180 36990 -12060
rect 37110 -12180 37155 -12060
rect 37275 -12180 37330 -12060
rect 37450 -12180 37495 -12060
rect 37615 -12180 37660 -12060
rect 37780 -12180 37825 -12060
rect 37945 -12180 38000 -12060
rect 38120 -12180 38165 -12060
rect 38285 -12180 38330 -12060
rect 38450 -12180 38495 -12060
rect 38615 -12180 38670 -12060
rect 38790 -12180 38835 -12060
rect 38955 -12180 39000 -12060
rect 39120 -12180 39165 -12060
rect 39285 -12180 39340 -12060
rect 39460 -12180 39505 -12060
rect 39625 -12180 39670 -12060
rect 39790 -12180 39835 -12060
rect 39955 -12180 40010 -12060
rect 40130 -12180 40175 -12060
rect 40295 -12180 40340 -12060
rect 40460 -12180 40505 -12060
rect 40625 -12180 40680 -12060
rect 40800 -12180 40845 -12060
rect 40965 -12180 41010 -12060
rect 41130 -12180 41175 -12060
rect 41295 -12180 41350 -12060
rect 41470 -12180 41515 -12060
rect 41635 -12180 41680 -12060
rect 41800 -12180 41845 -12060
rect 41965 -12180 41975 -12060
rect 36475 -12225 41975 -12180
rect 36475 -12345 36485 -12225
rect 36605 -12345 36660 -12225
rect 36780 -12345 36825 -12225
rect 36945 -12345 36990 -12225
rect 37110 -12345 37155 -12225
rect 37275 -12345 37330 -12225
rect 37450 -12345 37495 -12225
rect 37615 -12345 37660 -12225
rect 37780 -12345 37825 -12225
rect 37945 -12345 38000 -12225
rect 38120 -12345 38165 -12225
rect 38285 -12345 38330 -12225
rect 38450 -12345 38495 -12225
rect 38615 -12345 38670 -12225
rect 38790 -12345 38835 -12225
rect 38955 -12345 39000 -12225
rect 39120 -12345 39165 -12225
rect 39285 -12345 39340 -12225
rect 39460 -12345 39505 -12225
rect 39625 -12345 39670 -12225
rect 39790 -12345 39835 -12225
rect 39955 -12345 40010 -12225
rect 40130 -12345 40175 -12225
rect 40295 -12345 40340 -12225
rect 40460 -12345 40505 -12225
rect 40625 -12345 40680 -12225
rect 40800 -12345 40845 -12225
rect 40965 -12345 41010 -12225
rect 41130 -12345 41175 -12225
rect 41295 -12345 41350 -12225
rect 41470 -12345 41515 -12225
rect 41635 -12345 41680 -12225
rect 41800 -12345 41845 -12225
rect 41965 -12345 41975 -12225
rect 36475 -12390 41975 -12345
rect 36475 -12510 36485 -12390
rect 36605 -12510 36660 -12390
rect 36780 -12510 36825 -12390
rect 36945 -12510 36990 -12390
rect 37110 -12510 37155 -12390
rect 37275 -12510 37330 -12390
rect 37450 -12510 37495 -12390
rect 37615 -12510 37660 -12390
rect 37780 -12510 37825 -12390
rect 37945 -12510 38000 -12390
rect 38120 -12510 38165 -12390
rect 38285 -12510 38330 -12390
rect 38450 -12510 38495 -12390
rect 38615 -12510 38670 -12390
rect 38790 -12510 38835 -12390
rect 38955 -12510 39000 -12390
rect 39120 -12510 39165 -12390
rect 39285 -12510 39340 -12390
rect 39460 -12510 39505 -12390
rect 39625 -12510 39670 -12390
rect 39790 -12510 39835 -12390
rect 39955 -12510 40010 -12390
rect 40130 -12510 40175 -12390
rect 40295 -12510 40340 -12390
rect 40460 -12510 40505 -12390
rect 40625 -12510 40680 -12390
rect 40800 -12510 40845 -12390
rect 40965 -12510 41010 -12390
rect 41130 -12510 41175 -12390
rect 41295 -12510 41350 -12390
rect 41470 -12510 41515 -12390
rect 41635 -12510 41680 -12390
rect 41800 -12510 41845 -12390
rect 41965 -12510 41975 -12390
rect 36475 -12555 41975 -12510
rect 36475 -12675 36485 -12555
rect 36605 -12675 36660 -12555
rect 36780 -12675 36825 -12555
rect 36945 -12675 36990 -12555
rect 37110 -12675 37155 -12555
rect 37275 -12675 37330 -12555
rect 37450 -12675 37495 -12555
rect 37615 -12675 37660 -12555
rect 37780 -12675 37825 -12555
rect 37945 -12675 38000 -12555
rect 38120 -12675 38165 -12555
rect 38285 -12675 38330 -12555
rect 38450 -12675 38495 -12555
rect 38615 -12675 38670 -12555
rect 38790 -12675 38835 -12555
rect 38955 -12675 39000 -12555
rect 39120 -12675 39165 -12555
rect 39285 -12675 39340 -12555
rect 39460 -12675 39505 -12555
rect 39625 -12675 39670 -12555
rect 39790 -12675 39835 -12555
rect 39955 -12675 40010 -12555
rect 40130 -12675 40175 -12555
rect 40295 -12675 40340 -12555
rect 40460 -12675 40505 -12555
rect 40625 -12675 40680 -12555
rect 40800 -12675 40845 -12555
rect 40965 -12675 41010 -12555
rect 41130 -12675 41175 -12555
rect 41295 -12675 41350 -12555
rect 41470 -12675 41515 -12555
rect 41635 -12675 41680 -12555
rect 41800 -12675 41845 -12555
rect 41965 -12675 41975 -12555
rect 36475 -12730 41975 -12675
rect 36475 -12850 36485 -12730
rect 36605 -12850 36660 -12730
rect 36780 -12850 36825 -12730
rect 36945 -12850 36990 -12730
rect 37110 -12850 37155 -12730
rect 37275 -12850 37330 -12730
rect 37450 -12850 37495 -12730
rect 37615 -12850 37660 -12730
rect 37780 -12850 37825 -12730
rect 37945 -12850 38000 -12730
rect 38120 -12850 38165 -12730
rect 38285 -12850 38330 -12730
rect 38450 -12850 38495 -12730
rect 38615 -12850 38670 -12730
rect 38790 -12850 38835 -12730
rect 38955 -12850 39000 -12730
rect 39120 -12850 39165 -12730
rect 39285 -12850 39340 -12730
rect 39460 -12850 39505 -12730
rect 39625 -12850 39670 -12730
rect 39790 -12850 39835 -12730
rect 39955 -12850 40010 -12730
rect 40130 -12850 40175 -12730
rect 40295 -12850 40340 -12730
rect 40460 -12850 40505 -12730
rect 40625 -12850 40680 -12730
rect 40800 -12850 40845 -12730
rect 40965 -12850 41010 -12730
rect 41130 -12850 41175 -12730
rect 41295 -12850 41350 -12730
rect 41470 -12850 41515 -12730
rect 41635 -12850 41680 -12730
rect 41800 -12850 41845 -12730
rect 41965 -12850 41975 -12730
rect 36475 -12895 41975 -12850
rect 36475 -13015 36485 -12895
rect 36605 -13015 36660 -12895
rect 36780 -13015 36825 -12895
rect 36945 -13015 36990 -12895
rect 37110 -13015 37155 -12895
rect 37275 -13015 37330 -12895
rect 37450 -13015 37495 -12895
rect 37615 -13015 37660 -12895
rect 37780 -13015 37825 -12895
rect 37945 -13015 38000 -12895
rect 38120 -13015 38165 -12895
rect 38285 -13015 38330 -12895
rect 38450 -13015 38495 -12895
rect 38615 -13015 38670 -12895
rect 38790 -13015 38835 -12895
rect 38955 -13015 39000 -12895
rect 39120 -13015 39165 -12895
rect 39285 -13015 39340 -12895
rect 39460 -13015 39505 -12895
rect 39625 -13015 39670 -12895
rect 39790 -13015 39835 -12895
rect 39955 -13015 40010 -12895
rect 40130 -13015 40175 -12895
rect 40295 -13015 40340 -12895
rect 40460 -13015 40505 -12895
rect 40625 -13015 40680 -12895
rect 40800 -13015 40845 -12895
rect 40965 -13015 41010 -12895
rect 41130 -13015 41175 -12895
rect 41295 -13015 41350 -12895
rect 41470 -13015 41515 -12895
rect 41635 -13015 41680 -12895
rect 41800 -13015 41845 -12895
rect 41965 -13015 41975 -12895
rect 36475 -13060 41975 -13015
rect 36475 -13180 36485 -13060
rect 36605 -13180 36660 -13060
rect 36780 -13180 36825 -13060
rect 36945 -13180 36990 -13060
rect 37110 -13180 37155 -13060
rect 37275 -13180 37330 -13060
rect 37450 -13180 37495 -13060
rect 37615 -13180 37660 -13060
rect 37780 -13180 37825 -13060
rect 37945 -13180 38000 -13060
rect 38120 -13180 38165 -13060
rect 38285 -13180 38330 -13060
rect 38450 -13180 38495 -13060
rect 38615 -13180 38670 -13060
rect 38790 -13180 38835 -13060
rect 38955 -13180 39000 -13060
rect 39120 -13180 39165 -13060
rect 39285 -13180 39340 -13060
rect 39460 -13180 39505 -13060
rect 39625 -13180 39670 -13060
rect 39790 -13180 39835 -13060
rect 39955 -13180 40010 -13060
rect 40130 -13180 40175 -13060
rect 40295 -13180 40340 -13060
rect 40460 -13180 40505 -13060
rect 40625 -13180 40680 -13060
rect 40800 -13180 40845 -13060
rect 40965 -13180 41010 -13060
rect 41130 -13180 41175 -13060
rect 41295 -13180 41350 -13060
rect 41470 -13180 41515 -13060
rect 41635 -13180 41680 -13060
rect 41800 -13180 41845 -13060
rect 41965 -13180 41975 -13060
rect 36475 -13225 41975 -13180
rect 36475 -13345 36485 -13225
rect 36605 -13345 36660 -13225
rect 36780 -13345 36825 -13225
rect 36945 -13345 36990 -13225
rect 37110 -13345 37155 -13225
rect 37275 -13345 37330 -13225
rect 37450 -13345 37495 -13225
rect 37615 -13345 37660 -13225
rect 37780 -13345 37825 -13225
rect 37945 -13345 38000 -13225
rect 38120 -13345 38165 -13225
rect 38285 -13345 38330 -13225
rect 38450 -13345 38495 -13225
rect 38615 -13345 38670 -13225
rect 38790 -13345 38835 -13225
rect 38955 -13345 39000 -13225
rect 39120 -13345 39165 -13225
rect 39285 -13345 39340 -13225
rect 39460 -13345 39505 -13225
rect 39625 -13345 39670 -13225
rect 39790 -13345 39835 -13225
rect 39955 -13345 40010 -13225
rect 40130 -13345 40175 -13225
rect 40295 -13345 40340 -13225
rect 40460 -13345 40505 -13225
rect 40625 -13345 40680 -13225
rect 40800 -13345 40845 -13225
rect 40965 -13345 41010 -13225
rect 41130 -13345 41175 -13225
rect 41295 -13345 41350 -13225
rect 41470 -13345 41515 -13225
rect 41635 -13345 41680 -13225
rect 41800 -13345 41845 -13225
rect 41965 -13345 41975 -13225
rect 36475 -13400 41975 -13345
rect 36475 -13520 36485 -13400
rect 36605 -13520 36660 -13400
rect 36780 -13520 36825 -13400
rect 36945 -13520 36990 -13400
rect 37110 -13520 37155 -13400
rect 37275 -13520 37330 -13400
rect 37450 -13520 37495 -13400
rect 37615 -13520 37660 -13400
rect 37780 -13520 37825 -13400
rect 37945 -13520 38000 -13400
rect 38120 -13520 38165 -13400
rect 38285 -13520 38330 -13400
rect 38450 -13520 38495 -13400
rect 38615 -13520 38670 -13400
rect 38790 -13520 38835 -13400
rect 38955 -13520 39000 -13400
rect 39120 -13520 39165 -13400
rect 39285 -13520 39340 -13400
rect 39460 -13520 39505 -13400
rect 39625 -13520 39670 -13400
rect 39790 -13520 39835 -13400
rect 39955 -13520 40010 -13400
rect 40130 -13520 40175 -13400
rect 40295 -13520 40340 -13400
rect 40460 -13520 40505 -13400
rect 40625 -13520 40680 -13400
rect 40800 -13520 40845 -13400
rect 40965 -13520 41010 -13400
rect 41130 -13520 41175 -13400
rect 41295 -13520 41350 -13400
rect 41470 -13520 41515 -13400
rect 41635 -13520 41680 -13400
rect 41800 -13520 41845 -13400
rect 41965 -13520 41975 -13400
rect 36475 -13565 41975 -13520
rect 36475 -13685 36485 -13565
rect 36605 -13685 36660 -13565
rect 36780 -13685 36825 -13565
rect 36945 -13685 36990 -13565
rect 37110 -13685 37155 -13565
rect 37275 -13685 37330 -13565
rect 37450 -13685 37495 -13565
rect 37615 -13685 37660 -13565
rect 37780 -13685 37825 -13565
rect 37945 -13685 38000 -13565
rect 38120 -13685 38165 -13565
rect 38285 -13685 38330 -13565
rect 38450 -13685 38495 -13565
rect 38615 -13685 38670 -13565
rect 38790 -13685 38835 -13565
rect 38955 -13685 39000 -13565
rect 39120 -13685 39165 -13565
rect 39285 -13685 39340 -13565
rect 39460 -13685 39505 -13565
rect 39625 -13685 39670 -13565
rect 39790 -13685 39835 -13565
rect 39955 -13685 40010 -13565
rect 40130 -13685 40175 -13565
rect 40295 -13685 40340 -13565
rect 40460 -13685 40505 -13565
rect 40625 -13685 40680 -13565
rect 40800 -13685 40845 -13565
rect 40965 -13685 41010 -13565
rect 41130 -13685 41175 -13565
rect 41295 -13685 41350 -13565
rect 41470 -13685 41515 -13565
rect 41635 -13685 41680 -13565
rect 41800 -13685 41845 -13565
rect 41965 -13685 41975 -13565
rect 36475 -13730 41975 -13685
rect 36475 -13850 36485 -13730
rect 36605 -13850 36660 -13730
rect 36780 -13850 36825 -13730
rect 36945 -13850 36990 -13730
rect 37110 -13850 37155 -13730
rect 37275 -13850 37330 -13730
rect 37450 -13850 37495 -13730
rect 37615 -13850 37660 -13730
rect 37780 -13850 37825 -13730
rect 37945 -13850 38000 -13730
rect 38120 -13850 38165 -13730
rect 38285 -13850 38330 -13730
rect 38450 -13850 38495 -13730
rect 38615 -13850 38670 -13730
rect 38790 -13850 38835 -13730
rect 38955 -13850 39000 -13730
rect 39120 -13850 39165 -13730
rect 39285 -13850 39340 -13730
rect 39460 -13850 39505 -13730
rect 39625 -13850 39670 -13730
rect 39790 -13850 39835 -13730
rect 39955 -13850 40010 -13730
rect 40130 -13850 40175 -13730
rect 40295 -13850 40340 -13730
rect 40460 -13850 40505 -13730
rect 40625 -13850 40680 -13730
rect 40800 -13850 40845 -13730
rect 40965 -13850 41010 -13730
rect 41130 -13850 41175 -13730
rect 41295 -13850 41350 -13730
rect 41470 -13850 41515 -13730
rect 41635 -13850 41680 -13730
rect 41800 -13850 41845 -13730
rect 41965 -13850 41975 -13730
rect 36475 -13895 41975 -13850
rect 36475 -14015 36485 -13895
rect 36605 -14015 36660 -13895
rect 36780 -14015 36825 -13895
rect 36945 -14015 36990 -13895
rect 37110 -14015 37155 -13895
rect 37275 -14015 37330 -13895
rect 37450 -14015 37495 -13895
rect 37615 -14015 37660 -13895
rect 37780 -14015 37825 -13895
rect 37945 -14015 38000 -13895
rect 38120 -14015 38165 -13895
rect 38285 -14015 38330 -13895
rect 38450 -14015 38495 -13895
rect 38615 -14015 38670 -13895
rect 38790 -14015 38835 -13895
rect 38955 -14015 39000 -13895
rect 39120 -14015 39165 -13895
rect 39285 -14015 39340 -13895
rect 39460 -14015 39505 -13895
rect 39625 -14015 39670 -13895
rect 39790 -14015 39835 -13895
rect 39955 -14015 40010 -13895
rect 40130 -14015 40175 -13895
rect 40295 -14015 40340 -13895
rect 40460 -14015 40505 -13895
rect 40625 -14015 40680 -13895
rect 40800 -14015 40845 -13895
rect 40965 -14015 41010 -13895
rect 41130 -14015 41175 -13895
rect 41295 -14015 41350 -13895
rect 41470 -14015 41515 -13895
rect 41635 -14015 41680 -13895
rect 41800 -14015 41845 -13895
rect 41965 -14015 41975 -13895
rect 36475 -14070 41975 -14015
rect 36475 -14190 36485 -14070
rect 36605 -14190 36660 -14070
rect 36780 -14190 36825 -14070
rect 36945 -14190 36990 -14070
rect 37110 -14190 37155 -14070
rect 37275 -14190 37330 -14070
rect 37450 -14190 37495 -14070
rect 37615 -14190 37660 -14070
rect 37780 -14190 37825 -14070
rect 37945 -14190 38000 -14070
rect 38120 -14190 38165 -14070
rect 38285 -14190 38330 -14070
rect 38450 -14190 38495 -14070
rect 38615 -14190 38670 -14070
rect 38790 -14190 38835 -14070
rect 38955 -14190 39000 -14070
rect 39120 -14190 39165 -14070
rect 39285 -14190 39340 -14070
rect 39460 -14190 39505 -14070
rect 39625 -14190 39670 -14070
rect 39790 -14190 39835 -14070
rect 39955 -14190 40010 -14070
rect 40130 -14190 40175 -14070
rect 40295 -14190 40340 -14070
rect 40460 -14190 40505 -14070
rect 40625 -14190 40680 -14070
rect 40800 -14190 40845 -14070
rect 40965 -14190 41010 -14070
rect 41130 -14190 41175 -14070
rect 41295 -14190 41350 -14070
rect 41470 -14190 41515 -14070
rect 41635 -14190 41680 -14070
rect 41800 -14190 41845 -14070
rect 41965 -14190 41975 -14070
rect 36475 -14235 41975 -14190
rect 36475 -14355 36485 -14235
rect 36605 -14355 36660 -14235
rect 36780 -14355 36825 -14235
rect 36945 -14355 36990 -14235
rect 37110 -14355 37155 -14235
rect 37275 -14355 37330 -14235
rect 37450 -14355 37495 -14235
rect 37615 -14355 37660 -14235
rect 37780 -14355 37825 -14235
rect 37945 -14355 38000 -14235
rect 38120 -14355 38165 -14235
rect 38285 -14355 38330 -14235
rect 38450 -14355 38495 -14235
rect 38615 -14355 38670 -14235
rect 38790 -14355 38835 -14235
rect 38955 -14355 39000 -14235
rect 39120 -14355 39165 -14235
rect 39285 -14355 39340 -14235
rect 39460 -14355 39505 -14235
rect 39625 -14355 39670 -14235
rect 39790 -14355 39835 -14235
rect 39955 -14355 40010 -14235
rect 40130 -14355 40175 -14235
rect 40295 -14355 40340 -14235
rect 40460 -14355 40505 -14235
rect 40625 -14355 40680 -14235
rect 40800 -14355 40845 -14235
rect 40965 -14355 41010 -14235
rect 41130 -14355 41175 -14235
rect 41295 -14355 41350 -14235
rect 41470 -14355 41515 -14235
rect 41635 -14355 41680 -14235
rect 41800 -14355 41845 -14235
rect 41965 -14355 41975 -14235
rect 36475 -14400 41975 -14355
rect 36475 -14520 36485 -14400
rect 36605 -14520 36660 -14400
rect 36780 -14520 36825 -14400
rect 36945 -14520 36990 -14400
rect 37110 -14520 37155 -14400
rect 37275 -14520 37330 -14400
rect 37450 -14520 37495 -14400
rect 37615 -14520 37660 -14400
rect 37780 -14520 37825 -14400
rect 37945 -14520 38000 -14400
rect 38120 -14520 38165 -14400
rect 38285 -14520 38330 -14400
rect 38450 -14520 38495 -14400
rect 38615 -14520 38670 -14400
rect 38790 -14520 38835 -14400
rect 38955 -14520 39000 -14400
rect 39120 -14520 39165 -14400
rect 39285 -14520 39340 -14400
rect 39460 -14520 39505 -14400
rect 39625 -14520 39670 -14400
rect 39790 -14520 39835 -14400
rect 39955 -14520 40010 -14400
rect 40130 -14520 40175 -14400
rect 40295 -14520 40340 -14400
rect 40460 -14520 40505 -14400
rect 40625 -14520 40680 -14400
rect 40800 -14520 40845 -14400
rect 40965 -14520 41010 -14400
rect 41130 -14520 41175 -14400
rect 41295 -14520 41350 -14400
rect 41470 -14520 41515 -14400
rect 41635 -14520 41680 -14400
rect 41800 -14520 41845 -14400
rect 41965 -14520 41975 -14400
rect 36475 -14565 41975 -14520
rect 36475 -14685 36485 -14565
rect 36605 -14685 36660 -14565
rect 36780 -14685 36825 -14565
rect 36945 -14685 36990 -14565
rect 37110 -14685 37155 -14565
rect 37275 -14685 37330 -14565
rect 37450 -14685 37495 -14565
rect 37615 -14685 37660 -14565
rect 37780 -14685 37825 -14565
rect 37945 -14685 38000 -14565
rect 38120 -14685 38165 -14565
rect 38285 -14685 38330 -14565
rect 38450 -14685 38495 -14565
rect 38615 -14685 38670 -14565
rect 38790 -14685 38835 -14565
rect 38955 -14685 39000 -14565
rect 39120 -14685 39165 -14565
rect 39285 -14685 39340 -14565
rect 39460 -14685 39505 -14565
rect 39625 -14685 39670 -14565
rect 39790 -14685 39835 -14565
rect 39955 -14685 40010 -14565
rect 40130 -14685 40175 -14565
rect 40295 -14685 40340 -14565
rect 40460 -14685 40505 -14565
rect 40625 -14685 40680 -14565
rect 40800 -14685 40845 -14565
rect 40965 -14685 41010 -14565
rect 41130 -14685 41175 -14565
rect 41295 -14685 41350 -14565
rect 41470 -14685 41515 -14565
rect 41635 -14685 41680 -14565
rect 41800 -14685 41845 -14565
rect 41965 -14685 41975 -14565
rect 36475 -14740 41975 -14685
rect 36475 -14860 36485 -14740
rect 36605 -14860 36660 -14740
rect 36780 -14860 36825 -14740
rect 36945 -14860 36990 -14740
rect 37110 -14860 37155 -14740
rect 37275 -14860 37330 -14740
rect 37450 -14860 37495 -14740
rect 37615 -14860 37660 -14740
rect 37780 -14860 37825 -14740
rect 37945 -14860 38000 -14740
rect 38120 -14860 38165 -14740
rect 38285 -14860 38330 -14740
rect 38450 -14860 38495 -14740
rect 38615 -14860 38670 -14740
rect 38790 -14860 38835 -14740
rect 38955 -14860 39000 -14740
rect 39120 -14860 39165 -14740
rect 39285 -14860 39340 -14740
rect 39460 -14860 39505 -14740
rect 39625 -14860 39670 -14740
rect 39790 -14860 39835 -14740
rect 39955 -14860 40010 -14740
rect 40130 -14860 40175 -14740
rect 40295 -14860 40340 -14740
rect 40460 -14860 40505 -14740
rect 40625 -14860 40680 -14740
rect 40800 -14860 40845 -14740
rect 40965 -14860 41010 -14740
rect 41130 -14860 41175 -14740
rect 41295 -14860 41350 -14740
rect 41470 -14860 41515 -14740
rect 41635 -14860 41680 -14740
rect 41800 -14860 41845 -14740
rect 41965 -14860 41975 -14740
rect 36475 -14905 41975 -14860
rect 36475 -15025 36485 -14905
rect 36605 -15025 36660 -14905
rect 36780 -15025 36825 -14905
rect 36945 -15025 36990 -14905
rect 37110 -15025 37155 -14905
rect 37275 -15025 37330 -14905
rect 37450 -15025 37495 -14905
rect 37615 -15025 37660 -14905
rect 37780 -15025 37825 -14905
rect 37945 -15025 38000 -14905
rect 38120 -15025 38165 -14905
rect 38285 -15025 38330 -14905
rect 38450 -15025 38495 -14905
rect 38615 -15025 38670 -14905
rect 38790 -15025 38835 -14905
rect 38955 -15025 39000 -14905
rect 39120 -15025 39165 -14905
rect 39285 -15025 39340 -14905
rect 39460 -15025 39505 -14905
rect 39625 -15025 39670 -14905
rect 39790 -15025 39835 -14905
rect 39955 -15025 40010 -14905
rect 40130 -15025 40175 -14905
rect 40295 -15025 40340 -14905
rect 40460 -15025 40505 -14905
rect 40625 -15025 40680 -14905
rect 40800 -15025 40845 -14905
rect 40965 -15025 41010 -14905
rect 41130 -15025 41175 -14905
rect 41295 -15025 41350 -14905
rect 41470 -15025 41515 -14905
rect 41635 -15025 41680 -14905
rect 41800 -15025 41845 -14905
rect 41965 -15025 41975 -14905
rect 36475 -15070 41975 -15025
rect 36475 -15190 36485 -15070
rect 36605 -15190 36660 -15070
rect 36780 -15190 36825 -15070
rect 36945 -15190 36990 -15070
rect 37110 -15190 37155 -15070
rect 37275 -15190 37330 -15070
rect 37450 -15190 37495 -15070
rect 37615 -15190 37660 -15070
rect 37780 -15190 37825 -15070
rect 37945 -15190 38000 -15070
rect 38120 -15190 38165 -15070
rect 38285 -15190 38330 -15070
rect 38450 -15190 38495 -15070
rect 38615 -15190 38670 -15070
rect 38790 -15190 38835 -15070
rect 38955 -15190 39000 -15070
rect 39120 -15190 39165 -15070
rect 39285 -15190 39340 -15070
rect 39460 -15190 39505 -15070
rect 39625 -15190 39670 -15070
rect 39790 -15190 39835 -15070
rect 39955 -15190 40010 -15070
rect 40130 -15190 40175 -15070
rect 40295 -15190 40340 -15070
rect 40460 -15190 40505 -15070
rect 40625 -15190 40680 -15070
rect 40800 -15190 40845 -15070
rect 40965 -15190 41010 -15070
rect 41130 -15190 41175 -15070
rect 41295 -15190 41350 -15070
rect 41470 -15190 41515 -15070
rect 41635 -15190 41680 -15070
rect 41800 -15190 41845 -15070
rect 41965 -15190 41975 -15070
rect 36475 -15235 41975 -15190
rect 36475 -15355 36485 -15235
rect 36605 -15355 36660 -15235
rect 36780 -15355 36825 -15235
rect 36945 -15355 36990 -15235
rect 37110 -15355 37155 -15235
rect 37275 -15355 37330 -15235
rect 37450 -15355 37495 -15235
rect 37615 -15355 37660 -15235
rect 37780 -15355 37825 -15235
rect 37945 -15355 38000 -15235
rect 38120 -15355 38165 -15235
rect 38285 -15355 38330 -15235
rect 38450 -15355 38495 -15235
rect 38615 -15355 38670 -15235
rect 38790 -15355 38835 -15235
rect 38955 -15355 39000 -15235
rect 39120 -15355 39165 -15235
rect 39285 -15355 39340 -15235
rect 39460 -15355 39505 -15235
rect 39625 -15355 39670 -15235
rect 39790 -15355 39835 -15235
rect 39955 -15355 40010 -15235
rect 40130 -15355 40175 -15235
rect 40295 -15355 40340 -15235
rect 40460 -15355 40505 -15235
rect 40625 -15355 40680 -15235
rect 40800 -15355 40845 -15235
rect 40965 -15355 41010 -15235
rect 41130 -15355 41175 -15235
rect 41295 -15355 41350 -15235
rect 41470 -15355 41515 -15235
rect 41635 -15355 41680 -15235
rect 41800 -15355 41845 -15235
rect 41965 -15355 41975 -15235
rect 36475 -15410 41975 -15355
rect 36475 -15530 36485 -15410
rect 36605 -15530 36660 -15410
rect 36780 -15530 36825 -15410
rect 36945 -15530 36990 -15410
rect 37110 -15530 37155 -15410
rect 37275 -15530 37330 -15410
rect 37450 -15530 37495 -15410
rect 37615 -15530 37660 -15410
rect 37780 -15530 37825 -15410
rect 37945 -15530 38000 -15410
rect 38120 -15530 38165 -15410
rect 38285 -15530 38330 -15410
rect 38450 -15530 38495 -15410
rect 38615 -15530 38670 -15410
rect 38790 -15530 38835 -15410
rect 38955 -15530 39000 -15410
rect 39120 -15530 39165 -15410
rect 39285 -15530 39340 -15410
rect 39460 -15530 39505 -15410
rect 39625 -15530 39670 -15410
rect 39790 -15530 39835 -15410
rect 39955 -15530 40010 -15410
rect 40130 -15530 40175 -15410
rect 40295 -15530 40340 -15410
rect 40460 -15530 40505 -15410
rect 40625 -15530 40680 -15410
rect 40800 -15530 40845 -15410
rect 40965 -15530 41010 -15410
rect 41130 -15530 41175 -15410
rect 41295 -15530 41350 -15410
rect 41470 -15530 41515 -15410
rect 41635 -15530 41680 -15410
rect 41800 -15530 41845 -15410
rect 41965 -15530 41975 -15410
rect 36475 -15540 41975 -15530
rect 42165 -10050 47665 -10040
rect 42165 -10170 42175 -10050
rect 42295 -10170 42350 -10050
rect 42470 -10170 42515 -10050
rect 42635 -10170 42680 -10050
rect 42800 -10170 42845 -10050
rect 42965 -10170 43020 -10050
rect 43140 -10170 43185 -10050
rect 43305 -10170 43350 -10050
rect 43470 -10170 43515 -10050
rect 43635 -10170 43690 -10050
rect 43810 -10170 43855 -10050
rect 43975 -10170 44020 -10050
rect 44140 -10170 44185 -10050
rect 44305 -10170 44360 -10050
rect 44480 -10170 44525 -10050
rect 44645 -10170 44690 -10050
rect 44810 -10170 44855 -10050
rect 44975 -10170 45030 -10050
rect 45150 -10170 45195 -10050
rect 45315 -10170 45360 -10050
rect 45480 -10170 45525 -10050
rect 45645 -10170 45700 -10050
rect 45820 -10170 45865 -10050
rect 45985 -10170 46030 -10050
rect 46150 -10170 46195 -10050
rect 46315 -10170 46370 -10050
rect 46490 -10170 46535 -10050
rect 46655 -10170 46700 -10050
rect 46820 -10170 46865 -10050
rect 46985 -10170 47040 -10050
rect 47160 -10170 47205 -10050
rect 47325 -10170 47370 -10050
rect 47490 -10170 47535 -10050
rect 47655 -10170 47665 -10050
rect 42165 -10215 47665 -10170
rect 42165 -10335 42175 -10215
rect 42295 -10335 42350 -10215
rect 42470 -10335 42515 -10215
rect 42635 -10335 42680 -10215
rect 42800 -10335 42845 -10215
rect 42965 -10335 43020 -10215
rect 43140 -10335 43185 -10215
rect 43305 -10335 43350 -10215
rect 43470 -10335 43515 -10215
rect 43635 -10335 43690 -10215
rect 43810 -10335 43855 -10215
rect 43975 -10335 44020 -10215
rect 44140 -10335 44185 -10215
rect 44305 -10335 44360 -10215
rect 44480 -10335 44525 -10215
rect 44645 -10335 44690 -10215
rect 44810 -10335 44855 -10215
rect 44975 -10335 45030 -10215
rect 45150 -10335 45195 -10215
rect 45315 -10335 45360 -10215
rect 45480 -10335 45525 -10215
rect 45645 -10335 45700 -10215
rect 45820 -10335 45865 -10215
rect 45985 -10335 46030 -10215
rect 46150 -10335 46195 -10215
rect 46315 -10335 46370 -10215
rect 46490 -10335 46535 -10215
rect 46655 -10335 46700 -10215
rect 46820 -10335 46865 -10215
rect 46985 -10335 47040 -10215
rect 47160 -10335 47205 -10215
rect 47325 -10335 47370 -10215
rect 47490 -10335 47535 -10215
rect 47655 -10335 47665 -10215
rect 42165 -10380 47665 -10335
rect 42165 -10500 42175 -10380
rect 42295 -10500 42350 -10380
rect 42470 -10500 42515 -10380
rect 42635 -10500 42680 -10380
rect 42800 -10500 42845 -10380
rect 42965 -10500 43020 -10380
rect 43140 -10500 43185 -10380
rect 43305 -10500 43350 -10380
rect 43470 -10500 43515 -10380
rect 43635 -10500 43690 -10380
rect 43810 -10500 43855 -10380
rect 43975 -10500 44020 -10380
rect 44140 -10500 44185 -10380
rect 44305 -10500 44360 -10380
rect 44480 -10500 44525 -10380
rect 44645 -10500 44690 -10380
rect 44810 -10500 44855 -10380
rect 44975 -10500 45030 -10380
rect 45150 -10500 45195 -10380
rect 45315 -10500 45360 -10380
rect 45480 -10500 45525 -10380
rect 45645 -10500 45700 -10380
rect 45820 -10500 45865 -10380
rect 45985 -10500 46030 -10380
rect 46150 -10500 46195 -10380
rect 46315 -10500 46370 -10380
rect 46490 -10500 46535 -10380
rect 46655 -10500 46700 -10380
rect 46820 -10500 46865 -10380
rect 46985 -10500 47040 -10380
rect 47160 -10500 47205 -10380
rect 47325 -10500 47370 -10380
rect 47490 -10500 47535 -10380
rect 47655 -10500 47665 -10380
rect 42165 -10545 47665 -10500
rect 42165 -10665 42175 -10545
rect 42295 -10665 42350 -10545
rect 42470 -10665 42515 -10545
rect 42635 -10665 42680 -10545
rect 42800 -10665 42845 -10545
rect 42965 -10665 43020 -10545
rect 43140 -10665 43185 -10545
rect 43305 -10665 43350 -10545
rect 43470 -10665 43515 -10545
rect 43635 -10665 43690 -10545
rect 43810 -10665 43855 -10545
rect 43975 -10665 44020 -10545
rect 44140 -10665 44185 -10545
rect 44305 -10665 44360 -10545
rect 44480 -10665 44525 -10545
rect 44645 -10665 44690 -10545
rect 44810 -10665 44855 -10545
rect 44975 -10665 45030 -10545
rect 45150 -10665 45195 -10545
rect 45315 -10665 45360 -10545
rect 45480 -10665 45525 -10545
rect 45645 -10665 45700 -10545
rect 45820 -10665 45865 -10545
rect 45985 -10665 46030 -10545
rect 46150 -10665 46195 -10545
rect 46315 -10665 46370 -10545
rect 46490 -10665 46535 -10545
rect 46655 -10665 46700 -10545
rect 46820 -10665 46865 -10545
rect 46985 -10665 47040 -10545
rect 47160 -10665 47205 -10545
rect 47325 -10665 47370 -10545
rect 47490 -10665 47535 -10545
rect 47655 -10665 47665 -10545
rect 42165 -10720 47665 -10665
rect 42165 -10840 42175 -10720
rect 42295 -10840 42350 -10720
rect 42470 -10840 42515 -10720
rect 42635 -10840 42680 -10720
rect 42800 -10840 42845 -10720
rect 42965 -10840 43020 -10720
rect 43140 -10840 43185 -10720
rect 43305 -10840 43350 -10720
rect 43470 -10840 43515 -10720
rect 43635 -10840 43690 -10720
rect 43810 -10840 43855 -10720
rect 43975 -10840 44020 -10720
rect 44140 -10840 44185 -10720
rect 44305 -10840 44360 -10720
rect 44480 -10840 44525 -10720
rect 44645 -10840 44690 -10720
rect 44810 -10840 44855 -10720
rect 44975 -10840 45030 -10720
rect 45150 -10840 45195 -10720
rect 45315 -10840 45360 -10720
rect 45480 -10840 45525 -10720
rect 45645 -10840 45700 -10720
rect 45820 -10840 45865 -10720
rect 45985 -10840 46030 -10720
rect 46150 -10840 46195 -10720
rect 46315 -10840 46370 -10720
rect 46490 -10840 46535 -10720
rect 46655 -10840 46700 -10720
rect 46820 -10840 46865 -10720
rect 46985 -10840 47040 -10720
rect 47160 -10840 47205 -10720
rect 47325 -10840 47370 -10720
rect 47490 -10840 47535 -10720
rect 47655 -10840 47665 -10720
rect 42165 -10885 47665 -10840
rect 42165 -11005 42175 -10885
rect 42295 -11005 42350 -10885
rect 42470 -11005 42515 -10885
rect 42635 -11005 42680 -10885
rect 42800 -11005 42845 -10885
rect 42965 -11005 43020 -10885
rect 43140 -11005 43185 -10885
rect 43305 -11005 43350 -10885
rect 43470 -11005 43515 -10885
rect 43635 -11005 43690 -10885
rect 43810 -11005 43855 -10885
rect 43975 -11005 44020 -10885
rect 44140 -11005 44185 -10885
rect 44305 -11005 44360 -10885
rect 44480 -11005 44525 -10885
rect 44645 -11005 44690 -10885
rect 44810 -11005 44855 -10885
rect 44975 -11005 45030 -10885
rect 45150 -11005 45195 -10885
rect 45315 -11005 45360 -10885
rect 45480 -11005 45525 -10885
rect 45645 -11005 45700 -10885
rect 45820 -11005 45865 -10885
rect 45985 -11005 46030 -10885
rect 46150 -11005 46195 -10885
rect 46315 -11005 46370 -10885
rect 46490 -11005 46535 -10885
rect 46655 -11005 46700 -10885
rect 46820 -11005 46865 -10885
rect 46985 -11005 47040 -10885
rect 47160 -11005 47205 -10885
rect 47325 -11005 47370 -10885
rect 47490 -11005 47535 -10885
rect 47655 -11005 47665 -10885
rect 42165 -11050 47665 -11005
rect 42165 -11170 42175 -11050
rect 42295 -11170 42350 -11050
rect 42470 -11170 42515 -11050
rect 42635 -11170 42680 -11050
rect 42800 -11170 42845 -11050
rect 42965 -11170 43020 -11050
rect 43140 -11170 43185 -11050
rect 43305 -11170 43350 -11050
rect 43470 -11170 43515 -11050
rect 43635 -11170 43690 -11050
rect 43810 -11170 43855 -11050
rect 43975 -11170 44020 -11050
rect 44140 -11170 44185 -11050
rect 44305 -11170 44360 -11050
rect 44480 -11170 44525 -11050
rect 44645 -11170 44690 -11050
rect 44810 -11170 44855 -11050
rect 44975 -11170 45030 -11050
rect 45150 -11170 45195 -11050
rect 45315 -11170 45360 -11050
rect 45480 -11170 45525 -11050
rect 45645 -11170 45700 -11050
rect 45820 -11170 45865 -11050
rect 45985 -11170 46030 -11050
rect 46150 -11170 46195 -11050
rect 46315 -11170 46370 -11050
rect 46490 -11170 46535 -11050
rect 46655 -11170 46700 -11050
rect 46820 -11170 46865 -11050
rect 46985 -11170 47040 -11050
rect 47160 -11170 47205 -11050
rect 47325 -11170 47370 -11050
rect 47490 -11170 47535 -11050
rect 47655 -11170 47665 -11050
rect 42165 -11215 47665 -11170
rect 42165 -11335 42175 -11215
rect 42295 -11335 42350 -11215
rect 42470 -11335 42515 -11215
rect 42635 -11335 42680 -11215
rect 42800 -11335 42845 -11215
rect 42965 -11335 43020 -11215
rect 43140 -11335 43185 -11215
rect 43305 -11335 43350 -11215
rect 43470 -11335 43515 -11215
rect 43635 -11335 43690 -11215
rect 43810 -11335 43855 -11215
rect 43975 -11335 44020 -11215
rect 44140 -11335 44185 -11215
rect 44305 -11335 44360 -11215
rect 44480 -11335 44525 -11215
rect 44645 -11335 44690 -11215
rect 44810 -11335 44855 -11215
rect 44975 -11335 45030 -11215
rect 45150 -11335 45195 -11215
rect 45315 -11335 45360 -11215
rect 45480 -11335 45525 -11215
rect 45645 -11335 45700 -11215
rect 45820 -11335 45865 -11215
rect 45985 -11335 46030 -11215
rect 46150 -11335 46195 -11215
rect 46315 -11335 46370 -11215
rect 46490 -11335 46535 -11215
rect 46655 -11335 46700 -11215
rect 46820 -11335 46865 -11215
rect 46985 -11335 47040 -11215
rect 47160 -11335 47205 -11215
rect 47325 -11335 47370 -11215
rect 47490 -11335 47535 -11215
rect 47655 -11335 47665 -11215
rect 42165 -11390 47665 -11335
rect 42165 -11510 42175 -11390
rect 42295 -11510 42350 -11390
rect 42470 -11510 42515 -11390
rect 42635 -11510 42680 -11390
rect 42800 -11510 42845 -11390
rect 42965 -11510 43020 -11390
rect 43140 -11510 43185 -11390
rect 43305 -11510 43350 -11390
rect 43470 -11510 43515 -11390
rect 43635 -11510 43690 -11390
rect 43810 -11510 43855 -11390
rect 43975 -11510 44020 -11390
rect 44140 -11510 44185 -11390
rect 44305 -11510 44360 -11390
rect 44480 -11510 44525 -11390
rect 44645 -11510 44690 -11390
rect 44810 -11510 44855 -11390
rect 44975 -11510 45030 -11390
rect 45150 -11510 45195 -11390
rect 45315 -11510 45360 -11390
rect 45480 -11510 45525 -11390
rect 45645 -11510 45700 -11390
rect 45820 -11510 45865 -11390
rect 45985 -11510 46030 -11390
rect 46150 -11510 46195 -11390
rect 46315 -11510 46370 -11390
rect 46490 -11510 46535 -11390
rect 46655 -11510 46700 -11390
rect 46820 -11510 46865 -11390
rect 46985 -11510 47040 -11390
rect 47160 -11510 47205 -11390
rect 47325 -11510 47370 -11390
rect 47490 -11510 47535 -11390
rect 47655 -11510 47665 -11390
rect 42165 -11555 47665 -11510
rect 42165 -11675 42175 -11555
rect 42295 -11675 42350 -11555
rect 42470 -11675 42515 -11555
rect 42635 -11675 42680 -11555
rect 42800 -11675 42845 -11555
rect 42965 -11675 43020 -11555
rect 43140 -11675 43185 -11555
rect 43305 -11675 43350 -11555
rect 43470 -11675 43515 -11555
rect 43635 -11675 43690 -11555
rect 43810 -11675 43855 -11555
rect 43975 -11675 44020 -11555
rect 44140 -11675 44185 -11555
rect 44305 -11675 44360 -11555
rect 44480 -11675 44525 -11555
rect 44645 -11675 44690 -11555
rect 44810 -11675 44855 -11555
rect 44975 -11675 45030 -11555
rect 45150 -11675 45195 -11555
rect 45315 -11675 45360 -11555
rect 45480 -11675 45525 -11555
rect 45645 -11675 45700 -11555
rect 45820 -11675 45865 -11555
rect 45985 -11675 46030 -11555
rect 46150 -11675 46195 -11555
rect 46315 -11675 46370 -11555
rect 46490 -11675 46535 -11555
rect 46655 -11675 46700 -11555
rect 46820 -11675 46865 -11555
rect 46985 -11675 47040 -11555
rect 47160 -11675 47205 -11555
rect 47325 -11675 47370 -11555
rect 47490 -11675 47535 -11555
rect 47655 -11675 47665 -11555
rect 42165 -11720 47665 -11675
rect 42165 -11840 42175 -11720
rect 42295 -11840 42350 -11720
rect 42470 -11840 42515 -11720
rect 42635 -11840 42680 -11720
rect 42800 -11840 42845 -11720
rect 42965 -11840 43020 -11720
rect 43140 -11840 43185 -11720
rect 43305 -11840 43350 -11720
rect 43470 -11840 43515 -11720
rect 43635 -11840 43690 -11720
rect 43810 -11840 43855 -11720
rect 43975 -11840 44020 -11720
rect 44140 -11840 44185 -11720
rect 44305 -11840 44360 -11720
rect 44480 -11840 44525 -11720
rect 44645 -11840 44690 -11720
rect 44810 -11840 44855 -11720
rect 44975 -11840 45030 -11720
rect 45150 -11840 45195 -11720
rect 45315 -11840 45360 -11720
rect 45480 -11840 45525 -11720
rect 45645 -11840 45700 -11720
rect 45820 -11840 45865 -11720
rect 45985 -11840 46030 -11720
rect 46150 -11840 46195 -11720
rect 46315 -11840 46370 -11720
rect 46490 -11840 46535 -11720
rect 46655 -11840 46700 -11720
rect 46820 -11840 46865 -11720
rect 46985 -11840 47040 -11720
rect 47160 -11840 47205 -11720
rect 47325 -11840 47370 -11720
rect 47490 -11840 47535 -11720
rect 47655 -11840 47665 -11720
rect 42165 -11885 47665 -11840
rect 42165 -12005 42175 -11885
rect 42295 -12005 42350 -11885
rect 42470 -12005 42515 -11885
rect 42635 -12005 42680 -11885
rect 42800 -12005 42845 -11885
rect 42965 -12005 43020 -11885
rect 43140 -12005 43185 -11885
rect 43305 -12005 43350 -11885
rect 43470 -12005 43515 -11885
rect 43635 -12005 43690 -11885
rect 43810 -12005 43855 -11885
rect 43975 -12005 44020 -11885
rect 44140 -12005 44185 -11885
rect 44305 -12005 44360 -11885
rect 44480 -12005 44525 -11885
rect 44645 -12005 44690 -11885
rect 44810 -12005 44855 -11885
rect 44975 -12005 45030 -11885
rect 45150 -12005 45195 -11885
rect 45315 -12005 45360 -11885
rect 45480 -12005 45525 -11885
rect 45645 -12005 45700 -11885
rect 45820 -12005 45865 -11885
rect 45985 -12005 46030 -11885
rect 46150 -12005 46195 -11885
rect 46315 -12005 46370 -11885
rect 46490 -12005 46535 -11885
rect 46655 -12005 46700 -11885
rect 46820 -12005 46865 -11885
rect 46985 -12005 47040 -11885
rect 47160 -12005 47205 -11885
rect 47325 -12005 47370 -11885
rect 47490 -12005 47535 -11885
rect 47655 -12005 47665 -11885
rect 42165 -12060 47665 -12005
rect 42165 -12180 42175 -12060
rect 42295 -12180 42350 -12060
rect 42470 -12180 42515 -12060
rect 42635 -12180 42680 -12060
rect 42800 -12180 42845 -12060
rect 42965 -12180 43020 -12060
rect 43140 -12180 43185 -12060
rect 43305 -12180 43350 -12060
rect 43470 -12180 43515 -12060
rect 43635 -12180 43690 -12060
rect 43810 -12180 43855 -12060
rect 43975 -12180 44020 -12060
rect 44140 -12180 44185 -12060
rect 44305 -12180 44360 -12060
rect 44480 -12180 44525 -12060
rect 44645 -12180 44690 -12060
rect 44810 -12180 44855 -12060
rect 44975 -12180 45030 -12060
rect 45150 -12180 45195 -12060
rect 45315 -12180 45360 -12060
rect 45480 -12180 45525 -12060
rect 45645 -12180 45700 -12060
rect 45820 -12180 45865 -12060
rect 45985 -12180 46030 -12060
rect 46150 -12180 46195 -12060
rect 46315 -12180 46370 -12060
rect 46490 -12180 46535 -12060
rect 46655 -12180 46700 -12060
rect 46820 -12180 46865 -12060
rect 46985 -12180 47040 -12060
rect 47160 -12180 47205 -12060
rect 47325 -12180 47370 -12060
rect 47490 -12180 47535 -12060
rect 47655 -12180 47665 -12060
rect 42165 -12225 47665 -12180
rect 42165 -12345 42175 -12225
rect 42295 -12345 42350 -12225
rect 42470 -12345 42515 -12225
rect 42635 -12345 42680 -12225
rect 42800 -12345 42845 -12225
rect 42965 -12345 43020 -12225
rect 43140 -12345 43185 -12225
rect 43305 -12345 43350 -12225
rect 43470 -12345 43515 -12225
rect 43635 -12345 43690 -12225
rect 43810 -12345 43855 -12225
rect 43975 -12345 44020 -12225
rect 44140 -12345 44185 -12225
rect 44305 -12345 44360 -12225
rect 44480 -12345 44525 -12225
rect 44645 -12345 44690 -12225
rect 44810 -12345 44855 -12225
rect 44975 -12345 45030 -12225
rect 45150 -12345 45195 -12225
rect 45315 -12345 45360 -12225
rect 45480 -12345 45525 -12225
rect 45645 -12345 45700 -12225
rect 45820 -12345 45865 -12225
rect 45985 -12345 46030 -12225
rect 46150 -12345 46195 -12225
rect 46315 -12345 46370 -12225
rect 46490 -12345 46535 -12225
rect 46655 -12345 46700 -12225
rect 46820 -12345 46865 -12225
rect 46985 -12345 47040 -12225
rect 47160 -12345 47205 -12225
rect 47325 -12345 47370 -12225
rect 47490 -12345 47535 -12225
rect 47655 -12345 47665 -12225
rect 42165 -12390 47665 -12345
rect 42165 -12510 42175 -12390
rect 42295 -12510 42350 -12390
rect 42470 -12510 42515 -12390
rect 42635 -12510 42680 -12390
rect 42800 -12510 42845 -12390
rect 42965 -12510 43020 -12390
rect 43140 -12510 43185 -12390
rect 43305 -12510 43350 -12390
rect 43470 -12510 43515 -12390
rect 43635 -12510 43690 -12390
rect 43810 -12510 43855 -12390
rect 43975 -12510 44020 -12390
rect 44140 -12510 44185 -12390
rect 44305 -12510 44360 -12390
rect 44480 -12510 44525 -12390
rect 44645 -12510 44690 -12390
rect 44810 -12510 44855 -12390
rect 44975 -12510 45030 -12390
rect 45150 -12510 45195 -12390
rect 45315 -12510 45360 -12390
rect 45480 -12510 45525 -12390
rect 45645 -12510 45700 -12390
rect 45820 -12510 45865 -12390
rect 45985 -12510 46030 -12390
rect 46150 -12510 46195 -12390
rect 46315 -12510 46370 -12390
rect 46490 -12510 46535 -12390
rect 46655 -12510 46700 -12390
rect 46820 -12510 46865 -12390
rect 46985 -12510 47040 -12390
rect 47160 -12510 47205 -12390
rect 47325 -12510 47370 -12390
rect 47490 -12510 47535 -12390
rect 47655 -12510 47665 -12390
rect 42165 -12555 47665 -12510
rect 42165 -12675 42175 -12555
rect 42295 -12675 42350 -12555
rect 42470 -12675 42515 -12555
rect 42635 -12675 42680 -12555
rect 42800 -12675 42845 -12555
rect 42965 -12675 43020 -12555
rect 43140 -12675 43185 -12555
rect 43305 -12675 43350 -12555
rect 43470 -12675 43515 -12555
rect 43635 -12675 43690 -12555
rect 43810 -12675 43855 -12555
rect 43975 -12675 44020 -12555
rect 44140 -12675 44185 -12555
rect 44305 -12675 44360 -12555
rect 44480 -12675 44525 -12555
rect 44645 -12675 44690 -12555
rect 44810 -12675 44855 -12555
rect 44975 -12675 45030 -12555
rect 45150 -12675 45195 -12555
rect 45315 -12675 45360 -12555
rect 45480 -12675 45525 -12555
rect 45645 -12675 45700 -12555
rect 45820 -12675 45865 -12555
rect 45985 -12675 46030 -12555
rect 46150 -12675 46195 -12555
rect 46315 -12675 46370 -12555
rect 46490 -12675 46535 -12555
rect 46655 -12675 46700 -12555
rect 46820 -12675 46865 -12555
rect 46985 -12675 47040 -12555
rect 47160 -12675 47205 -12555
rect 47325 -12675 47370 -12555
rect 47490 -12675 47535 -12555
rect 47655 -12675 47665 -12555
rect 42165 -12730 47665 -12675
rect 42165 -12850 42175 -12730
rect 42295 -12850 42350 -12730
rect 42470 -12850 42515 -12730
rect 42635 -12850 42680 -12730
rect 42800 -12850 42845 -12730
rect 42965 -12850 43020 -12730
rect 43140 -12850 43185 -12730
rect 43305 -12850 43350 -12730
rect 43470 -12850 43515 -12730
rect 43635 -12850 43690 -12730
rect 43810 -12850 43855 -12730
rect 43975 -12850 44020 -12730
rect 44140 -12850 44185 -12730
rect 44305 -12850 44360 -12730
rect 44480 -12850 44525 -12730
rect 44645 -12850 44690 -12730
rect 44810 -12850 44855 -12730
rect 44975 -12850 45030 -12730
rect 45150 -12850 45195 -12730
rect 45315 -12850 45360 -12730
rect 45480 -12850 45525 -12730
rect 45645 -12850 45700 -12730
rect 45820 -12850 45865 -12730
rect 45985 -12850 46030 -12730
rect 46150 -12850 46195 -12730
rect 46315 -12850 46370 -12730
rect 46490 -12850 46535 -12730
rect 46655 -12850 46700 -12730
rect 46820 -12850 46865 -12730
rect 46985 -12850 47040 -12730
rect 47160 -12850 47205 -12730
rect 47325 -12850 47370 -12730
rect 47490 -12850 47535 -12730
rect 47655 -12850 47665 -12730
rect 42165 -12895 47665 -12850
rect 42165 -13015 42175 -12895
rect 42295 -13015 42350 -12895
rect 42470 -13015 42515 -12895
rect 42635 -13015 42680 -12895
rect 42800 -13015 42845 -12895
rect 42965 -13015 43020 -12895
rect 43140 -13015 43185 -12895
rect 43305 -13015 43350 -12895
rect 43470 -13015 43515 -12895
rect 43635 -13015 43690 -12895
rect 43810 -13015 43855 -12895
rect 43975 -13015 44020 -12895
rect 44140 -13015 44185 -12895
rect 44305 -13015 44360 -12895
rect 44480 -13015 44525 -12895
rect 44645 -13015 44690 -12895
rect 44810 -13015 44855 -12895
rect 44975 -13015 45030 -12895
rect 45150 -13015 45195 -12895
rect 45315 -13015 45360 -12895
rect 45480 -13015 45525 -12895
rect 45645 -13015 45700 -12895
rect 45820 -13015 45865 -12895
rect 45985 -13015 46030 -12895
rect 46150 -13015 46195 -12895
rect 46315 -13015 46370 -12895
rect 46490 -13015 46535 -12895
rect 46655 -13015 46700 -12895
rect 46820 -13015 46865 -12895
rect 46985 -13015 47040 -12895
rect 47160 -13015 47205 -12895
rect 47325 -13015 47370 -12895
rect 47490 -13015 47535 -12895
rect 47655 -13015 47665 -12895
rect 42165 -13060 47665 -13015
rect 42165 -13180 42175 -13060
rect 42295 -13180 42350 -13060
rect 42470 -13180 42515 -13060
rect 42635 -13180 42680 -13060
rect 42800 -13180 42845 -13060
rect 42965 -13180 43020 -13060
rect 43140 -13180 43185 -13060
rect 43305 -13180 43350 -13060
rect 43470 -13180 43515 -13060
rect 43635 -13180 43690 -13060
rect 43810 -13180 43855 -13060
rect 43975 -13180 44020 -13060
rect 44140 -13180 44185 -13060
rect 44305 -13180 44360 -13060
rect 44480 -13180 44525 -13060
rect 44645 -13180 44690 -13060
rect 44810 -13180 44855 -13060
rect 44975 -13180 45030 -13060
rect 45150 -13180 45195 -13060
rect 45315 -13180 45360 -13060
rect 45480 -13180 45525 -13060
rect 45645 -13180 45700 -13060
rect 45820 -13180 45865 -13060
rect 45985 -13180 46030 -13060
rect 46150 -13180 46195 -13060
rect 46315 -13180 46370 -13060
rect 46490 -13180 46535 -13060
rect 46655 -13180 46700 -13060
rect 46820 -13180 46865 -13060
rect 46985 -13180 47040 -13060
rect 47160 -13180 47205 -13060
rect 47325 -13180 47370 -13060
rect 47490 -13180 47535 -13060
rect 47655 -13180 47665 -13060
rect 42165 -13225 47665 -13180
rect 42165 -13345 42175 -13225
rect 42295 -13345 42350 -13225
rect 42470 -13345 42515 -13225
rect 42635 -13345 42680 -13225
rect 42800 -13345 42845 -13225
rect 42965 -13345 43020 -13225
rect 43140 -13345 43185 -13225
rect 43305 -13345 43350 -13225
rect 43470 -13345 43515 -13225
rect 43635 -13345 43690 -13225
rect 43810 -13345 43855 -13225
rect 43975 -13345 44020 -13225
rect 44140 -13345 44185 -13225
rect 44305 -13345 44360 -13225
rect 44480 -13345 44525 -13225
rect 44645 -13345 44690 -13225
rect 44810 -13345 44855 -13225
rect 44975 -13345 45030 -13225
rect 45150 -13345 45195 -13225
rect 45315 -13345 45360 -13225
rect 45480 -13345 45525 -13225
rect 45645 -13345 45700 -13225
rect 45820 -13345 45865 -13225
rect 45985 -13345 46030 -13225
rect 46150 -13345 46195 -13225
rect 46315 -13345 46370 -13225
rect 46490 -13345 46535 -13225
rect 46655 -13345 46700 -13225
rect 46820 -13345 46865 -13225
rect 46985 -13345 47040 -13225
rect 47160 -13345 47205 -13225
rect 47325 -13345 47370 -13225
rect 47490 -13345 47535 -13225
rect 47655 -13345 47665 -13225
rect 42165 -13400 47665 -13345
rect 42165 -13520 42175 -13400
rect 42295 -13520 42350 -13400
rect 42470 -13520 42515 -13400
rect 42635 -13520 42680 -13400
rect 42800 -13520 42845 -13400
rect 42965 -13520 43020 -13400
rect 43140 -13520 43185 -13400
rect 43305 -13520 43350 -13400
rect 43470 -13520 43515 -13400
rect 43635 -13520 43690 -13400
rect 43810 -13520 43855 -13400
rect 43975 -13520 44020 -13400
rect 44140 -13520 44185 -13400
rect 44305 -13520 44360 -13400
rect 44480 -13520 44525 -13400
rect 44645 -13520 44690 -13400
rect 44810 -13520 44855 -13400
rect 44975 -13520 45030 -13400
rect 45150 -13520 45195 -13400
rect 45315 -13520 45360 -13400
rect 45480 -13520 45525 -13400
rect 45645 -13520 45700 -13400
rect 45820 -13520 45865 -13400
rect 45985 -13520 46030 -13400
rect 46150 -13520 46195 -13400
rect 46315 -13520 46370 -13400
rect 46490 -13520 46535 -13400
rect 46655 -13520 46700 -13400
rect 46820 -13520 46865 -13400
rect 46985 -13520 47040 -13400
rect 47160 -13520 47205 -13400
rect 47325 -13520 47370 -13400
rect 47490 -13520 47535 -13400
rect 47655 -13520 47665 -13400
rect 42165 -13565 47665 -13520
rect 42165 -13685 42175 -13565
rect 42295 -13685 42350 -13565
rect 42470 -13685 42515 -13565
rect 42635 -13685 42680 -13565
rect 42800 -13685 42845 -13565
rect 42965 -13685 43020 -13565
rect 43140 -13685 43185 -13565
rect 43305 -13685 43350 -13565
rect 43470 -13685 43515 -13565
rect 43635 -13685 43690 -13565
rect 43810 -13685 43855 -13565
rect 43975 -13685 44020 -13565
rect 44140 -13685 44185 -13565
rect 44305 -13685 44360 -13565
rect 44480 -13685 44525 -13565
rect 44645 -13685 44690 -13565
rect 44810 -13685 44855 -13565
rect 44975 -13685 45030 -13565
rect 45150 -13685 45195 -13565
rect 45315 -13685 45360 -13565
rect 45480 -13685 45525 -13565
rect 45645 -13685 45700 -13565
rect 45820 -13685 45865 -13565
rect 45985 -13685 46030 -13565
rect 46150 -13685 46195 -13565
rect 46315 -13685 46370 -13565
rect 46490 -13685 46535 -13565
rect 46655 -13685 46700 -13565
rect 46820 -13685 46865 -13565
rect 46985 -13685 47040 -13565
rect 47160 -13685 47205 -13565
rect 47325 -13685 47370 -13565
rect 47490 -13685 47535 -13565
rect 47655 -13685 47665 -13565
rect 42165 -13730 47665 -13685
rect 42165 -13850 42175 -13730
rect 42295 -13850 42350 -13730
rect 42470 -13850 42515 -13730
rect 42635 -13850 42680 -13730
rect 42800 -13850 42845 -13730
rect 42965 -13850 43020 -13730
rect 43140 -13850 43185 -13730
rect 43305 -13850 43350 -13730
rect 43470 -13850 43515 -13730
rect 43635 -13850 43690 -13730
rect 43810 -13850 43855 -13730
rect 43975 -13850 44020 -13730
rect 44140 -13850 44185 -13730
rect 44305 -13850 44360 -13730
rect 44480 -13850 44525 -13730
rect 44645 -13850 44690 -13730
rect 44810 -13850 44855 -13730
rect 44975 -13850 45030 -13730
rect 45150 -13850 45195 -13730
rect 45315 -13850 45360 -13730
rect 45480 -13850 45525 -13730
rect 45645 -13850 45700 -13730
rect 45820 -13850 45865 -13730
rect 45985 -13850 46030 -13730
rect 46150 -13850 46195 -13730
rect 46315 -13850 46370 -13730
rect 46490 -13850 46535 -13730
rect 46655 -13850 46700 -13730
rect 46820 -13850 46865 -13730
rect 46985 -13850 47040 -13730
rect 47160 -13850 47205 -13730
rect 47325 -13850 47370 -13730
rect 47490 -13850 47535 -13730
rect 47655 -13850 47665 -13730
rect 42165 -13895 47665 -13850
rect 42165 -14015 42175 -13895
rect 42295 -14015 42350 -13895
rect 42470 -14015 42515 -13895
rect 42635 -14015 42680 -13895
rect 42800 -14015 42845 -13895
rect 42965 -14015 43020 -13895
rect 43140 -14015 43185 -13895
rect 43305 -14015 43350 -13895
rect 43470 -14015 43515 -13895
rect 43635 -14015 43690 -13895
rect 43810 -14015 43855 -13895
rect 43975 -14015 44020 -13895
rect 44140 -14015 44185 -13895
rect 44305 -14015 44360 -13895
rect 44480 -14015 44525 -13895
rect 44645 -14015 44690 -13895
rect 44810 -14015 44855 -13895
rect 44975 -14015 45030 -13895
rect 45150 -14015 45195 -13895
rect 45315 -14015 45360 -13895
rect 45480 -14015 45525 -13895
rect 45645 -14015 45700 -13895
rect 45820 -14015 45865 -13895
rect 45985 -14015 46030 -13895
rect 46150 -14015 46195 -13895
rect 46315 -14015 46370 -13895
rect 46490 -14015 46535 -13895
rect 46655 -14015 46700 -13895
rect 46820 -14015 46865 -13895
rect 46985 -14015 47040 -13895
rect 47160 -14015 47205 -13895
rect 47325 -14015 47370 -13895
rect 47490 -14015 47535 -13895
rect 47655 -14015 47665 -13895
rect 42165 -14070 47665 -14015
rect 42165 -14190 42175 -14070
rect 42295 -14190 42350 -14070
rect 42470 -14190 42515 -14070
rect 42635 -14190 42680 -14070
rect 42800 -14190 42845 -14070
rect 42965 -14190 43020 -14070
rect 43140 -14190 43185 -14070
rect 43305 -14190 43350 -14070
rect 43470 -14190 43515 -14070
rect 43635 -14190 43690 -14070
rect 43810 -14190 43855 -14070
rect 43975 -14190 44020 -14070
rect 44140 -14190 44185 -14070
rect 44305 -14190 44360 -14070
rect 44480 -14190 44525 -14070
rect 44645 -14190 44690 -14070
rect 44810 -14190 44855 -14070
rect 44975 -14190 45030 -14070
rect 45150 -14190 45195 -14070
rect 45315 -14190 45360 -14070
rect 45480 -14190 45525 -14070
rect 45645 -14190 45700 -14070
rect 45820 -14190 45865 -14070
rect 45985 -14190 46030 -14070
rect 46150 -14190 46195 -14070
rect 46315 -14190 46370 -14070
rect 46490 -14190 46535 -14070
rect 46655 -14190 46700 -14070
rect 46820 -14190 46865 -14070
rect 46985 -14190 47040 -14070
rect 47160 -14190 47205 -14070
rect 47325 -14190 47370 -14070
rect 47490 -14190 47535 -14070
rect 47655 -14190 47665 -14070
rect 42165 -14235 47665 -14190
rect 42165 -14355 42175 -14235
rect 42295 -14355 42350 -14235
rect 42470 -14355 42515 -14235
rect 42635 -14355 42680 -14235
rect 42800 -14355 42845 -14235
rect 42965 -14355 43020 -14235
rect 43140 -14355 43185 -14235
rect 43305 -14355 43350 -14235
rect 43470 -14355 43515 -14235
rect 43635 -14355 43690 -14235
rect 43810 -14355 43855 -14235
rect 43975 -14355 44020 -14235
rect 44140 -14355 44185 -14235
rect 44305 -14355 44360 -14235
rect 44480 -14355 44525 -14235
rect 44645 -14355 44690 -14235
rect 44810 -14355 44855 -14235
rect 44975 -14355 45030 -14235
rect 45150 -14355 45195 -14235
rect 45315 -14355 45360 -14235
rect 45480 -14355 45525 -14235
rect 45645 -14355 45700 -14235
rect 45820 -14355 45865 -14235
rect 45985 -14355 46030 -14235
rect 46150 -14355 46195 -14235
rect 46315 -14355 46370 -14235
rect 46490 -14355 46535 -14235
rect 46655 -14355 46700 -14235
rect 46820 -14355 46865 -14235
rect 46985 -14355 47040 -14235
rect 47160 -14355 47205 -14235
rect 47325 -14355 47370 -14235
rect 47490 -14355 47535 -14235
rect 47655 -14355 47665 -14235
rect 42165 -14400 47665 -14355
rect 42165 -14520 42175 -14400
rect 42295 -14520 42350 -14400
rect 42470 -14520 42515 -14400
rect 42635 -14520 42680 -14400
rect 42800 -14520 42845 -14400
rect 42965 -14520 43020 -14400
rect 43140 -14520 43185 -14400
rect 43305 -14520 43350 -14400
rect 43470 -14520 43515 -14400
rect 43635 -14520 43690 -14400
rect 43810 -14520 43855 -14400
rect 43975 -14520 44020 -14400
rect 44140 -14520 44185 -14400
rect 44305 -14520 44360 -14400
rect 44480 -14520 44525 -14400
rect 44645 -14520 44690 -14400
rect 44810 -14520 44855 -14400
rect 44975 -14520 45030 -14400
rect 45150 -14520 45195 -14400
rect 45315 -14520 45360 -14400
rect 45480 -14520 45525 -14400
rect 45645 -14520 45700 -14400
rect 45820 -14520 45865 -14400
rect 45985 -14520 46030 -14400
rect 46150 -14520 46195 -14400
rect 46315 -14520 46370 -14400
rect 46490 -14520 46535 -14400
rect 46655 -14520 46700 -14400
rect 46820 -14520 46865 -14400
rect 46985 -14520 47040 -14400
rect 47160 -14520 47205 -14400
rect 47325 -14520 47370 -14400
rect 47490 -14520 47535 -14400
rect 47655 -14520 47665 -14400
rect 42165 -14565 47665 -14520
rect 42165 -14685 42175 -14565
rect 42295 -14685 42350 -14565
rect 42470 -14685 42515 -14565
rect 42635 -14685 42680 -14565
rect 42800 -14685 42845 -14565
rect 42965 -14685 43020 -14565
rect 43140 -14685 43185 -14565
rect 43305 -14685 43350 -14565
rect 43470 -14685 43515 -14565
rect 43635 -14685 43690 -14565
rect 43810 -14685 43855 -14565
rect 43975 -14685 44020 -14565
rect 44140 -14685 44185 -14565
rect 44305 -14685 44360 -14565
rect 44480 -14685 44525 -14565
rect 44645 -14685 44690 -14565
rect 44810 -14685 44855 -14565
rect 44975 -14685 45030 -14565
rect 45150 -14685 45195 -14565
rect 45315 -14685 45360 -14565
rect 45480 -14685 45525 -14565
rect 45645 -14685 45700 -14565
rect 45820 -14685 45865 -14565
rect 45985 -14685 46030 -14565
rect 46150 -14685 46195 -14565
rect 46315 -14685 46370 -14565
rect 46490 -14685 46535 -14565
rect 46655 -14685 46700 -14565
rect 46820 -14685 46865 -14565
rect 46985 -14685 47040 -14565
rect 47160 -14685 47205 -14565
rect 47325 -14685 47370 -14565
rect 47490 -14685 47535 -14565
rect 47655 -14685 47665 -14565
rect 42165 -14740 47665 -14685
rect 42165 -14860 42175 -14740
rect 42295 -14860 42350 -14740
rect 42470 -14860 42515 -14740
rect 42635 -14860 42680 -14740
rect 42800 -14860 42845 -14740
rect 42965 -14860 43020 -14740
rect 43140 -14860 43185 -14740
rect 43305 -14860 43350 -14740
rect 43470 -14860 43515 -14740
rect 43635 -14860 43690 -14740
rect 43810 -14860 43855 -14740
rect 43975 -14860 44020 -14740
rect 44140 -14860 44185 -14740
rect 44305 -14860 44360 -14740
rect 44480 -14860 44525 -14740
rect 44645 -14860 44690 -14740
rect 44810 -14860 44855 -14740
rect 44975 -14860 45030 -14740
rect 45150 -14860 45195 -14740
rect 45315 -14860 45360 -14740
rect 45480 -14860 45525 -14740
rect 45645 -14860 45700 -14740
rect 45820 -14860 45865 -14740
rect 45985 -14860 46030 -14740
rect 46150 -14860 46195 -14740
rect 46315 -14860 46370 -14740
rect 46490 -14860 46535 -14740
rect 46655 -14860 46700 -14740
rect 46820 -14860 46865 -14740
rect 46985 -14860 47040 -14740
rect 47160 -14860 47205 -14740
rect 47325 -14860 47370 -14740
rect 47490 -14860 47535 -14740
rect 47655 -14860 47665 -14740
rect 42165 -14905 47665 -14860
rect 42165 -15025 42175 -14905
rect 42295 -15025 42350 -14905
rect 42470 -15025 42515 -14905
rect 42635 -15025 42680 -14905
rect 42800 -15025 42845 -14905
rect 42965 -15025 43020 -14905
rect 43140 -15025 43185 -14905
rect 43305 -15025 43350 -14905
rect 43470 -15025 43515 -14905
rect 43635 -15025 43690 -14905
rect 43810 -15025 43855 -14905
rect 43975 -15025 44020 -14905
rect 44140 -15025 44185 -14905
rect 44305 -15025 44360 -14905
rect 44480 -15025 44525 -14905
rect 44645 -15025 44690 -14905
rect 44810 -15025 44855 -14905
rect 44975 -15025 45030 -14905
rect 45150 -15025 45195 -14905
rect 45315 -15025 45360 -14905
rect 45480 -15025 45525 -14905
rect 45645 -15025 45700 -14905
rect 45820 -15025 45865 -14905
rect 45985 -15025 46030 -14905
rect 46150 -15025 46195 -14905
rect 46315 -15025 46370 -14905
rect 46490 -15025 46535 -14905
rect 46655 -15025 46700 -14905
rect 46820 -15025 46865 -14905
rect 46985 -15025 47040 -14905
rect 47160 -15025 47205 -14905
rect 47325 -15025 47370 -14905
rect 47490 -15025 47535 -14905
rect 47655 -15025 47665 -14905
rect 42165 -15070 47665 -15025
rect 42165 -15190 42175 -15070
rect 42295 -15190 42350 -15070
rect 42470 -15190 42515 -15070
rect 42635 -15190 42680 -15070
rect 42800 -15190 42845 -15070
rect 42965 -15190 43020 -15070
rect 43140 -15190 43185 -15070
rect 43305 -15190 43350 -15070
rect 43470 -15190 43515 -15070
rect 43635 -15190 43690 -15070
rect 43810 -15190 43855 -15070
rect 43975 -15190 44020 -15070
rect 44140 -15190 44185 -15070
rect 44305 -15190 44360 -15070
rect 44480 -15190 44525 -15070
rect 44645 -15190 44690 -15070
rect 44810 -15190 44855 -15070
rect 44975 -15190 45030 -15070
rect 45150 -15190 45195 -15070
rect 45315 -15190 45360 -15070
rect 45480 -15190 45525 -15070
rect 45645 -15190 45700 -15070
rect 45820 -15190 45865 -15070
rect 45985 -15190 46030 -15070
rect 46150 -15190 46195 -15070
rect 46315 -15190 46370 -15070
rect 46490 -15190 46535 -15070
rect 46655 -15190 46700 -15070
rect 46820 -15190 46865 -15070
rect 46985 -15190 47040 -15070
rect 47160 -15190 47205 -15070
rect 47325 -15190 47370 -15070
rect 47490 -15190 47535 -15070
rect 47655 -15190 47665 -15070
rect 42165 -15235 47665 -15190
rect 42165 -15355 42175 -15235
rect 42295 -15355 42350 -15235
rect 42470 -15355 42515 -15235
rect 42635 -15355 42680 -15235
rect 42800 -15355 42845 -15235
rect 42965 -15355 43020 -15235
rect 43140 -15355 43185 -15235
rect 43305 -15355 43350 -15235
rect 43470 -15355 43515 -15235
rect 43635 -15355 43690 -15235
rect 43810 -15355 43855 -15235
rect 43975 -15355 44020 -15235
rect 44140 -15355 44185 -15235
rect 44305 -15355 44360 -15235
rect 44480 -15355 44525 -15235
rect 44645 -15355 44690 -15235
rect 44810 -15355 44855 -15235
rect 44975 -15355 45030 -15235
rect 45150 -15355 45195 -15235
rect 45315 -15355 45360 -15235
rect 45480 -15355 45525 -15235
rect 45645 -15355 45700 -15235
rect 45820 -15355 45865 -15235
rect 45985 -15355 46030 -15235
rect 46150 -15355 46195 -15235
rect 46315 -15355 46370 -15235
rect 46490 -15355 46535 -15235
rect 46655 -15355 46700 -15235
rect 46820 -15355 46865 -15235
rect 46985 -15355 47040 -15235
rect 47160 -15355 47205 -15235
rect 47325 -15355 47370 -15235
rect 47490 -15355 47535 -15235
rect 47655 -15355 47665 -15235
rect 42165 -15410 47665 -15355
rect 42165 -15530 42175 -15410
rect 42295 -15530 42350 -15410
rect 42470 -15530 42515 -15410
rect 42635 -15530 42680 -15410
rect 42800 -15530 42845 -15410
rect 42965 -15530 43020 -15410
rect 43140 -15530 43185 -15410
rect 43305 -15530 43350 -15410
rect 43470 -15530 43515 -15410
rect 43635 -15530 43690 -15410
rect 43810 -15530 43855 -15410
rect 43975 -15530 44020 -15410
rect 44140 -15530 44185 -15410
rect 44305 -15530 44360 -15410
rect 44480 -15530 44525 -15410
rect 44645 -15530 44690 -15410
rect 44810 -15530 44855 -15410
rect 44975 -15530 45030 -15410
rect 45150 -15530 45195 -15410
rect 45315 -15530 45360 -15410
rect 45480 -15530 45525 -15410
rect 45645 -15530 45700 -15410
rect 45820 -15530 45865 -15410
rect 45985 -15530 46030 -15410
rect 46150 -15530 46195 -15410
rect 46315 -15530 46370 -15410
rect 46490 -15530 46535 -15410
rect 46655 -15530 46700 -15410
rect 46820 -15530 46865 -15410
rect 46985 -15530 47040 -15410
rect 47160 -15530 47205 -15410
rect 47325 -15530 47370 -15410
rect 47490 -15530 47535 -15410
rect 47655 -15530 47665 -15410
rect 42165 -15540 47665 -15530
rect 47855 -10050 53355 -10040
rect 47855 -10170 47865 -10050
rect 47985 -10170 48040 -10050
rect 48160 -10170 48205 -10050
rect 48325 -10170 48370 -10050
rect 48490 -10170 48535 -10050
rect 48655 -10170 48710 -10050
rect 48830 -10170 48875 -10050
rect 48995 -10170 49040 -10050
rect 49160 -10170 49205 -10050
rect 49325 -10170 49380 -10050
rect 49500 -10170 49545 -10050
rect 49665 -10170 49710 -10050
rect 49830 -10170 49875 -10050
rect 49995 -10170 50050 -10050
rect 50170 -10170 50215 -10050
rect 50335 -10170 50380 -10050
rect 50500 -10170 50545 -10050
rect 50665 -10170 50720 -10050
rect 50840 -10170 50885 -10050
rect 51005 -10170 51050 -10050
rect 51170 -10170 51215 -10050
rect 51335 -10170 51390 -10050
rect 51510 -10170 51555 -10050
rect 51675 -10170 51720 -10050
rect 51840 -10170 51885 -10050
rect 52005 -10170 52060 -10050
rect 52180 -10170 52225 -10050
rect 52345 -10170 52390 -10050
rect 52510 -10170 52555 -10050
rect 52675 -10170 52730 -10050
rect 52850 -10170 52895 -10050
rect 53015 -10170 53060 -10050
rect 53180 -10170 53225 -10050
rect 53345 -10170 53355 -10050
rect 47855 -10215 53355 -10170
rect 47855 -10335 47865 -10215
rect 47985 -10335 48040 -10215
rect 48160 -10335 48205 -10215
rect 48325 -10335 48370 -10215
rect 48490 -10335 48535 -10215
rect 48655 -10335 48710 -10215
rect 48830 -10335 48875 -10215
rect 48995 -10335 49040 -10215
rect 49160 -10335 49205 -10215
rect 49325 -10335 49380 -10215
rect 49500 -10335 49545 -10215
rect 49665 -10335 49710 -10215
rect 49830 -10335 49875 -10215
rect 49995 -10335 50050 -10215
rect 50170 -10335 50215 -10215
rect 50335 -10335 50380 -10215
rect 50500 -10335 50545 -10215
rect 50665 -10335 50720 -10215
rect 50840 -10335 50885 -10215
rect 51005 -10335 51050 -10215
rect 51170 -10335 51215 -10215
rect 51335 -10335 51390 -10215
rect 51510 -10335 51555 -10215
rect 51675 -10335 51720 -10215
rect 51840 -10335 51885 -10215
rect 52005 -10335 52060 -10215
rect 52180 -10335 52225 -10215
rect 52345 -10335 52390 -10215
rect 52510 -10335 52555 -10215
rect 52675 -10335 52730 -10215
rect 52850 -10335 52895 -10215
rect 53015 -10335 53060 -10215
rect 53180 -10335 53225 -10215
rect 53345 -10335 53355 -10215
rect 47855 -10380 53355 -10335
rect 47855 -10500 47865 -10380
rect 47985 -10500 48040 -10380
rect 48160 -10500 48205 -10380
rect 48325 -10500 48370 -10380
rect 48490 -10500 48535 -10380
rect 48655 -10500 48710 -10380
rect 48830 -10500 48875 -10380
rect 48995 -10500 49040 -10380
rect 49160 -10500 49205 -10380
rect 49325 -10500 49380 -10380
rect 49500 -10500 49545 -10380
rect 49665 -10500 49710 -10380
rect 49830 -10500 49875 -10380
rect 49995 -10500 50050 -10380
rect 50170 -10500 50215 -10380
rect 50335 -10500 50380 -10380
rect 50500 -10500 50545 -10380
rect 50665 -10500 50720 -10380
rect 50840 -10500 50885 -10380
rect 51005 -10500 51050 -10380
rect 51170 -10500 51215 -10380
rect 51335 -10500 51390 -10380
rect 51510 -10500 51555 -10380
rect 51675 -10500 51720 -10380
rect 51840 -10500 51885 -10380
rect 52005 -10500 52060 -10380
rect 52180 -10500 52225 -10380
rect 52345 -10500 52390 -10380
rect 52510 -10500 52555 -10380
rect 52675 -10500 52730 -10380
rect 52850 -10500 52895 -10380
rect 53015 -10500 53060 -10380
rect 53180 -10500 53225 -10380
rect 53345 -10500 53355 -10380
rect 47855 -10545 53355 -10500
rect 47855 -10665 47865 -10545
rect 47985 -10665 48040 -10545
rect 48160 -10665 48205 -10545
rect 48325 -10665 48370 -10545
rect 48490 -10665 48535 -10545
rect 48655 -10665 48710 -10545
rect 48830 -10665 48875 -10545
rect 48995 -10665 49040 -10545
rect 49160 -10665 49205 -10545
rect 49325 -10665 49380 -10545
rect 49500 -10665 49545 -10545
rect 49665 -10665 49710 -10545
rect 49830 -10665 49875 -10545
rect 49995 -10665 50050 -10545
rect 50170 -10665 50215 -10545
rect 50335 -10665 50380 -10545
rect 50500 -10665 50545 -10545
rect 50665 -10665 50720 -10545
rect 50840 -10665 50885 -10545
rect 51005 -10665 51050 -10545
rect 51170 -10665 51215 -10545
rect 51335 -10665 51390 -10545
rect 51510 -10665 51555 -10545
rect 51675 -10665 51720 -10545
rect 51840 -10665 51885 -10545
rect 52005 -10665 52060 -10545
rect 52180 -10665 52225 -10545
rect 52345 -10665 52390 -10545
rect 52510 -10665 52555 -10545
rect 52675 -10665 52730 -10545
rect 52850 -10665 52895 -10545
rect 53015 -10665 53060 -10545
rect 53180 -10665 53225 -10545
rect 53345 -10665 53355 -10545
rect 47855 -10720 53355 -10665
rect 47855 -10840 47865 -10720
rect 47985 -10840 48040 -10720
rect 48160 -10840 48205 -10720
rect 48325 -10840 48370 -10720
rect 48490 -10840 48535 -10720
rect 48655 -10840 48710 -10720
rect 48830 -10840 48875 -10720
rect 48995 -10840 49040 -10720
rect 49160 -10840 49205 -10720
rect 49325 -10840 49380 -10720
rect 49500 -10840 49545 -10720
rect 49665 -10840 49710 -10720
rect 49830 -10840 49875 -10720
rect 49995 -10840 50050 -10720
rect 50170 -10840 50215 -10720
rect 50335 -10840 50380 -10720
rect 50500 -10840 50545 -10720
rect 50665 -10840 50720 -10720
rect 50840 -10840 50885 -10720
rect 51005 -10840 51050 -10720
rect 51170 -10840 51215 -10720
rect 51335 -10840 51390 -10720
rect 51510 -10840 51555 -10720
rect 51675 -10840 51720 -10720
rect 51840 -10840 51885 -10720
rect 52005 -10840 52060 -10720
rect 52180 -10840 52225 -10720
rect 52345 -10840 52390 -10720
rect 52510 -10840 52555 -10720
rect 52675 -10840 52730 -10720
rect 52850 -10840 52895 -10720
rect 53015 -10840 53060 -10720
rect 53180 -10840 53225 -10720
rect 53345 -10840 53355 -10720
rect 47855 -10885 53355 -10840
rect 47855 -11005 47865 -10885
rect 47985 -11005 48040 -10885
rect 48160 -11005 48205 -10885
rect 48325 -11005 48370 -10885
rect 48490 -11005 48535 -10885
rect 48655 -11005 48710 -10885
rect 48830 -11005 48875 -10885
rect 48995 -11005 49040 -10885
rect 49160 -11005 49205 -10885
rect 49325 -11005 49380 -10885
rect 49500 -11005 49545 -10885
rect 49665 -11005 49710 -10885
rect 49830 -11005 49875 -10885
rect 49995 -11005 50050 -10885
rect 50170 -11005 50215 -10885
rect 50335 -11005 50380 -10885
rect 50500 -11005 50545 -10885
rect 50665 -11005 50720 -10885
rect 50840 -11005 50885 -10885
rect 51005 -11005 51050 -10885
rect 51170 -11005 51215 -10885
rect 51335 -11005 51390 -10885
rect 51510 -11005 51555 -10885
rect 51675 -11005 51720 -10885
rect 51840 -11005 51885 -10885
rect 52005 -11005 52060 -10885
rect 52180 -11005 52225 -10885
rect 52345 -11005 52390 -10885
rect 52510 -11005 52555 -10885
rect 52675 -11005 52730 -10885
rect 52850 -11005 52895 -10885
rect 53015 -11005 53060 -10885
rect 53180 -11005 53225 -10885
rect 53345 -11005 53355 -10885
rect 47855 -11050 53355 -11005
rect 47855 -11170 47865 -11050
rect 47985 -11170 48040 -11050
rect 48160 -11170 48205 -11050
rect 48325 -11170 48370 -11050
rect 48490 -11170 48535 -11050
rect 48655 -11170 48710 -11050
rect 48830 -11170 48875 -11050
rect 48995 -11170 49040 -11050
rect 49160 -11170 49205 -11050
rect 49325 -11170 49380 -11050
rect 49500 -11170 49545 -11050
rect 49665 -11170 49710 -11050
rect 49830 -11170 49875 -11050
rect 49995 -11170 50050 -11050
rect 50170 -11170 50215 -11050
rect 50335 -11170 50380 -11050
rect 50500 -11170 50545 -11050
rect 50665 -11170 50720 -11050
rect 50840 -11170 50885 -11050
rect 51005 -11170 51050 -11050
rect 51170 -11170 51215 -11050
rect 51335 -11170 51390 -11050
rect 51510 -11170 51555 -11050
rect 51675 -11170 51720 -11050
rect 51840 -11170 51885 -11050
rect 52005 -11170 52060 -11050
rect 52180 -11170 52225 -11050
rect 52345 -11170 52390 -11050
rect 52510 -11170 52555 -11050
rect 52675 -11170 52730 -11050
rect 52850 -11170 52895 -11050
rect 53015 -11170 53060 -11050
rect 53180 -11170 53225 -11050
rect 53345 -11170 53355 -11050
rect 47855 -11215 53355 -11170
rect 47855 -11335 47865 -11215
rect 47985 -11335 48040 -11215
rect 48160 -11335 48205 -11215
rect 48325 -11335 48370 -11215
rect 48490 -11335 48535 -11215
rect 48655 -11335 48710 -11215
rect 48830 -11335 48875 -11215
rect 48995 -11335 49040 -11215
rect 49160 -11335 49205 -11215
rect 49325 -11335 49380 -11215
rect 49500 -11335 49545 -11215
rect 49665 -11335 49710 -11215
rect 49830 -11335 49875 -11215
rect 49995 -11335 50050 -11215
rect 50170 -11335 50215 -11215
rect 50335 -11335 50380 -11215
rect 50500 -11335 50545 -11215
rect 50665 -11335 50720 -11215
rect 50840 -11335 50885 -11215
rect 51005 -11335 51050 -11215
rect 51170 -11335 51215 -11215
rect 51335 -11335 51390 -11215
rect 51510 -11335 51555 -11215
rect 51675 -11335 51720 -11215
rect 51840 -11335 51885 -11215
rect 52005 -11335 52060 -11215
rect 52180 -11335 52225 -11215
rect 52345 -11335 52390 -11215
rect 52510 -11335 52555 -11215
rect 52675 -11335 52730 -11215
rect 52850 -11335 52895 -11215
rect 53015 -11335 53060 -11215
rect 53180 -11335 53225 -11215
rect 53345 -11335 53355 -11215
rect 47855 -11390 53355 -11335
rect 47855 -11510 47865 -11390
rect 47985 -11510 48040 -11390
rect 48160 -11510 48205 -11390
rect 48325 -11510 48370 -11390
rect 48490 -11510 48535 -11390
rect 48655 -11510 48710 -11390
rect 48830 -11510 48875 -11390
rect 48995 -11510 49040 -11390
rect 49160 -11510 49205 -11390
rect 49325 -11510 49380 -11390
rect 49500 -11510 49545 -11390
rect 49665 -11510 49710 -11390
rect 49830 -11510 49875 -11390
rect 49995 -11510 50050 -11390
rect 50170 -11510 50215 -11390
rect 50335 -11510 50380 -11390
rect 50500 -11510 50545 -11390
rect 50665 -11510 50720 -11390
rect 50840 -11510 50885 -11390
rect 51005 -11510 51050 -11390
rect 51170 -11510 51215 -11390
rect 51335 -11510 51390 -11390
rect 51510 -11510 51555 -11390
rect 51675 -11510 51720 -11390
rect 51840 -11510 51885 -11390
rect 52005 -11510 52060 -11390
rect 52180 -11510 52225 -11390
rect 52345 -11510 52390 -11390
rect 52510 -11510 52555 -11390
rect 52675 -11510 52730 -11390
rect 52850 -11510 52895 -11390
rect 53015 -11510 53060 -11390
rect 53180 -11510 53225 -11390
rect 53345 -11510 53355 -11390
rect 47855 -11555 53355 -11510
rect 47855 -11675 47865 -11555
rect 47985 -11675 48040 -11555
rect 48160 -11675 48205 -11555
rect 48325 -11675 48370 -11555
rect 48490 -11675 48535 -11555
rect 48655 -11675 48710 -11555
rect 48830 -11675 48875 -11555
rect 48995 -11675 49040 -11555
rect 49160 -11675 49205 -11555
rect 49325 -11675 49380 -11555
rect 49500 -11675 49545 -11555
rect 49665 -11675 49710 -11555
rect 49830 -11675 49875 -11555
rect 49995 -11675 50050 -11555
rect 50170 -11675 50215 -11555
rect 50335 -11675 50380 -11555
rect 50500 -11675 50545 -11555
rect 50665 -11675 50720 -11555
rect 50840 -11675 50885 -11555
rect 51005 -11675 51050 -11555
rect 51170 -11675 51215 -11555
rect 51335 -11675 51390 -11555
rect 51510 -11675 51555 -11555
rect 51675 -11675 51720 -11555
rect 51840 -11675 51885 -11555
rect 52005 -11675 52060 -11555
rect 52180 -11675 52225 -11555
rect 52345 -11675 52390 -11555
rect 52510 -11675 52555 -11555
rect 52675 -11675 52730 -11555
rect 52850 -11675 52895 -11555
rect 53015 -11675 53060 -11555
rect 53180 -11675 53225 -11555
rect 53345 -11675 53355 -11555
rect 47855 -11720 53355 -11675
rect 47855 -11840 47865 -11720
rect 47985 -11840 48040 -11720
rect 48160 -11840 48205 -11720
rect 48325 -11840 48370 -11720
rect 48490 -11840 48535 -11720
rect 48655 -11840 48710 -11720
rect 48830 -11840 48875 -11720
rect 48995 -11840 49040 -11720
rect 49160 -11840 49205 -11720
rect 49325 -11840 49380 -11720
rect 49500 -11840 49545 -11720
rect 49665 -11840 49710 -11720
rect 49830 -11840 49875 -11720
rect 49995 -11840 50050 -11720
rect 50170 -11840 50215 -11720
rect 50335 -11840 50380 -11720
rect 50500 -11840 50545 -11720
rect 50665 -11840 50720 -11720
rect 50840 -11840 50885 -11720
rect 51005 -11840 51050 -11720
rect 51170 -11840 51215 -11720
rect 51335 -11840 51390 -11720
rect 51510 -11840 51555 -11720
rect 51675 -11840 51720 -11720
rect 51840 -11840 51885 -11720
rect 52005 -11840 52060 -11720
rect 52180 -11840 52225 -11720
rect 52345 -11840 52390 -11720
rect 52510 -11840 52555 -11720
rect 52675 -11840 52730 -11720
rect 52850 -11840 52895 -11720
rect 53015 -11840 53060 -11720
rect 53180 -11840 53225 -11720
rect 53345 -11840 53355 -11720
rect 47855 -11885 53355 -11840
rect 47855 -12005 47865 -11885
rect 47985 -12005 48040 -11885
rect 48160 -12005 48205 -11885
rect 48325 -12005 48370 -11885
rect 48490 -12005 48535 -11885
rect 48655 -12005 48710 -11885
rect 48830 -12005 48875 -11885
rect 48995 -12005 49040 -11885
rect 49160 -12005 49205 -11885
rect 49325 -12005 49380 -11885
rect 49500 -12005 49545 -11885
rect 49665 -12005 49710 -11885
rect 49830 -12005 49875 -11885
rect 49995 -12005 50050 -11885
rect 50170 -12005 50215 -11885
rect 50335 -12005 50380 -11885
rect 50500 -12005 50545 -11885
rect 50665 -12005 50720 -11885
rect 50840 -12005 50885 -11885
rect 51005 -12005 51050 -11885
rect 51170 -12005 51215 -11885
rect 51335 -12005 51390 -11885
rect 51510 -12005 51555 -11885
rect 51675 -12005 51720 -11885
rect 51840 -12005 51885 -11885
rect 52005 -12005 52060 -11885
rect 52180 -12005 52225 -11885
rect 52345 -12005 52390 -11885
rect 52510 -12005 52555 -11885
rect 52675 -12005 52730 -11885
rect 52850 -12005 52895 -11885
rect 53015 -12005 53060 -11885
rect 53180 -12005 53225 -11885
rect 53345 -12005 53355 -11885
rect 47855 -12060 53355 -12005
rect 47855 -12180 47865 -12060
rect 47985 -12180 48040 -12060
rect 48160 -12180 48205 -12060
rect 48325 -12180 48370 -12060
rect 48490 -12180 48535 -12060
rect 48655 -12180 48710 -12060
rect 48830 -12180 48875 -12060
rect 48995 -12180 49040 -12060
rect 49160 -12180 49205 -12060
rect 49325 -12180 49380 -12060
rect 49500 -12180 49545 -12060
rect 49665 -12180 49710 -12060
rect 49830 -12180 49875 -12060
rect 49995 -12180 50050 -12060
rect 50170 -12180 50215 -12060
rect 50335 -12180 50380 -12060
rect 50500 -12180 50545 -12060
rect 50665 -12180 50720 -12060
rect 50840 -12180 50885 -12060
rect 51005 -12180 51050 -12060
rect 51170 -12180 51215 -12060
rect 51335 -12180 51390 -12060
rect 51510 -12180 51555 -12060
rect 51675 -12180 51720 -12060
rect 51840 -12180 51885 -12060
rect 52005 -12180 52060 -12060
rect 52180 -12180 52225 -12060
rect 52345 -12180 52390 -12060
rect 52510 -12180 52555 -12060
rect 52675 -12180 52730 -12060
rect 52850 -12180 52895 -12060
rect 53015 -12180 53060 -12060
rect 53180 -12180 53225 -12060
rect 53345 -12180 53355 -12060
rect 47855 -12225 53355 -12180
rect 47855 -12345 47865 -12225
rect 47985 -12345 48040 -12225
rect 48160 -12345 48205 -12225
rect 48325 -12345 48370 -12225
rect 48490 -12345 48535 -12225
rect 48655 -12345 48710 -12225
rect 48830 -12345 48875 -12225
rect 48995 -12345 49040 -12225
rect 49160 -12345 49205 -12225
rect 49325 -12345 49380 -12225
rect 49500 -12345 49545 -12225
rect 49665 -12345 49710 -12225
rect 49830 -12345 49875 -12225
rect 49995 -12345 50050 -12225
rect 50170 -12345 50215 -12225
rect 50335 -12345 50380 -12225
rect 50500 -12345 50545 -12225
rect 50665 -12345 50720 -12225
rect 50840 -12345 50885 -12225
rect 51005 -12345 51050 -12225
rect 51170 -12345 51215 -12225
rect 51335 -12345 51390 -12225
rect 51510 -12345 51555 -12225
rect 51675 -12345 51720 -12225
rect 51840 -12345 51885 -12225
rect 52005 -12345 52060 -12225
rect 52180 -12345 52225 -12225
rect 52345 -12345 52390 -12225
rect 52510 -12345 52555 -12225
rect 52675 -12345 52730 -12225
rect 52850 -12345 52895 -12225
rect 53015 -12345 53060 -12225
rect 53180 -12345 53225 -12225
rect 53345 -12345 53355 -12225
rect 47855 -12390 53355 -12345
rect 47855 -12510 47865 -12390
rect 47985 -12510 48040 -12390
rect 48160 -12510 48205 -12390
rect 48325 -12510 48370 -12390
rect 48490 -12510 48535 -12390
rect 48655 -12510 48710 -12390
rect 48830 -12510 48875 -12390
rect 48995 -12510 49040 -12390
rect 49160 -12510 49205 -12390
rect 49325 -12510 49380 -12390
rect 49500 -12510 49545 -12390
rect 49665 -12510 49710 -12390
rect 49830 -12510 49875 -12390
rect 49995 -12510 50050 -12390
rect 50170 -12510 50215 -12390
rect 50335 -12510 50380 -12390
rect 50500 -12510 50545 -12390
rect 50665 -12510 50720 -12390
rect 50840 -12510 50885 -12390
rect 51005 -12510 51050 -12390
rect 51170 -12510 51215 -12390
rect 51335 -12510 51390 -12390
rect 51510 -12510 51555 -12390
rect 51675 -12510 51720 -12390
rect 51840 -12510 51885 -12390
rect 52005 -12510 52060 -12390
rect 52180 -12510 52225 -12390
rect 52345 -12510 52390 -12390
rect 52510 -12510 52555 -12390
rect 52675 -12510 52730 -12390
rect 52850 -12510 52895 -12390
rect 53015 -12510 53060 -12390
rect 53180 -12510 53225 -12390
rect 53345 -12510 53355 -12390
rect 47855 -12555 53355 -12510
rect 47855 -12675 47865 -12555
rect 47985 -12675 48040 -12555
rect 48160 -12675 48205 -12555
rect 48325 -12675 48370 -12555
rect 48490 -12675 48535 -12555
rect 48655 -12675 48710 -12555
rect 48830 -12675 48875 -12555
rect 48995 -12675 49040 -12555
rect 49160 -12675 49205 -12555
rect 49325 -12675 49380 -12555
rect 49500 -12675 49545 -12555
rect 49665 -12675 49710 -12555
rect 49830 -12675 49875 -12555
rect 49995 -12675 50050 -12555
rect 50170 -12675 50215 -12555
rect 50335 -12675 50380 -12555
rect 50500 -12675 50545 -12555
rect 50665 -12675 50720 -12555
rect 50840 -12675 50885 -12555
rect 51005 -12675 51050 -12555
rect 51170 -12675 51215 -12555
rect 51335 -12675 51390 -12555
rect 51510 -12675 51555 -12555
rect 51675 -12675 51720 -12555
rect 51840 -12675 51885 -12555
rect 52005 -12675 52060 -12555
rect 52180 -12675 52225 -12555
rect 52345 -12675 52390 -12555
rect 52510 -12675 52555 -12555
rect 52675 -12675 52730 -12555
rect 52850 -12675 52895 -12555
rect 53015 -12675 53060 -12555
rect 53180 -12675 53225 -12555
rect 53345 -12675 53355 -12555
rect 47855 -12730 53355 -12675
rect 47855 -12850 47865 -12730
rect 47985 -12850 48040 -12730
rect 48160 -12850 48205 -12730
rect 48325 -12850 48370 -12730
rect 48490 -12850 48535 -12730
rect 48655 -12850 48710 -12730
rect 48830 -12850 48875 -12730
rect 48995 -12850 49040 -12730
rect 49160 -12850 49205 -12730
rect 49325 -12850 49380 -12730
rect 49500 -12850 49545 -12730
rect 49665 -12850 49710 -12730
rect 49830 -12850 49875 -12730
rect 49995 -12850 50050 -12730
rect 50170 -12850 50215 -12730
rect 50335 -12850 50380 -12730
rect 50500 -12850 50545 -12730
rect 50665 -12850 50720 -12730
rect 50840 -12850 50885 -12730
rect 51005 -12850 51050 -12730
rect 51170 -12850 51215 -12730
rect 51335 -12850 51390 -12730
rect 51510 -12850 51555 -12730
rect 51675 -12850 51720 -12730
rect 51840 -12850 51885 -12730
rect 52005 -12850 52060 -12730
rect 52180 -12850 52225 -12730
rect 52345 -12850 52390 -12730
rect 52510 -12850 52555 -12730
rect 52675 -12850 52730 -12730
rect 52850 -12850 52895 -12730
rect 53015 -12850 53060 -12730
rect 53180 -12850 53225 -12730
rect 53345 -12850 53355 -12730
rect 47855 -12895 53355 -12850
rect 47855 -13015 47865 -12895
rect 47985 -13015 48040 -12895
rect 48160 -13015 48205 -12895
rect 48325 -13015 48370 -12895
rect 48490 -13015 48535 -12895
rect 48655 -13015 48710 -12895
rect 48830 -13015 48875 -12895
rect 48995 -13015 49040 -12895
rect 49160 -13015 49205 -12895
rect 49325 -13015 49380 -12895
rect 49500 -13015 49545 -12895
rect 49665 -13015 49710 -12895
rect 49830 -13015 49875 -12895
rect 49995 -13015 50050 -12895
rect 50170 -13015 50215 -12895
rect 50335 -13015 50380 -12895
rect 50500 -13015 50545 -12895
rect 50665 -13015 50720 -12895
rect 50840 -13015 50885 -12895
rect 51005 -13015 51050 -12895
rect 51170 -13015 51215 -12895
rect 51335 -13015 51390 -12895
rect 51510 -13015 51555 -12895
rect 51675 -13015 51720 -12895
rect 51840 -13015 51885 -12895
rect 52005 -13015 52060 -12895
rect 52180 -13015 52225 -12895
rect 52345 -13015 52390 -12895
rect 52510 -13015 52555 -12895
rect 52675 -13015 52730 -12895
rect 52850 -13015 52895 -12895
rect 53015 -13015 53060 -12895
rect 53180 -13015 53225 -12895
rect 53345 -13015 53355 -12895
rect 47855 -13060 53355 -13015
rect 47855 -13180 47865 -13060
rect 47985 -13180 48040 -13060
rect 48160 -13180 48205 -13060
rect 48325 -13180 48370 -13060
rect 48490 -13180 48535 -13060
rect 48655 -13180 48710 -13060
rect 48830 -13180 48875 -13060
rect 48995 -13180 49040 -13060
rect 49160 -13180 49205 -13060
rect 49325 -13180 49380 -13060
rect 49500 -13180 49545 -13060
rect 49665 -13180 49710 -13060
rect 49830 -13180 49875 -13060
rect 49995 -13180 50050 -13060
rect 50170 -13180 50215 -13060
rect 50335 -13180 50380 -13060
rect 50500 -13180 50545 -13060
rect 50665 -13180 50720 -13060
rect 50840 -13180 50885 -13060
rect 51005 -13180 51050 -13060
rect 51170 -13180 51215 -13060
rect 51335 -13180 51390 -13060
rect 51510 -13180 51555 -13060
rect 51675 -13180 51720 -13060
rect 51840 -13180 51885 -13060
rect 52005 -13180 52060 -13060
rect 52180 -13180 52225 -13060
rect 52345 -13180 52390 -13060
rect 52510 -13180 52555 -13060
rect 52675 -13180 52730 -13060
rect 52850 -13180 52895 -13060
rect 53015 -13180 53060 -13060
rect 53180 -13180 53225 -13060
rect 53345 -13180 53355 -13060
rect 47855 -13225 53355 -13180
rect 47855 -13345 47865 -13225
rect 47985 -13345 48040 -13225
rect 48160 -13345 48205 -13225
rect 48325 -13345 48370 -13225
rect 48490 -13345 48535 -13225
rect 48655 -13345 48710 -13225
rect 48830 -13345 48875 -13225
rect 48995 -13345 49040 -13225
rect 49160 -13345 49205 -13225
rect 49325 -13345 49380 -13225
rect 49500 -13345 49545 -13225
rect 49665 -13345 49710 -13225
rect 49830 -13345 49875 -13225
rect 49995 -13345 50050 -13225
rect 50170 -13345 50215 -13225
rect 50335 -13345 50380 -13225
rect 50500 -13345 50545 -13225
rect 50665 -13345 50720 -13225
rect 50840 -13345 50885 -13225
rect 51005 -13345 51050 -13225
rect 51170 -13345 51215 -13225
rect 51335 -13345 51390 -13225
rect 51510 -13345 51555 -13225
rect 51675 -13345 51720 -13225
rect 51840 -13345 51885 -13225
rect 52005 -13345 52060 -13225
rect 52180 -13345 52225 -13225
rect 52345 -13345 52390 -13225
rect 52510 -13345 52555 -13225
rect 52675 -13345 52730 -13225
rect 52850 -13345 52895 -13225
rect 53015 -13345 53060 -13225
rect 53180 -13345 53225 -13225
rect 53345 -13345 53355 -13225
rect 47855 -13400 53355 -13345
rect 47855 -13520 47865 -13400
rect 47985 -13520 48040 -13400
rect 48160 -13520 48205 -13400
rect 48325 -13520 48370 -13400
rect 48490 -13520 48535 -13400
rect 48655 -13520 48710 -13400
rect 48830 -13520 48875 -13400
rect 48995 -13520 49040 -13400
rect 49160 -13520 49205 -13400
rect 49325 -13520 49380 -13400
rect 49500 -13520 49545 -13400
rect 49665 -13520 49710 -13400
rect 49830 -13520 49875 -13400
rect 49995 -13520 50050 -13400
rect 50170 -13520 50215 -13400
rect 50335 -13520 50380 -13400
rect 50500 -13520 50545 -13400
rect 50665 -13520 50720 -13400
rect 50840 -13520 50885 -13400
rect 51005 -13520 51050 -13400
rect 51170 -13520 51215 -13400
rect 51335 -13520 51390 -13400
rect 51510 -13520 51555 -13400
rect 51675 -13520 51720 -13400
rect 51840 -13520 51885 -13400
rect 52005 -13520 52060 -13400
rect 52180 -13520 52225 -13400
rect 52345 -13520 52390 -13400
rect 52510 -13520 52555 -13400
rect 52675 -13520 52730 -13400
rect 52850 -13520 52895 -13400
rect 53015 -13520 53060 -13400
rect 53180 -13520 53225 -13400
rect 53345 -13520 53355 -13400
rect 47855 -13565 53355 -13520
rect 47855 -13685 47865 -13565
rect 47985 -13685 48040 -13565
rect 48160 -13685 48205 -13565
rect 48325 -13685 48370 -13565
rect 48490 -13685 48535 -13565
rect 48655 -13685 48710 -13565
rect 48830 -13685 48875 -13565
rect 48995 -13685 49040 -13565
rect 49160 -13685 49205 -13565
rect 49325 -13685 49380 -13565
rect 49500 -13685 49545 -13565
rect 49665 -13685 49710 -13565
rect 49830 -13685 49875 -13565
rect 49995 -13685 50050 -13565
rect 50170 -13685 50215 -13565
rect 50335 -13685 50380 -13565
rect 50500 -13685 50545 -13565
rect 50665 -13685 50720 -13565
rect 50840 -13685 50885 -13565
rect 51005 -13685 51050 -13565
rect 51170 -13685 51215 -13565
rect 51335 -13685 51390 -13565
rect 51510 -13685 51555 -13565
rect 51675 -13685 51720 -13565
rect 51840 -13685 51885 -13565
rect 52005 -13685 52060 -13565
rect 52180 -13685 52225 -13565
rect 52345 -13685 52390 -13565
rect 52510 -13685 52555 -13565
rect 52675 -13685 52730 -13565
rect 52850 -13685 52895 -13565
rect 53015 -13685 53060 -13565
rect 53180 -13685 53225 -13565
rect 53345 -13685 53355 -13565
rect 47855 -13730 53355 -13685
rect 47855 -13850 47865 -13730
rect 47985 -13850 48040 -13730
rect 48160 -13850 48205 -13730
rect 48325 -13850 48370 -13730
rect 48490 -13850 48535 -13730
rect 48655 -13850 48710 -13730
rect 48830 -13850 48875 -13730
rect 48995 -13850 49040 -13730
rect 49160 -13850 49205 -13730
rect 49325 -13850 49380 -13730
rect 49500 -13850 49545 -13730
rect 49665 -13850 49710 -13730
rect 49830 -13850 49875 -13730
rect 49995 -13850 50050 -13730
rect 50170 -13850 50215 -13730
rect 50335 -13850 50380 -13730
rect 50500 -13850 50545 -13730
rect 50665 -13850 50720 -13730
rect 50840 -13850 50885 -13730
rect 51005 -13850 51050 -13730
rect 51170 -13850 51215 -13730
rect 51335 -13850 51390 -13730
rect 51510 -13850 51555 -13730
rect 51675 -13850 51720 -13730
rect 51840 -13850 51885 -13730
rect 52005 -13850 52060 -13730
rect 52180 -13850 52225 -13730
rect 52345 -13850 52390 -13730
rect 52510 -13850 52555 -13730
rect 52675 -13850 52730 -13730
rect 52850 -13850 52895 -13730
rect 53015 -13850 53060 -13730
rect 53180 -13850 53225 -13730
rect 53345 -13850 53355 -13730
rect 47855 -13895 53355 -13850
rect 47855 -14015 47865 -13895
rect 47985 -14015 48040 -13895
rect 48160 -14015 48205 -13895
rect 48325 -14015 48370 -13895
rect 48490 -14015 48535 -13895
rect 48655 -14015 48710 -13895
rect 48830 -14015 48875 -13895
rect 48995 -14015 49040 -13895
rect 49160 -14015 49205 -13895
rect 49325 -14015 49380 -13895
rect 49500 -14015 49545 -13895
rect 49665 -14015 49710 -13895
rect 49830 -14015 49875 -13895
rect 49995 -14015 50050 -13895
rect 50170 -14015 50215 -13895
rect 50335 -14015 50380 -13895
rect 50500 -14015 50545 -13895
rect 50665 -14015 50720 -13895
rect 50840 -14015 50885 -13895
rect 51005 -14015 51050 -13895
rect 51170 -14015 51215 -13895
rect 51335 -14015 51390 -13895
rect 51510 -14015 51555 -13895
rect 51675 -14015 51720 -13895
rect 51840 -14015 51885 -13895
rect 52005 -14015 52060 -13895
rect 52180 -14015 52225 -13895
rect 52345 -14015 52390 -13895
rect 52510 -14015 52555 -13895
rect 52675 -14015 52730 -13895
rect 52850 -14015 52895 -13895
rect 53015 -14015 53060 -13895
rect 53180 -14015 53225 -13895
rect 53345 -14015 53355 -13895
rect 47855 -14070 53355 -14015
rect 47855 -14190 47865 -14070
rect 47985 -14190 48040 -14070
rect 48160 -14190 48205 -14070
rect 48325 -14190 48370 -14070
rect 48490 -14190 48535 -14070
rect 48655 -14190 48710 -14070
rect 48830 -14190 48875 -14070
rect 48995 -14190 49040 -14070
rect 49160 -14190 49205 -14070
rect 49325 -14190 49380 -14070
rect 49500 -14190 49545 -14070
rect 49665 -14190 49710 -14070
rect 49830 -14190 49875 -14070
rect 49995 -14190 50050 -14070
rect 50170 -14190 50215 -14070
rect 50335 -14190 50380 -14070
rect 50500 -14190 50545 -14070
rect 50665 -14190 50720 -14070
rect 50840 -14190 50885 -14070
rect 51005 -14190 51050 -14070
rect 51170 -14190 51215 -14070
rect 51335 -14190 51390 -14070
rect 51510 -14190 51555 -14070
rect 51675 -14190 51720 -14070
rect 51840 -14190 51885 -14070
rect 52005 -14190 52060 -14070
rect 52180 -14190 52225 -14070
rect 52345 -14190 52390 -14070
rect 52510 -14190 52555 -14070
rect 52675 -14190 52730 -14070
rect 52850 -14190 52895 -14070
rect 53015 -14190 53060 -14070
rect 53180 -14190 53225 -14070
rect 53345 -14190 53355 -14070
rect 47855 -14235 53355 -14190
rect 47855 -14355 47865 -14235
rect 47985 -14355 48040 -14235
rect 48160 -14355 48205 -14235
rect 48325 -14355 48370 -14235
rect 48490 -14355 48535 -14235
rect 48655 -14355 48710 -14235
rect 48830 -14355 48875 -14235
rect 48995 -14355 49040 -14235
rect 49160 -14355 49205 -14235
rect 49325 -14355 49380 -14235
rect 49500 -14355 49545 -14235
rect 49665 -14355 49710 -14235
rect 49830 -14355 49875 -14235
rect 49995 -14355 50050 -14235
rect 50170 -14355 50215 -14235
rect 50335 -14355 50380 -14235
rect 50500 -14355 50545 -14235
rect 50665 -14355 50720 -14235
rect 50840 -14355 50885 -14235
rect 51005 -14355 51050 -14235
rect 51170 -14355 51215 -14235
rect 51335 -14355 51390 -14235
rect 51510 -14355 51555 -14235
rect 51675 -14355 51720 -14235
rect 51840 -14355 51885 -14235
rect 52005 -14355 52060 -14235
rect 52180 -14355 52225 -14235
rect 52345 -14355 52390 -14235
rect 52510 -14355 52555 -14235
rect 52675 -14355 52730 -14235
rect 52850 -14355 52895 -14235
rect 53015 -14355 53060 -14235
rect 53180 -14355 53225 -14235
rect 53345 -14355 53355 -14235
rect 47855 -14400 53355 -14355
rect 47855 -14520 47865 -14400
rect 47985 -14520 48040 -14400
rect 48160 -14520 48205 -14400
rect 48325 -14520 48370 -14400
rect 48490 -14520 48535 -14400
rect 48655 -14520 48710 -14400
rect 48830 -14520 48875 -14400
rect 48995 -14520 49040 -14400
rect 49160 -14520 49205 -14400
rect 49325 -14520 49380 -14400
rect 49500 -14520 49545 -14400
rect 49665 -14520 49710 -14400
rect 49830 -14520 49875 -14400
rect 49995 -14520 50050 -14400
rect 50170 -14520 50215 -14400
rect 50335 -14520 50380 -14400
rect 50500 -14520 50545 -14400
rect 50665 -14520 50720 -14400
rect 50840 -14520 50885 -14400
rect 51005 -14520 51050 -14400
rect 51170 -14520 51215 -14400
rect 51335 -14520 51390 -14400
rect 51510 -14520 51555 -14400
rect 51675 -14520 51720 -14400
rect 51840 -14520 51885 -14400
rect 52005 -14520 52060 -14400
rect 52180 -14520 52225 -14400
rect 52345 -14520 52390 -14400
rect 52510 -14520 52555 -14400
rect 52675 -14520 52730 -14400
rect 52850 -14520 52895 -14400
rect 53015 -14520 53060 -14400
rect 53180 -14520 53225 -14400
rect 53345 -14520 53355 -14400
rect 47855 -14565 53355 -14520
rect 47855 -14685 47865 -14565
rect 47985 -14685 48040 -14565
rect 48160 -14685 48205 -14565
rect 48325 -14685 48370 -14565
rect 48490 -14685 48535 -14565
rect 48655 -14685 48710 -14565
rect 48830 -14685 48875 -14565
rect 48995 -14685 49040 -14565
rect 49160 -14685 49205 -14565
rect 49325 -14685 49380 -14565
rect 49500 -14685 49545 -14565
rect 49665 -14685 49710 -14565
rect 49830 -14685 49875 -14565
rect 49995 -14685 50050 -14565
rect 50170 -14685 50215 -14565
rect 50335 -14685 50380 -14565
rect 50500 -14685 50545 -14565
rect 50665 -14685 50720 -14565
rect 50840 -14685 50885 -14565
rect 51005 -14685 51050 -14565
rect 51170 -14685 51215 -14565
rect 51335 -14685 51390 -14565
rect 51510 -14685 51555 -14565
rect 51675 -14685 51720 -14565
rect 51840 -14685 51885 -14565
rect 52005 -14685 52060 -14565
rect 52180 -14685 52225 -14565
rect 52345 -14685 52390 -14565
rect 52510 -14685 52555 -14565
rect 52675 -14685 52730 -14565
rect 52850 -14685 52895 -14565
rect 53015 -14685 53060 -14565
rect 53180 -14685 53225 -14565
rect 53345 -14685 53355 -14565
rect 47855 -14740 53355 -14685
rect 47855 -14860 47865 -14740
rect 47985 -14860 48040 -14740
rect 48160 -14860 48205 -14740
rect 48325 -14860 48370 -14740
rect 48490 -14860 48535 -14740
rect 48655 -14860 48710 -14740
rect 48830 -14860 48875 -14740
rect 48995 -14860 49040 -14740
rect 49160 -14860 49205 -14740
rect 49325 -14860 49380 -14740
rect 49500 -14860 49545 -14740
rect 49665 -14860 49710 -14740
rect 49830 -14860 49875 -14740
rect 49995 -14860 50050 -14740
rect 50170 -14860 50215 -14740
rect 50335 -14860 50380 -14740
rect 50500 -14860 50545 -14740
rect 50665 -14860 50720 -14740
rect 50840 -14860 50885 -14740
rect 51005 -14860 51050 -14740
rect 51170 -14860 51215 -14740
rect 51335 -14860 51390 -14740
rect 51510 -14860 51555 -14740
rect 51675 -14860 51720 -14740
rect 51840 -14860 51885 -14740
rect 52005 -14860 52060 -14740
rect 52180 -14860 52225 -14740
rect 52345 -14860 52390 -14740
rect 52510 -14860 52555 -14740
rect 52675 -14860 52730 -14740
rect 52850 -14860 52895 -14740
rect 53015 -14860 53060 -14740
rect 53180 -14860 53225 -14740
rect 53345 -14860 53355 -14740
rect 47855 -14905 53355 -14860
rect 47855 -15025 47865 -14905
rect 47985 -15025 48040 -14905
rect 48160 -15025 48205 -14905
rect 48325 -15025 48370 -14905
rect 48490 -15025 48535 -14905
rect 48655 -15025 48710 -14905
rect 48830 -15025 48875 -14905
rect 48995 -15025 49040 -14905
rect 49160 -15025 49205 -14905
rect 49325 -15025 49380 -14905
rect 49500 -15025 49545 -14905
rect 49665 -15025 49710 -14905
rect 49830 -15025 49875 -14905
rect 49995 -15025 50050 -14905
rect 50170 -15025 50215 -14905
rect 50335 -15025 50380 -14905
rect 50500 -15025 50545 -14905
rect 50665 -15025 50720 -14905
rect 50840 -15025 50885 -14905
rect 51005 -15025 51050 -14905
rect 51170 -15025 51215 -14905
rect 51335 -15025 51390 -14905
rect 51510 -15025 51555 -14905
rect 51675 -15025 51720 -14905
rect 51840 -15025 51885 -14905
rect 52005 -15025 52060 -14905
rect 52180 -15025 52225 -14905
rect 52345 -15025 52390 -14905
rect 52510 -15025 52555 -14905
rect 52675 -15025 52730 -14905
rect 52850 -15025 52895 -14905
rect 53015 -15025 53060 -14905
rect 53180 -15025 53225 -14905
rect 53345 -15025 53355 -14905
rect 47855 -15070 53355 -15025
rect 47855 -15190 47865 -15070
rect 47985 -15190 48040 -15070
rect 48160 -15190 48205 -15070
rect 48325 -15190 48370 -15070
rect 48490 -15190 48535 -15070
rect 48655 -15190 48710 -15070
rect 48830 -15190 48875 -15070
rect 48995 -15190 49040 -15070
rect 49160 -15190 49205 -15070
rect 49325 -15190 49380 -15070
rect 49500 -15190 49545 -15070
rect 49665 -15190 49710 -15070
rect 49830 -15190 49875 -15070
rect 49995 -15190 50050 -15070
rect 50170 -15190 50215 -15070
rect 50335 -15190 50380 -15070
rect 50500 -15190 50545 -15070
rect 50665 -15190 50720 -15070
rect 50840 -15190 50885 -15070
rect 51005 -15190 51050 -15070
rect 51170 -15190 51215 -15070
rect 51335 -15190 51390 -15070
rect 51510 -15190 51555 -15070
rect 51675 -15190 51720 -15070
rect 51840 -15190 51885 -15070
rect 52005 -15190 52060 -15070
rect 52180 -15190 52225 -15070
rect 52345 -15190 52390 -15070
rect 52510 -15190 52555 -15070
rect 52675 -15190 52730 -15070
rect 52850 -15190 52895 -15070
rect 53015 -15190 53060 -15070
rect 53180 -15190 53225 -15070
rect 53345 -15190 53355 -15070
rect 47855 -15235 53355 -15190
rect 47855 -15355 47865 -15235
rect 47985 -15355 48040 -15235
rect 48160 -15355 48205 -15235
rect 48325 -15355 48370 -15235
rect 48490 -15355 48535 -15235
rect 48655 -15355 48710 -15235
rect 48830 -15355 48875 -15235
rect 48995 -15355 49040 -15235
rect 49160 -15355 49205 -15235
rect 49325 -15355 49380 -15235
rect 49500 -15355 49545 -15235
rect 49665 -15355 49710 -15235
rect 49830 -15355 49875 -15235
rect 49995 -15355 50050 -15235
rect 50170 -15355 50215 -15235
rect 50335 -15355 50380 -15235
rect 50500 -15355 50545 -15235
rect 50665 -15355 50720 -15235
rect 50840 -15355 50885 -15235
rect 51005 -15355 51050 -15235
rect 51170 -15355 51215 -15235
rect 51335 -15355 51390 -15235
rect 51510 -15355 51555 -15235
rect 51675 -15355 51720 -15235
rect 51840 -15355 51885 -15235
rect 52005 -15355 52060 -15235
rect 52180 -15355 52225 -15235
rect 52345 -15355 52390 -15235
rect 52510 -15355 52555 -15235
rect 52675 -15355 52730 -15235
rect 52850 -15355 52895 -15235
rect 53015 -15355 53060 -15235
rect 53180 -15355 53225 -15235
rect 53345 -15355 53355 -15235
rect 47855 -15410 53355 -15355
rect 47855 -15530 47865 -15410
rect 47985 -15530 48040 -15410
rect 48160 -15530 48205 -15410
rect 48325 -15530 48370 -15410
rect 48490 -15530 48535 -15410
rect 48655 -15530 48710 -15410
rect 48830 -15530 48875 -15410
rect 48995 -15530 49040 -15410
rect 49160 -15530 49205 -15410
rect 49325 -15530 49380 -15410
rect 49500 -15530 49545 -15410
rect 49665 -15530 49710 -15410
rect 49830 -15530 49875 -15410
rect 49995 -15530 50050 -15410
rect 50170 -15530 50215 -15410
rect 50335 -15530 50380 -15410
rect 50500 -15530 50545 -15410
rect 50665 -15530 50720 -15410
rect 50840 -15530 50885 -15410
rect 51005 -15530 51050 -15410
rect 51170 -15530 51215 -15410
rect 51335 -15530 51390 -15410
rect 51510 -15530 51555 -15410
rect 51675 -15530 51720 -15410
rect 51840 -15530 51885 -15410
rect 52005 -15530 52060 -15410
rect 52180 -15530 52225 -15410
rect 52345 -15530 52390 -15410
rect 52510 -15530 52555 -15410
rect 52675 -15530 52730 -15410
rect 52850 -15530 52895 -15410
rect 53015 -15530 53060 -15410
rect 53180 -15530 53225 -15410
rect 53345 -15530 53355 -15410
rect 47855 -15540 53355 -15530
<< mimcap2contact >>
rect 30795 7080 30915 7200
rect 30960 7080 31080 7200
rect 31125 7080 31245 7200
rect 31290 7080 31410 7200
rect 31465 7080 31585 7200
rect 31630 7080 31750 7200
rect 31795 7080 31915 7200
rect 31960 7080 32080 7200
rect 32135 7080 32255 7200
rect 32300 7080 32420 7200
rect 32465 7080 32585 7200
rect 32630 7080 32750 7200
rect 32805 7080 32925 7200
rect 32970 7080 33090 7200
rect 33135 7080 33255 7200
rect 33300 7080 33420 7200
rect 33475 7080 33595 7200
rect 33640 7080 33760 7200
rect 33805 7080 33925 7200
rect 33970 7080 34090 7200
rect 34145 7080 34265 7200
rect 34310 7080 34430 7200
rect 34475 7080 34595 7200
rect 34640 7080 34760 7200
rect 34815 7080 34935 7200
rect 34980 7080 35100 7200
rect 35145 7080 35265 7200
rect 35310 7080 35430 7200
rect 35485 7080 35605 7200
rect 35650 7080 35770 7200
rect 35815 7080 35935 7200
rect 35980 7080 36100 7200
rect 36155 7080 36275 7200
rect 30795 6905 30915 7025
rect 30960 6905 31080 7025
rect 31125 6905 31245 7025
rect 31290 6905 31410 7025
rect 31465 6905 31585 7025
rect 31630 6905 31750 7025
rect 31795 6905 31915 7025
rect 31960 6905 32080 7025
rect 32135 6905 32255 7025
rect 32300 6905 32420 7025
rect 32465 6905 32585 7025
rect 32630 6905 32750 7025
rect 32805 6905 32925 7025
rect 32970 6905 33090 7025
rect 33135 6905 33255 7025
rect 33300 6905 33420 7025
rect 33475 6905 33595 7025
rect 33640 6905 33760 7025
rect 33805 6905 33925 7025
rect 33970 6905 34090 7025
rect 34145 6905 34265 7025
rect 34310 6905 34430 7025
rect 34475 6905 34595 7025
rect 34640 6905 34760 7025
rect 34815 6905 34935 7025
rect 34980 6905 35100 7025
rect 35145 6905 35265 7025
rect 35310 6905 35430 7025
rect 35485 6905 35605 7025
rect 35650 6905 35770 7025
rect 35815 6905 35935 7025
rect 35980 6905 36100 7025
rect 36155 6905 36275 7025
rect 30795 6740 30915 6860
rect 30960 6740 31080 6860
rect 31125 6740 31245 6860
rect 31290 6740 31410 6860
rect 31465 6740 31585 6860
rect 31630 6740 31750 6860
rect 31795 6740 31915 6860
rect 31960 6740 32080 6860
rect 32135 6740 32255 6860
rect 32300 6740 32420 6860
rect 32465 6740 32585 6860
rect 32630 6740 32750 6860
rect 32805 6740 32925 6860
rect 32970 6740 33090 6860
rect 33135 6740 33255 6860
rect 33300 6740 33420 6860
rect 33475 6740 33595 6860
rect 33640 6740 33760 6860
rect 33805 6740 33925 6860
rect 33970 6740 34090 6860
rect 34145 6740 34265 6860
rect 34310 6740 34430 6860
rect 34475 6740 34595 6860
rect 34640 6740 34760 6860
rect 34815 6740 34935 6860
rect 34980 6740 35100 6860
rect 35145 6740 35265 6860
rect 35310 6740 35430 6860
rect 35485 6740 35605 6860
rect 35650 6740 35770 6860
rect 35815 6740 35935 6860
rect 35980 6740 36100 6860
rect 36155 6740 36275 6860
rect 30795 6575 30915 6695
rect 30960 6575 31080 6695
rect 31125 6575 31245 6695
rect 31290 6575 31410 6695
rect 31465 6575 31585 6695
rect 31630 6575 31750 6695
rect 31795 6575 31915 6695
rect 31960 6575 32080 6695
rect 32135 6575 32255 6695
rect 32300 6575 32420 6695
rect 32465 6575 32585 6695
rect 32630 6575 32750 6695
rect 32805 6575 32925 6695
rect 32970 6575 33090 6695
rect 33135 6575 33255 6695
rect 33300 6575 33420 6695
rect 33475 6575 33595 6695
rect 33640 6575 33760 6695
rect 33805 6575 33925 6695
rect 33970 6575 34090 6695
rect 34145 6575 34265 6695
rect 34310 6575 34430 6695
rect 34475 6575 34595 6695
rect 34640 6575 34760 6695
rect 34815 6575 34935 6695
rect 34980 6575 35100 6695
rect 35145 6575 35265 6695
rect 35310 6575 35430 6695
rect 35485 6575 35605 6695
rect 35650 6575 35770 6695
rect 35815 6575 35935 6695
rect 35980 6575 36100 6695
rect 36155 6575 36275 6695
rect 30795 6410 30915 6530
rect 30960 6410 31080 6530
rect 31125 6410 31245 6530
rect 31290 6410 31410 6530
rect 31465 6410 31585 6530
rect 31630 6410 31750 6530
rect 31795 6410 31915 6530
rect 31960 6410 32080 6530
rect 32135 6410 32255 6530
rect 32300 6410 32420 6530
rect 32465 6410 32585 6530
rect 32630 6410 32750 6530
rect 32805 6410 32925 6530
rect 32970 6410 33090 6530
rect 33135 6410 33255 6530
rect 33300 6410 33420 6530
rect 33475 6410 33595 6530
rect 33640 6410 33760 6530
rect 33805 6410 33925 6530
rect 33970 6410 34090 6530
rect 34145 6410 34265 6530
rect 34310 6410 34430 6530
rect 34475 6410 34595 6530
rect 34640 6410 34760 6530
rect 34815 6410 34935 6530
rect 34980 6410 35100 6530
rect 35145 6410 35265 6530
rect 35310 6410 35430 6530
rect 35485 6410 35605 6530
rect 35650 6410 35770 6530
rect 35815 6410 35935 6530
rect 35980 6410 36100 6530
rect 36155 6410 36275 6530
rect 30795 6235 30915 6355
rect 30960 6235 31080 6355
rect 31125 6235 31245 6355
rect 31290 6235 31410 6355
rect 31465 6235 31585 6355
rect 31630 6235 31750 6355
rect 31795 6235 31915 6355
rect 31960 6235 32080 6355
rect 32135 6235 32255 6355
rect 32300 6235 32420 6355
rect 32465 6235 32585 6355
rect 32630 6235 32750 6355
rect 32805 6235 32925 6355
rect 32970 6235 33090 6355
rect 33135 6235 33255 6355
rect 33300 6235 33420 6355
rect 33475 6235 33595 6355
rect 33640 6235 33760 6355
rect 33805 6235 33925 6355
rect 33970 6235 34090 6355
rect 34145 6235 34265 6355
rect 34310 6235 34430 6355
rect 34475 6235 34595 6355
rect 34640 6235 34760 6355
rect 34815 6235 34935 6355
rect 34980 6235 35100 6355
rect 35145 6235 35265 6355
rect 35310 6235 35430 6355
rect 35485 6235 35605 6355
rect 35650 6235 35770 6355
rect 35815 6235 35935 6355
rect 35980 6235 36100 6355
rect 36155 6235 36275 6355
rect 30795 6070 30915 6190
rect 30960 6070 31080 6190
rect 31125 6070 31245 6190
rect 31290 6070 31410 6190
rect 31465 6070 31585 6190
rect 31630 6070 31750 6190
rect 31795 6070 31915 6190
rect 31960 6070 32080 6190
rect 32135 6070 32255 6190
rect 32300 6070 32420 6190
rect 32465 6070 32585 6190
rect 32630 6070 32750 6190
rect 32805 6070 32925 6190
rect 32970 6070 33090 6190
rect 33135 6070 33255 6190
rect 33300 6070 33420 6190
rect 33475 6070 33595 6190
rect 33640 6070 33760 6190
rect 33805 6070 33925 6190
rect 33970 6070 34090 6190
rect 34145 6070 34265 6190
rect 34310 6070 34430 6190
rect 34475 6070 34595 6190
rect 34640 6070 34760 6190
rect 34815 6070 34935 6190
rect 34980 6070 35100 6190
rect 35145 6070 35265 6190
rect 35310 6070 35430 6190
rect 35485 6070 35605 6190
rect 35650 6070 35770 6190
rect 35815 6070 35935 6190
rect 35980 6070 36100 6190
rect 36155 6070 36275 6190
rect 30795 5905 30915 6025
rect 30960 5905 31080 6025
rect 31125 5905 31245 6025
rect 31290 5905 31410 6025
rect 31465 5905 31585 6025
rect 31630 5905 31750 6025
rect 31795 5905 31915 6025
rect 31960 5905 32080 6025
rect 32135 5905 32255 6025
rect 32300 5905 32420 6025
rect 32465 5905 32585 6025
rect 32630 5905 32750 6025
rect 32805 5905 32925 6025
rect 32970 5905 33090 6025
rect 33135 5905 33255 6025
rect 33300 5905 33420 6025
rect 33475 5905 33595 6025
rect 33640 5905 33760 6025
rect 33805 5905 33925 6025
rect 33970 5905 34090 6025
rect 34145 5905 34265 6025
rect 34310 5905 34430 6025
rect 34475 5905 34595 6025
rect 34640 5905 34760 6025
rect 34815 5905 34935 6025
rect 34980 5905 35100 6025
rect 35145 5905 35265 6025
rect 35310 5905 35430 6025
rect 35485 5905 35605 6025
rect 35650 5905 35770 6025
rect 35815 5905 35935 6025
rect 35980 5905 36100 6025
rect 36155 5905 36275 6025
rect 30795 5740 30915 5860
rect 30960 5740 31080 5860
rect 31125 5740 31245 5860
rect 31290 5740 31410 5860
rect 31465 5740 31585 5860
rect 31630 5740 31750 5860
rect 31795 5740 31915 5860
rect 31960 5740 32080 5860
rect 32135 5740 32255 5860
rect 32300 5740 32420 5860
rect 32465 5740 32585 5860
rect 32630 5740 32750 5860
rect 32805 5740 32925 5860
rect 32970 5740 33090 5860
rect 33135 5740 33255 5860
rect 33300 5740 33420 5860
rect 33475 5740 33595 5860
rect 33640 5740 33760 5860
rect 33805 5740 33925 5860
rect 33970 5740 34090 5860
rect 34145 5740 34265 5860
rect 34310 5740 34430 5860
rect 34475 5740 34595 5860
rect 34640 5740 34760 5860
rect 34815 5740 34935 5860
rect 34980 5740 35100 5860
rect 35145 5740 35265 5860
rect 35310 5740 35430 5860
rect 35485 5740 35605 5860
rect 35650 5740 35770 5860
rect 35815 5740 35935 5860
rect 35980 5740 36100 5860
rect 36155 5740 36275 5860
rect 30795 5565 30915 5685
rect 30960 5565 31080 5685
rect 31125 5565 31245 5685
rect 31290 5565 31410 5685
rect 31465 5565 31585 5685
rect 31630 5565 31750 5685
rect 31795 5565 31915 5685
rect 31960 5565 32080 5685
rect 32135 5565 32255 5685
rect 32300 5565 32420 5685
rect 32465 5565 32585 5685
rect 32630 5565 32750 5685
rect 32805 5565 32925 5685
rect 32970 5565 33090 5685
rect 33135 5565 33255 5685
rect 33300 5565 33420 5685
rect 33475 5565 33595 5685
rect 33640 5565 33760 5685
rect 33805 5565 33925 5685
rect 33970 5565 34090 5685
rect 34145 5565 34265 5685
rect 34310 5565 34430 5685
rect 34475 5565 34595 5685
rect 34640 5565 34760 5685
rect 34815 5565 34935 5685
rect 34980 5565 35100 5685
rect 35145 5565 35265 5685
rect 35310 5565 35430 5685
rect 35485 5565 35605 5685
rect 35650 5565 35770 5685
rect 35815 5565 35935 5685
rect 35980 5565 36100 5685
rect 36155 5565 36275 5685
rect 30795 5400 30915 5520
rect 30960 5400 31080 5520
rect 31125 5400 31245 5520
rect 31290 5400 31410 5520
rect 31465 5400 31585 5520
rect 31630 5400 31750 5520
rect 31795 5400 31915 5520
rect 31960 5400 32080 5520
rect 32135 5400 32255 5520
rect 32300 5400 32420 5520
rect 32465 5400 32585 5520
rect 32630 5400 32750 5520
rect 32805 5400 32925 5520
rect 32970 5400 33090 5520
rect 33135 5400 33255 5520
rect 33300 5400 33420 5520
rect 33475 5400 33595 5520
rect 33640 5400 33760 5520
rect 33805 5400 33925 5520
rect 33970 5400 34090 5520
rect 34145 5400 34265 5520
rect 34310 5400 34430 5520
rect 34475 5400 34595 5520
rect 34640 5400 34760 5520
rect 34815 5400 34935 5520
rect 34980 5400 35100 5520
rect 35145 5400 35265 5520
rect 35310 5400 35430 5520
rect 35485 5400 35605 5520
rect 35650 5400 35770 5520
rect 35815 5400 35935 5520
rect 35980 5400 36100 5520
rect 36155 5400 36275 5520
rect 30795 5235 30915 5355
rect 30960 5235 31080 5355
rect 31125 5235 31245 5355
rect 31290 5235 31410 5355
rect 31465 5235 31585 5355
rect 31630 5235 31750 5355
rect 31795 5235 31915 5355
rect 31960 5235 32080 5355
rect 32135 5235 32255 5355
rect 32300 5235 32420 5355
rect 32465 5235 32585 5355
rect 32630 5235 32750 5355
rect 32805 5235 32925 5355
rect 32970 5235 33090 5355
rect 33135 5235 33255 5355
rect 33300 5235 33420 5355
rect 33475 5235 33595 5355
rect 33640 5235 33760 5355
rect 33805 5235 33925 5355
rect 33970 5235 34090 5355
rect 34145 5235 34265 5355
rect 34310 5235 34430 5355
rect 34475 5235 34595 5355
rect 34640 5235 34760 5355
rect 34815 5235 34935 5355
rect 34980 5235 35100 5355
rect 35145 5235 35265 5355
rect 35310 5235 35430 5355
rect 35485 5235 35605 5355
rect 35650 5235 35770 5355
rect 35815 5235 35935 5355
rect 35980 5235 36100 5355
rect 36155 5235 36275 5355
rect 30795 5070 30915 5190
rect 30960 5070 31080 5190
rect 31125 5070 31245 5190
rect 31290 5070 31410 5190
rect 31465 5070 31585 5190
rect 31630 5070 31750 5190
rect 31795 5070 31915 5190
rect 31960 5070 32080 5190
rect 32135 5070 32255 5190
rect 32300 5070 32420 5190
rect 32465 5070 32585 5190
rect 32630 5070 32750 5190
rect 32805 5070 32925 5190
rect 32970 5070 33090 5190
rect 33135 5070 33255 5190
rect 33300 5070 33420 5190
rect 33475 5070 33595 5190
rect 33640 5070 33760 5190
rect 33805 5070 33925 5190
rect 33970 5070 34090 5190
rect 34145 5070 34265 5190
rect 34310 5070 34430 5190
rect 34475 5070 34595 5190
rect 34640 5070 34760 5190
rect 34815 5070 34935 5190
rect 34980 5070 35100 5190
rect 35145 5070 35265 5190
rect 35310 5070 35430 5190
rect 35485 5070 35605 5190
rect 35650 5070 35770 5190
rect 35815 5070 35935 5190
rect 35980 5070 36100 5190
rect 36155 5070 36275 5190
rect 30795 4895 30915 5015
rect 30960 4895 31080 5015
rect 31125 4895 31245 5015
rect 31290 4895 31410 5015
rect 31465 4895 31585 5015
rect 31630 4895 31750 5015
rect 31795 4895 31915 5015
rect 31960 4895 32080 5015
rect 32135 4895 32255 5015
rect 32300 4895 32420 5015
rect 32465 4895 32585 5015
rect 32630 4895 32750 5015
rect 32805 4895 32925 5015
rect 32970 4895 33090 5015
rect 33135 4895 33255 5015
rect 33300 4895 33420 5015
rect 33475 4895 33595 5015
rect 33640 4895 33760 5015
rect 33805 4895 33925 5015
rect 33970 4895 34090 5015
rect 34145 4895 34265 5015
rect 34310 4895 34430 5015
rect 34475 4895 34595 5015
rect 34640 4895 34760 5015
rect 34815 4895 34935 5015
rect 34980 4895 35100 5015
rect 35145 4895 35265 5015
rect 35310 4895 35430 5015
rect 35485 4895 35605 5015
rect 35650 4895 35770 5015
rect 35815 4895 35935 5015
rect 35980 4895 36100 5015
rect 36155 4895 36275 5015
rect 30795 4730 30915 4850
rect 30960 4730 31080 4850
rect 31125 4730 31245 4850
rect 31290 4730 31410 4850
rect 31465 4730 31585 4850
rect 31630 4730 31750 4850
rect 31795 4730 31915 4850
rect 31960 4730 32080 4850
rect 32135 4730 32255 4850
rect 32300 4730 32420 4850
rect 32465 4730 32585 4850
rect 32630 4730 32750 4850
rect 32805 4730 32925 4850
rect 32970 4730 33090 4850
rect 33135 4730 33255 4850
rect 33300 4730 33420 4850
rect 33475 4730 33595 4850
rect 33640 4730 33760 4850
rect 33805 4730 33925 4850
rect 33970 4730 34090 4850
rect 34145 4730 34265 4850
rect 34310 4730 34430 4850
rect 34475 4730 34595 4850
rect 34640 4730 34760 4850
rect 34815 4730 34935 4850
rect 34980 4730 35100 4850
rect 35145 4730 35265 4850
rect 35310 4730 35430 4850
rect 35485 4730 35605 4850
rect 35650 4730 35770 4850
rect 35815 4730 35935 4850
rect 35980 4730 36100 4850
rect 36155 4730 36275 4850
rect 30795 4565 30915 4685
rect 30960 4565 31080 4685
rect 31125 4565 31245 4685
rect 31290 4565 31410 4685
rect 31465 4565 31585 4685
rect 31630 4565 31750 4685
rect 31795 4565 31915 4685
rect 31960 4565 32080 4685
rect 32135 4565 32255 4685
rect 32300 4565 32420 4685
rect 32465 4565 32585 4685
rect 32630 4565 32750 4685
rect 32805 4565 32925 4685
rect 32970 4565 33090 4685
rect 33135 4565 33255 4685
rect 33300 4565 33420 4685
rect 33475 4565 33595 4685
rect 33640 4565 33760 4685
rect 33805 4565 33925 4685
rect 33970 4565 34090 4685
rect 34145 4565 34265 4685
rect 34310 4565 34430 4685
rect 34475 4565 34595 4685
rect 34640 4565 34760 4685
rect 34815 4565 34935 4685
rect 34980 4565 35100 4685
rect 35145 4565 35265 4685
rect 35310 4565 35430 4685
rect 35485 4565 35605 4685
rect 35650 4565 35770 4685
rect 35815 4565 35935 4685
rect 35980 4565 36100 4685
rect 36155 4565 36275 4685
rect 30795 4400 30915 4520
rect 30960 4400 31080 4520
rect 31125 4400 31245 4520
rect 31290 4400 31410 4520
rect 31465 4400 31585 4520
rect 31630 4400 31750 4520
rect 31795 4400 31915 4520
rect 31960 4400 32080 4520
rect 32135 4400 32255 4520
rect 32300 4400 32420 4520
rect 32465 4400 32585 4520
rect 32630 4400 32750 4520
rect 32805 4400 32925 4520
rect 32970 4400 33090 4520
rect 33135 4400 33255 4520
rect 33300 4400 33420 4520
rect 33475 4400 33595 4520
rect 33640 4400 33760 4520
rect 33805 4400 33925 4520
rect 33970 4400 34090 4520
rect 34145 4400 34265 4520
rect 34310 4400 34430 4520
rect 34475 4400 34595 4520
rect 34640 4400 34760 4520
rect 34815 4400 34935 4520
rect 34980 4400 35100 4520
rect 35145 4400 35265 4520
rect 35310 4400 35430 4520
rect 35485 4400 35605 4520
rect 35650 4400 35770 4520
rect 35815 4400 35935 4520
rect 35980 4400 36100 4520
rect 36155 4400 36275 4520
rect 30795 4225 30915 4345
rect 30960 4225 31080 4345
rect 31125 4225 31245 4345
rect 31290 4225 31410 4345
rect 31465 4225 31585 4345
rect 31630 4225 31750 4345
rect 31795 4225 31915 4345
rect 31960 4225 32080 4345
rect 32135 4225 32255 4345
rect 32300 4225 32420 4345
rect 32465 4225 32585 4345
rect 32630 4225 32750 4345
rect 32805 4225 32925 4345
rect 32970 4225 33090 4345
rect 33135 4225 33255 4345
rect 33300 4225 33420 4345
rect 33475 4225 33595 4345
rect 33640 4225 33760 4345
rect 33805 4225 33925 4345
rect 33970 4225 34090 4345
rect 34145 4225 34265 4345
rect 34310 4225 34430 4345
rect 34475 4225 34595 4345
rect 34640 4225 34760 4345
rect 34815 4225 34935 4345
rect 34980 4225 35100 4345
rect 35145 4225 35265 4345
rect 35310 4225 35430 4345
rect 35485 4225 35605 4345
rect 35650 4225 35770 4345
rect 35815 4225 35935 4345
rect 35980 4225 36100 4345
rect 36155 4225 36275 4345
rect 30795 4060 30915 4180
rect 30960 4060 31080 4180
rect 31125 4060 31245 4180
rect 31290 4060 31410 4180
rect 31465 4060 31585 4180
rect 31630 4060 31750 4180
rect 31795 4060 31915 4180
rect 31960 4060 32080 4180
rect 32135 4060 32255 4180
rect 32300 4060 32420 4180
rect 32465 4060 32585 4180
rect 32630 4060 32750 4180
rect 32805 4060 32925 4180
rect 32970 4060 33090 4180
rect 33135 4060 33255 4180
rect 33300 4060 33420 4180
rect 33475 4060 33595 4180
rect 33640 4060 33760 4180
rect 33805 4060 33925 4180
rect 33970 4060 34090 4180
rect 34145 4060 34265 4180
rect 34310 4060 34430 4180
rect 34475 4060 34595 4180
rect 34640 4060 34760 4180
rect 34815 4060 34935 4180
rect 34980 4060 35100 4180
rect 35145 4060 35265 4180
rect 35310 4060 35430 4180
rect 35485 4060 35605 4180
rect 35650 4060 35770 4180
rect 35815 4060 35935 4180
rect 35980 4060 36100 4180
rect 36155 4060 36275 4180
rect 30795 3895 30915 4015
rect 30960 3895 31080 4015
rect 31125 3895 31245 4015
rect 31290 3895 31410 4015
rect 31465 3895 31585 4015
rect 31630 3895 31750 4015
rect 31795 3895 31915 4015
rect 31960 3895 32080 4015
rect 32135 3895 32255 4015
rect 32300 3895 32420 4015
rect 32465 3895 32585 4015
rect 32630 3895 32750 4015
rect 32805 3895 32925 4015
rect 32970 3895 33090 4015
rect 33135 3895 33255 4015
rect 33300 3895 33420 4015
rect 33475 3895 33595 4015
rect 33640 3895 33760 4015
rect 33805 3895 33925 4015
rect 33970 3895 34090 4015
rect 34145 3895 34265 4015
rect 34310 3895 34430 4015
rect 34475 3895 34595 4015
rect 34640 3895 34760 4015
rect 34815 3895 34935 4015
rect 34980 3895 35100 4015
rect 35145 3895 35265 4015
rect 35310 3895 35430 4015
rect 35485 3895 35605 4015
rect 35650 3895 35770 4015
rect 35815 3895 35935 4015
rect 35980 3895 36100 4015
rect 36155 3895 36275 4015
rect 30795 3730 30915 3850
rect 30960 3730 31080 3850
rect 31125 3730 31245 3850
rect 31290 3730 31410 3850
rect 31465 3730 31585 3850
rect 31630 3730 31750 3850
rect 31795 3730 31915 3850
rect 31960 3730 32080 3850
rect 32135 3730 32255 3850
rect 32300 3730 32420 3850
rect 32465 3730 32585 3850
rect 32630 3730 32750 3850
rect 32805 3730 32925 3850
rect 32970 3730 33090 3850
rect 33135 3730 33255 3850
rect 33300 3730 33420 3850
rect 33475 3730 33595 3850
rect 33640 3730 33760 3850
rect 33805 3730 33925 3850
rect 33970 3730 34090 3850
rect 34145 3730 34265 3850
rect 34310 3730 34430 3850
rect 34475 3730 34595 3850
rect 34640 3730 34760 3850
rect 34815 3730 34935 3850
rect 34980 3730 35100 3850
rect 35145 3730 35265 3850
rect 35310 3730 35430 3850
rect 35485 3730 35605 3850
rect 35650 3730 35770 3850
rect 35815 3730 35935 3850
rect 35980 3730 36100 3850
rect 36155 3730 36275 3850
rect 30795 3555 30915 3675
rect 30960 3555 31080 3675
rect 31125 3555 31245 3675
rect 31290 3555 31410 3675
rect 31465 3555 31585 3675
rect 31630 3555 31750 3675
rect 31795 3555 31915 3675
rect 31960 3555 32080 3675
rect 32135 3555 32255 3675
rect 32300 3555 32420 3675
rect 32465 3555 32585 3675
rect 32630 3555 32750 3675
rect 32805 3555 32925 3675
rect 32970 3555 33090 3675
rect 33135 3555 33255 3675
rect 33300 3555 33420 3675
rect 33475 3555 33595 3675
rect 33640 3555 33760 3675
rect 33805 3555 33925 3675
rect 33970 3555 34090 3675
rect 34145 3555 34265 3675
rect 34310 3555 34430 3675
rect 34475 3555 34595 3675
rect 34640 3555 34760 3675
rect 34815 3555 34935 3675
rect 34980 3555 35100 3675
rect 35145 3555 35265 3675
rect 35310 3555 35430 3675
rect 35485 3555 35605 3675
rect 35650 3555 35770 3675
rect 35815 3555 35935 3675
rect 35980 3555 36100 3675
rect 36155 3555 36275 3675
rect 30795 3390 30915 3510
rect 30960 3390 31080 3510
rect 31125 3390 31245 3510
rect 31290 3390 31410 3510
rect 31465 3390 31585 3510
rect 31630 3390 31750 3510
rect 31795 3390 31915 3510
rect 31960 3390 32080 3510
rect 32135 3390 32255 3510
rect 32300 3390 32420 3510
rect 32465 3390 32585 3510
rect 32630 3390 32750 3510
rect 32805 3390 32925 3510
rect 32970 3390 33090 3510
rect 33135 3390 33255 3510
rect 33300 3390 33420 3510
rect 33475 3390 33595 3510
rect 33640 3390 33760 3510
rect 33805 3390 33925 3510
rect 33970 3390 34090 3510
rect 34145 3390 34265 3510
rect 34310 3390 34430 3510
rect 34475 3390 34595 3510
rect 34640 3390 34760 3510
rect 34815 3390 34935 3510
rect 34980 3390 35100 3510
rect 35145 3390 35265 3510
rect 35310 3390 35430 3510
rect 35485 3390 35605 3510
rect 35650 3390 35770 3510
rect 35815 3390 35935 3510
rect 35980 3390 36100 3510
rect 36155 3390 36275 3510
rect 30795 3225 30915 3345
rect 30960 3225 31080 3345
rect 31125 3225 31245 3345
rect 31290 3225 31410 3345
rect 31465 3225 31585 3345
rect 31630 3225 31750 3345
rect 31795 3225 31915 3345
rect 31960 3225 32080 3345
rect 32135 3225 32255 3345
rect 32300 3225 32420 3345
rect 32465 3225 32585 3345
rect 32630 3225 32750 3345
rect 32805 3225 32925 3345
rect 32970 3225 33090 3345
rect 33135 3225 33255 3345
rect 33300 3225 33420 3345
rect 33475 3225 33595 3345
rect 33640 3225 33760 3345
rect 33805 3225 33925 3345
rect 33970 3225 34090 3345
rect 34145 3225 34265 3345
rect 34310 3225 34430 3345
rect 34475 3225 34595 3345
rect 34640 3225 34760 3345
rect 34815 3225 34935 3345
rect 34980 3225 35100 3345
rect 35145 3225 35265 3345
rect 35310 3225 35430 3345
rect 35485 3225 35605 3345
rect 35650 3225 35770 3345
rect 35815 3225 35935 3345
rect 35980 3225 36100 3345
rect 36155 3225 36275 3345
rect 30795 3060 30915 3180
rect 30960 3060 31080 3180
rect 31125 3060 31245 3180
rect 31290 3060 31410 3180
rect 31465 3060 31585 3180
rect 31630 3060 31750 3180
rect 31795 3060 31915 3180
rect 31960 3060 32080 3180
rect 32135 3060 32255 3180
rect 32300 3060 32420 3180
rect 32465 3060 32585 3180
rect 32630 3060 32750 3180
rect 32805 3060 32925 3180
rect 32970 3060 33090 3180
rect 33135 3060 33255 3180
rect 33300 3060 33420 3180
rect 33475 3060 33595 3180
rect 33640 3060 33760 3180
rect 33805 3060 33925 3180
rect 33970 3060 34090 3180
rect 34145 3060 34265 3180
rect 34310 3060 34430 3180
rect 34475 3060 34595 3180
rect 34640 3060 34760 3180
rect 34815 3060 34935 3180
rect 34980 3060 35100 3180
rect 35145 3060 35265 3180
rect 35310 3060 35430 3180
rect 35485 3060 35605 3180
rect 35650 3060 35770 3180
rect 35815 3060 35935 3180
rect 35980 3060 36100 3180
rect 36155 3060 36275 3180
rect 30795 2885 30915 3005
rect 30960 2885 31080 3005
rect 31125 2885 31245 3005
rect 31290 2885 31410 3005
rect 31465 2885 31585 3005
rect 31630 2885 31750 3005
rect 31795 2885 31915 3005
rect 31960 2885 32080 3005
rect 32135 2885 32255 3005
rect 32300 2885 32420 3005
rect 32465 2885 32585 3005
rect 32630 2885 32750 3005
rect 32805 2885 32925 3005
rect 32970 2885 33090 3005
rect 33135 2885 33255 3005
rect 33300 2885 33420 3005
rect 33475 2885 33595 3005
rect 33640 2885 33760 3005
rect 33805 2885 33925 3005
rect 33970 2885 34090 3005
rect 34145 2885 34265 3005
rect 34310 2885 34430 3005
rect 34475 2885 34595 3005
rect 34640 2885 34760 3005
rect 34815 2885 34935 3005
rect 34980 2885 35100 3005
rect 35145 2885 35265 3005
rect 35310 2885 35430 3005
rect 35485 2885 35605 3005
rect 35650 2885 35770 3005
rect 35815 2885 35935 3005
rect 35980 2885 36100 3005
rect 36155 2885 36275 3005
rect 30795 2720 30915 2840
rect 30960 2720 31080 2840
rect 31125 2720 31245 2840
rect 31290 2720 31410 2840
rect 31465 2720 31585 2840
rect 31630 2720 31750 2840
rect 31795 2720 31915 2840
rect 31960 2720 32080 2840
rect 32135 2720 32255 2840
rect 32300 2720 32420 2840
rect 32465 2720 32585 2840
rect 32630 2720 32750 2840
rect 32805 2720 32925 2840
rect 32970 2720 33090 2840
rect 33135 2720 33255 2840
rect 33300 2720 33420 2840
rect 33475 2720 33595 2840
rect 33640 2720 33760 2840
rect 33805 2720 33925 2840
rect 33970 2720 34090 2840
rect 34145 2720 34265 2840
rect 34310 2720 34430 2840
rect 34475 2720 34595 2840
rect 34640 2720 34760 2840
rect 34815 2720 34935 2840
rect 34980 2720 35100 2840
rect 35145 2720 35265 2840
rect 35310 2720 35430 2840
rect 35485 2720 35605 2840
rect 35650 2720 35770 2840
rect 35815 2720 35935 2840
rect 35980 2720 36100 2840
rect 36155 2720 36275 2840
rect 30795 2555 30915 2675
rect 30960 2555 31080 2675
rect 31125 2555 31245 2675
rect 31290 2555 31410 2675
rect 31465 2555 31585 2675
rect 31630 2555 31750 2675
rect 31795 2555 31915 2675
rect 31960 2555 32080 2675
rect 32135 2555 32255 2675
rect 32300 2555 32420 2675
rect 32465 2555 32585 2675
rect 32630 2555 32750 2675
rect 32805 2555 32925 2675
rect 32970 2555 33090 2675
rect 33135 2555 33255 2675
rect 33300 2555 33420 2675
rect 33475 2555 33595 2675
rect 33640 2555 33760 2675
rect 33805 2555 33925 2675
rect 33970 2555 34090 2675
rect 34145 2555 34265 2675
rect 34310 2555 34430 2675
rect 34475 2555 34595 2675
rect 34640 2555 34760 2675
rect 34815 2555 34935 2675
rect 34980 2555 35100 2675
rect 35145 2555 35265 2675
rect 35310 2555 35430 2675
rect 35485 2555 35605 2675
rect 35650 2555 35770 2675
rect 35815 2555 35935 2675
rect 35980 2555 36100 2675
rect 36155 2555 36275 2675
rect 30795 2390 30915 2510
rect 30960 2390 31080 2510
rect 31125 2390 31245 2510
rect 31290 2390 31410 2510
rect 31465 2390 31585 2510
rect 31630 2390 31750 2510
rect 31795 2390 31915 2510
rect 31960 2390 32080 2510
rect 32135 2390 32255 2510
rect 32300 2390 32420 2510
rect 32465 2390 32585 2510
rect 32630 2390 32750 2510
rect 32805 2390 32925 2510
rect 32970 2390 33090 2510
rect 33135 2390 33255 2510
rect 33300 2390 33420 2510
rect 33475 2390 33595 2510
rect 33640 2390 33760 2510
rect 33805 2390 33925 2510
rect 33970 2390 34090 2510
rect 34145 2390 34265 2510
rect 34310 2390 34430 2510
rect 34475 2390 34595 2510
rect 34640 2390 34760 2510
rect 34815 2390 34935 2510
rect 34980 2390 35100 2510
rect 35145 2390 35265 2510
rect 35310 2390 35430 2510
rect 35485 2390 35605 2510
rect 35650 2390 35770 2510
rect 35815 2390 35935 2510
rect 35980 2390 36100 2510
rect 36155 2390 36275 2510
rect 30795 2215 30915 2335
rect 30960 2215 31080 2335
rect 31125 2215 31245 2335
rect 31290 2215 31410 2335
rect 31465 2215 31585 2335
rect 31630 2215 31750 2335
rect 31795 2215 31915 2335
rect 31960 2215 32080 2335
rect 32135 2215 32255 2335
rect 32300 2215 32420 2335
rect 32465 2215 32585 2335
rect 32630 2215 32750 2335
rect 32805 2215 32925 2335
rect 32970 2215 33090 2335
rect 33135 2215 33255 2335
rect 33300 2215 33420 2335
rect 33475 2215 33595 2335
rect 33640 2215 33760 2335
rect 33805 2215 33925 2335
rect 33970 2215 34090 2335
rect 34145 2215 34265 2335
rect 34310 2215 34430 2335
rect 34475 2215 34595 2335
rect 34640 2215 34760 2335
rect 34815 2215 34935 2335
rect 34980 2215 35100 2335
rect 35145 2215 35265 2335
rect 35310 2215 35430 2335
rect 35485 2215 35605 2335
rect 35650 2215 35770 2335
rect 35815 2215 35935 2335
rect 35980 2215 36100 2335
rect 36155 2215 36275 2335
rect 30795 2050 30915 2170
rect 30960 2050 31080 2170
rect 31125 2050 31245 2170
rect 31290 2050 31410 2170
rect 31465 2050 31585 2170
rect 31630 2050 31750 2170
rect 31795 2050 31915 2170
rect 31960 2050 32080 2170
rect 32135 2050 32255 2170
rect 32300 2050 32420 2170
rect 32465 2050 32585 2170
rect 32630 2050 32750 2170
rect 32805 2050 32925 2170
rect 32970 2050 33090 2170
rect 33135 2050 33255 2170
rect 33300 2050 33420 2170
rect 33475 2050 33595 2170
rect 33640 2050 33760 2170
rect 33805 2050 33925 2170
rect 33970 2050 34090 2170
rect 34145 2050 34265 2170
rect 34310 2050 34430 2170
rect 34475 2050 34595 2170
rect 34640 2050 34760 2170
rect 34815 2050 34935 2170
rect 34980 2050 35100 2170
rect 35145 2050 35265 2170
rect 35310 2050 35430 2170
rect 35485 2050 35605 2170
rect 35650 2050 35770 2170
rect 35815 2050 35935 2170
rect 35980 2050 36100 2170
rect 36155 2050 36275 2170
rect 30795 1885 30915 2005
rect 30960 1885 31080 2005
rect 31125 1885 31245 2005
rect 31290 1885 31410 2005
rect 31465 1885 31585 2005
rect 31630 1885 31750 2005
rect 31795 1885 31915 2005
rect 31960 1885 32080 2005
rect 32135 1885 32255 2005
rect 32300 1885 32420 2005
rect 32465 1885 32585 2005
rect 32630 1885 32750 2005
rect 32805 1885 32925 2005
rect 32970 1885 33090 2005
rect 33135 1885 33255 2005
rect 33300 1885 33420 2005
rect 33475 1885 33595 2005
rect 33640 1885 33760 2005
rect 33805 1885 33925 2005
rect 33970 1885 34090 2005
rect 34145 1885 34265 2005
rect 34310 1885 34430 2005
rect 34475 1885 34595 2005
rect 34640 1885 34760 2005
rect 34815 1885 34935 2005
rect 34980 1885 35100 2005
rect 35145 1885 35265 2005
rect 35310 1885 35430 2005
rect 35485 1885 35605 2005
rect 35650 1885 35770 2005
rect 35815 1885 35935 2005
rect 35980 1885 36100 2005
rect 36155 1885 36275 2005
rect 30795 1720 30915 1840
rect 30960 1720 31080 1840
rect 31125 1720 31245 1840
rect 31290 1720 31410 1840
rect 31465 1720 31585 1840
rect 31630 1720 31750 1840
rect 31795 1720 31915 1840
rect 31960 1720 32080 1840
rect 32135 1720 32255 1840
rect 32300 1720 32420 1840
rect 32465 1720 32585 1840
rect 32630 1720 32750 1840
rect 32805 1720 32925 1840
rect 32970 1720 33090 1840
rect 33135 1720 33255 1840
rect 33300 1720 33420 1840
rect 33475 1720 33595 1840
rect 33640 1720 33760 1840
rect 33805 1720 33925 1840
rect 33970 1720 34090 1840
rect 34145 1720 34265 1840
rect 34310 1720 34430 1840
rect 34475 1720 34595 1840
rect 34640 1720 34760 1840
rect 34815 1720 34935 1840
rect 34980 1720 35100 1840
rect 35145 1720 35265 1840
rect 35310 1720 35430 1840
rect 35485 1720 35605 1840
rect 35650 1720 35770 1840
rect 35815 1720 35935 1840
rect 35980 1720 36100 1840
rect 36155 1720 36275 1840
rect 36485 7080 36605 7200
rect 36650 7080 36770 7200
rect 36815 7080 36935 7200
rect 36980 7080 37100 7200
rect 37155 7080 37275 7200
rect 37320 7080 37440 7200
rect 37485 7080 37605 7200
rect 37650 7080 37770 7200
rect 37825 7080 37945 7200
rect 37990 7080 38110 7200
rect 38155 7080 38275 7200
rect 38320 7080 38440 7200
rect 38495 7080 38615 7200
rect 38660 7080 38780 7200
rect 38825 7080 38945 7200
rect 38990 7080 39110 7200
rect 39165 7080 39285 7200
rect 39330 7080 39450 7200
rect 39495 7080 39615 7200
rect 39660 7080 39780 7200
rect 39835 7080 39955 7200
rect 40000 7080 40120 7200
rect 40165 7080 40285 7200
rect 40330 7080 40450 7200
rect 40505 7080 40625 7200
rect 40670 7080 40790 7200
rect 40835 7080 40955 7200
rect 41000 7080 41120 7200
rect 41175 7080 41295 7200
rect 41340 7080 41460 7200
rect 41505 7080 41625 7200
rect 41670 7080 41790 7200
rect 41845 7080 41965 7200
rect 36485 6905 36605 7025
rect 36650 6905 36770 7025
rect 36815 6905 36935 7025
rect 36980 6905 37100 7025
rect 37155 6905 37275 7025
rect 37320 6905 37440 7025
rect 37485 6905 37605 7025
rect 37650 6905 37770 7025
rect 37825 6905 37945 7025
rect 37990 6905 38110 7025
rect 38155 6905 38275 7025
rect 38320 6905 38440 7025
rect 38495 6905 38615 7025
rect 38660 6905 38780 7025
rect 38825 6905 38945 7025
rect 38990 6905 39110 7025
rect 39165 6905 39285 7025
rect 39330 6905 39450 7025
rect 39495 6905 39615 7025
rect 39660 6905 39780 7025
rect 39835 6905 39955 7025
rect 40000 6905 40120 7025
rect 40165 6905 40285 7025
rect 40330 6905 40450 7025
rect 40505 6905 40625 7025
rect 40670 6905 40790 7025
rect 40835 6905 40955 7025
rect 41000 6905 41120 7025
rect 41175 6905 41295 7025
rect 41340 6905 41460 7025
rect 41505 6905 41625 7025
rect 41670 6905 41790 7025
rect 41845 6905 41965 7025
rect 36485 6740 36605 6860
rect 36650 6740 36770 6860
rect 36815 6740 36935 6860
rect 36980 6740 37100 6860
rect 37155 6740 37275 6860
rect 37320 6740 37440 6860
rect 37485 6740 37605 6860
rect 37650 6740 37770 6860
rect 37825 6740 37945 6860
rect 37990 6740 38110 6860
rect 38155 6740 38275 6860
rect 38320 6740 38440 6860
rect 38495 6740 38615 6860
rect 38660 6740 38780 6860
rect 38825 6740 38945 6860
rect 38990 6740 39110 6860
rect 39165 6740 39285 6860
rect 39330 6740 39450 6860
rect 39495 6740 39615 6860
rect 39660 6740 39780 6860
rect 39835 6740 39955 6860
rect 40000 6740 40120 6860
rect 40165 6740 40285 6860
rect 40330 6740 40450 6860
rect 40505 6740 40625 6860
rect 40670 6740 40790 6860
rect 40835 6740 40955 6860
rect 41000 6740 41120 6860
rect 41175 6740 41295 6860
rect 41340 6740 41460 6860
rect 41505 6740 41625 6860
rect 41670 6740 41790 6860
rect 41845 6740 41965 6860
rect 36485 6575 36605 6695
rect 36650 6575 36770 6695
rect 36815 6575 36935 6695
rect 36980 6575 37100 6695
rect 37155 6575 37275 6695
rect 37320 6575 37440 6695
rect 37485 6575 37605 6695
rect 37650 6575 37770 6695
rect 37825 6575 37945 6695
rect 37990 6575 38110 6695
rect 38155 6575 38275 6695
rect 38320 6575 38440 6695
rect 38495 6575 38615 6695
rect 38660 6575 38780 6695
rect 38825 6575 38945 6695
rect 38990 6575 39110 6695
rect 39165 6575 39285 6695
rect 39330 6575 39450 6695
rect 39495 6575 39615 6695
rect 39660 6575 39780 6695
rect 39835 6575 39955 6695
rect 40000 6575 40120 6695
rect 40165 6575 40285 6695
rect 40330 6575 40450 6695
rect 40505 6575 40625 6695
rect 40670 6575 40790 6695
rect 40835 6575 40955 6695
rect 41000 6575 41120 6695
rect 41175 6575 41295 6695
rect 41340 6575 41460 6695
rect 41505 6575 41625 6695
rect 41670 6575 41790 6695
rect 41845 6575 41965 6695
rect 36485 6410 36605 6530
rect 36650 6410 36770 6530
rect 36815 6410 36935 6530
rect 36980 6410 37100 6530
rect 37155 6410 37275 6530
rect 37320 6410 37440 6530
rect 37485 6410 37605 6530
rect 37650 6410 37770 6530
rect 37825 6410 37945 6530
rect 37990 6410 38110 6530
rect 38155 6410 38275 6530
rect 38320 6410 38440 6530
rect 38495 6410 38615 6530
rect 38660 6410 38780 6530
rect 38825 6410 38945 6530
rect 38990 6410 39110 6530
rect 39165 6410 39285 6530
rect 39330 6410 39450 6530
rect 39495 6410 39615 6530
rect 39660 6410 39780 6530
rect 39835 6410 39955 6530
rect 40000 6410 40120 6530
rect 40165 6410 40285 6530
rect 40330 6410 40450 6530
rect 40505 6410 40625 6530
rect 40670 6410 40790 6530
rect 40835 6410 40955 6530
rect 41000 6410 41120 6530
rect 41175 6410 41295 6530
rect 41340 6410 41460 6530
rect 41505 6410 41625 6530
rect 41670 6410 41790 6530
rect 41845 6410 41965 6530
rect 36485 6235 36605 6355
rect 36650 6235 36770 6355
rect 36815 6235 36935 6355
rect 36980 6235 37100 6355
rect 37155 6235 37275 6355
rect 37320 6235 37440 6355
rect 37485 6235 37605 6355
rect 37650 6235 37770 6355
rect 37825 6235 37945 6355
rect 37990 6235 38110 6355
rect 38155 6235 38275 6355
rect 38320 6235 38440 6355
rect 38495 6235 38615 6355
rect 38660 6235 38780 6355
rect 38825 6235 38945 6355
rect 38990 6235 39110 6355
rect 39165 6235 39285 6355
rect 39330 6235 39450 6355
rect 39495 6235 39615 6355
rect 39660 6235 39780 6355
rect 39835 6235 39955 6355
rect 40000 6235 40120 6355
rect 40165 6235 40285 6355
rect 40330 6235 40450 6355
rect 40505 6235 40625 6355
rect 40670 6235 40790 6355
rect 40835 6235 40955 6355
rect 41000 6235 41120 6355
rect 41175 6235 41295 6355
rect 41340 6235 41460 6355
rect 41505 6235 41625 6355
rect 41670 6235 41790 6355
rect 41845 6235 41965 6355
rect 36485 6070 36605 6190
rect 36650 6070 36770 6190
rect 36815 6070 36935 6190
rect 36980 6070 37100 6190
rect 37155 6070 37275 6190
rect 37320 6070 37440 6190
rect 37485 6070 37605 6190
rect 37650 6070 37770 6190
rect 37825 6070 37945 6190
rect 37990 6070 38110 6190
rect 38155 6070 38275 6190
rect 38320 6070 38440 6190
rect 38495 6070 38615 6190
rect 38660 6070 38780 6190
rect 38825 6070 38945 6190
rect 38990 6070 39110 6190
rect 39165 6070 39285 6190
rect 39330 6070 39450 6190
rect 39495 6070 39615 6190
rect 39660 6070 39780 6190
rect 39835 6070 39955 6190
rect 40000 6070 40120 6190
rect 40165 6070 40285 6190
rect 40330 6070 40450 6190
rect 40505 6070 40625 6190
rect 40670 6070 40790 6190
rect 40835 6070 40955 6190
rect 41000 6070 41120 6190
rect 41175 6070 41295 6190
rect 41340 6070 41460 6190
rect 41505 6070 41625 6190
rect 41670 6070 41790 6190
rect 41845 6070 41965 6190
rect 36485 5905 36605 6025
rect 36650 5905 36770 6025
rect 36815 5905 36935 6025
rect 36980 5905 37100 6025
rect 37155 5905 37275 6025
rect 37320 5905 37440 6025
rect 37485 5905 37605 6025
rect 37650 5905 37770 6025
rect 37825 5905 37945 6025
rect 37990 5905 38110 6025
rect 38155 5905 38275 6025
rect 38320 5905 38440 6025
rect 38495 5905 38615 6025
rect 38660 5905 38780 6025
rect 38825 5905 38945 6025
rect 38990 5905 39110 6025
rect 39165 5905 39285 6025
rect 39330 5905 39450 6025
rect 39495 5905 39615 6025
rect 39660 5905 39780 6025
rect 39835 5905 39955 6025
rect 40000 5905 40120 6025
rect 40165 5905 40285 6025
rect 40330 5905 40450 6025
rect 40505 5905 40625 6025
rect 40670 5905 40790 6025
rect 40835 5905 40955 6025
rect 41000 5905 41120 6025
rect 41175 5905 41295 6025
rect 41340 5905 41460 6025
rect 41505 5905 41625 6025
rect 41670 5905 41790 6025
rect 41845 5905 41965 6025
rect 36485 5740 36605 5860
rect 36650 5740 36770 5860
rect 36815 5740 36935 5860
rect 36980 5740 37100 5860
rect 37155 5740 37275 5860
rect 37320 5740 37440 5860
rect 37485 5740 37605 5860
rect 37650 5740 37770 5860
rect 37825 5740 37945 5860
rect 37990 5740 38110 5860
rect 38155 5740 38275 5860
rect 38320 5740 38440 5860
rect 38495 5740 38615 5860
rect 38660 5740 38780 5860
rect 38825 5740 38945 5860
rect 38990 5740 39110 5860
rect 39165 5740 39285 5860
rect 39330 5740 39450 5860
rect 39495 5740 39615 5860
rect 39660 5740 39780 5860
rect 39835 5740 39955 5860
rect 40000 5740 40120 5860
rect 40165 5740 40285 5860
rect 40330 5740 40450 5860
rect 40505 5740 40625 5860
rect 40670 5740 40790 5860
rect 40835 5740 40955 5860
rect 41000 5740 41120 5860
rect 41175 5740 41295 5860
rect 41340 5740 41460 5860
rect 41505 5740 41625 5860
rect 41670 5740 41790 5860
rect 41845 5740 41965 5860
rect 36485 5565 36605 5685
rect 36650 5565 36770 5685
rect 36815 5565 36935 5685
rect 36980 5565 37100 5685
rect 37155 5565 37275 5685
rect 37320 5565 37440 5685
rect 37485 5565 37605 5685
rect 37650 5565 37770 5685
rect 37825 5565 37945 5685
rect 37990 5565 38110 5685
rect 38155 5565 38275 5685
rect 38320 5565 38440 5685
rect 38495 5565 38615 5685
rect 38660 5565 38780 5685
rect 38825 5565 38945 5685
rect 38990 5565 39110 5685
rect 39165 5565 39285 5685
rect 39330 5565 39450 5685
rect 39495 5565 39615 5685
rect 39660 5565 39780 5685
rect 39835 5565 39955 5685
rect 40000 5565 40120 5685
rect 40165 5565 40285 5685
rect 40330 5565 40450 5685
rect 40505 5565 40625 5685
rect 40670 5565 40790 5685
rect 40835 5565 40955 5685
rect 41000 5565 41120 5685
rect 41175 5565 41295 5685
rect 41340 5565 41460 5685
rect 41505 5565 41625 5685
rect 41670 5565 41790 5685
rect 41845 5565 41965 5685
rect 36485 5400 36605 5520
rect 36650 5400 36770 5520
rect 36815 5400 36935 5520
rect 36980 5400 37100 5520
rect 37155 5400 37275 5520
rect 37320 5400 37440 5520
rect 37485 5400 37605 5520
rect 37650 5400 37770 5520
rect 37825 5400 37945 5520
rect 37990 5400 38110 5520
rect 38155 5400 38275 5520
rect 38320 5400 38440 5520
rect 38495 5400 38615 5520
rect 38660 5400 38780 5520
rect 38825 5400 38945 5520
rect 38990 5400 39110 5520
rect 39165 5400 39285 5520
rect 39330 5400 39450 5520
rect 39495 5400 39615 5520
rect 39660 5400 39780 5520
rect 39835 5400 39955 5520
rect 40000 5400 40120 5520
rect 40165 5400 40285 5520
rect 40330 5400 40450 5520
rect 40505 5400 40625 5520
rect 40670 5400 40790 5520
rect 40835 5400 40955 5520
rect 41000 5400 41120 5520
rect 41175 5400 41295 5520
rect 41340 5400 41460 5520
rect 41505 5400 41625 5520
rect 41670 5400 41790 5520
rect 41845 5400 41965 5520
rect 36485 5235 36605 5355
rect 36650 5235 36770 5355
rect 36815 5235 36935 5355
rect 36980 5235 37100 5355
rect 37155 5235 37275 5355
rect 37320 5235 37440 5355
rect 37485 5235 37605 5355
rect 37650 5235 37770 5355
rect 37825 5235 37945 5355
rect 37990 5235 38110 5355
rect 38155 5235 38275 5355
rect 38320 5235 38440 5355
rect 38495 5235 38615 5355
rect 38660 5235 38780 5355
rect 38825 5235 38945 5355
rect 38990 5235 39110 5355
rect 39165 5235 39285 5355
rect 39330 5235 39450 5355
rect 39495 5235 39615 5355
rect 39660 5235 39780 5355
rect 39835 5235 39955 5355
rect 40000 5235 40120 5355
rect 40165 5235 40285 5355
rect 40330 5235 40450 5355
rect 40505 5235 40625 5355
rect 40670 5235 40790 5355
rect 40835 5235 40955 5355
rect 41000 5235 41120 5355
rect 41175 5235 41295 5355
rect 41340 5235 41460 5355
rect 41505 5235 41625 5355
rect 41670 5235 41790 5355
rect 41845 5235 41965 5355
rect 36485 5070 36605 5190
rect 36650 5070 36770 5190
rect 36815 5070 36935 5190
rect 36980 5070 37100 5190
rect 37155 5070 37275 5190
rect 37320 5070 37440 5190
rect 37485 5070 37605 5190
rect 37650 5070 37770 5190
rect 37825 5070 37945 5190
rect 37990 5070 38110 5190
rect 38155 5070 38275 5190
rect 38320 5070 38440 5190
rect 38495 5070 38615 5190
rect 38660 5070 38780 5190
rect 38825 5070 38945 5190
rect 38990 5070 39110 5190
rect 39165 5070 39285 5190
rect 39330 5070 39450 5190
rect 39495 5070 39615 5190
rect 39660 5070 39780 5190
rect 39835 5070 39955 5190
rect 40000 5070 40120 5190
rect 40165 5070 40285 5190
rect 40330 5070 40450 5190
rect 40505 5070 40625 5190
rect 40670 5070 40790 5190
rect 40835 5070 40955 5190
rect 41000 5070 41120 5190
rect 41175 5070 41295 5190
rect 41340 5070 41460 5190
rect 41505 5070 41625 5190
rect 41670 5070 41790 5190
rect 41845 5070 41965 5190
rect 36485 4895 36605 5015
rect 36650 4895 36770 5015
rect 36815 4895 36935 5015
rect 36980 4895 37100 5015
rect 37155 4895 37275 5015
rect 37320 4895 37440 5015
rect 37485 4895 37605 5015
rect 37650 4895 37770 5015
rect 37825 4895 37945 5015
rect 37990 4895 38110 5015
rect 38155 4895 38275 5015
rect 38320 4895 38440 5015
rect 38495 4895 38615 5015
rect 38660 4895 38780 5015
rect 38825 4895 38945 5015
rect 38990 4895 39110 5015
rect 39165 4895 39285 5015
rect 39330 4895 39450 5015
rect 39495 4895 39615 5015
rect 39660 4895 39780 5015
rect 39835 4895 39955 5015
rect 40000 4895 40120 5015
rect 40165 4895 40285 5015
rect 40330 4895 40450 5015
rect 40505 4895 40625 5015
rect 40670 4895 40790 5015
rect 40835 4895 40955 5015
rect 41000 4895 41120 5015
rect 41175 4895 41295 5015
rect 41340 4895 41460 5015
rect 41505 4895 41625 5015
rect 41670 4895 41790 5015
rect 41845 4895 41965 5015
rect 36485 4730 36605 4850
rect 36650 4730 36770 4850
rect 36815 4730 36935 4850
rect 36980 4730 37100 4850
rect 37155 4730 37275 4850
rect 37320 4730 37440 4850
rect 37485 4730 37605 4850
rect 37650 4730 37770 4850
rect 37825 4730 37945 4850
rect 37990 4730 38110 4850
rect 38155 4730 38275 4850
rect 38320 4730 38440 4850
rect 38495 4730 38615 4850
rect 38660 4730 38780 4850
rect 38825 4730 38945 4850
rect 38990 4730 39110 4850
rect 39165 4730 39285 4850
rect 39330 4730 39450 4850
rect 39495 4730 39615 4850
rect 39660 4730 39780 4850
rect 39835 4730 39955 4850
rect 40000 4730 40120 4850
rect 40165 4730 40285 4850
rect 40330 4730 40450 4850
rect 40505 4730 40625 4850
rect 40670 4730 40790 4850
rect 40835 4730 40955 4850
rect 41000 4730 41120 4850
rect 41175 4730 41295 4850
rect 41340 4730 41460 4850
rect 41505 4730 41625 4850
rect 41670 4730 41790 4850
rect 41845 4730 41965 4850
rect 36485 4565 36605 4685
rect 36650 4565 36770 4685
rect 36815 4565 36935 4685
rect 36980 4565 37100 4685
rect 37155 4565 37275 4685
rect 37320 4565 37440 4685
rect 37485 4565 37605 4685
rect 37650 4565 37770 4685
rect 37825 4565 37945 4685
rect 37990 4565 38110 4685
rect 38155 4565 38275 4685
rect 38320 4565 38440 4685
rect 38495 4565 38615 4685
rect 38660 4565 38780 4685
rect 38825 4565 38945 4685
rect 38990 4565 39110 4685
rect 39165 4565 39285 4685
rect 39330 4565 39450 4685
rect 39495 4565 39615 4685
rect 39660 4565 39780 4685
rect 39835 4565 39955 4685
rect 40000 4565 40120 4685
rect 40165 4565 40285 4685
rect 40330 4565 40450 4685
rect 40505 4565 40625 4685
rect 40670 4565 40790 4685
rect 40835 4565 40955 4685
rect 41000 4565 41120 4685
rect 41175 4565 41295 4685
rect 41340 4565 41460 4685
rect 41505 4565 41625 4685
rect 41670 4565 41790 4685
rect 41845 4565 41965 4685
rect 36485 4400 36605 4520
rect 36650 4400 36770 4520
rect 36815 4400 36935 4520
rect 36980 4400 37100 4520
rect 37155 4400 37275 4520
rect 37320 4400 37440 4520
rect 37485 4400 37605 4520
rect 37650 4400 37770 4520
rect 37825 4400 37945 4520
rect 37990 4400 38110 4520
rect 38155 4400 38275 4520
rect 38320 4400 38440 4520
rect 38495 4400 38615 4520
rect 38660 4400 38780 4520
rect 38825 4400 38945 4520
rect 38990 4400 39110 4520
rect 39165 4400 39285 4520
rect 39330 4400 39450 4520
rect 39495 4400 39615 4520
rect 39660 4400 39780 4520
rect 39835 4400 39955 4520
rect 40000 4400 40120 4520
rect 40165 4400 40285 4520
rect 40330 4400 40450 4520
rect 40505 4400 40625 4520
rect 40670 4400 40790 4520
rect 40835 4400 40955 4520
rect 41000 4400 41120 4520
rect 41175 4400 41295 4520
rect 41340 4400 41460 4520
rect 41505 4400 41625 4520
rect 41670 4400 41790 4520
rect 41845 4400 41965 4520
rect 36485 4225 36605 4345
rect 36650 4225 36770 4345
rect 36815 4225 36935 4345
rect 36980 4225 37100 4345
rect 37155 4225 37275 4345
rect 37320 4225 37440 4345
rect 37485 4225 37605 4345
rect 37650 4225 37770 4345
rect 37825 4225 37945 4345
rect 37990 4225 38110 4345
rect 38155 4225 38275 4345
rect 38320 4225 38440 4345
rect 38495 4225 38615 4345
rect 38660 4225 38780 4345
rect 38825 4225 38945 4345
rect 38990 4225 39110 4345
rect 39165 4225 39285 4345
rect 39330 4225 39450 4345
rect 39495 4225 39615 4345
rect 39660 4225 39780 4345
rect 39835 4225 39955 4345
rect 40000 4225 40120 4345
rect 40165 4225 40285 4345
rect 40330 4225 40450 4345
rect 40505 4225 40625 4345
rect 40670 4225 40790 4345
rect 40835 4225 40955 4345
rect 41000 4225 41120 4345
rect 41175 4225 41295 4345
rect 41340 4225 41460 4345
rect 41505 4225 41625 4345
rect 41670 4225 41790 4345
rect 41845 4225 41965 4345
rect 36485 4060 36605 4180
rect 36650 4060 36770 4180
rect 36815 4060 36935 4180
rect 36980 4060 37100 4180
rect 37155 4060 37275 4180
rect 37320 4060 37440 4180
rect 37485 4060 37605 4180
rect 37650 4060 37770 4180
rect 37825 4060 37945 4180
rect 37990 4060 38110 4180
rect 38155 4060 38275 4180
rect 38320 4060 38440 4180
rect 38495 4060 38615 4180
rect 38660 4060 38780 4180
rect 38825 4060 38945 4180
rect 38990 4060 39110 4180
rect 39165 4060 39285 4180
rect 39330 4060 39450 4180
rect 39495 4060 39615 4180
rect 39660 4060 39780 4180
rect 39835 4060 39955 4180
rect 40000 4060 40120 4180
rect 40165 4060 40285 4180
rect 40330 4060 40450 4180
rect 40505 4060 40625 4180
rect 40670 4060 40790 4180
rect 40835 4060 40955 4180
rect 41000 4060 41120 4180
rect 41175 4060 41295 4180
rect 41340 4060 41460 4180
rect 41505 4060 41625 4180
rect 41670 4060 41790 4180
rect 41845 4060 41965 4180
rect 36485 3895 36605 4015
rect 36650 3895 36770 4015
rect 36815 3895 36935 4015
rect 36980 3895 37100 4015
rect 37155 3895 37275 4015
rect 37320 3895 37440 4015
rect 37485 3895 37605 4015
rect 37650 3895 37770 4015
rect 37825 3895 37945 4015
rect 37990 3895 38110 4015
rect 38155 3895 38275 4015
rect 38320 3895 38440 4015
rect 38495 3895 38615 4015
rect 38660 3895 38780 4015
rect 38825 3895 38945 4015
rect 38990 3895 39110 4015
rect 39165 3895 39285 4015
rect 39330 3895 39450 4015
rect 39495 3895 39615 4015
rect 39660 3895 39780 4015
rect 39835 3895 39955 4015
rect 40000 3895 40120 4015
rect 40165 3895 40285 4015
rect 40330 3895 40450 4015
rect 40505 3895 40625 4015
rect 40670 3895 40790 4015
rect 40835 3895 40955 4015
rect 41000 3895 41120 4015
rect 41175 3895 41295 4015
rect 41340 3895 41460 4015
rect 41505 3895 41625 4015
rect 41670 3895 41790 4015
rect 41845 3895 41965 4015
rect 36485 3730 36605 3850
rect 36650 3730 36770 3850
rect 36815 3730 36935 3850
rect 36980 3730 37100 3850
rect 37155 3730 37275 3850
rect 37320 3730 37440 3850
rect 37485 3730 37605 3850
rect 37650 3730 37770 3850
rect 37825 3730 37945 3850
rect 37990 3730 38110 3850
rect 38155 3730 38275 3850
rect 38320 3730 38440 3850
rect 38495 3730 38615 3850
rect 38660 3730 38780 3850
rect 38825 3730 38945 3850
rect 38990 3730 39110 3850
rect 39165 3730 39285 3850
rect 39330 3730 39450 3850
rect 39495 3730 39615 3850
rect 39660 3730 39780 3850
rect 39835 3730 39955 3850
rect 40000 3730 40120 3850
rect 40165 3730 40285 3850
rect 40330 3730 40450 3850
rect 40505 3730 40625 3850
rect 40670 3730 40790 3850
rect 40835 3730 40955 3850
rect 41000 3730 41120 3850
rect 41175 3730 41295 3850
rect 41340 3730 41460 3850
rect 41505 3730 41625 3850
rect 41670 3730 41790 3850
rect 41845 3730 41965 3850
rect 36485 3555 36605 3675
rect 36650 3555 36770 3675
rect 36815 3555 36935 3675
rect 36980 3555 37100 3675
rect 37155 3555 37275 3675
rect 37320 3555 37440 3675
rect 37485 3555 37605 3675
rect 37650 3555 37770 3675
rect 37825 3555 37945 3675
rect 37990 3555 38110 3675
rect 38155 3555 38275 3675
rect 38320 3555 38440 3675
rect 38495 3555 38615 3675
rect 38660 3555 38780 3675
rect 38825 3555 38945 3675
rect 38990 3555 39110 3675
rect 39165 3555 39285 3675
rect 39330 3555 39450 3675
rect 39495 3555 39615 3675
rect 39660 3555 39780 3675
rect 39835 3555 39955 3675
rect 40000 3555 40120 3675
rect 40165 3555 40285 3675
rect 40330 3555 40450 3675
rect 40505 3555 40625 3675
rect 40670 3555 40790 3675
rect 40835 3555 40955 3675
rect 41000 3555 41120 3675
rect 41175 3555 41295 3675
rect 41340 3555 41460 3675
rect 41505 3555 41625 3675
rect 41670 3555 41790 3675
rect 41845 3555 41965 3675
rect 36485 3390 36605 3510
rect 36650 3390 36770 3510
rect 36815 3390 36935 3510
rect 36980 3390 37100 3510
rect 37155 3390 37275 3510
rect 37320 3390 37440 3510
rect 37485 3390 37605 3510
rect 37650 3390 37770 3510
rect 37825 3390 37945 3510
rect 37990 3390 38110 3510
rect 38155 3390 38275 3510
rect 38320 3390 38440 3510
rect 38495 3390 38615 3510
rect 38660 3390 38780 3510
rect 38825 3390 38945 3510
rect 38990 3390 39110 3510
rect 39165 3390 39285 3510
rect 39330 3390 39450 3510
rect 39495 3390 39615 3510
rect 39660 3390 39780 3510
rect 39835 3390 39955 3510
rect 40000 3390 40120 3510
rect 40165 3390 40285 3510
rect 40330 3390 40450 3510
rect 40505 3390 40625 3510
rect 40670 3390 40790 3510
rect 40835 3390 40955 3510
rect 41000 3390 41120 3510
rect 41175 3390 41295 3510
rect 41340 3390 41460 3510
rect 41505 3390 41625 3510
rect 41670 3390 41790 3510
rect 41845 3390 41965 3510
rect 36485 3225 36605 3345
rect 36650 3225 36770 3345
rect 36815 3225 36935 3345
rect 36980 3225 37100 3345
rect 37155 3225 37275 3345
rect 37320 3225 37440 3345
rect 37485 3225 37605 3345
rect 37650 3225 37770 3345
rect 37825 3225 37945 3345
rect 37990 3225 38110 3345
rect 38155 3225 38275 3345
rect 38320 3225 38440 3345
rect 38495 3225 38615 3345
rect 38660 3225 38780 3345
rect 38825 3225 38945 3345
rect 38990 3225 39110 3345
rect 39165 3225 39285 3345
rect 39330 3225 39450 3345
rect 39495 3225 39615 3345
rect 39660 3225 39780 3345
rect 39835 3225 39955 3345
rect 40000 3225 40120 3345
rect 40165 3225 40285 3345
rect 40330 3225 40450 3345
rect 40505 3225 40625 3345
rect 40670 3225 40790 3345
rect 40835 3225 40955 3345
rect 41000 3225 41120 3345
rect 41175 3225 41295 3345
rect 41340 3225 41460 3345
rect 41505 3225 41625 3345
rect 41670 3225 41790 3345
rect 41845 3225 41965 3345
rect 36485 3060 36605 3180
rect 36650 3060 36770 3180
rect 36815 3060 36935 3180
rect 36980 3060 37100 3180
rect 37155 3060 37275 3180
rect 37320 3060 37440 3180
rect 37485 3060 37605 3180
rect 37650 3060 37770 3180
rect 37825 3060 37945 3180
rect 37990 3060 38110 3180
rect 38155 3060 38275 3180
rect 38320 3060 38440 3180
rect 38495 3060 38615 3180
rect 38660 3060 38780 3180
rect 38825 3060 38945 3180
rect 38990 3060 39110 3180
rect 39165 3060 39285 3180
rect 39330 3060 39450 3180
rect 39495 3060 39615 3180
rect 39660 3060 39780 3180
rect 39835 3060 39955 3180
rect 40000 3060 40120 3180
rect 40165 3060 40285 3180
rect 40330 3060 40450 3180
rect 40505 3060 40625 3180
rect 40670 3060 40790 3180
rect 40835 3060 40955 3180
rect 41000 3060 41120 3180
rect 41175 3060 41295 3180
rect 41340 3060 41460 3180
rect 41505 3060 41625 3180
rect 41670 3060 41790 3180
rect 41845 3060 41965 3180
rect 36485 2885 36605 3005
rect 36650 2885 36770 3005
rect 36815 2885 36935 3005
rect 36980 2885 37100 3005
rect 37155 2885 37275 3005
rect 37320 2885 37440 3005
rect 37485 2885 37605 3005
rect 37650 2885 37770 3005
rect 37825 2885 37945 3005
rect 37990 2885 38110 3005
rect 38155 2885 38275 3005
rect 38320 2885 38440 3005
rect 38495 2885 38615 3005
rect 38660 2885 38780 3005
rect 38825 2885 38945 3005
rect 38990 2885 39110 3005
rect 39165 2885 39285 3005
rect 39330 2885 39450 3005
rect 39495 2885 39615 3005
rect 39660 2885 39780 3005
rect 39835 2885 39955 3005
rect 40000 2885 40120 3005
rect 40165 2885 40285 3005
rect 40330 2885 40450 3005
rect 40505 2885 40625 3005
rect 40670 2885 40790 3005
rect 40835 2885 40955 3005
rect 41000 2885 41120 3005
rect 41175 2885 41295 3005
rect 41340 2885 41460 3005
rect 41505 2885 41625 3005
rect 41670 2885 41790 3005
rect 41845 2885 41965 3005
rect 36485 2720 36605 2840
rect 36650 2720 36770 2840
rect 36815 2720 36935 2840
rect 36980 2720 37100 2840
rect 37155 2720 37275 2840
rect 37320 2720 37440 2840
rect 37485 2720 37605 2840
rect 37650 2720 37770 2840
rect 37825 2720 37945 2840
rect 37990 2720 38110 2840
rect 38155 2720 38275 2840
rect 38320 2720 38440 2840
rect 38495 2720 38615 2840
rect 38660 2720 38780 2840
rect 38825 2720 38945 2840
rect 38990 2720 39110 2840
rect 39165 2720 39285 2840
rect 39330 2720 39450 2840
rect 39495 2720 39615 2840
rect 39660 2720 39780 2840
rect 39835 2720 39955 2840
rect 40000 2720 40120 2840
rect 40165 2720 40285 2840
rect 40330 2720 40450 2840
rect 40505 2720 40625 2840
rect 40670 2720 40790 2840
rect 40835 2720 40955 2840
rect 41000 2720 41120 2840
rect 41175 2720 41295 2840
rect 41340 2720 41460 2840
rect 41505 2720 41625 2840
rect 41670 2720 41790 2840
rect 41845 2720 41965 2840
rect 36485 2555 36605 2675
rect 36650 2555 36770 2675
rect 36815 2555 36935 2675
rect 36980 2555 37100 2675
rect 37155 2555 37275 2675
rect 37320 2555 37440 2675
rect 37485 2555 37605 2675
rect 37650 2555 37770 2675
rect 37825 2555 37945 2675
rect 37990 2555 38110 2675
rect 38155 2555 38275 2675
rect 38320 2555 38440 2675
rect 38495 2555 38615 2675
rect 38660 2555 38780 2675
rect 38825 2555 38945 2675
rect 38990 2555 39110 2675
rect 39165 2555 39285 2675
rect 39330 2555 39450 2675
rect 39495 2555 39615 2675
rect 39660 2555 39780 2675
rect 39835 2555 39955 2675
rect 40000 2555 40120 2675
rect 40165 2555 40285 2675
rect 40330 2555 40450 2675
rect 40505 2555 40625 2675
rect 40670 2555 40790 2675
rect 40835 2555 40955 2675
rect 41000 2555 41120 2675
rect 41175 2555 41295 2675
rect 41340 2555 41460 2675
rect 41505 2555 41625 2675
rect 41670 2555 41790 2675
rect 41845 2555 41965 2675
rect 36485 2390 36605 2510
rect 36650 2390 36770 2510
rect 36815 2390 36935 2510
rect 36980 2390 37100 2510
rect 37155 2390 37275 2510
rect 37320 2390 37440 2510
rect 37485 2390 37605 2510
rect 37650 2390 37770 2510
rect 37825 2390 37945 2510
rect 37990 2390 38110 2510
rect 38155 2390 38275 2510
rect 38320 2390 38440 2510
rect 38495 2390 38615 2510
rect 38660 2390 38780 2510
rect 38825 2390 38945 2510
rect 38990 2390 39110 2510
rect 39165 2390 39285 2510
rect 39330 2390 39450 2510
rect 39495 2390 39615 2510
rect 39660 2390 39780 2510
rect 39835 2390 39955 2510
rect 40000 2390 40120 2510
rect 40165 2390 40285 2510
rect 40330 2390 40450 2510
rect 40505 2390 40625 2510
rect 40670 2390 40790 2510
rect 40835 2390 40955 2510
rect 41000 2390 41120 2510
rect 41175 2390 41295 2510
rect 41340 2390 41460 2510
rect 41505 2390 41625 2510
rect 41670 2390 41790 2510
rect 41845 2390 41965 2510
rect 36485 2215 36605 2335
rect 36650 2215 36770 2335
rect 36815 2215 36935 2335
rect 36980 2215 37100 2335
rect 37155 2215 37275 2335
rect 37320 2215 37440 2335
rect 37485 2215 37605 2335
rect 37650 2215 37770 2335
rect 37825 2215 37945 2335
rect 37990 2215 38110 2335
rect 38155 2215 38275 2335
rect 38320 2215 38440 2335
rect 38495 2215 38615 2335
rect 38660 2215 38780 2335
rect 38825 2215 38945 2335
rect 38990 2215 39110 2335
rect 39165 2215 39285 2335
rect 39330 2215 39450 2335
rect 39495 2215 39615 2335
rect 39660 2215 39780 2335
rect 39835 2215 39955 2335
rect 40000 2215 40120 2335
rect 40165 2215 40285 2335
rect 40330 2215 40450 2335
rect 40505 2215 40625 2335
rect 40670 2215 40790 2335
rect 40835 2215 40955 2335
rect 41000 2215 41120 2335
rect 41175 2215 41295 2335
rect 41340 2215 41460 2335
rect 41505 2215 41625 2335
rect 41670 2215 41790 2335
rect 41845 2215 41965 2335
rect 36485 2050 36605 2170
rect 36650 2050 36770 2170
rect 36815 2050 36935 2170
rect 36980 2050 37100 2170
rect 37155 2050 37275 2170
rect 37320 2050 37440 2170
rect 37485 2050 37605 2170
rect 37650 2050 37770 2170
rect 37825 2050 37945 2170
rect 37990 2050 38110 2170
rect 38155 2050 38275 2170
rect 38320 2050 38440 2170
rect 38495 2050 38615 2170
rect 38660 2050 38780 2170
rect 38825 2050 38945 2170
rect 38990 2050 39110 2170
rect 39165 2050 39285 2170
rect 39330 2050 39450 2170
rect 39495 2050 39615 2170
rect 39660 2050 39780 2170
rect 39835 2050 39955 2170
rect 40000 2050 40120 2170
rect 40165 2050 40285 2170
rect 40330 2050 40450 2170
rect 40505 2050 40625 2170
rect 40670 2050 40790 2170
rect 40835 2050 40955 2170
rect 41000 2050 41120 2170
rect 41175 2050 41295 2170
rect 41340 2050 41460 2170
rect 41505 2050 41625 2170
rect 41670 2050 41790 2170
rect 41845 2050 41965 2170
rect 36485 1885 36605 2005
rect 36650 1885 36770 2005
rect 36815 1885 36935 2005
rect 36980 1885 37100 2005
rect 37155 1885 37275 2005
rect 37320 1885 37440 2005
rect 37485 1885 37605 2005
rect 37650 1885 37770 2005
rect 37825 1885 37945 2005
rect 37990 1885 38110 2005
rect 38155 1885 38275 2005
rect 38320 1885 38440 2005
rect 38495 1885 38615 2005
rect 38660 1885 38780 2005
rect 38825 1885 38945 2005
rect 38990 1885 39110 2005
rect 39165 1885 39285 2005
rect 39330 1885 39450 2005
rect 39495 1885 39615 2005
rect 39660 1885 39780 2005
rect 39835 1885 39955 2005
rect 40000 1885 40120 2005
rect 40165 1885 40285 2005
rect 40330 1885 40450 2005
rect 40505 1885 40625 2005
rect 40670 1885 40790 2005
rect 40835 1885 40955 2005
rect 41000 1885 41120 2005
rect 41175 1885 41295 2005
rect 41340 1885 41460 2005
rect 41505 1885 41625 2005
rect 41670 1885 41790 2005
rect 41845 1885 41965 2005
rect 36485 1720 36605 1840
rect 36650 1720 36770 1840
rect 36815 1720 36935 1840
rect 36980 1720 37100 1840
rect 37155 1720 37275 1840
rect 37320 1720 37440 1840
rect 37485 1720 37605 1840
rect 37650 1720 37770 1840
rect 37825 1720 37945 1840
rect 37990 1720 38110 1840
rect 38155 1720 38275 1840
rect 38320 1720 38440 1840
rect 38495 1720 38615 1840
rect 38660 1720 38780 1840
rect 38825 1720 38945 1840
rect 38990 1720 39110 1840
rect 39165 1720 39285 1840
rect 39330 1720 39450 1840
rect 39495 1720 39615 1840
rect 39660 1720 39780 1840
rect 39835 1720 39955 1840
rect 40000 1720 40120 1840
rect 40165 1720 40285 1840
rect 40330 1720 40450 1840
rect 40505 1720 40625 1840
rect 40670 1720 40790 1840
rect 40835 1720 40955 1840
rect 41000 1720 41120 1840
rect 41175 1720 41295 1840
rect 41340 1720 41460 1840
rect 41505 1720 41625 1840
rect 41670 1720 41790 1840
rect 41845 1720 41965 1840
rect 42175 7080 42295 7200
rect 42340 7080 42460 7200
rect 42505 7080 42625 7200
rect 42670 7080 42790 7200
rect 42845 7080 42965 7200
rect 43010 7080 43130 7200
rect 43175 7080 43295 7200
rect 43340 7080 43460 7200
rect 43515 7080 43635 7200
rect 43680 7080 43800 7200
rect 43845 7080 43965 7200
rect 44010 7080 44130 7200
rect 44185 7080 44305 7200
rect 44350 7080 44470 7200
rect 44515 7080 44635 7200
rect 44680 7080 44800 7200
rect 44855 7080 44975 7200
rect 45020 7080 45140 7200
rect 45185 7080 45305 7200
rect 45350 7080 45470 7200
rect 45525 7080 45645 7200
rect 45690 7080 45810 7200
rect 45855 7080 45975 7200
rect 46020 7080 46140 7200
rect 46195 7080 46315 7200
rect 46360 7080 46480 7200
rect 46525 7080 46645 7200
rect 46690 7080 46810 7200
rect 46865 7080 46985 7200
rect 47030 7080 47150 7200
rect 47195 7080 47315 7200
rect 47360 7080 47480 7200
rect 47535 7080 47655 7200
rect 42175 6905 42295 7025
rect 42340 6905 42460 7025
rect 42505 6905 42625 7025
rect 42670 6905 42790 7025
rect 42845 6905 42965 7025
rect 43010 6905 43130 7025
rect 43175 6905 43295 7025
rect 43340 6905 43460 7025
rect 43515 6905 43635 7025
rect 43680 6905 43800 7025
rect 43845 6905 43965 7025
rect 44010 6905 44130 7025
rect 44185 6905 44305 7025
rect 44350 6905 44470 7025
rect 44515 6905 44635 7025
rect 44680 6905 44800 7025
rect 44855 6905 44975 7025
rect 45020 6905 45140 7025
rect 45185 6905 45305 7025
rect 45350 6905 45470 7025
rect 45525 6905 45645 7025
rect 45690 6905 45810 7025
rect 45855 6905 45975 7025
rect 46020 6905 46140 7025
rect 46195 6905 46315 7025
rect 46360 6905 46480 7025
rect 46525 6905 46645 7025
rect 46690 6905 46810 7025
rect 46865 6905 46985 7025
rect 47030 6905 47150 7025
rect 47195 6905 47315 7025
rect 47360 6905 47480 7025
rect 47535 6905 47655 7025
rect 42175 6740 42295 6860
rect 42340 6740 42460 6860
rect 42505 6740 42625 6860
rect 42670 6740 42790 6860
rect 42845 6740 42965 6860
rect 43010 6740 43130 6860
rect 43175 6740 43295 6860
rect 43340 6740 43460 6860
rect 43515 6740 43635 6860
rect 43680 6740 43800 6860
rect 43845 6740 43965 6860
rect 44010 6740 44130 6860
rect 44185 6740 44305 6860
rect 44350 6740 44470 6860
rect 44515 6740 44635 6860
rect 44680 6740 44800 6860
rect 44855 6740 44975 6860
rect 45020 6740 45140 6860
rect 45185 6740 45305 6860
rect 45350 6740 45470 6860
rect 45525 6740 45645 6860
rect 45690 6740 45810 6860
rect 45855 6740 45975 6860
rect 46020 6740 46140 6860
rect 46195 6740 46315 6860
rect 46360 6740 46480 6860
rect 46525 6740 46645 6860
rect 46690 6740 46810 6860
rect 46865 6740 46985 6860
rect 47030 6740 47150 6860
rect 47195 6740 47315 6860
rect 47360 6740 47480 6860
rect 47535 6740 47655 6860
rect 42175 6575 42295 6695
rect 42340 6575 42460 6695
rect 42505 6575 42625 6695
rect 42670 6575 42790 6695
rect 42845 6575 42965 6695
rect 43010 6575 43130 6695
rect 43175 6575 43295 6695
rect 43340 6575 43460 6695
rect 43515 6575 43635 6695
rect 43680 6575 43800 6695
rect 43845 6575 43965 6695
rect 44010 6575 44130 6695
rect 44185 6575 44305 6695
rect 44350 6575 44470 6695
rect 44515 6575 44635 6695
rect 44680 6575 44800 6695
rect 44855 6575 44975 6695
rect 45020 6575 45140 6695
rect 45185 6575 45305 6695
rect 45350 6575 45470 6695
rect 45525 6575 45645 6695
rect 45690 6575 45810 6695
rect 45855 6575 45975 6695
rect 46020 6575 46140 6695
rect 46195 6575 46315 6695
rect 46360 6575 46480 6695
rect 46525 6575 46645 6695
rect 46690 6575 46810 6695
rect 46865 6575 46985 6695
rect 47030 6575 47150 6695
rect 47195 6575 47315 6695
rect 47360 6575 47480 6695
rect 47535 6575 47655 6695
rect 42175 6410 42295 6530
rect 42340 6410 42460 6530
rect 42505 6410 42625 6530
rect 42670 6410 42790 6530
rect 42845 6410 42965 6530
rect 43010 6410 43130 6530
rect 43175 6410 43295 6530
rect 43340 6410 43460 6530
rect 43515 6410 43635 6530
rect 43680 6410 43800 6530
rect 43845 6410 43965 6530
rect 44010 6410 44130 6530
rect 44185 6410 44305 6530
rect 44350 6410 44470 6530
rect 44515 6410 44635 6530
rect 44680 6410 44800 6530
rect 44855 6410 44975 6530
rect 45020 6410 45140 6530
rect 45185 6410 45305 6530
rect 45350 6410 45470 6530
rect 45525 6410 45645 6530
rect 45690 6410 45810 6530
rect 45855 6410 45975 6530
rect 46020 6410 46140 6530
rect 46195 6410 46315 6530
rect 46360 6410 46480 6530
rect 46525 6410 46645 6530
rect 46690 6410 46810 6530
rect 46865 6410 46985 6530
rect 47030 6410 47150 6530
rect 47195 6410 47315 6530
rect 47360 6410 47480 6530
rect 47535 6410 47655 6530
rect 42175 6235 42295 6355
rect 42340 6235 42460 6355
rect 42505 6235 42625 6355
rect 42670 6235 42790 6355
rect 42845 6235 42965 6355
rect 43010 6235 43130 6355
rect 43175 6235 43295 6355
rect 43340 6235 43460 6355
rect 43515 6235 43635 6355
rect 43680 6235 43800 6355
rect 43845 6235 43965 6355
rect 44010 6235 44130 6355
rect 44185 6235 44305 6355
rect 44350 6235 44470 6355
rect 44515 6235 44635 6355
rect 44680 6235 44800 6355
rect 44855 6235 44975 6355
rect 45020 6235 45140 6355
rect 45185 6235 45305 6355
rect 45350 6235 45470 6355
rect 45525 6235 45645 6355
rect 45690 6235 45810 6355
rect 45855 6235 45975 6355
rect 46020 6235 46140 6355
rect 46195 6235 46315 6355
rect 46360 6235 46480 6355
rect 46525 6235 46645 6355
rect 46690 6235 46810 6355
rect 46865 6235 46985 6355
rect 47030 6235 47150 6355
rect 47195 6235 47315 6355
rect 47360 6235 47480 6355
rect 47535 6235 47655 6355
rect 42175 6070 42295 6190
rect 42340 6070 42460 6190
rect 42505 6070 42625 6190
rect 42670 6070 42790 6190
rect 42845 6070 42965 6190
rect 43010 6070 43130 6190
rect 43175 6070 43295 6190
rect 43340 6070 43460 6190
rect 43515 6070 43635 6190
rect 43680 6070 43800 6190
rect 43845 6070 43965 6190
rect 44010 6070 44130 6190
rect 44185 6070 44305 6190
rect 44350 6070 44470 6190
rect 44515 6070 44635 6190
rect 44680 6070 44800 6190
rect 44855 6070 44975 6190
rect 45020 6070 45140 6190
rect 45185 6070 45305 6190
rect 45350 6070 45470 6190
rect 45525 6070 45645 6190
rect 45690 6070 45810 6190
rect 45855 6070 45975 6190
rect 46020 6070 46140 6190
rect 46195 6070 46315 6190
rect 46360 6070 46480 6190
rect 46525 6070 46645 6190
rect 46690 6070 46810 6190
rect 46865 6070 46985 6190
rect 47030 6070 47150 6190
rect 47195 6070 47315 6190
rect 47360 6070 47480 6190
rect 47535 6070 47655 6190
rect 42175 5905 42295 6025
rect 42340 5905 42460 6025
rect 42505 5905 42625 6025
rect 42670 5905 42790 6025
rect 42845 5905 42965 6025
rect 43010 5905 43130 6025
rect 43175 5905 43295 6025
rect 43340 5905 43460 6025
rect 43515 5905 43635 6025
rect 43680 5905 43800 6025
rect 43845 5905 43965 6025
rect 44010 5905 44130 6025
rect 44185 5905 44305 6025
rect 44350 5905 44470 6025
rect 44515 5905 44635 6025
rect 44680 5905 44800 6025
rect 44855 5905 44975 6025
rect 45020 5905 45140 6025
rect 45185 5905 45305 6025
rect 45350 5905 45470 6025
rect 45525 5905 45645 6025
rect 45690 5905 45810 6025
rect 45855 5905 45975 6025
rect 46020 5905 46140 6025
rect 46195 5905 46315 6025
rect 46360 5905 46480 6025
rect 46525 5905 46645 6025
rect 46690 5905 46810 6025
rect 46865 5905 46985 6025
rect 47030 5905 47150 6025
rect 47195 5905 47315 6025
rect 47360 5905 47480 6025
rect 47535 5905 47655 6025
rect 42175 5740 42295 5860
rect 42340 5740 42460 5860
rect 42505 5740 42625 5860
rect 42670 5740 42790 5860
rect 42845 5740 42965 5860
rect 43010 5740 43130 5860
rect 43175 5740 43295 5860
rect 43340 5740 43460 5860
rect 43515 5740 43635 5860
rect 43680 5740 43800 5860
rect 43845 5740 43965 5860
rect 44010 5740 44130 5860
rect 44185 5740 44305 5860
rect 44350 5740 44470 5860
rect 44515 5740 44635 5860
rect 44680 5740 44800 5860
rect 44855 5740 44975 5860
rect 45020 5740 45140 5860
rect 45185 5740 45305 5860
rect 45350 5740 45470 5860
rect 45525 5740 45645 5860
rect 45690 5740 45810 5860
rect 45855 5740 45975 5860
rect 46020 5740 46140 5860
rect 46195 5740 46315 5860
rect 46360 5740 46480 5860
rect 46525 5740 46645 5860
rect 46690 5740 46810 5860
rect 46865 5740 46985 5860
rect 47030 5740 47150 5860
rect 47195 5740 47315 5860
rect 47360 5740 47480 5860
rect 47535 5740 47655 5860
rect 42175 5565 42295 5685
rect 42340 5565 42460 5685
rect 42505 5565 42625 5685
rect 42670 5565 42790 5685
rect 42845 5565 42965 5685
rect 43010 5565 43130 5685
rect 43175 5565 43295 5685
rect 43340 5565 43460 5685
rect 43515 5565 43635 5685
rect 43680 5565 43800 5685
rect 43845 5565 43965 5685
rect 44010 5565 44130 5685
rect 44185 5565 44305 5685
rect 44350 5565 44470 5685
rect 44515 5565 44635 5685
rect 44680 5565 44800 5685
rect 44855 5565 44975 5685
rect 45020 5565 45140 5685
rect 45185 5565 45305 5685
rect 45350 5565 45470 5685
rect 45525 5565 45645 5685
rect 45690 5565 45810 5685
rect 45855 5565 45975 5685
rect 46020 5565 46140 5685
rect 46195 5565 46315 5685
rect 46360 5565 46480 5685
rect 46525 5565 46645 5685
rect 46690 5565 46810 5685
rect 46865 5565 46985 5685
rect 47030 5565 47150 5685
rect 47195 5565 47315 5685
rect 47360 5565 47480 5685
rect 47535 5565 47655 5685
rect 42175 5400 42295 5520
rect 42340 5400 42460 5520
rect 42505 5400 42625 5520
rect 42670 5400 42790 5520
rect 42845 5400 42965 5520
rect 43010 5400 43130 5520
rect 43175 5400 43295 5520
rect 43340 5400 43460 5520
rect 43515 5400 43635 5520
rect 43680 5400 43800 5520
rect 43845 5400 43965 5520
rect 44010 5400 44130 5520
rect 44185 5400 44305 5520
rect 44350 5400 44470 5520
rect 44515 5400 44635 5520
rect 44680 5400 44800 5520
rect 44855 5400 44975 5520
rect 45020 5400 45140 5520
rect 45185 5400 45305 5520
rect 45350 5400 45470 5520
rect 45525 5400 45645 5520
rect 45690 5400 45810 5520
rect 45855 5400 45975 5520
rect 46020 5400 46140 5520
rect 46195 5400 46315 5520
rect 46360 5400 46480 5520
rect 46525 5400 46645 5520
rect 46690 5400 46810 5520
rect 46865 5400 46985 5520
rect 47030 5400 47150 5520
rect 47195 5400 47315 5520
rect 47360 5400 47480 5520
rect 47535 5400 47655 5520
rect 42175 5235 42295 5355
rect 42340 5235 42460 5355
rect 42505 5235 42625 5355
rect 42670 5235 42790 5355
rect 42845 5235 42965 5355
rect 43010 5235 43130 5355
rect 43175 5235 43295 5355
rect 43340 5235 43460 5355
rect 43515 5235 43635 5355
rect 43680 5235 43800 5355
rect 43845 5235 43965 5355
rect 44010 5235 44130 5355
rect 44185 5235 44305 5355
rect 44350 5235 44470 5355
rect 44515 5235 44635 5355
rect 44680 5235 44800 5355
rect 44855 5235 44975 5355
rect 45020 5235 45140 5355
rect 45185 5235 45305 5355
rect 45350 5235 45470 5355
rect 45525 5235 45645 5355
rect 45690 5235 45810 5355
rect 45855 5235 45975 5355
rect 46020 5235 46140 5355
rect 46195 5235 46315 5355
rect 46360 5235 46480 5355
rect 46525 5235 46645 5355
rect 46690 5235 46810 5355
rect 46865 5235 46985 5355
rect 47030 5235 47150 5355
rect 47195 5235 47315 5355
rect 47360 5235 47480 5355
rect 47535 5235 47655 5355
rect 42175 5070 42295 5190
rect 42340 5070 42460 5190
rect 42505 5070 42625 5190
rect 42670 5070 42790 5190
rect 42845 5070 42965 5190
rect 43010 5070 43130 5190
rect 43175 5070 43295 5190
rect 43340 5070 43460 5190
rect 43515 5070 43635 5190
rect 43680 5070 43800 5190
rect 43845 5070 43965 5190
rect 44010 5070 44130 5190
rect 44185 5070 44305 5190
rect 44350 5070 44470 5190
rect 44515 5070 44635 5190
rect 44680 5070 44800 5190
rect 44855 5070 44975 5190
rect 45020 5070 45140 5190
rect 45185 5070 45305 5190
rect 45350 5070 45470 5190
rect 45525 5070 45645 5190
rect 45690 5070 45810 5190
rect 45855 5070 45975 5190
rect 46020 5070 46140 5190
rect 46195 5070 46315 5190
rect 46360 5070 46480 5190
rect 46525 5070 46645 5190
rect 46690 5070 46810 5190
rect 46865 5070 46985 5190
rect 47030 5070 47150 5190
rect 47195 5070 47315 5190
rect 47360 5070 47480 5190
rect 47535 5070 47655 5190
rect 42175 4895 42295 5015
rect 42340 4895 42460 5015
rect 42505 4895 42625 5015
rect 42670 4895 42790 5015
rect 42845 4895 42965 5015
rect 43010 4895 43130 5015
rect 43175 4895 43295 5015
rect 43340 4895 43460 5015
rect 43515 4895 43635 5015
rect 43680 4895 43800 5015
rect 43845 4895 43965 5015
rect 44010 4895 44130 5015
rect 44185 4895 44305 5015
rect 44350 4895 44470 5015
rect 44515 4895 44635 5015
rect 44680 4895 44800 5015
rect 44855 4895 44975 5015
rect 45020 4895 45140 5015
rect 45185 4895 45305 5015
rect 45350 4895 45470 5015
rect 45525 4895 45645 5015
rect 45690 4895 45810 5015
rect 45855 4895 45975 5015
rect 46020 4895 46140 5015
rect 46195 4895 46315 5015
rect 46360 4895 46480 5015
rect 46525 4895 46645 5015
rect 46690 4895 46810 5015
rect 46865 4895 46985 5015
rect 47030 4895 47150 5015
rect 47195 4895 47315 5015
rect 47360 4895 47480 5015
rect 47535 4895 47655 5015
rect 42175 4730 42295 4850
rect 42340 4730 42460 4850
rect 42505 4730 42625 4850
rect 42670 4730 42790 4850
rect 42845 4730 42965 4850
rect 43010 4730 43130 4850
rect 43175 4730 43295 4850
rect 43340 4730 43460 4850
rect 43515 4730 43635 4850
rect 43680 4730 43800 4850
rect 43845 4730 43965 4850
rect 44010 4730 44130 4850
rect 44185 4730 44305 4850
rect 44350 4730 44470 4850
rect 44515 4730 44635 4850
rect 44680 4730 44800 4850
rect 44855 4730 44975 4850
rect 45020 4730 45140 4850
rect 45185 4730 45305 4850
rect 45350 4730 45470 4850
rect 45525 4730 45645 4850
rect 45690 4730 45810 4850
rect 45855 4730 45975 4850
rect 46020 4730 46140 4850
rect 46195 4730 46315 4850
rect 46360 4730 46480 4850
rect 46525 4730 46645 4850
rect 46690 4730 46810 4850
rect 46865 4730 46985 4850
rect 47030 4730 47150 4850
rect 47195 4730 47315 4850
rect 47360 4730 47480 4850
rect 47535 4730 47655 4850
rect 42175 4565 42295 4685
rect 42340 4565 42460 4685
rect 42505 4565 42625 4685
rect 42670 4565 42790 4685
rect 42845 4565 42965 4685
rect 43010 4565 43130 4685
rect 43175 4565 43295 4685
rect 43340 4565 43460 4685
rect 43515 4565 43635 4685
rect 43680 4565 43800 4685
rect 43845 4565 43965 4685
rect 44010 4565 44130 4685
rect 44185 4565 44305 4685
rect 44350 4565 44470 4685
rect 44515 4565 44635 4685
rect 44680 4565 44800 4685
rect 44855 4565 44975 4685
rect 45020 4565 45140 4685
rect 45185 4565 45305 4685
rect 45350 4565 45470 4685
rect 45525 4565 45645 4685
rect 45690 4565 45810 4685
rect 45855 4565 45975 4685
rect 46020 4565 46140 4685
rect 46195 4565 46315 4685
rect 46360 4565 46480 4685
rect 46525 4565 46645 4685
rect 46690 4565 46810 4685
rect 46865 4565 46985 4685
rect 47030 4565 47150 4685
rect 47195 4565 47315 4685
rect 47360 4565 47480 4685
rect 47535 4565 47655 4685
rect 42175 4400 42295 4520
rect 42340 4400 42460 4520
rect 42505 4400 42625 4520
rect 42670 4400 42790 4520
rect 42845 4400 42965 4520
rect 43010 4400 43130 4520
rect 43175 4400 43295 4520
rect 43340 4400 43460 4520
rect 43515 4400 43635 4520
rect 43680 4400 43800 4520
rect 43845 4400 43965 4520
rect 44010 4400 44130 4520
rect 44185 4400 44305 4520
rect 44350 4400 44470 4520
rect 44515 4400 44635 4520
rect 44680 4400 44800 4520
rect 44855 4400 44975 4520
rect 45020 4400 45140 4520
rect 45185 4400 45305 4520
rect 45350 4400 45470 4520
rect 45525 4400 45645 4520
rect 45690 4400 45810 4520
rect 45855 4400 45975 4520
rect 46020 4400 46140 4520
rect 46195 4400 46315 4520
rect 46360 4400 46480 4520
rect 46525 4400 46645 4520
rect 46690 4400 46810 4520
rect 46865 4400 46985 4520
rect 47030 4400 47150 4520
rect 47195 4400 47315 4520
rect 47360 4400 47480 4520
rect 47535 4400 47655 4520
rect 42175 4225 42295 4345
rect 42340 4225 42460 4345
rect 42505 4225 42625 4345
rect 42670 4225 42790 4345
rect 42845 4225 42965 4345
rect 43010 4225 43130 4345
rect 43175 4225 43295 4345
rect 43340 4225 43460 4345
rect 43515 4225 43635 4345
rect 43680 4225 43800 4345
rect 43845 4225 43965 4345
rect 44010 4225 44130 4345
rect 44185 4225 44305 4345
rect 44350 4225 44470 4345
rect 44515 4225 44635 4345
rect 44680 4225 44800 4345
rect 44855 4225 44975 4345
rect 45020 4225 45140 4345
rect 45185 4225 45305 4345
rect 45350 4225 45470 4345
rect 45525 4225 45645 4345
rect 45690 4225 45810 4345
rect 45855 4225 45975 4345
rect 46020 4225 46140 4345
rect 46195 4225 46315 4345
rect 46360 4225 46480 4345
rect 46525 4225 46645 4345
rect 46690 4225 46810 4345
rect 46865 4225 46985 4345
rect 47030 4225 47150 4345
rect 47195 4225 47315 4345
rect 47360 4225 47480 4345
rect 47535 4225 47655 4345
rect 42175 4060 42295 4180
rect 42340 4060 42460 4180
rect 42505 4060 42625 4180
rect 42670 4060 42790 4180
rect 42845 4060 42965 4180
rect 43010 4060 43130 4180
rect 43175 4060 43295 4180
rect 43340 4060 43460 4180
rect 43515 4060 43635 4180
rect 43680 4060 43800 4180
rect 43845 4060 43965 4180
rect 44010 4060 44130 4180
rect 44185 4060 44305 4180
rect 44350 4060 44470 4180
rect 44515 4060 44635 4180
rect 44680 4060 44800 4180
rect 44855 4060 44975 4180
rect 45020 4060 45140 4180
rect 45185 4060 45305 4180
rect 45350 4060 45470 4180
rect 45525 4060 45645 4180
rect 45690 4060 45810 4180
rect 45855 4060 45975 4180
rect 46020 4060 46140 4180
rect 46195 4060 46315 4180
rect 46360 4060 46480 4180
rect 46525 4060 46645 4180
rect 46690 4060 46810 4180
rect 46865 4060 46985 4180
rect 47030 4060 47150 4180
rect 47195 4060 47315 4180
rect 47360 4060 47480 4180
rect 47535 4060 47655 4180
rect 42175 3895 42295 4015
rect 42340 3895 42460 4015
rect 42505 3895 42625 4015
rect 42670 3895 42790 4015
rect 42845 3895 42965 4015
rect 43010 3895 43130 4015
rect 43175 3895 43295 4015
rect 43340 3895 43460 4015
rect 43515 3895 43635 4015
rect 43680 3895 43800 4015
rect 43845 3895 43965 4015
rect 44010 3895 44130 4015
rect 44185 3895 44305 4015
rect 44350 3895 44470 4015
rect 44515 3895 44635 4015
rect 44680 3895 44800 4015
rect 44855 3895 44975 4015
rect 45020 3895 45140 4015
rect 45185 3895 45305 4015
rect 45350 3895 45470 4015
rect 45525 3895 45645 4015
rect 45690 3895 45810 4015
rect 45855 3895 45975 4015
rect 46020 3895 46140 4015
rect 46195 3895 46315 4015
rect 46360 3895 46480 4015
rect 46525 3895 46645 4015
rect 46690 3895 46810 4015
rect 46865 3895 46985 4015
rect 47030 3895 47150 4015
rect 47195 3895 47315 4015
rect 47360 3895 47480 4015
rect 47535 3895 47655 4015
rect 42175 3730 42295 3850
rect 42340 3730 42460 3850
rect 42505 3730 42625 3850
rect 42670 3730 42790 3850
rect 42845 3730 42965 3850
rect 43010 3730 43130 3850
rect 43175 3730 43295 3850
rect 43340 3730 43460 3850
rect 43515 3730 43635 3850
rect 43680 3730 43800 3850
rect 43845 3730 43965 3850
rect 44010 3730 44130 3850
rect 44185 3730 44305 3850
rect 44350 3730 44470 3850
rect 44515 3730 44635 3850
rect 44680 3730 44800 3850
rect 44855 3730 44975 3850
rect 45020 3730 45140 3850
rect 45185 3730 45305 3850
rect 45350 3730 45470 3850
rect 45525 3730 45645 3850
rect 45690 3730 45810 3850
rect 45855 3730 45975 3850
rect 46020 3730 46140 3850
rect 46195 3730 46315 3850
rect 46360 3730 46480 3850
rect 46525 3730 46645 3850
rect 46690 3730 46810 3850
rect 46865 3730 46985 3850
rect 47030 3730 47150 3850
rect 47195 3730 47315 3850
rect 47360 3730 47480 3850
rect 47535 3730 47655 3850
rect 42175 3555 42295 3675
rect 42340 3555 42460 3675
rect 42505 3555 42625 3675
rect 42670 3555 42790 3675
rect 42845 3555 42965 3675
rect 43010 3555 43130 3675
rect 43175 3555 43295 3675
rect 43340 3555 43460 3675
rect 43515 3555 43635 3675
rect 43680 3555 43800 3675
rect 43845 3555 43965 3675
rect 44010 3555 44130 3675
rect 44185 3555 44305 3675
rect 44350 3555 44470 3675
rect 44515 3555 44635 3675
rect 44680 3555 44800 3675
rect 44855 3555 44975 3675
rect 45020 3555 45140 3675
rect 45185 3555 45305 3675
rect 45350 3555 45470 3675
rect 45525 3555 45645 3675
rect 45690 3555 45810 3675
rect 45855 3555 45975 3675
rect 46020 3555 46140 3675
rect 46195 3555 46315 3675
rect 46360 3555 46480 3675
rect 46525 3555 46645 3675
rect 46690 3555 46810 3675
rect 46865 3555 46985 3675
rect 47030 3555 47150 3675
rect 47195 3555 47315 3675
rect 47360 3555 47480 3675
rect 47535 3555 47655 3675
rect 42175 3390 42295 3510
rect 42340 3390 42460 3510
rect 42505 3390 42625 3510
rect 42670 3390 42790 3510
rect 42845 3390 42965 3510
rect 43010 3390 43130 3510
rect 43175 3390 43295 3510
rect 43340 3390 43460 3510
rect 43515 3390 43635 3510
rect 43680 3390 43800 3510
rect 43845 3390 43965 3510
rect 44010 3390 44130 3510
rect 44185 3390 44305 3510
rect 44350 3390 44470 3510
rect 44515 3390 44635 3510
rect 44680 3390 44800 3510
rect 44855 3390 44975 3510
rect 45020 3390 45140 3510
rect 45185 3390 45305 3510
rect 45350 3390 45470 3510
rect 45525 3390 45645 3510
rect 45690 3390 45810 3510
rect 45855 3390 45975 3510
rect 46020 3390 46140 3510
rect 46195 3390 46315 3510
rect 46360 3390 46480 3510
rect 46525 3390 46645 3510
rect 46690 3390 46810 3510
rect 46865 3390 46985 3510
rect 47030 3390 47150 3510
rect 47195 3390 47315 3510
rect 47360 3390 47480 3510
rect 47535 3390 47655 3510
rect 42175 3225 42295 3345
rect 42340 3225 42460 3345
rect 42505 3225 42625 3345
rect 42670 3225 42790 3345
rect 42845 3225 42965 3345
rect 43010 3225 43130 3345
rect 43175 3225 43295 3345
rect 43340 3225 43460 3345
rect 43515 3225 43635 3345
rect 43680 3225 43800 3345
rect 43845 3225 43965 3345
rect 44010 3225 44130 3345
rect 44185 3225 44305 3345
rect 44350 3225 44470 3345
rect 44515 3225 44635 3345
rect 44680 3225 44800 3345
rect 44855 3225 44975 3345
rect 45020 3225 45140 3345
rect 45185 3225 45305 3345
rect 45350 3225 45470 3345
rect 45525 3225 45645 3345
rect 45690 3225 45810 3345
rect 45855 3225 45975 3345
rect 46020 3225 46140 3345
rect 46195 3225 46315 3345
rect 46360 3225 46480 3345
rect 46525 3225 46645 3345
rect 46690 3225 46810 3345
rect 46865 3225 46985 3345
rect 47030 3225 47150 3345
rect 47195 3225 47315 3345
rect 47360 3225 47480 3345
rect 47535 3225 47655 3345
rect 42175 3060 42295 3180
rect 42340 3060 42460 3180
rect 42505 3060 42625 3180
rect 42670 3060 42790 3180
rect 42845 3060 42965 3180
rect 43010 3060 43130 3180
rect 43175 3060 43295 3180
rect 43340 3060 43460 3180
rect 43515 3060 43635 3180
rect 43680 3060 43800 3180
rect 43845 3060 43965 3180
rect 44010 3060 44130 3180
rect 44185 3060 44305 3180
rect 44350 3060 44470 3180
rect 44515 3060 44635 3180
rect 44680 3060 44800 3180
rect 44855 3060 44975 3180
rect 45020 3060 45140 3180
rect 45185 3060 45305 3180
rect 45350 3060 45470 3180
rect 45525 3060 45645 3180
rect 45690 3060 45810 3180
rect 45855 3060 45975 3180
rect 46020 3060 46140 3180
rect 46195 3060 46315 3180
rect 46360 3060 46480 3180
rect 46525 3060 46645 3180
rect 46690 3060 46810 3180
rect 46865 3060 46985 3180
rect 47030 3060 47150 3180
rect 47195 3060 47315 3180
rect 47360 3060 47480 3180
rect 47535 3060 47655 3180
rect 42175 2885 42295 3005
rect 42340 2885 42460 3005
rect 42505 2885 42625 3005
rect 42670 2885 42790 3005
rect 42845 2885 42965 3005
rect 43010 2885 43130 3005
rect 43175 2885 43295 3005
rect 43340 2885 43460 3005
rect 43515 2885 43635 3005
rect 43680 2885 43800 3005
rect 43845 2885 43965 3005
rect 44010 2885 44130 3005
rect 44185 2885 44305 3005
rect 44350 2885 44470 3005
rect 44515 2885 44635 3005
rect 44680 2885 44800 3005
rect 44855 2885 44975 3005
rect 45020 2885 45140 3005
rect 45185 2885 45305 3005
rect 45350 2885 45470 3005
rect 45525 2885 45645 3005
rect 45690 2885 45810 3005
rect 45855 2885 45975 3005
rect 46020 2885 46140 3005
rect 46195 2885 46315 3005
rect 46360 2885 46480 3005
rect 46525 2885 46645 3005
rect 46690 2885 46810 3005
rect 46865 2885 46985 3005
rect 47030 2885 47150 3005
rect 47195 2885 47315 3005
rect 47360 2885 47480 3005
rect 47535 2885 47655 3005
rect 42175 2720 42295 2840
rect 42340 2720 42460 2840
rect 42505 2720 42625 2840
rect 42670 2720 42790 2840
rect 42845 2720 42965 2840
rect 43010 2720 43130 2840
rect 43175 2720 43295 2840
rect 43340 2720 43460 2840
rect 43515 2720 43635 2840
rect 43680 2720 43800 2840
rect 43845 2720 43965 2840
rect 44010 2720 44130 2840
rect 44185 2720 44305 2840
rect 44350 2720 44470 2840
rect 44515 2720 44635 2840
rect 44680 2720 44800 2840
rect 44855 2720 44975 2840
rect 45020 2720 45140 2840
rect 45185 2720 45305 2840
rect 45350 2720 45470 2840
rect 45525 2720 45645 2840
rect 45690 2720 45810 2840
rect 45855 2720 45975 2840
rect 46020 2720 46140 2840
rect 46195 2720 46315 2840
rect 46360 2720 46480 2840
rect 46525 2720 46645 2840
rect 46690 2720 46810 2840
rect 46865 2720 46985 2840
rect 47030 2720 47150 2840
rect 47195 2720 47315 2840
rect 47360 2720 47480 2840
rect 47535 2720 47655 2840
rect 42175 2555 42295 2675
rect 42340 2555 42460 2675
rect 42505 2555 42625 2675
rect 42670 2555 42790 2675
rect 42845 2555 42965 2675
rect 43010 2555 43130 2675
rect 43175 2555 43295 2675
rect 43340 2555 43460 2675
rect 43515 2555 43635 2675
rect 43680 2555 43800 2675
rect 43845 2555 43965 2675
rect 44010 2555 44130 2675
rect 44185 2555 44305 2675
rect 44350 2555 44470 2675
rect 44515 2555 44635 2675
rect 44680 2555 44800 2675
rect 44855 2555 44975 2675
rect 45020 2555 45140 2675
rect 45185 2555 45305 2675
rect 45350 2555 45470 2675
rect 45525 2555 45645 2675
rect 45690 2555 45810 2675
rect 45855 2555 45975 2675
rect 46020 2555 46140 2675
rect 46195 2555 46315 2675
rect 46360 2555 46480 2675
rect 46525 2555 46645 2675
rect 46690 2555 46810 2675
rect 46865 2555 46985 2675
rect 47030 2555 47150 2675
rect 47195 2555 47315 2675
rect 47360 2555 47480 2675
rect 47535 2555 47655 2675
rect 42175 2390 42295 2510
rect 42340 2390 42460 2510
rect 42505 2390 42625 2510
rect 42670 2390 42790 2510
rect 42845 2390 42965 2510
rect 43010 2390 43130 2510
rect 43175 2390 43295 2510
rect 43340 2390 43460 2510
rect 43515 2390 43635 2510
rect 43680 2390 43800 2510
rect 43845 2390 43965 2510
rect 44010 2390 44130 2510
rect 44185 2390 44305 2510
rect 44350 2390 44470 2510
rect 44515 2390 44635 2510
rect 44680 2390 44800 2510
rect 44855 2390 44975 2510
rect 45020 2390 45140 2510
rect 45185 2390 45305 2510
rect 45350 2390 45470 2510
rect 45525 2390 45645 2510
rect 45690 2390 45810 2510
rect 45855 2390 45975 2510
rect 46020 2390 46140 2510
rect 46195 2390 46315 2510
rect 46360 2390 46480 2510
rect 46525 2390 46645 2510
rect 46690 2390 46810 2510
rect 46865 2390 46985 2510
rect 47030 2390 47150 2510
rect 47195 2390 47315 2510
rect 47360 2390 47480 2510
rect 47535 2390 47655 2510
rect 42175 2215 42295 2335
rect 42340 2215 42460 2335
rect 42505 2215 42625 2335
rect 42670 2215 42790 2335
rect 42845 2215 42965 2335
rect 43010 2215 43130 2335
rect 43175 2215 43295 2335
rect 43340 2215 43460 2335
rect 43515 2215 43635 2335
rect 43680 2215 43800 2335
rect 43845 2215 43965 2335
rect 44010 2215 44130 2335
rect 44185 2215 44305 2335
rect 44350 2215 44470 2335
rect 44515 2215 44635 2335
rect 44680 2215 44800 2335
rect 44855 2215 44975 2335
rect 45020 2215 45140 2335
rect 45185 2215 45305 2335
rect 45350 2215 45470 2335
rect 45525 2215 45645 2335
rect 45690 2215 45810 2335
rect 45855 2215 45975 2335
rect 46020 2215 46140 2335
rect 46195 2215 46315 2335
rect 46360 2215 46480 2335
rect 46525 2215 46645 2335
rect 46690 2215 46810 2335
rect 46865 2215 46985 2335
rect 47030 2215 47150 2335
rect 47195 2215 47315 2335
rect 47360 2215 47480 2335
rect 47535 2215 47655 2335
rect 42175 2050 42295 2170
rect 42340 2050 42460 2170
rect 42505 2050 42625 2170
rect 42670 2050 42790 2170
rect 42845 2050 42965 2170
rect 43010 2050 43130 2170
rect 43175 2050 43295 2170
rect 43340 2050 43460 2170
rect 43515 2050 43635 2170
rect 43680 2050 43800 2170
rect 43845 2050 43965 2170
rect 44010 2050 44130 2170
rect 44185 2050 44305 2170
rect 44350 2050 44470 2170
rect 44515 2050 44635 2170
rect 44680 2050 44800 2170
rect 44855 2050 44975 2170
rect 45020 2050 45140 2170
rect 45185 2050 45305 2170
rect 45350 2050 45470 2170
rect 45525 2050 45645 2170
rect 45690 2050 45810 2170
rect 45855 2050 45975 2170
rect 46020 2050 46140 2170
rect 46195 2050 46315 2170
rect 46360 2050 46480 2170
rect 46525 2050 46645 2170
rect 46690 2050 46810 2170
rect 46865 2050 46985 2170
rect 47030 2050 47150 2170
rect 47195 2050 47315 2170
rect 47360 2050 47480 2170
rect 47535 2050 47655 2170
rect 42175 1885 42295 2005
rect 42340 1885 42460 2005
rect 42505 1885 42625 2005
rect 42670 1885 42790 2005
rect 42845 1885 42965 2005
rect 43010 1885 43130 2005
rect 43175 1885 43295 2005
rect 43340 1885 43460 2005
rect 43515 1885 43635 2005
rect 43680 1885 43800 2005
rect 43845 1885 43965 2005
rect 44010 1885 44130 2005
rect 44185 1885 44305 2005
rect 44350 1885 44470 2005
rect 44515 1885 44635 2005
rect 44680 1885 44800 2005
rect 44855 1885 44975 2005
rect 45020 1885 45140 2005
rect 45185 1885 45305 2005
rect 45350 1885 45470 2005
rect 45525 1885 45645 2005
rect 45690 1885 45810 2005
rect 45855 1885 45975 2005
rect 46020 1885 46140 2005
rect 46195 1885 46315 2005
rect 46360 1885 46480 2005
rect 46525 1885 46645 2005
rect 46690 1885 46810 2005
rect 46865 1885 46985 2005
rect 47030 1885 47150 2005
rect 47195 1885 47315 2005
rect 47360 1885 47480 2005
rect 47535 1885 47655 2005
rect 42175 1720 42295 1840
rect 42340 1720 42460 1840
rect 42505 1720 42625 1840
rect 42670 1720 42790 1840
rect 42845 1720 42965 1840
rect 43010 1720 43130 1840
rect 43175 1720 43295 1840
rect 43340 1720 43460 1840
rect 43515 1720 43635 1840
rect 43680 1720 43800 1840
rect 43845 1720 43965 1840
rect 44010 1720 44130 1840
rect 44185 1720 44305 1840
rect 44350 1720 44470 1840
rect 44515 1720 44635 1840
rect 44680 1720 44800 1840
rect 44855 1720 44975 1840
rect 45020 1720 45140 1840
rect 45185 1720 45305 1840
rect 45350 1720 45470 1840
rect 45525 1720 45645 1840
rect 45690 1720 45810 1840
rect 45855 1720 45975 1840
rect 46020 1720 46140 1840
rect 46195 1720 46315 1840
rect 46360 1720 46480 1840
rect 46525 1720 46645 1840
rect 46690 1720 46810 1840
rect 46865 1720 46985 1840
rect 47030 1720 47150 1840
rect 47195 1720 47315 1840
rect 47360 1720 47480 1840
rect 47535 1720 47655 1840
rect 47865 7080 47985 7200
rect 48030 7080 48150 7200
rect 48195 7080 48315 7200
rect 48360 7080 48480 7200
rect 48535 7080 48655 7200
rect 48700 7080 48820 7200
rect 48865 7080 48985 7200
rect 49030 7080 49150 7200
rect 49205 7080 49325 7200
rect 49370 7080 49490 7200
rect 49535 7080 49655 7200
rect 49700 7080 49820 7200
rect 49875 7080 49995 7200
rect 50040 7080 50160 7200
rect 50205 7080 50325 7200
rect 50370 7080 50490 7200
rect 50545 7080 50665 7200
rect 50710 7080 50830 7200
rect 50875 7080 50995 7200
rect 51040 7080 51160 7200
rect 51215 7080 51335 7200
rect 51380 7080 51500 7200
rect 51545 7080 51665 7200
rect 51710 7080 51830 7200
rect 51885 7080 52005 7200
rect 52050 7080 52170 7200
rect 52215 7080 52335 7200
rect 52380 7080 52500 7200
rect 52555 7080 52675 7200
rect 52720 7080 52840 7200
rect 52885 7080 53005 7200
rect 53050 7080 53170 7200
rect 53225 7080 53345 7200
rect 47865 6905 47985 7025
rect 48030 6905 48150 7025
rect 48195 6905 48315 7025
rect 48360 6905 48480 7025
rect 48535 6905 48655 7025
rect 48700 6905 48820 7025
rect 48865 6905 48985 7025
rect 49030 6905 49150 7025
rect 49205 6905 49325 7025
rect 49370 6905 49490 7025
rect 49535 6905 49655 7025
rect 49700 6905 49820 7025
rect 49875 6905 49995 7025
rect 50040 6905 50160 7025
rect 50205 6905 50325 7025
rect 50370 6905 50490 7025
rect 50545 6905 50665 7025
rect 50710 6905 50830 7025
rect 50875 6905 50995 7025
rect 51040 6905 51160 7025
rect 51215 6905 51335 7025
rect 51380 6905 51500 7025
rect 51545 6905 51665 7025
rect 51710 6905 51830 7025
rect 51885 6905 52005 7025
rect 52050 6905 52170 7025
rect 52215 6905 52335 7025
rect 52380 6905 52500 7025
rect 52555 6905 52675 7025
rect 52720 6905 52840 7025
rect 52885 6905 53005 7025
rect 53050 6905 53170 7025
rect 53225 6905 53345 7025
rect 47865 6740 47985 6860
rect 48030 6740 48150 6860
rect 48195 6740 48315 6860
rect 48360 6740 48480 6860
rect 48535 6740 48655 6860
rect 48700 6740 48820 6860
rect 48865 6740 48985 6860
rect 49030 6740 49150 6860
rect 49205 6740 49325 6860
rect 49370 6740 49490 6860
rect 49535 6740 49655 6860
rect 49700 6740 49820 6860
rect 49875 6740 49995 6860
rect 50040 6740 50160 6860
rect 50205 6740 50325 6860
rect 50370 6740 50490 6860
rect 50545 6740 50665 6860
rect 50710 6740 50830 6860
rect 50875 6740 50995 6860
rect 51040 6740 51160 6860
rect 51215 6740 51335 6860
rect 51380 6740 51500 6860
rect 51545 6740 51665 6860
rect 51710 6740 51830 6860
rect 51885 6740 52005 6860
rect 52050 6740 52170 6860
rect 52215 6740 52335 6860
rect 52380 6740 52500 6860
rect 52555 6740 52675 6860
rect 52720 6740 52840 6860
rect 52885 6740 53005 6860
rect 53050 6740 53170 6860
rect 53225 6740 53345 6860
rect 47865 6575 47985 6695
rect 48030 6575 48150 6695
rect 48195 6575 48315 6695
rect 48360 6575 48480 6695
rect 48535 6575 48655 6695
rect 48700 6575 48820 6695
rect 48865 6575 48985 6695
rect 49030 6575 49150 6695
rect 49205 6575 49325 6695
rect 49370 6575 49490 6695
rect 49535 6575 49655 6695
rect 49700 6575 49820 6695
rect 49875 6575 49995 6695
rect 50040 6575 50160 6695
rect 50205 6575 50325 6695
rect 50370 6575 50490 6695
rect 50545 6575 50665 6695
rect 50710 6575 50830 6695
rect 50875 6575 50995 6695
rect 51040 6575 51160 6695
rect 51215 6575 51335 6695
rect 51380 6575 51500 6695
rect 51545 6575 51665 6695
rect 51710 6575 51830 6695
rect 51885 6575 52005 6695
rect 52050 6575 52170 6695
rect 52215 6575 52335 6695
rect 52380 6575 52500 6695
rect 52555 6575 52675 6695
rect 52720 6575 52840 6695
rect 52885 6575 53005 6695
rect 53050 6575 53170 6695
rect 53225 6575 53345 6695
rect 47865 6410 47985 6530
rect 48030 6410 48150 6530
rect 48195 6410 48315 6530
rect 48360 6410 48480 6530
rect 48535 6410 48655 6530
rect 48700 6410 48820 6530
rect 48865 6410 48985 6530
rect 49030 6410 49150 6530
rect 49205 6410 49325 6530
rect 49370 6410 49490 6530
rect 49535 6410 49655 6530
rect 49700 6410 49820 6530
rect 49875 6410 49995 6530
rect 50040 6410 50160 6530
rect 50205 6410 50325 6530
rect 50370 6410 50490 6530
rect 50545 6410 50665 6530
rect 50710 6410 50830 6530
rect 50875 6410 50995 6530
rect 51040 6410 51160 6530
rect 51215 6410 51335 6530
rect 51380 6410 51500 6530
rect 51545 6410 51665 6530
rect 51710 6410 51830 6530
rect 51885 6410 52005 6530
rect 52050 6410 52170 6530
rect 52215 6410 52335 6530
rect 52380 6410 52500 6530
rect 52555 6410 52675 6530
rect 52720 6410 52840 6530
rect 52885 6410 53005 6530
rect 53050 6410 53170 6530
rect 53225 6410 53345 6530
rect 47865 6235 47985 6355
rect 48030 6235 48150 6355
rect 48195 6235 48315 6355
rect 48360 6235 48480 6355
rect 48535 6235 48655 6355
rect 48700 6235 48820 6355
rect 48865 6235 48985 6355
rect 49030 6235 49150 6355
rect 49205 6235 49325 6355
rect 49370 6235 49490 6355
rect 49535 6235 49655 6355
rect 49700 6235 49820 6355
rect 49875 6235 49995 6355
rect 50040 6235 50160 6355
rect 50205 6235 50325 6355
rect 50370 6235 50490 6355
rect 50545 6235 50665 6355
rect 50710 6235 50830 6355
rect 50875 6235 50995 6355
rect 51040 6235 51160 6355
rect 51215 6235 51335 6355
rect 51380 6235 51500 6355
rect 51545 6235 51665 6355
rect 51710 6235 51830 6355
rect 51885 6235 52005 6355
rect 52050 6235 52170 6355
rect 52215 6235 52335 6355
rect 52380 6235 52500 6355
rect 52555 6235 52675 6355
rect 52720 6235 52840 6355
rect 52885 6235 53005 6355
rect 53050 6235 53170 6355
rect 53225 6235 53345 6355
rect 47865 6070 47985 6190
rect 48030 6070 48150 6190
rect 48195 6070 48315 6190
rect 48360 6070 48480 6190
rect 48535 6070 48655 6190
rect 48700 6070 48820 6190
rect 48865 6070 48985 6190
rect 49030 6070 49150 6190
rect 49205 6070 49325 6190
rect 49370 6070 49490 6190
rect 49535 6070 49655 6190
rect 49700 6070 49820 6190
rect 49875 6070 49995 6190
rect 50040 6070 50160 6190
rect 50205 6070 50325 6190
rect 50370 6070 50490 6190
rect 50545 6070 50665 6190
rect 50710 6070 50830 6190
rect 50875 6070 50995 6190
rect 51040 6070 51160 6190
rect 51215 6070 51335 6190
rect 51380 6070 51500 6190
rect 51545 6070 51665 6190
rect 51710 6070 51830 6190
rect 51885 6070 52005 6190
rect 52050 6070 52170 6190
rect 52215 6070 52335 6190
rect 52380 6070 52500 6190
rect 52555 6070 52675 6190
rect 52720 6070 52840 6190
rect 52885 6070 53005 6190
rect 53050 6070 53170 6190
rect 53225 6070 53345 6190
rect 47865 5905 47985 6025
rect 48030 5905 48150 6025
rect 48195 5905 48315 6025
rect 48360 5905 48480 6025
rect 48535 5905 48655 6025
rect 48700 5905 48820 6025
rect 48865 5905 48985 6025
rect 49030 5905 49150 6025
rect 49205 5905 49325 6025
rect 49370 5905 49490 6025
rect 49535 5905 49655 6025
rect 49700 5905 49820 6025
rect 49875 5905 49995 6025
rect 50040 5905 50160 6025
rect 50205 5905 50325 6025
rect 50370 5905 50490 6025
rect 50545 5905 50665 6025
rect 50710 5905 50830 6025
rect 50875 5905 50995 6025
rect 51040 5905 51160 6025
rect 51215 5905 51335 6025
rect 51380 5905 51500 6025
rect 51545 5905 51665 6025
rect 51710 5905 51830 6025
rect 51885 5905 52005 6025
rect 52050 5905 52170 6025
rect 52215 5905 52335 6025
rect 52380 5905 52500 6025
rect 52555 5905 52675 6025
rect 52720 5905 52840 6025
rect 52885 5905 53005 6025
rect 53050 5905 53170 6025
rect 53225 5905 53345 6025
rect 47865 5740 47985 5860
rect 48030 5740 48150 5860
rect 48195 5740 48315 5860
rect 48360 5740 48480 5860
rect 48535 5740 48655 5860
rect 48700 5740 48820 5860
rect 48865 5740 48985 5860
rect 49030 5740 49150 5860
rect 49205 5740 49325 5860
rect 49370 5740 49490 5860
rect 49535 5740 49655 5860
rect 49700 5740 49820 5860
rect 49875 5740 49995 5860
rect 50040 5740 50160 5860
rect 50205 5740 50325 5860
rect 50370 5740 50490 5860
rect 50545 5740 50665 5860
rect 50710 5740 50830 5860
rect 50875 5740 50995 5860
rect 51040 5740 51160 5860
rect 51215 5740 51335 5860
rect 51380 5740 51500 5860
rect 51545 5740 51665 5860
rect 51710 5740 51830 5860
rect 51885 5740 52005 5860
rect 52050 5740 52170 5860
rect 52215 5740 52335 5860
rect 52380 5740 52500 5860
rect 52555 5740 52675 5860
rect 52720 5740 52840 5860
rect 52885 5740 53005 5860
rect 53050 5740 53170 5860
rect 53225 5740 53345 5860
rect 47865 5565 47985 5685
rect 48030 5565 48150 5685
rect 48195 5565 48315 5685
rect 48360 5565 48480 5685
rect 48535 5565 48655 5685
rect 48700 5565 48820 5685
rect 48865 5565 48985 5685
rect 49030 5565 49150 5685
rect 49205 5565 49325 5685
rect 49370 5565 49490 5685
rect 49535 5565 49655 5685
rect 49700 5565 49820 5685
rect 49875 5565 49995 5685
rect 50040 5565 50160 5685
rect 50205 5565 50325 5685
rect 50370 5565 50490 5685
rect 50545 5565 50665 5685
rect 50710 5565 50830 5685
rect 50875 5565 50995 5685
rect 51040 5565 51160 5685
rect 51215 5565 51335 5685
rect 51380 5565 51500 5685
rect 51545 5565 51665 5685
rect 51710 5565 51830 5685
rect 51885 5565 52005 5685
rect 52050 5565 52170 5685
rect 52215 5565 52335 5685
rect 52380 5565 52500 5685
rect 52555 5565 52675 5685
rect 52720 5565 52840 5685
rect 52885 5565 53005 5685
rect 53050 5565 53170 5685
rect 53225 5565 53345 5685
rect 47865 5400 47985 5520
rect 48030 5400 48150 5520
rect 48195 5400 48315 5520
rect 48360 5400 48480 5520
rect 48535 5400 48655 5520
rect 48700 5400 48820 5520
rect 48865 5400 48985 5520
rect 49030 5400 49150 5520
rect 49205 5400 49325 5520
rect 49370 5400 49490 5520
rect 49535 5400 49655 5520
rect 49700 5400 49820 5520
rect 49875 5400 49995 5520
rect 50040 5400 50160 5520
rect 50205 5400 50325 5520
rect 50370 5400 50490 5520
rect 50545 5400 50665 5520
rect 50710 5400 50830 5520
rect 50875 5400 50995 5520
rect 51040 5400 51160 5520
rect 51215 5400 51335 5520
rect 51380 5400 51500 5520
rect 51545 5400 51665 5520
rect 51710 5400 51830 5520
rect 51885 5400 52005 5520
rect 52050 5400 52170 5520
rect 52215 5400 52335 5520
rect 52380 5400 52500 5520
rect 52555 5400 52675 5520
rect 52720 5400 52840 5520
rect 52885 5400 53005 5520
rect 53050 5400 53170 5520
rect 53225 5400 53345 5520
rect 47865 5235 47985 5355
rect 48030 5235 48150 5355
rect 48195 5235 48315 5355
rect 48360 5235 48480 5355
rect 48535 5235 48655 5355
rect 48700 5235 48820 5355
rect 48865 5235 48985 5355
rect 49030 5235 49150 5355
rect 49205 5235 49325 5355
rect 49370 5235 49490 5355
rect 49535 5235 49655 5355
rect 49700 5235 49820 5355
rect 49875 5235 49995 5355
rect 50040 5235 50160 5355
rect 50205 5235 50325 5355
rect 50370 5235 50490 5355
rect 50545 5235 50665 5355
rect 50710 5235 50830 5355
rect 50875 5235 50995 5355
rect 51040 5235 51160 5355
rect 51215 5235 51335 5355
rect 51380 5235 51500 5355
rect 51545 5235 51665 5355
rect 51710 5235 51830 5355
rect 51885 5235 52005 5355
rect 52050 5235 52170 5355
rect 52215 5235 52335 5355
rect 52380 5235 52500 5355
rect 52555 5235 52675 5355
rect 52720 5235 52840 5355
rect 52885 5235 53005 5355
rect 53050 5235 53170 5355
rect 53225 5235 53345 5355
rect 47865 5070 47985 5190
rect 48030 5070 48150 5190
rect 48195 5070 48315 5190
rect 48360 5070 48480 5190
rect 48535 5070 48655 5190
rect 48700 5070 48820 5190
rect 48865 5070 48985 5190
rect 49030 5070 49150 5190
rect 49205 5070 49325 5190
rect 49370 5070 49490 5190
rect 49535 5070 49655 5190
rect 49700 5070 49820 5190
rect 49875 5070 49995 5190
rect 50040 5070 50160 5190
rect 50205 5070 50325 5190
rect 50370 5070 50490 5190
rect 50545 5070 50665 5190
rect 50710 5070 50830 5190
rect 50875 5070 50995 5190
rect 51040 5070 51160 5190
rect 51215 5070 51335 5190
rect 51380 5070 51500 5190
rect 51545 5070 51665 5190
rect 51710 5070 51830 5190
rect 51885 5070 52005 5190
rect 52050 5070 52170 5190
rect 52215 5070 52335 5190
rect 52380 5070 52500 5190
rect 52555 5070 52675 5190
rect 52720 5070 52840 5190
rect 52885 5070 53005 5190
rect 53050 5070 53170 5190
rect 53225 5070 53345 5190
rect 47865 4895 47985 5015
rect 48030 4895 48150 5015
rect 48195 4895 48315 5015
rect 48360 4895 48480 5015
rect 48535 4895 48655 5015
rect 48700 4895 48820 5015
rect 48865 4895 48985 5015
rect 49030 4895 49150 5015
rect 49205 4895 49325 5015
rect 49370 4895 49490 5015
rect 49535 4895 49655 5015
rect 49700 4895 49820 5015
rect 49875 4895 49995 5015
rect 50040 4895 50160 5015
rect 50205 4895 50325 5015
rect 50370 4895 50490 5015
rect 50545 4895 50665 5015
rect 50710 4895 50830 5015
rect 50875 4895 50995 5015
rect 51040 4895 51160 5015
rect 51215 4895 51335 5015
rect 51380 4895 51500 5015
rect 51545 4895 51665 5015
rect 51710 4895 51830 5015
rect 51885 4895 52005 5015
rect 52050 4895 52170 5015
rect 52215 4895 52335 5015
rect 52380 4895 52500 5015
rect 52555 4895 52675 5015
rect 52720 4895 52840 5015
rect 52885 4895 53005 5015
rect 53050 4895 53170 5015
rect 53225 4895 53345 5015
rect 47865 4730 47985 4850
rect 48030 4730 48150 4850
rect 48195 4730 48315 4850
rect 48360 4730 48480 4850
rect 48535 4730 48655 4850
rect 48700 4730 48820 4850
rect 48865 4730 48985 4850
rect 49030 4730 49150 4850
rect 49205 4730 49325 4850
rect 49370 4730 49490 4850
rect 49535 4730 49655 4850
rect 49700 4730 49820 4850
rect 49875 4730 49995 4850
rect 50040 4730 50160 4850
rect 50205 4730 50325 4850
rect 50370 4730 50490 4850
rect 50545 4730 50665 4850
rect 50710 4730 50830 4850
rect 50875 4730 50995 4850
rect 51040 4730 51160 4850
rect 51215 4730 51335 4850
rect 51380 4730 51500 4850
rect 51545 4730 51665 4850
rect 51710 4730 51830 4850
rect 51885 4730 52005 4850
rect 52050 4730 52170 4850
rect 52215 4730 52335 4850
rect 52380 4730 52500 4850
rect 52555 4730 52675 4850
rect 52720 4730 52840 4850
rect 52885 4730 53005 4850
rect 53050 4730 53170 4850
rect 53225 4730 53345 4850
rect 47865 4565 47985 4685
rect 48030 4565 48150 4685
rect 48195 4565 48315 4685
rect 48360 4565 48480 4685
rect 48535 4565 48655 4685
rect 48700 4565 48820 4685
rect 48865 4565 48985 4685
rect 49030 4565 49150 4685
rect 49205 4565 49325 4685
rect 49370 4565 49490 4685
rect 49535 4565 49655 4685
rect 49700 4565 49820 4685
rect 49875 4565 49995 4685
rect 50040 4565 50160 4685
rect 50205 4565 50325 4685
rect 50370 4565 50490 4685
rect 50545 4565 50665 4685
rect 50710 4565 50830 4685
rect 50875 4565 50995 4685
rect 51040 4565 51160 4685
rect 51215 4565 51335 4685
rect 51380 4565 51500 4685
rect 51545 4565 51665 4685
rect 51710 4565 51830 4685
rect 51885 4565 52005 4685
rect 52050 4565 52170 4685
rect 52215 4565 52335 4685
rect 52380 4565 52500 4685
rect 52555 4565 52675 4685
rect 52720 4565 52840 4685
rect 52885 4565 53005 4685
rect 53050 4565 53170 4685
rect 53225 4565 53345 4685
rect 47865 4400 47985 4520
rect 48030 4400 48150 4520
rect 48195 4400 48315 4520
rect 48360 4400 48480 4520
rect 48535 4400 48655 4520
rect 48700 4400 48820 4520
rect 48865 4400 48985 4520
rect 49030 4400 49150 4520
rect 49205 4400 49325 4520
rect 49370 4400 49490 4520
rect 49535 4400 49655 4520
rect 49700 4400 49820 4520
rect 49875 4400 49995 4520
rect 50040 4400 50160 4520
rect 50205 4400 50325 4520
rect 50370 4400 50490 4520
rect 50545 4400 50665 4520
rect 50710 4400 50830 4520
rect 50875 4400 50995 4520
rect 51040 4400 51160 4520
rect 51215 4400 51335 4520
rect 51380 4400 51500 4520
rect 51545 4400 51665 4520
rect 51710 4400 51830 4520
rect 51885 4400 52005 4520
rect 52050 4400 52170 4520
rect 52215 4400 52335 4520
rect 52380 4400 52500 4520
rect 52555 4400 52675 4520
rect 52720 4400 52840 4520
rect 52885 4400 53005 4520
rect 53050 4400 53170 4520
rect 53225 4400 53345 4520
rect 47865 4225 47985 4345
rect 48030 4225 48150 4345
rect 48195 4225 48315 4345
rect 48360 4225 48480 4345
rect 48535 4225 48655 4345
rect 48700 4225 48820 4345
rect 48865 4225 48985 4345
rect 49030 4225 49150 4345
rect 49205 4225 49325 4345
rect 49370 4225 49490 4345
rect 49535 4225 49655 4345
rect 49700 4225 49820 4345
rect 49875 4225 49995 4345
rect 50040 4225 50160 4345
rect 50205 4225 50325 4345
rect 50370 4225 50490 4345
rect 50545 4225 50665 4345
rect 50710 4225 50830 4345
rect 50875 4225 50995 4345
rect 51040 4225 51160 4345
rect 51215 4225 51335 4345
rect 51380 4225 51500 4345
rect 51545 4225 51665 4345
rect 51710 4225 51830 4345
rect 51885 4225 52005 4345
rect 52050 4225 52170 4345
rect 52215 4225 52335 4345
rect 52380 4225 52500 4345
rect 52555 4225 52675 4345
rect 52720 4225 52840 4345
rect 52885 4225 53005 4345
rect 53050 4225 53170 4345
rect 53225 4225 53345 4345
rect 47865 4060 47985 4180
rect 48030 4060 48150 4180
rect 48195 4060 48315 4180
rect 48360 4060 48480 4180
rect 48535 4060 48655 4180
rect 48700 4060 48820 4180
rect 48865 4060 48985 4180
rect 49030 4060 49150 4180
rect 49205 4060 49325 4180
rect 49370 4060 49490 4180
rect 49535 4060 49655 4180
rect 49700 4060 49820 4180
rect 49875 4060 49995 4180
rect 50040 4060 50160 4180
rect 50205 4060 50325 4180
rect 50370 4060 50490 4180
rect 50545 4060 50665 4180
rect 50710 4060 50830 4180
rect 50875 4060 50995 4180
rect 51040 4060 51160 4180
rect 51215 4060 51335 4180
rect 51380 4060 51500 4180
rect 51545 4060 51665 4180
rect 51710 4060 51830 4180
rect 51885 4060 52005 4180
rect 52050 4060 52170 4180
rect 52215 4060 52335 4180
rect 52380 4060 52500 4180
rect 52555 4060 52675 4180
rect 52720 4060 52840 4180
rect 52885 4060 53005 4180
rect 53050 4060 53170 4180
rect 53225 4060 53345 4180
rect 47865 3895 47985 4015
rect 48030 3895 48150 4015
rect 48195 3895 48315 4015
rect 48360 3895 48480 4015
rect 48535 3895 48655 4015
rect 48700 3895 48820 4015
rect 48865 3895 48985 4015
rect 49030 3895 49150 4015
rect 49205 3895 49325 4015
rect 49370 3895 49490 4015
rect 49535 3895 49655 4015
rect 49700 3895 49820 4015
rect 49875 3895 49995 4015
rect 50040 3895 50160 4015
rect 50205 3895 50325 4015
rect 50370 3895 50490 4015
rect 50545 3895 50665 4015
rect 50710 3895 50830 4015
rect 50875 3895 50995 4015
rect 51040 3895 51160 4015
rect 51215 3895 51335 4015
rect 51380 3895 51500 4015
rect 51545 3895 51665 4015
rect 51710 3895 51830 4015
rect 51885 3895 52005 4015
rect 52050 3895 52170 4015
rect 52215 3895 52335 4015
rect 52380 3895 52500 4015
rect 52555 3895 52675 4015
rect 52720 3895 52840 4015
rect 52885 3895 53005 4015
rect 53050 3895 53170 4015
rect 53225 3895 53345 4015
rect 47865 3730 47985 3850
rect 48030 3730 48150 3850
rect 48195 3730 48315 3850
rect 48360 3730 48480 3850
rect 48535 3730 48655 3850
rect 48700 3730 48820 3850
rect 48865 3730 48985 3850
rect 49030 3730 49150 3850
rect 49205 3730 49325 3850
rect 49370 3730 49490 3850
rect 49535 3730 49655 3850
rect 49700 3730 49820 3850
rect 49875 3730 49995 3850
rect 50040 3730 50160 3850
rect 50205 3730 50325 3850
rect 50370 3730 50490 3850
rect 50545 3730 50665 3850
rect 50710 3730 50830 3850
rect 50875 3730 50995 3850
rect 51040 3730 51160 3850
rect 51215 3730 51335 3850
rect 51380 3730 51500 3850
rect 51545 3730 51665 3850
rect 51710 3730 51830 3850
rect 51885 3730 52005 3850
rect 52050 3730 52170 3850
rect 52215 3730 52335 3850
rect 52380 3730 52500 3850
rect 52555 3730 52675 3850
rect 52720 3730 52840 3850
rect 52885 3730 53005 3850
rect 53050 3730 53170 3850
rect 53225 3730 53345 3850
rect 47865 3555 47985 3675
rect 48030 3555 48150 3675
rect 48195 3555 48315 3675
rect 48360 3555 48480 3675
rect 48535 3555 48655 3675
rect 48700 3555 48820 3675
rect 48865 3555 48985 3675
rect 49030 3555 49150 3675
rect 49205 3555 49325 3675
rect 49370 3555 49490 3675
rect 49535 3555 49655 3675
rect 49700 3555 49820 3675
rect 49875 3555 49995 3675
rect 50040 3555 50160 3675
rect 50205 3555 50325 3675
rect 50370 3555 50490 3675
rect 50545 3555 50665 3675
rect 50710 3555 50830 3675
rect 50875 3555 50995 3675
rect 51040 3555 51160 3675
rect 51215 3555 51335 3675
rect 51380 3555 51500 3675
rect 51545 3555 51665 3675
rect 51710 3555 51830 3675
rect 51885 3555 52005 3675
rect 52050 3555 52170 3675
rect 52215 3555 52335 3675
rect 52380 3555 52500 3675
rect 52555 3555 52675 3675
rect 52720 3555 52840 3675
rect 52885 3555 53005 3675
rect 53050 3555 53170 3675
rect 53225 3555 53345 3675
rect 47865 3390 47985 3510
rect 48030 3390 48150 3510
rect 48195 3390 48315 3510
rect 48360 3390 48480 3510
rect 48535 3390 48655 3510
rect 48700 3390 48820 3510
rect 48865 3390 48985 3510
rect 49030 3390 49150 3510
rect 49205 3390 49325 3510
rect 49370 3390 49490 3510
rect 49535 3390 49655 3510
rect 49700 3390 49820 3510
rect 49875 3390 49995 3510
rect 50040 3390 50160 3510
rect 50205 3390 50325 3510
rect 50370 3390 50490 3510
rect 50545 3390 50665 3510
rect 50710 3390 50830 3510
rect 50875 3390 50995 3510
rect 51040 3390 51160 3510
rect 51215 3390 51335 3510
rect 51380 3390 51500 3510
rect 51545 3390 51665 3510
rect 51710 3390 51830 3510
rect 51885 3390 52005 3510
rect 52050 3390 52170 3510
rect 52215 3390 52335 3510
rect 52380 3390 52500 3510
rect 52555 3390 52675 3510
rect 52720 3390 52840 3510
rect 52885 3390 53005 3510
rect 53050 3390 53170 3510
rect 53225 3390 53345 3510
rect 47865 3225 47985 3345
rect 48030 3225 48150 3345
rect 48195 3225 48315 3345
rect 48360 3225 48480 3345
rect 48535 3225 48655 3345
rect 48700 3225 48820 3345
rect 48865 3225 48985 3345
rect 49030 3225 49150 3345
rect 49205 3225 49325 3345
rect 49370 3225 49490 3345
rect 49535 3225 49655 3345
rect 49700 3225 49820 3345
rect 49875 3225 49995 3345
rect 50040 3225 50160 3345
rect 50205 3225 50325 3345
rect 50370 3225 50490 3345
rect 50545 3225 50665 3345
rect 50710 3225 50830 3345
rect 50875 3225 50995 3345
rect 51040 3225 51160 3345
rect 51215 3225 51335 3345
rect 51380 3225 51500 3345
rect 51545 3225 51665 3345
rect 51710 3225 51830 3345
rect 51885 3225 52005 3345
rect 52050 3225 52170 3345
rect 52215 3225 52335 3345
rect 52380 3225 52500 3345
rect 52555 3225 52675 3345
rect 52720 3225 52840 3345
rect 52885 3225 53005 3345
rect 53050 3225 53170 3345
rect 53225 3225 53345 3345
rect 47865 3060 47985 3180
rect 48030 3060 48150 3180
rect 48195 3060 48315 3180
rect 48360 3060 48480 3180
rect 48535 3060 48655 3180
rect 48700 3060 48820 3180
rect 48865 3060 48985 3180
rect 49030 3060 49150 3180
rect 49205 3060 49325 3180
rect 49370 3060 49490 3180
rect 49535 3060 49655 3180
rect 49700 3060 49820 3180
rect 49875 3060 49995 3180
rect 50040 3060 50160 3180
rect 50205 3060 50325 3180
rect 50370 3060 50490 3180
rect 50545 3060 50665 3180
rect 50710 3060 50830 3180
rect 50875 3060 50995 3180
rect 51040 3060 51160 3180
rect 51215 3060 51335 3180
rect 51380 3060 51500 3180
rect 51545 3060 51665 3180
rect 51710 3060 51830 3180
rect 51885 3060 52005 3180
rect 52050 3060 52170 3180
rect 52215 3060 52335 3180
rect 52380 3060 52500 3180
rect 52555 3060 52675 3180
rect 52720 3060 52840 3180
rect 52885 3060 53005 3180
rect 53050 3060 53170 3180
rect 53225 3060 53345 3180
rect 47865 2885 47985 3005
rect 48030 2885 48150 3005
rect 48195 2885 48315 3005
rect 48360 2885 48480 3005
rect 48535 2885 48655 3005
rect 48700 2885 48820 3005
rect 48865 2885 48985 3005
rect 49030 2885 49150 3005
rect 49205 2885 49325 3005
rect 49370 2885 49490 3005
rect 49535 2885 49655 3005
rect 49700 2885 49820 3005
rect 49875 2885 49995 3005
rect 50040 2885 50160 3005
rect 50205 2885 50325 3005
rect 50370 2885 50490 3005
rect 50545 2885 50665 3005
rect 50710 2885 50830 3005
rect 50875 2885 50995 3005
rect 51040 2885 51160 3005
rect 51215 2885 51335 3005
rect 51380 2885 51500 3005
rect 51545 2885 51665 3005
rect 51710 2885 51830 3005
rect 51885 2885 52005 3005
rect 52050 2885 52170 3005
rect 52215 2885 52335 3005
rect 52380 2885 52500 3005
rect 52555 2885 52675 3005
rect 52720 2885 52840 3005
rect 52885 2885 53005 3005
rect 53050 2885 53170 3005
rect 53225 2885 53345 3005
rect 47865 2720 47985 2840
rect 48030 2720 48150 2840
rect 48195 2720 48315 2840
rect 48360 2720 48480 2840
rect 48535 2720 48655 2840
rect 48700 2720 48820 2840
rect 48865 2720 48985 2840
rect 49030 2720 49150 2840
rect 49205 2720 49325 2840
rect 49370 2720 49490 2840
rect 49535 2720 49655 2840
rect 49700 2720 49820 2840
rect 49875 2720 49995 2840
rect 50040 2720 50160 2840
rect 50205 2720 50325 2840
rect 50370 2720 50490 2840
rect 50545 2720 50665 2840
rect 50710 2720 50830 2840
rect 50875 2720 50995 2840
rect 51040 2720 51160 2840
rect 51215 2720 51335 2840
rect 51380 2720 51500 2840
rect 51545 2720 51665 2840
rect 51710 2720 51830 2840
rect 51885 2720 52005 2840
rect 52050 2720 52170 2840
rect 52215 2720 52335 2840
rect 52380 2720 52500 2840
rect 52555 2720 52675 2840
rect 52720 2720 52840 2840
rect 52885 2720 53005 2840
rect 53050 2720 53170 2840
rect 53225 2720 53345 2840
rect 47865 2555 47985 2675
rect 48030 2555 48150 2675
rect 48195 2555 48315 2675
rect 48360 2555 48480 2675
rect 48535 2555 48655 2675
rect 48700 2555 48820 2675
rect 48865 2555 48985 2675
rect 49030 2555 49150 2675
rect 49205 2555 49325 2675
rect 49370 2555 49490 2675
rect 49535 2555 49655 2675
rect 49700 2555 49820 2675
rect 49875 2555 49995 2675
rect 50040 2555 50160 2675
rect 50205 2555 50325 2675
rect 50370 2555 50490 2675
rect 50545 2555 50665 2675
rect 50710 2555 50830 2675
rect 50875 2555 50995 2675
rect 51040 2555 51160 2675
rect 51215 2555 51335 2675
rect 51380 2555 51500 2675
rect 51545 2555 51665 2675
rect 51710 2555 51830 2675
rect 51885 2555 52005 2675
rect 52050 2555 52170 2675
rect 52215 2555 52335 2675
rect 52380 2555 52500 2675
rect 52555 2555 52675 2675
rect 52720 2555 52840 2675
rect 52885 2555 53005 2675
rect 53050 2555 53170 2675
rect 53225 2555 53345 2675
rect 47865 2390 47985 2510
rect 48030 2390 48150 2510
rect 48195 2390 48315 2510
rect 48360 2390 48480 2510
rect 48535 2390 48655 2510
rect 48700 2390 48820 2510
rect 48865 2390 48985 2510
rect 49030 2390 49150 2510
rect 49205 2390 49325 2510
rect 49370 2390 49490 2510
rect 49535 2390 49655 2510
rect 49700 2390 49820 2510
rect 49875 2390 49995 2510
rect 50040 2390 50160 2510
rect 50205 2390 50325 2510
rect 50370 2390 50490 2510
rect 50545 2390 50665 2510
rect 50710 2390 50830 2510
rect 50875 2390 50995 2510
rect 51040 2390 51160 2510
rect 51215 2390 51335 2510
rect 51380 2390 51500 2510
rect 51545 2390 51665 2510
rect 51710 2390 51830 2510
rect 51885 2390 52005 2510
rect 52050 2390 52170 2510
rect 52215 2390 52335 2510
rect 52380 2390 52500 2510
rect 52555 2390 52675 2510
rect 52720 2390 52840 2510
rect 52885 2390 53005 2510
rect 53050 2390 53170 2510
rect 53225 2390 53345 2510
rect 47865 2215 47985 2335
rect 48030 2215 48150 2335
rect 48195 2215 48315 2335
rect 48360 2215 48480 2335
rect 48535 2215 48655 2335
rect 48700 2215 48820 2335
rect 48865 2215 48985 2335
rect 49030 2215 49150 2335
rect 49205 2215 49325 2335
rect 49370 2215 49490 2335
rect 49535 2215 49655 2335
rect 49700 2215 49820 2335
rect 49875 2215 49995 2335
rect 50040 2215 50160 2335
rect 50205 2215 50325 2335
rect 50370 2215 50490 2335
rect 50545 2215 50665 2335
rect 50710 2215 50830 2335
rect 50875 2215 50995 2335
rect 51040 2215 51160 2335
rect 51215 2215 51335 2335
rect 51380 2215 51500 2335
rect 51545 2215 51665 2335
rect 51710 2215 51830 2335
rect 51885 2215 52005 2335
rect 52050 2215 52170 2335
rect 52215 2215 52335 2335
rect 52380 2215 52500 2335
rect 52555 2215 52675 2335
rect 52720 2215 52840 2335
rect 52885 2215 53005 2335
rect 53050 2215 53170 2335
rect 53225 2215 53345 2335
rect 47865 2050 47985 2170
rect 48030 2050 48150 2170
rect 48195 2050 48315 2170
rect 48360 2050 48480 2170
rect 48535 2050 48655 2170
rect 48700 2050 48820 2170
rect 48865 2050 48985 2170
rect 49030 2050 49150 2170
rect 49205 2050 49325 2170
rect 49370 2050 49490 2170
rect 49535 2050 49655 2170
rect 49700 2050 49820 2170
rect 49875 2050 49995 2170
rect 50040 2050 50160 2170
rect 50205 2050 50325 2170
rect 50370 2050 50490 2170
rect 50545 2050 50665 2170
rect 50710 2050 50830 2170
rect 50875 2050 50995 2170
rect 51040 2050 51160 2170
rect 51215 2050 51335 2170
rect 51380 2050 51500 2170
rect 51545 2050 51665 2170
rect 51710 2050 51830 2170
rect 51885 2050 52005 2170
rect 52050 2050 52170 2170
rect 52215 2050 52335 2170
rect 52380 2050 52500 2170
rect 52555 2050 52675 2170
rect 52720 2050 52840 2170
rect 52885 2050 53005 2170
rect 53050 2050 53170 2170
rect 53225 2050 53345 2170
rect 47865 1885 47985 2005
rect 48030 1885 48150 2005
rect 48195 1885 48315 2005
rect 48360 1885 48480 2005
rect 48535 1885 48655 2005
rect 48700 1885 48820 2005
rect 48865 1885 48985 2005
rect 49030 1885 49150 2005
rect 49205 1885 49325 2005
rect 49370 1885 49490 2005
rect 49535 1885 49655 2005
rect 49700 1885 49820 2005
rect 49875 1885 49995 2005
rect 50040 1885 50160 2005
rect 50205 1885 50325 2005
rect 50370 1885 50490 2005
rect 50545 1885 50665 2005
rect 50710 1885 50830 2005
rect 50875 1885 50995 2005
rect 51040 1885 51160 2005
rect 51215 1885 51335 2005
rect 51380 1885 51500 2005
rect 51545 1885 51665 2005
rect 51710 1885 51830 2005
rect 51885 1885 52005 2005
rect 52050 1885 52170 2005
rect 52215 1885 52335 2005
rect 52380 1885 52500 2005
rect 52555 1885 52675 2005
rect 52720 1885 52840 2005
rect 52885 1885 53005 2005
rect 53050 1885 53170 2005
rect 53225 1885 53345 2005
rect 47865 1720 47985 1840
rect 48030 1720 48150 1840
rect 48195 1720 48315 1840
rect 48360 1720 48480 1840
rect 48535 1720 48655 1840
rect 48700 1720 48820 1840
rect 48865 1720 48985 1840
rect 49030 1720 49150 1840
rect 49205 1720 49325 1840
rect 49370 1720 49490 1840
rect 49535 1720 49655 1840
rect 49700 1720 49820 1840
rect 49875 1720 49995 1840
rect 50040 1720 50160 1840
rect 50205 1720 50325 1840
rect 50370 1720 50490 1840
rect 50545 1720 50665 1840
rect 50710 1720 50830 1840
rect 50875 1720 50995 1840
rect 51040 1720 51160 1840
rect 51215 1720 51335 1840
rect 51380 1720 51500 1840
rect 51545 1720 51665 1840
rect 51710 1720 51830 1840
rect 51885 1720 52005 1840
rect 52050 1720 52170 1840
rect 52215 1720 52335 1840
rect 52380 1720 52500 1840
rect 52555 1720 52675 1840
rect 52720 1720 52840 1840
rect 52885 1720 53005 1840
rect 53050 1720 53170 1840
rect 53225 1720 53345 1840
rect 30795 1300 30915 1420
rect 30970 1300 31090 1420
rect 31135 1300 31255 1420
rect 31300 1300 31420 1420
rect 31465 1300 31585 1420
rect 31640 1300 31760 1420
rect 31805 1300 31925 1420
rect 31970 1300 32090 1420
rect 32135 1300 32255 1420
rect 32310 1300 32430 1420
rect 32475 1300 32595 1420
rect 32640 1300 32760 1420
rect 32805 1300 32925 1420
rect 32980 1300 33100 1420
rect 33145 1300 33265 1420
rect 33310 1300 33430 1420
rect 33475 1300 33595 1420
rect 33650 1300 33770 1420
rect 33815 1300 33935 1420
rect 33980 1300 34100 1420
rect 34145 1300 34265 1420
rect 34320 1300 34440 1420
rect 34485 1300 34605 1420
rect 34650 1300 34770 1420
rect 34815 1300 34935 1420
rect 34990 1300 35110 1420
rect 35155 1300 35275 1420
rect 35320 1300 35440 1420
rect 35485 1300 35605 1420
rect 35660 1300 35780 1420
rect 35825 1300 35945 1420
rect 35990 1300 36110 1420
rect 36155 1300 36275 1420
rect 30795 1135 30915 1255
rect 30970 1135 31090 1255
rect 31135 1135 31255 1255
rect 31300 1135 31420 1255
rect 31465 1135 31585 1255
rect 31640 1135 31760 1255
rect 31805 1135 31925 1255
rect 31970 1135 32090 1255
rect 32135 1135 32255 1255
rect 32310 1135 32430 1255
rect 32475 1135 32595 1255
rect 32640 1135 32760 1255
rect 32805 1135 32925 1255
rect 32980 1135 33100 1255
rect 33145 1135 33265 1255
rect 33310 1135 33430 1255
rect 33475 1135 33595 1255
rect 33650 1135 33770 1255
rect 33815 1135 33935 1255
rect 33980 1135 34100 1255
rect 34145 1135 34265 1255
rect 34320 1135 34440 1255
rect 34485 1135 34605 1255
rect 34650 1135 34770 1255
rect 34815 1135 34935 1255
rect 34990 1135 35110 1255
rect 35155 1135 35275 1255
rect 35320 1135 35440 1255
rect 35485 1135 35605 1255
rect 35660 1135 35780 1255
rect 35825 1135 35945 1255
rect 35990 1135 36110 1255
rect 36155 1135 36275 1255
rect 30795 970 30915 1090
rect 30970 970 31090 1090
rect 31135 970 31255 1090
rect 31300 970 31420 1090
rect 31465 970 31585 1090
rect 31640 970 31760 1090
rect 31805 970 31925 1090
rect 31970 970 32090 1090
rect 32135 970 32255 1090
rect 32310 970 32430 1090
rect 32475 970 32595 1090
rect 32640 970 32760 1090
rect 32805 970 32925 1090
rect 32980 970 33100 1090
rect 33145 970 33265 1090
rect 33310 970 33430 1090
rect 33475 970 33595 1090
rect 33650 970 33770 1090
rect 33815 970 33935 1090
rect 33980 970 34100 1090
rect 34145 970 34265 1090
rect 34320 970 34440 1090
rect 34485 970 34605 1090
rect 34650 970 34770 1090
rect 34815 970 34935 1090
rect 34990 970 35110 1090
rect 35155 970 35275 1090
rect 35320 970 35440 1090
rect 35485 970 35605 1090
rect 35660 970 35780 1090
rect 35825 970 35945 1090
rect 35990 970 36110 1090
rect 36155 970 36275 1090
rect 30795 805 30915 925
rect 30970 805 31090 925
rect 31135 805 31255 925
rect 31300 805 31420 925
rect 31465 805 31585 925
rect 31640 805 31760 925
rect 31805 805 31925 925
rect 31970 805 32090 925
rect 32135 805 32255 925
rect 32310 805 32430 925
rect 32475 805 32595 925
rect 32640 805 32760 925
rect 32805 805 32925 925
rect 32980 805 33100 925
rect 33145 805 33265 925
rect 33310 805 33430 925
rect 33475 805 33595 925
rect 33650 805 33770 925
rect 33815 805 33935 925
rect 33980 805 34100 925
rect 34145 805 34265 925
rect 34320 805 34440 925
rect 34485 805 34605 925
rect 34650 805 34770 925
rect 34815 805 34935 925
rect 34990 805 35110 925
rect 35155 805 35275 925
rect 35320 805 35440 925
rect 35485 805 35605 925
rect 35660 805 35780 925
rect 35825 805 35945 925
rect 35990 805 36110 925
rect 36155 805 36275 925
rect 30795 630 30915 750
rect 30970 630 31090 750
rect 31135 630 31255 750
rect 31300 630 31420 750
rect 31465 630 31585 750
rect 31640 630 31760 750
rect 31805 630 31925 750
rect 31970 630 32090 750
rect 32135 630 32255 750
rect 32310 630 32430 750
rect 32475 630 32595 750
rect 32640 630 32760 750
rect 32805 630 32925 750
rect 32980 630 33100 750
rect 33145 630 33265 750
rect 33310 630 33430 750
rect 33475 630 33595 750
rect 33650 630 33770 750
rect 33815 630 33935 750
rect 33980 630 34100 750
rect 34145 630 34265 750
rect 34320 630 34440 750
rect 34485 630 34605 750
rect 34650 630 34770 750
rect 34815 630 34935 750
rect 34990 630 35110 750
rect 35155 630 35275 750
rect 35320 630 35440 750
rect 35485 630 35605 750
rect 35660 630 35780 750
rect 35825 630 35945 750
rect 35990 630 36110 750
rect 36155 630 36275 750
rect 30795 465 30915 585
rect 30970 465 31090 585
rect 31135 465 31255 585
rect 31300 465 31420 585
rect 31465 465 31585 585
rect 31640 465 31760 585
rect 31805 465 31925 585
rect 31970 465 32090 585
rect 32135 465 32255 585
rect 32310 465 32430 585
rect 32475 465 32595 585
rect 32640 465 32760 585
rect 32805 465 32925 585
rect 32980 465 33100 585
rect 33145 465 33265 585
rect 33310 465 33430 585
rect 33475 465 33595 585
rect 33650 465 33770 585
rect 33815 465 33935 585
rect 33980 465 34100 585
rect 34145 465 34265 585
rect 34320 465 34440 585
rect 34485 465 34605 585
rect 34650 465 34770 585
rect 34815 465 34935 585
rect 34990 465 35110 585
rect 35155 465 35275 585
rect 35320 465 35440 585
rect 35485 465 35605 585
rect 35660 465 35780 585
rect 35825 465 35945 585
rect 35990 465 36110 585
rect 36155 465 36275 585
rect 30795 300 30915 420
rect 30970 300 31090 420
rect 31135 300 31255 420
rect 31300 300 31420 420
rect 31465 300 31585 420
rect 31640 300 31760 420
rect 31805 300 31925 420
rect 31970 300 32090 420
rect 32135 300 32255 420
rect 32310 300 32430 420
rect 32475 300 32595 420
rect 32640 300 32760 420
rect 32805 300 32925 420
rect 32980 300 33100 420
rect 33145 300 33265 420
rect 33310 300 33430 420
rect 33475 300 33595 420
rect 33650 300 33770 420
rect 33815 300 33935 420
rect 33980 300 34100 420
rect 34145 300 34265 420
rect 34320 300 34440 420
rect 34485 300 34605 420
rect 34650 300 34770 420
rect 34815 300 34935 420
rect 34990 300 35110 420
rect 35155 300 35275 420
rect 35320 300 35440 420
rect 35485 300 35605 420
rect 35660 300 35780 420
rect 35825 300 35945 420
rect 35990 300 36110 420
rect 36155 300 36275 420
rect 30795 135 30915 255
rect 30970 135 31090 255
rect 31135 135 31255 255
rect 31300 135 31420 255
rect 31465 135 31585 255
rect 31640 135 31760 255
rect 31805 135 31925 255
rect 31970 135 32090 255
rect 32135 135 32255 255
rect 32310 135 32430 255
rect 32475 135 32595 255
rect 32640 135 32760 255
rect 32805 135 32925 255
rect 32980 135 33100 255
rect 33145 135 33265 255
rect 33310 135 33430 255
rect 33475 135 33595 255
rect 33650 135 33770 255
rect 33815 135 33935 255
rect 33980 135 34100 255
rect 34145 135 34265 255
rect 34320 135 34440 255
rect 34485 135 34605 255
rect 34650 135 34770 255
rect 34815 135 34935 255
rect 34990 135 35110 255
rect 35155 135 35275 255
rect 35320 135 35440 255
rect 35485 135 35605 255
rect 35660 135 35780 255
rect 35825 135 35945 255
rect 35990 135 36110 255
rect 36155 135 36275 255
rect 30795 -40 30915 80
rect 30970 -40 31090 80
rect 31135 -40 31255 80
rect 31300 -40 31420 80
rect 31465 -40 31585 80
rect 31640 -40 31760 80
rect 31805 -40 31925 80
rect 31970 -40 32090 80
rect 32135 -40 32255 80
rect 32310 -40 32430 80
rect 32475 -40 32595 80
rect 32640 -40 32760 80
rect 32805 -40 32925 80
rect 32980 -40 33100 80
rect 33145 -40 33265 80
rect 33310 -40 33430 80
rect 33475 -40 33595 80
rect 33650 -40 33770 80
rect 33815 -40 33935 80
rect 33980 -40 34100 80
rect 34145 -40 34265 80
rect 34320 -40 34440 80
rect 34485 -40 34605 80
rect 34650 -40 34770 80
rect 34815 -40 34935 80
rect 34990 -40 35110 80
rect 35155 -40 35275 80
rect 35320 -40 35440 80
rect 35485 -40 35605 80
rect 35660 -40 35780 80
rect 35825 -40 35945 80
rect 35990 -40 36110 80
rect 36155 -40 36275 80
rect 30795 -205 30915 -85
rect 30970 -205 31090 -85
rect 31135 -205 31255 -85
rect 31300 -205 31420 -85
rect 31465 -205 31585 -85
rect 31640 -205 31760 -85
rect 31805 -205 31925 -85
rect 31970 -205 32090 -85
rect 32135 -205 32255 -85
rect 32310 -205 32430 -85
rect 32475 -205 32595 -85
rect 32640 -205 32760 -85
rect 32805 -205 32925 -85
rect 32980 -205 33100 -85
rect 33145 -205 33265 -85
rect 33310 -205 33430 -85
rect 33475 -205 33595 -85
rect 33650 -205 33770 -85
rect 33815 -205 33935 -85
rect 33980 -205 34100 -85
rect 34145 -205 34265 -85
rect 34320 -205 34440 -85
rect 34485 -205 34605 -85
rect 34650 -205 34770 -85
rect 34815 -205 34935 -85
rect 34990 -205 35110 -85
rect 35155 -205 35275 -85
rect 35320 -205 35440 -85
rect 35485 -205 35605 -85
rect 35660 -205 35780 -85
rect 35825 -205 35945 -85
rect 35990 -205 36110 -85
rect 36155 -205 36275 -85
rect 30795 -370 30915 -250
rect 30970 -370 31090 -250
rect 31135 -370 31255 -250
rect 31300 -370 31420 -250
rect 31465 -370 31585 -250
rect 31640 -370 31760 -250
rect 31805 -370 31925 -250
rect 31970 -370 32090 -250
rect 32135 -370 32255 -250
rect 32310 -370 32430 -250
rect 32475 -370 32595 -250
rect 32640 -370 32760 -250
rect 32805 -370 32925 -250
rect 32980 -370 33100 -250
rect 33145 -370 33265 -250
rect 33310 -370 33430 -250
rect 33475 -370 33595 -250
rect 33650 -370 33770 -250
rect 33815 -370 33935 -250
rect 33980 -370 34100 -250
rect 34145 -370 34265 -250
rect 34320 -370 34440 -250
rect 34485 -370 34605 -250
rect 34650 -370 34770 -250
rect 34815 -370 34935 -250
rect 34990 -370 35110 -250
rect 35155 -370 35275 -250
rect 35320 -370 35440 -250
rect 35485 -370 35605 -250
rect 35660 -370 35780 -250
rect 35825 -370 35945 -250
rect 35990 -370 36110 -250
rect 36155 -370 36275 -250
rect 30795 -535 30915 -415
rect 30970 -535 31090 -415
rect 31135 -535 31255 -415
rect 31300 -535 31420 -415
rect 31465 -535 31585 -415
rect 31640 -535 31760 -415
rect 31805 -535 31925 -415
rect 31970 -535 32090 -415
rect 32135 -535 32255 -415
rect 32310 -535 32430 -415
rect 32475 -535 32595 -415
rect 32640 -535 32760 -415
rect 32805 -535 32925 -415
rect 32980 -535 33100 -415
rect 33145 -535 33265 -415
rect 33310 -535 33430 -415
rect 33475 -535 33595 -415
rect 33650 -535 33770 -415
rect 33815 -535 33935 -415
rect 33980 -535 34100 -415
rect 34145 -535 34265 -415
rect 34320 -535 34440 -415
rect 34485 -535 34605 -415
rect 34650 -535 34770 -415
rect 34815 -535 34935 -415
rect 34990 -535 35110 -415
rect 35155 -535 35275 -415
rect 35320 -535 35440 -415
rect 35485 -535 35605 -415
rect 35660 -535 35780 -415
rect 35825 -535 35945 -415
rect 35990 -535 36110 -415
rect 36155 -535 36275 -415
rect 30795 -710 30915 -590
rect 30970 -710 31090 -590
rect 31135 -710 31255 -590
rect 31300 -710 31420 -590
rect 31465 -710 31585 -590
rect 31640 -710 31760 -590
rect 31805 -710 31925 -590
rect 31970 -710 32090 -590
rect 32135 -710 32255 -590
rect 32310 -710 32430 -590
rect 32475 -710 32595 -590
rect 32640 -710 32760 -590
rect 32805 -710 32925 -590
rect 32980 -710 33100 -590
rect 33145 -710 33265 -590
rect 33310 -710 33430 -590
rect 33475 -710 33595 -590
rect 33650 -710 33770 -590
rect 33815 -710 33935 -590
rect 33980 -710 34100 -590
rect 34145 -710 34265 -590
rect 34320 -710 34440 -590
rect 34485 -710 34605 -590
rect 34650 -710 34770 -590
rect 34815 -710 34935 -590
rect 34990 -710 35110 -590
rect 35155 -710 35275 -590
rect 35320 -710 35440 -590
rect 35485 -710 35605 -590
rect 35660 -710 35780 -590
rect 35825 -710 35945 -590
rect 35990 -710 36110 -590
rect 36155 -710 36275 -590
rect 30795 -875 30915 -755
rect 30970 -875 31090 -755
rect 31135 -875 31255 -755
rect 31300 -875 31420 -755
rect 31465 -875 31585 -755
rect 31640 -875 31760 -755
rect 31805 -875 31925 -755
rect 31970 -875 32090 -755
rect 32135 -875 32255 -755
rect 32310 -875 32430 -755
rect 32475 -875 32595 -755
rect 32640 -875 32760 -755
rect 32805 -875 32925 -755
rect 32980 -875 33100 -755
rect 33145 -875 33265 -755
rect 33310 -875 33430 -755
rect 33475 -875 33595 -755
rect 33650 -875 33770 -755
rect 33815 -875 33935 -755
rect 33980 -875 34100 -755
rect 34145 -875 34265 -755
rect 34320 -875 34440 -755
rect 34485 -875 34605 -755
rect 34650 -875 34770 -755
rect 34815 -875 34935 -755
rect 34990 -875 35110 -755
rect 35155 -875 35275 -755
rect 35320 -875 35440 -755
rect 35485 -875 35605 -755
rect 35660 -875 35780 -755
rect 35825 -875 35945 -755
rect 35990 -875 36110 -755
rect 36155 -875 36275 -755
rect 30795 -1040 30915 -920
rect 30970 -1040 31090 -920
rect 31135 -1040 31255 -920
rect 31300 -1040 31420 -920
rect 31465 -1040 31585 -920
rect 31640 -1040 31760 -920
rect 31805 -1040 31925 -920
rect 31970 -1040 32090 -920
rect 32135 -1040 32255 -920
rect 32310 -1040 32430 -920
rect 32475 -1040 32595 -920
rect 32640 -1040 32760 -920
rect 32805 -1040 32925 -920
rect 32980 -1040 33100 -920
rect 33145 -1040 33265 -920
rect 33310 -1040 33430 -920
rect 33475 -1040 33595 -920
rect 33650 -1040 33770 -920
rect 33815 -1040 33935 -920
rect 33980 -1040 34100 -920
rect 34145 -1040 34265 -920
rect 34320 -1040 34440 -920
rect 34485 -1040 34605 -920
rect 34650 -1040 34770 -920
rect 34815 -1040 34935 -920
rect 34990 -1040 35110 -920
rect 35155 -1040 35275 -920
rect 35320 -1040 35440 -920
rect 35485 -1040 35605 -920
rect 35660 -1040 35780 -920
rect 35825 -1040 35945 -920
rect 35990 -1040 36110 -920
rect 36155 -1040 36275 -920
rect 30795 -1205 30915 -1085
rect 30970 -1205 31090 -1085
rect 31135 -1205 31255 -1085
rect 31300 -1205 31420 -1085
rect 31465 -1205 31585 -1085
rect 31640 -1205 31760 -1085
rect 31805 -1205 31925 -1085
rect 31970 -1205 32090 -1085
rect 32135 -1205 32255 -1085
rect 32310 -1205 32430 -1085
rect 32475 -1205 32595 -1085
rect 32640 -1205 32760 -1085
rect 32805 -1205 32925 -1085
rect 32980 -1205 33100 -1085
rect 33145 -1205 33265 -1085
rect 33310 -1205 33430 -1085
rect 33475 -1205 33595 -1085
rect 33650 -1205 33770 -1085
rect 33815 -1205 33935 -1085
rect 33980 -1205 34100 -1085
rect 34145 -1205 34265 -1085
rect 34320 -1205 34440 -1085
rect 34485 -1205 34605 -1085
rect 34650 -1205 34770 -1085
rect 34815 -1205 34935 -1085
rect 34990 -1205 35110 -1085
rect 35155 -1205 35275 -1085
rect 35320 -1205 35440 -1085
rect 35485 -1205 35605 -1085
rect 35660 -1205 35780 -1085
rect 35825 -1205 35945 -1085
rect 35990 -1205 36110 -1085
rect 36155 -1205 36275 -1085
rect 30795 -1380 30915 -1260
rect 30970 -1380 31090 -1260
rect 31135 -1380 31255 -1260
rect 31300 -1380 31420 -1260
rect 31465 -1380 31585 -1260
rect 31640 -1380 31760 -1260
rect 31805 -1380 31925 -1260
rect 31970 -1380 32090 -1260
rect 32135 -1380 32255 -1260
rect 32310 -1380 32430 -1260
rect 32475 -1380 32595 -1260
rect 32640 -1380 32760 -1260
rect 32805 -1380 32925 -1260
rect 32980 -1380 33100 -1260
rect 33145 -1380 33265 -1260
rect 33310 -1380 33430 -1260
rect 33475 -1380 33595 -1260
rect 33650 -1380 33770 -1260
rect 33815 -1380 33935 -1260
rect 33980 -1380 34100 -1260
rect 34145 -1380 34265 -1260
rect 34320 -1380 34440 -1260
rect 34485 -1380 34605 -1260
rect 34650 -1380 34770 -1260
rect 34815 -1380 34935 -1260
rect 34990 -1380 35110 -1260
rect 35155 -1380 35275 -1260
rect 35320 -1380 35440 -1260
rect 35485 -1380 35605 -1260
rect 35660 -1380 35780 -1260
rect 35825 -1380 35945 -1260
rect 35990 -1380 36110 -1260
rect 36155 -1380 36275 -1260
rect 30795 -1545 30915 -1425
rect 30970 -1545 31090 -1425
rect 31135 -1545 31255 -1425
rect 31300 -1545 31420 -1425
rect 31465 -1545 31585 -1425
rect 31640 -1545 31760 -1425
rect 31805 -1545 31925 -1425
rect 31970 -1545 32090 -1425
rect 32135 -1545 32255 -1425
rect 32310 -1545 32430 -1425
rect 32475 -1545 32595 -1425
rect 32640 -1545 32760 -1425
rect 32805 -1545 32925 -1425
rect 32980 -1545 33100 -1425
rect 33145 -1545 33265 -1425
rect 33310 -1545 33430 -1425
rect 33475 -1545 33595 -1425
rect 33650 -1545 33770 -1425
rect 33815 -1545 33935 -1425
rect 33980 -1545 34100 -1425
rect 34145 -1545 34265 -1425
rect 34320 -1545 34440 -1425
rect 34485 -1545 34605 -1425
rect 34650 -1545 34770 -1425
rect 34815 -1545 34935 -1425
rect 34990 -1545 35110 -1425
rect 35155 -1545 35275 -1425
rect 35320 -1545 35440 -1425
rect 35485 -1545 35605 -1425
rect 35660 -1545 35780 -1425
rect 35825 -1545 35945 -1425
rect 35990 -1545 36110 -1425
rect 36155 -1545 36275 -1425
rect 30795 -1710 30915 -1590
rect 30970 -1710 31090 -1590
rect 31135 -1710 31255 -1590
rect 31300 -1710 31420 -1590
rect 31465 -1710 31585 -1590
rect 31640 -1710 31760 -1590
rect 31805 -1710 31925 -1590
rect 31970 -1710 32090 -1590
rect 32135 -1710 32255 -1590
rect 32310 -1710 32430 -1590
rect 32475 -1710 32595 -1590
rect 32640 -1710 32760 -1590
rect 32805 -1710 32925 -1590
rect 32980 -1710 33100 -1590
rect 33145 -1710 33265 -1590
rect 33310 -1710 33430 -1590
rect 33475 -1710 33595 -1590
rect 33650 -1710 33770 -1590
rect 33815 -1710 33935 -1590
rect 33980 -1710 34100 -1590
rect 34145 -1710 34265 -1590
rect 34320 -1710 34440 -1590
rect 34485 -1710 34605 -1590
rect 34650 -1710 34770 -1590
rect 34815 -1710 34935 -1590
rect 34990 -1710 35110 -1590
rect 35155 -1710 35275 -1590
rect 35320 -1710 35440 -1590
rect 35485 -1710 35605 -1590
rect 35660 -1710 35780 -1590
rect 35825 -1710 35945 -1590
rect 35990 -1710 36110 -1590
rect 36155 -1710 36275 -1590
rect 30795 -1875 30915 -1755
rect 30970 -1875 31090 -1755
rect 31135 -1875 31255 -1755
rect 31300 -1875 31420 -1755
rect 31465 -1875 31585 -1755
rect 31640 -1875 31760 -1755
rect 31805 -1875 31925 -1755
rect 31970 -1875 32090 -1755
rect 32135 -1875 32255 -1755
rect 32310 -1875 32430 -1755
rect 32475 -1875 32595 -1755
rect 32640 -1875 32760 -1755
rect 32805 -1875 32925 -1755
rect 32980 -1875 33100 -1755
rect 33145 -1875 33265 -1755
rect 33310 -1875 33430 -1755
rect 33475 -1875 33595 -1755
rect 33650 -1875 33770 -1755
rect 33815 -1875 33935 -1755
rect 33980 -1875 34100 -1755
rect 34145 -1875 34265 -1755
rect 34320 -1875 34440 -1755
rect 34485 -1875 34605 -1755
rect 34650 -1875 34770 -1755
rect 34815 -1875 34935 -1755
rect 34990 -1875 35110 -1755
rect 35155 -1875 35275 -1755
rect 35320 -1875 35440 -1755
rect 35485 -1875 35605 -1755
rect 35660 -1875 35780 -1755
rect 35825 -1875 35945 -1755
rect 35990 -1875 36110 -1755
rect 36155 -1875 36275 -1755
rect 30795 -2050 30915 -1930
rect 30970 -2050 31090 -1930
rect 31135 -2050 31255 -1930
rect 31300 -2050 31420 -1930
rect 31465 -2050 31585 -1930
rect 31640 -2050 31760 -1930
rect 31805 -2050 31925 -1930
rect 31970 -2050 32090 -1930
rect 32135 -2050 32255 -1930
rect 32310 -2050 32430 -1930
rect 32475 -2050 32595 -1930
rect 32640 -2050 32760 -1930
rect 32805 -2050 32925 -1930
rect 32980 -2050 33100 -1930
rect 33145 -2050 33265 -1930
rect 33310 -2050 33430 -1930
rect 33475 -2050 33595 -1930
rect 33650 -2050 33770 -1930
rect 33815 -2050 33935 -1930
rect 33980 -2050 34100 -1930
rect 34145 -2050 34265 -1930
rect 34320 -2050 34440 -1930
rect 34485 -2050 34605 -1930
rect 34650 -2050 34770 -1930
rect 34815 -2050 34935 -1930
rect 34990 -2050 35110 -1930
rect 35155 -2050 35275 -1930
rect 35320 -2050 35440 -1930
rect 35485 -2050 35605 -1930
rect 35660 -2050 35780 -1930
rect 35825 -2050 35945 -1930
rect 35990 -2050 36110 -1930
rect 36155 -2050 36275 -1930
rect 30795 -2215 30915 -2095
rect 30970 -2215 31090 -2095
rect 31135 -2215 31255 -2095
rect 31300 -2215 31420 -2095
rect 31465 -2215 31585 -2095
rect 31640 -2215 31760 -2095
rect 31805 -2215 31925 -2095
rect 31970 -2215 32090 -2095
rect 32135 -2215 32255 -2095
rect 32310 -2215 32430 -2095
rect 32475 -2215 32595 -2095
rect 32640 -2215 32760 -2095
rect 32805 -2215 32925 -2095
rect 32980 -2215 33100 -2095
rect 33145 -2215 33265 -2095
rect 33310 -2215 33430 -2095
rect 33475 -2215 33595 -2095
rect 33650 -2215 33770 -2095
rect 33815 -2215 33935 -2095
rect 33980 -2215 34100 -2095
rect 34145 -2215 34265 -2095
rect 34320 -2215 34440 -2095
rect 34485 -2215 34605 -2095
rect 34650 -2215 34770 -2095
rect 34815 -2215 34935 -2095
rect 34990 -2215 35110 -2095
rect 35155 -2215 35275 -2095
rect 35320 -2215 35440 -2095
rect 35485 -2215 35605 -2095
rect 35660 -2215 35780 -2095
rect 35825 -2215 35945 -2095
rect 35990 -2215 36110 -2095
rect 36155 -2215 36275 -2095
rect 30795 -2380 30915 -2260
rect 30970 -2380 31090 -2260
rect 31135 -2380 31255 -2260
rect 31300 -2380 31420 -2260
rect 31465 -2380 31585 -2260
rect 31640 -2380 31760 -2260
rect 31805 -2380 31925 -2260
rect 31970 -2380 32090 -2260
rect 32135 -2380 32255 -2260
rect 32310 -2380 32430 -2260
rect 32475 -2380 32595 -2260
rect 32640 -2380 32760 -2260
rect 32805 -2380 32925 -2260
rect 32980 -2380 33100 -2260
rect 33145 -2380 33265 -2260
rect 33310 -2380 33430 -2260
rect 33475 -2380 33595 -2260
rect 33650 -2380 33770 -2260
rect 33815 -2380 33935 -2260
rect 33980 -2380 34100 -2260
rect 34145 -2380 34265 -2260
rect 34320 -2380 34440 -2260
rect 34485 -2380 34605 -2260
rect 34650 -2380 34770 -2260
rect 34815 -2380 34935 -2260
rect 34990 -2380 35110 -2260
rect 35155 -2380 35275 -2260
rect 35320 -2380 35440 -2260
rect 35485 -2380 35605 -2260
rect 35660 -2380 35780 -2260
rect 35825 -2380 35945 -2260
rect 35990 -2380 36110 -2260
rect 36155 -2380 36275 -2260
rect 30795 -2545 30915 -2425
rect 30970 -2545 31090 -2425
rect 31135 -2545 31255 -2425
rect 31300 -2545 31420 -2425
rect 31465 -2545 31585 -2425
rect 31640 -2545 31760 -2425
rect 31805 -2545 31925 -2425
rect 31970 -2545 32090 -2425
rect 32135 -2545 32255 -2425
rect 32310 -2545 32430 -2425
rect 32475 -2545 32595 -2425
rect 32640 -2545 32760 -2425
rect 32805 -2545 32925 -2425
rect 32980 -2545 33100 -2425
rect 33145 -2545 33265 -2425
rect 33310 -2545 33430 -2425
rect 33475 -2545 33595 -2425
rect 33650 -2545 33770 -2425
rect 33815 -2545 33935 -2425
rect 33980 -2545 34100 -2425
rect 34145 -2545 34265 -2425
rect 34320 -2545 34440 -2425
rect 34485 -2545 34605 -2425
rect 34650 -2545 34770 -2425
rect 34815 -2545 34935 -2425
rect 34990 -2545 35110 -2425
rect 35155 -2545 35275 -2425
rect 35320 -2545 35440 -2425
rect 35485 -2545 35605 -2425
rect 35660 -2545 35780 -2425
rect 35825 -2545 35945 -2425
rect 35990 -2545 36110 -2425
rect 36155 -2545 36275 -2425
rect 30795 -2720 30915 -2600
rect 30970 -2720 31090 -2600
rect 31135 -2720 31255 -2600
rect 31300 -2720 31420 -2600
rect 31465 -2720 31585 -2600
rect 31640 -2720 31760 -2600
rect 31805 -2720 31925 -2600
rect 31970 -2720 32090 -2600
rect 32135 -2720 32255 -2600
rect 32310 -2720 32430 -2600
rect 32475 -2720 32595 -2600
rect 32640 -2720 32760 -2600
rect 32805 -2720 32925 -2600
rect 32980 -2720 33100 -2600
rect 33145 -2720 33265 -2600
rect 33310 -2720 33430 -2600
rect 33475 -2720 33595 -2600
rect 33650 -2720 33770 -2600
rect 33815 -2720 33935 -2600
rect 33980 -2720 34100 -2600
rect 34145 -2720 34265 -2600
rect 34320 -2720 34440 -2600
rect 34485 -2720 34605 -2600
rect 34650 -2720 34770 -2600
rect 34815 -2720 34935 -2600
rect 34990 -2720 35110 -2600
rect 35155 -2720 35275 -2600
rect 35320 -2720 35440 -2600
rect 35485 -2720 35605 -2600
rect 35660 -2720 35780 -2600
rect 35825 -2720 35945 -2600
rect 35990 -2720 36110 -2600
rect 36155 -2720 36275 -2600
rect 30795 -2885 30915 -2765
rect 30970 -2885 31090 -2765
rect 31135 -2885 31255 -2765
rect 31300 -2885 31420 -2765
rect 31465 -2885 31585 -2765
rect 31640 -2885 31760 -2765
rect 31805 -2885 31925 -2765
rect 31970 -2885 32090 -2765
rect 32135 -2885 32255 -2765
rect 32310 -2885 32430 -2765
rect 32475 -2885 32595 -2765
rect 32640 -2885 32760 -2765
rect 32805 -2885 32925 -2765
rect 32980 -2885 33100 -2765
rect 33145 -2885 33265 -2765
rect 33310 -2885 33430 -2765
rect 33475 -2885 33595 -2765
rect 33650 -2885 33770 -2765
rect 33815 -2885 33935 -2765
rect 33980 -2885 34100 -2765
rect 34145 -2885 34265 -2765
rect 34320 -2885 34440 -2765
rect 34485 -2885 34605 -2765
rect 34650 -2885 34770 -2765
rect 34815 -2885 34935 -2765
rect 34990 -2885 35110 -2765
rect 35155 -2885 35275 -2765
rect 35320 -2885 35440 -2765
rect 35485 -2885 35605 -2765
rect 35660 -2885 35780 -2765
rect 35825 -2885 35945 -2765
rect 35990 -2885 36110 -2765
rect 36155 -2885 36275 -2765
rect 30795 -3050 30915 -2930
rect 30970 -3050 31090 -2930
rect 31135 -3050 31255 -2930
rect 31300 -3050 31420 -2930
rect 31465 -3050 31585 -2930
rect 31640 -3050 31760 -2930
rect 31805 -3050 31925 -2930
rect 31970 -3050 32090 -2930
rect 32135 -3050 32255 -2930
rect 32310 -3050 32430 -2930
rect 32475 -3050 32595 -2930
rect 32640 -3050 32760 -2930
rect 32805 -3050 32925 -2930
rect 32980 -3050 33100 -2930
rect 33145 -3050 33265 -2930
rect 33310 -3050 33430 -2930
rect 33475 -3050 33595 -2930
rect 33650 -3050 33770 -2930
rect 33815 -3050 33935 -2930
rect 33980 -3050 34100 -2930
rect 34145 -3050 34265 -2930
rect 34320 -3050 34440 -2930
rect 34485 -3050 34605 -2930
rect 34650 -3050 34770 -2930
rect 34815 -3050 34935 -2930
rect 34990 -3050 35110 -2930
rect 35155 -3050 35275 -2930
rect 35320 -3050 35440 -2930
rect 35485 -3050 35605 -2930
rect 35660 -3050 35780 -2930
rect 35825 -3050 35945 -2930
rect 35990 -3050 36110 -2930
rect 36155 -3050 36275 -2930
rect 30795 -3215 30915 -3095
rect 30970 -3215 31090 -3095
rect 31135 -3215 31255 -3095
rect 31300 -3215 31420 -3095
rect 31465 -3215 31585 -3095
rect 31640 -3215 31760 -3095
rect 31805 -3215 31925 -3095
rect 31970 -3215 32090 -3095
rect 32135 -3215 32255 -3095
rect 32310 -3215 32430 -3095
rect 32475 -3215 32595 -3095
rect 32640 -3215 32760 -3095
rect 32805 -3215 32925 -3095
rect 32980 -3215 33100 -3095
rect 33145 -3215 33265 -3095
rect 33310 -3215 33430 -3095
rect 33475 -3215 33595 -3095
rect 33650 -3215 33770 -3095
rect 33815 -3215 33935 -3095
rect 33980 -3215 34100 -3095
rect 34145 -3215 34265 -3095
rect 34320 -3215 34440 -3095
rect 34485 -3215 34605 -3095
rect 34650 -3215 34770 -3095
rect 34815 -3215 34935 -3095
rect 34990 -3215 35110 -3095
rect 35155 -3215 35275 -3095
rect 35320 -3215 35440 -3095
rect 35485 -3215 35605 -3095
rect 35660 -3215 35780 -3095
rect 35825 -3215 35945 -3095
rect 35990 -3215 36110 -3095
rect 36155 -3215 36275 -3095
rect 30795 -3390 30915 -3270
rect 30970 -3390 31090 -3270
rect 31135 -3390 31255 -3270
rect 31300 -3390 31420 -3270
rect 31465 -3390 31585 -3270
rect 31640 -3390 31760 -3270
rect 31805 -3390 31925 -3270
rect 31970 -3390 32090 -3270
rect 32135 -3390 32255 -3270
rect 32310 -3390 32430 -3270
rect 32475 -3390 32595 -3270
rect 32640 -3390 32760 -3270
rect 32805 -3390 32925 -3270
rect 32980 -3390 33100 -3270
rect 33145 -3390 33265 -3270
rect 33310 -3390 33430 -3270
rect 33475 -3390 33595 -3270
rect 33650 -3390 33770 -3270
rect 33815 -3390 33935 -3270
rect 33980 -3390 34100 -3270
rect 34145 -3390 34265 -3270
rect 34320 -3390 34440 -3270
rect 34485 -3390 34605 -3270
rect 34650 -3390 34770 -3270
rect 34815 -3390 34935 -3270
rect 34990 -3390 35110 -3270
rect 35155 -3390 35275 -3270
rect 35320 -3390 35440 -3270
rect 35485 -3390 35605 -3270
rect 35660 -3390 35780 -3270
rect 35825 -3390 35945 -3270
rect 35990 -3390 36110 -3270
rect 36155 -3390 36275 -3270
rect 30795 -3555 30915 -3435
rect 30970 -3555 31090 -3435
rect 31135 -3555 31255 -3435
rect 31300 -3555 31420 -3435
rect 31465 -3555 31585 -3435
rect 31640 -3555 31760 -3435
rect 31805 -3555 31925 -3435
rect 31970 -3555 32090 -3435
rect 32135 -3555 32255 -3435
rect 32310 -3555 32430 -3435
rect 32475 -3555 32595 -3435
rect 32640 -3555 32760 -3435
rect 32805 -3555 32925 -3435
rect 32980 -3555 33100 -3435
rect 33145 -3555 33265 -3435
rect 33310 -3555 33430 -3435
rect 33475 -3555 33595 -3435
rect 33650 -3555 33770 -3435
rect 33815 -3555 33935 -3435
rect 33980 -3555 34100 -3435
rect 34145 -3555 34265 -3435
rect 34320 -3555 34440 -3435
rect 34485 -3555 34605 -3435
rect 34650 -3555 34770 -3435
rect 34815 -3555 34935 -3435
rect 34990 -3555 35110 -3435
rect 35155 -3555 35275 -3435
rect 35320 -3555 35440 -3435
rect 35485 -3555 35605 -3435
rect 35660 -3555 35780 -3435
rect 35825 -3555 35945 -3435
rect 35990 -3555 36110 -3435
rect 36155 -3555 36275 -3435
rect 30795 -3720 30915 -3600
rect 30970 -3720 31090 -3600
rect 31135 -3720 31255 -3600
rect 31300 -3720 31420 -3600
rect 31465 -3720 31585 -3600
rect 31640 -3720 31760 -3600
rect 31805 -3720 31925 -3600
rect 31970 -3720 32090 -3600
rect 32135 -3720 32255 -3600
rect 32310 -3720 32430 -3600
rect 32475 -3720 32595 -3600
rect 32640 -3720 32760 -3600
rect 32805 -3720 32925 -3600
rect 32980 -3720 33100 -3600
rect 33145 -3720 33265 -3600
rect 33310 -3720 33430 -3600
rect 33475 -3720 33595 -3600
rect 33650 -3720 33770 -3600
rect 33815 -3720 33935 -3600
rect 33980 -3720 34100 -3600
rect 34145 -3720 34265 -3600
rect 34320 -3720 34440 -3600
rect 34485 -3720 34605 -3600
rect 34650 -3720 34770 -3600
rect 34815 -3720 34935 -3600
rect 34990 -3720 35110 -3600
rect 35155 -3720 35275 -3600
rect 35320 -3720 35440 -3600
rect 35485 -3720 35605 -3600
rect 35660 -3720 35780 -3600
rect 35825 -3720 35945 -3600
rect 35990 -3720 36110 -3600
rect 36155 -3720 36275 -3600
rect 30795 -3885 30915 -3765
rect 30970 -3885 31090 -3765
rect 31135 -3885 31255 -3765
rect 31300 -3885 31420 -3765
rect 31465 -3885 31585 -3765
rect 31640 -3885 31760 -3765
rect 31805 -3885 31925 -3765
rect 31970 -3885 32090 -3765
rect 32135 -3885 32255 -3765
rect 32310 -3885 32430 -3765
rect 32475 -3885 32595 -3765
rect 32640 -3885 32760 -3765
rect 32805 -3885 32925 -3765
rect 32980 -3885 33100 -3765
rect 33145 -3885 33265 -3765
rect 33310 -3885 33430 -3765
rect 33475 -3885 33595 -3765
rect 33650 -3885 33770 -3765
rect 33815 -3885 33935 -3765
rect 33980 -3885 34100 -3765
rect 34145 -3885 34265 -3765
rect 34320 -3885 34440 -3765
rect 34485 -3885 34605 -3765
rect 34650 -3885 34770 -3765
rect 34815 -3885 34935 -3765
rect 34990 -3885 35110 -3765
rect 35155 -3885 35275 -3765
rect 35320 -3885 35440 -3765
rect 35485 -3885 35605 -3765
rect 35660 -3885 35780 -3765
rect 35825 -3885 35945 -3765
rect 35990 -3885 36110 -3765
rect 36155 -3885 36275 -3765
rect 30795 -4060 30915 -3940
rect 30970 -4060 31090 -3940
rect 31135 -4060 31255 -3940
rect 31300 -4060 31420 -3940
rect 31465 -4060 31585 -3940
rect 31640 -4060 31760 -3940
rect 31805 -4060 31925 -3940
rect 31970 -4060 32090 -3940
rect 32135 -4060 32255 -3940
rect 32310 -4060 32430 -3940
rect 32475 -4060 32595 -3940
rect 32640 -4060 32760 -3940
rect 32805 -4060 32925 -3940
rect 32980 -4060 33100 -3940
rect 33145 -4060 33265 -3940
rect 33310 -4060 33430 -3940
rect 33475 -4060 33595 -3940
rect 33650 -4060 33770 -3940
rect 33815 -4060 33935 -3940
rect 33980 -4060 34100 -3940
rect 34145 -4060 34265 -3940
rect 34320 -4060 34440 -3940
rect 34485 -4060 34605 -3940
rect 34650 -4060 34770 -3940
rect 34815 -4060 34935 -3940
rect 34990 -4060 35110 -3940
rect 35155 -4060 35275 -3940
rect 35320 -4060 35440 -3940
rect 35485 -4060 35605 -3940
rect 35660 -4060 35780 -3940
rect 35825 -4060 35945 -3940
rect 35990 -4060 36110 -3940
rect 36155 -4060 36275 -3940
rect 36485 1300 36605 1420
rect 36660 1300 36780 1420
rect 36825 1300 36945 1420
rect 36990 1300 37110 1420
rect 37155 1300 37275 1420
rect 37330 1300 37450 1420
rect 37495 1300 37615 1420
rect 37660 1300 37780 1420
rect 37825 1300 37945 1420
rect 38000 1300 38120 1420
rect 38165 1300 38285 1420
rect 38330 1300 38450 1420
rect 38495 1300 38615 1420
rect 38670 1300 38790 1420
rect 38835 1300 38955 1420
rect 39000 1300 39120 1420
rect 39165 1300 39285 1420
rect 39340 1300 39460 1420
rect 39505 1300 39625 1420
rect 39670 1300 39790 1420
rect 39835 1300 39955 1420
rect 40010 1300 40130 1420
rect 40175 1300 40295 1420
rect 40340 1300 40460 1420
rect 40505 1300 40625 1420
rect 40680 1300 40800 1420
rect 40845 1300 40965 1420
rect 41010 1300 41130 1420
rect 41175 1300 41295 1420
rect 41350 1300 41470 1420
rect 41515 1300 41635 1420
rect 41680 1300 41800 1420
rect 41845 1300 41965 1420
rect 36485 1135 36605 1255
rect 36660 1135 36780 1255
rect 36825 1135 36945 1255
rect 36990 1135 37110 1255
rect 37155 1135 37275 1255
rect 37330 1135 37450 1255
rect 37495 1135 37615 1255
rect 37660 1135 37780 1255
rect 37825 1135 37945 1255
rect 38000 1135 38120 1255
rect 38165 1135 38285 1255
rect 38330 1135 38450 1255
rect 38495 1135 38615 1255
rect 38670 1135 38790 1255
rect 38835 1135 38955 1255
rect 39000 1135 39120 1255
rect 39165 1135 39285 1255
rect 39340 1135 39460 1255
rect 39505 1135 39625 1255
rect 39670 1135 39790 1255
rect 39835 1135 39955 1255
rect 40010 1135 40130 1255
rect 40175 1135 40295 1255
rect 40340 1135 40460 1255
rect 40505 1135 40625 1255
rect 40680 1135 40800 1255
rect 40845 1135 40965 1255
rect 41010 1135 41130 1255
rect 41175 1135 41295 1255
rect 41350 1135 41470 1255
rect 41515 1135 41635 1255
rect 41680 1135 41800 1255
rect 41845 1135 41965 1255
rect 36485 970 36605 1090
rect 36660 970 36780 1090
rect 36825 970 36945 1090
rect 36990 970 37110 1090
rect 37155 970 37275 1090
rect 37330 970 37450 1090
rect 37495 970 37615 1090
rect 37660 970 37780 1090
rect 37825 970 37945 1090
rect 38000 970 38120 1090
rect 38165 970 38285 1090
rect 38330 970 38450 1090
rect 38495 970 38615 1090
rect 38670 970 38790 1090
rect 38835 970 38955 1090
rect 39000 970 39120 1090
rect 39165 970 39285 1090
rect 39340 970 39460 1090
rect 39505 970 39625 1090
rect 39670 970 39790 1090
rect 39835 970 39955 1090
rect 40010 970 40130 1090
rect 40175 970 40295 1090
rect 40340 970 40460 1090
rect 40505 970 40625 1090
rect 40680 970 40800 1090
rect 40845 970 40965 1090
rect 41010 970 41130 1090
rect 41175 970 41295 1090
rect 41350 970 41470 1090
rect 41515 970 41635 1090
rect 41680 970 41800 1090
rect 41845 970 41965 1090
rect 36485 805 36605 925
rect 36660 805 36780 925
rect 36825 805 36945 925
rect 36990 805 37110 925
rect 37155 805 37275 925
rect 37330 805 37450 925
rect 37495 805 37615 925
rect 37660 805 37780 925
rect 37825 805 37945 925
rect 38000 805 38120 925
rect 38165 805 38285 925
rect 38330 805 38450 925
rect 38495 805 38615 925
rect 38670 805 38790 925
rect 38835 805 38955 925
rect 39000 805 39120 925
rect 39165 805 39285 925
rect 39340 805 39460 925
rect 39505 805 39625 925
rect 39670 805 39790 925
rect 39835 805 39955 925
rect 40010 805 40130 925
rect 40175 805 40295 925
rect 40340 805 40460 925
rect 40505 805 40625 925
rect 40680 805 40800 925
rect 40845 805 40965 925
rect 41010 805 41130 925
rect 41175 805 41295 925
rect 41350 805 41470 925
rect 41515 805 41635 925
rect 41680 805 41800 925
rect 41845 805 41965 925
rect 36485 630 36605 750
rect 36660 630 36780 750
rect 36825 630 36945 750
rect 36990 630 37110 750
rect 37155 630 37275 750
rect 37330 630 37450 750
rect 37495 630 37615 750
rect 37660 630 37780 750
rect 37825 630 37945 750
rect 38000 630 38120 750
rect 38165 630 38285 750
rect 38330 630 38450 750
rect 38495 630 38615 750
rect 38670 630 38790 750
rect 38835 630 38955 750
rect 39000 630 39120 750
rect 39165 630 39285 750
rect 39340 630 39460 750
rect 39505 630 39625 750
rect 39670 630 39790 750
rect 39835 630 39955 750
rect 40010 630 40130 750
rect 40175 630 40295 750
rect 40340 630 40460 750
rect 40505 630 40625 750
rect 40680 630 40800 750
rect 40845 630 40965 750
rect 41010 630 41130 750
rect 41175 630 41295 750
rect 41350 630 41470 750
rect 41515 630 41635 750
rect 41680 630 41800 750
rect 41845 630 41965 750
rect 36485 465 36605 585
rect 36660 465 36780 585
rect 36825 465 36945 585
rect 36990 465 37110 585
rect 37155 465 37275 585
rect 37330 465 37450 585
rect 37495 465 37615 585
rect 37660 465 37780 585
rect 37825 465 37945 585
rect 38000 465 38120 585
rect 38165 465 38285 585
rect 38330 465 38450 585
rect 38495 465 38615 585
rect 38670 465 38790 585
rect 38835 465 38955 585
rect 39000 465 39120 585
rect 39165 465 39285 585
rect 39340 465 39460 585
rect 39505 465 39625 585
rect 39670 465 39790 585
rect 39835 465 39955 585
rect 40010 465 40130 585
rect 40175 465 40295 585
rect 40340 465 40460 585
rect 40505 465 40625 585
rect 40680 465 40800 585
rect 40845 465 40965 585
rect 41010 465 41130 585
rect 41175 465 41295 585
rect 41350 465 41470 585
rect 41515 465 41635 585
rect 41680 465 41800 585
rect 41845 465 41965 585
rect 36485 300 36605 420
rect 36660 300 36780 420
rect 36825 300 36945 420
rect 36990 300 37110 420
rect 37155 300 37275 420
rect 37330 300 37450 420
rect 37495 300 37615 420
rect 37660 300 37780 420
rect 37825 300 37945 420
rect 38000 300 38120 420
rect 38165 300 38285 420
rect 38330 300 38450 420
rect 38495 300 38615 420
rect 38670 300 38790 420
rect 38835 300 38955 420
rect 39000 300 39120 420
rect 39165 300 39285 420
rect 39340 300 39460 420
rect 39505 300 39625 420
rect 39670 300 39790 420
rect 39835 300 39955 420
rect 40010 300 40130 420
rect 40175 300 40295 420
rect 40340 300 40460 420
rect 40505 300 40625 420
rect 40680 300 40800 420
rect 40845 300 40965 420
rect 41010 300 41130 420
rect 41175 300 41295 420
rect 41350 300 41470 420
rect 41515 300 41635 420
rect 41680 300 41800 420
rect 41845 300 41965 420
rect 36485 135 36605 255
rect 36660 135 36780 255
rect 36825 135 36945 255
rect 36990 135 37110 255
rect 37155 135 37275 255
rect 37330 135 37450 255
rect 37495 135 37615 255
rect 37660 135 37780 255
rect 37825 135 37945 255
rect 38000 135 38120 255
rect 38165 135 38285 255
rect 38330 135 38450 255
rect 38495 135 38615 255
rect 38670 135 38790 255
rect 38835 135 38955 255
rect 39000 135 39120 255
rect 39165 135 39285 255
rect 39340 135 39460 255
rect 39505 135 39625 255
rect 39670 135 39790 255
rect 39835 135 39955 255
rect 40010 135 40130 255
rect 40175 135 40295 255
rect 40340 135 40460 255
rect 40505 135 40625 255
rect 40680 135 40800 255
rect 40845 135 40965 255
rect 41010 135 41130 255
rect 41175 135 41295 255
rect 41350 135 41470 255
rect 41515 135 41635 255
rect 41680 135 41800 255
rect 41845 135 41965 255
rect 36485 -40 36605 80
rect 36660 -40 36780 80
rect 36825 -40 36945 80
rect 36990 -40 37110 80
rect 37155 -40 37275 80
rect 37330 -40 37450 80
rect 37495 -40 37615 80
rect 37660 -40 37780 80
rect 37825 -40 37945 80
rect 38000 -40 38120 80
rect 38165 -40 38285 80
rect 38330 -40 38450 80
rect 38495 -40 38615 80
rect 38670 -40 38790 80
rect 38835 -40 38955 80
rect 39000 -40 39120 80
rect 39165 -40 39285 80
rect 39340 -40 39460 80
rect 39505 -40 39625 80
rect 39670 -40 39790 80
rect 39835 -40 39955 80
rect 40010 -40 40130 80
rect 40175 -40 40295 80
rect 40340 -40 40460 80
rect 40505 -40 40625 80
rect 40680 -40 40800 80
rect 40845 -40 40965 80
rect 41010 -40 41130 80
rect 41175 -40 41295 80
rect 41350 -40 41470 80
rect 41515 -40 41635 80
rect 41680 -40 41800 80
rect 41845 -40 41965 80
rect 36485 -205 36605 -85
rect 36660 -205 36780 -85
rect 36825 -205 36945 -85
rect 36990 -205 37110 -85
rect 37155 -205 37275 -85
rect 37330 -205 37450 -85
rect 37495 -205 37615 -85
rect 37660 -205 37780 -85
rect 37825 -205 37945 -85
rect 38000 -205 38120 -85
rect 38165 -205 38285 -85
rect 38330 -205 38450 -85
rect 38495 -205 38615 -85
rect 38670 -205 38790 -85
rect 38835 -205 38955 -85
rect 39000 -205 39120 -85
rect 39165 -205 39285 -85
rect 39340 -205 39460 -85
rect 39505 -205 39625 -85
rect 39670 -205 39790 -85
rect 39835 -205 39955 -85
rect 40010 -205 40130 -85
rect 40175 -205 40295 -85
rect 40340 -205 40460 -85
rect 40505 -205 40625 -85
rect 40680 -205 40800 -85
rect 40845 -205 40965 -85
rect 41010 -205 41130 -85
rect 41175 -205 41295 -85
rect 41350 -205 41470 -85
rect 41515 -205 41635 -85
rect 41680 -205 41800 -85
rect 41845 -205 41965 -85
rect 36485 -370 36605 -250
rect 36660 -370 36780 -250
rect 36825 -370 36945 -250
rect 36990 -370 37110 -250
rect 37155 -370 37275 -250
rect 37330 -370 37450 -250
rect 37495 -370 37615 -250
rect 37660 -370 37780 -250
rect 37825 -370 37945 -250
rect 38000 -370 38120 -250
rect 38165 -370 38285 -250
rect 38330 -370 38450 -250
rect 38495 -370 38615 -250
rect 38670 -370 38790 -250
rect 38835 -370 38955 -250
rect 39000 -370 39120 -250
rect 39165 -370 39285 -250
rect 39340 -370 39460 -250
rect 39505 -370 39625 -250
rect 39670 -370 39790 -250
rect 39835 -370 39955 -250
rect 40010 -370 40130 -250
rect 40175 -370 40295 -250
rect 40340 -370 40460 -250
rect 40505 -370 40625 -250
rect 40680 -370 40800 -250
rect 40845 -370 40965 -250
rect 41010 -370 41130 -250
rect 41175 -370 41295 -250
rect 41350 -370 41470 -250
rect 41515 -370 41635 -250
rect 41680 -370 41800 -250
rect 41845 -370 41965 -250
rect 36485 -535 36605 -415
rect 36660 -535 36780 -415
rect 36825 -535 36945 -415
rect 36990 -535 37110 -415
rect 37155 -535 37275 -415
rect 37330 -535 37450 -415
rect 37495 -535 37615 -415
rect 37660 -535 37780 -415
rect 37825 -535 37945 -415
rect 38000 -535 38120 -415
rect 38165 -535 38285 -415
rect 38330 -535 38450 -415
rect 38495 -535 38615 -415
rect 38670 -535 38790 -415
rect 38835 -535 38955 -415
rect 39000 -535 39120 -415
rect 39165 -535 39285 -415
rect 39340 -535 39460 -415
rect 39505 -535 39625 -415
rect 39670 -535 39790 -415
rect 39835 -535 39955 -415
rect 40010 -535 40130 -415
rect 40175 -535 40295 -415
rect 40340 -535 40460 -415
rect 40505 -535 40625 -415
rect 40680 -535 40800 -415
rect 40845 -535 40965 -415
rect 41010 -535 41130 -415
rect 41175 -535 41295 -415
rect 41350 -535 41470 -415
rect 41515 -535 41635 -415
rect 41680 -535 41800 -415
rect 41845 -535 41965 -415
rect 36485 -710 36605 -590
rect 36660 -710 36780 -590
rect 36825 -710 36945 -590
rect 36990 -710 37110 -590
rect 37155 -710 37275 -590
rect 37330 -710 37450 -590
rect 37495 -710 37615 -590
rect 37660 -710 37780 -590
rect 37825 -710 37945 -590
rect 38000 -710 38120 -590
rect 38165 -710 38285 -590
rect 38330 -710 38450 -590
rect 38495 -710 38615 -590
rect 38670 -710 38790 -590
rect 38835 -710 38955 -590
rect 39000 -710 39120 -590
rect 39165 -710 39285 -590
rect 39340 -710 39460 -590
rect 39505 -710 39625 -590
rect 39670 -710 39790 -590
rect 39835 -710 39955 -590
rect 40010 -710 40130 -590
rect 40175 -710 40295 -590
rect 40340 -710 40460 -590
rect 40505 -710 40625 -590
rect 40680 -710 40800 -590
rect 40845 -710 40965 -590
rect 41010 -710 41130 -590
rect 41175 -710 41295 -590
rect 41350 -710 41470 -590
rect 41515 -710 41635 -590
rect 41680 -710 41800 -590
rect 41845 -710 41965 -590
rect 36485 -875 36605 -755
rect 36660 -875 36780 -755
rect 36825 -875 36945 -755
rect 36990 -875 37110 -755
rect 37155 -875 37275 -755
rect 37330 -875 37450 -755
rect 37495 -875 37615 -755
rect 37660 -875 37780 -755
rect 37825 -875 37945 -755
rect 38000 -875 38120 -755
rect 38165 -875 38285 -755
rect 38330 -875 38450 -755
rect 38495 -875 38615 -755
rect 38670 -875 38790 -755
rect 38835 -875 38955 -755
rect 39000 -875 39120 -755
rect 39165 -875 39285 -755
rect 39340 -875 39460 -755
rect 39505 -875 39625 -755
rect 39670 -875 39790 -755
rect 39835 -875 39955 -755
rect 40010 -875 40130 -755
rect 40175 -875 40295 -755
rect 40340 -875 40460 -755
rect 40505 -875 40625 -755
rect 40680 -875 40800 -755
rect 40845 -875 40965 -755
rect 41010 -875 41130 -755
rect 41175 -875 41295 -755
rect 41350 -875 41470 -755
rect 41515 -875 41635 -755
rect 41680 -875 41800 -755
rect 41845 -875 41965 -755
rect 36485 -1040 36605 -920
rect 36660 -1040 36780 -920
rect 36825 -1040 36945 -920
rect 36990 -1040 37110 -920
rect 37155 -1040 37275 -920
rect 37330 -1040 37450 -920
rect 37495 -1040 37615 -920
rect 37660 -1040 37780 -920
rect 37825 -1040 37945 -920
rect 38000 -1040 38120 -920
rect 38165 -1040 38285 -920
rect 38330 -1040 38450 -920
rect 38495 -1040 38615 -920
rect 38670 -1040 38790 -920
rect 38835 -1040 38955 -920
rect 39000 -1040 39120 -920
rect 39165 -1040 39285 -920
rect 39340 -1040 39460 -920
rect 39505 -1040 39625 -920
rect 39670 -1040 39790 -920
rect 39835 -1040 39955 -920
rect 40010 -1040 40130 -920
rect 40175 -1040 40295 -920
rect 40340 -1040 40460 -920
rect 40505 -1040 40625 -920
rect 40680 -1040 40800 -920
rect 40845 -1040 40965 -920
rect 41010 -1040 41130 -920
rect 41175 -1040 41295 -920
rect 41350 -1040 41470 -920
rect 41515 -1040 41635 -920
rect 41680 -1040 41800 -920
rect 41845 -1040 41965 -920
rect 36485 -1205 36605 -1085
rect 36660 -1205 36780 -1085
rect 36825 -1205 36945 -1085
rect 36990 -1205 37110 -1085
rect 37155 -1205 37275 -1085
rect 37330 -1205 37450 -1085
rect 37495 -1205 37615 -1085
rect 37660 -1205 37780 -1085
rect 37825 -1205 37945 -1085
rect 38000 -1205 38120 -1085
rect 38165 -1205 38285 -1085
rect 38330 -1205 38450 -1085
rect 38495 -1205 38615 -1085
rect 38670 -1205 38790 -1085
rect 38835 -1205 38955 -1085
rect 39000 -1205 39120 -1085
rect 39165 -1205 39285 -1085
rect 39340 -1205 39460 -1085
rect 39505 -1205 39625 -1085
rect 39670 -1205 39790 -1085
rect 39835 -1205 39955 -1085
rect 40010 -1205 40130 -1085
rect 40175 -1205 40295 -1085
rect 40340 -1205 40460 -1085
rect 40505 -1205 40625 -1085
rect 40680 -1205 40800 -1085
rect 40845 -1205 40965 -1085
rect 41010 -1205 41130 -1085
rect 41175 -1205 41295 -1085
rect 41350 -1205 41470 -1085
rect 41515 -1205 41635 -1085
rect 41680 -1205 41800 -1085
rect 41845 -1205 41965 -1085
rect 36485 -1380 36605 -1260
rect 36660 -1380 36780 -1260
rect 36825 -1380 36945 -1260
rect 36990 -1380 37110 -1260
rect 37155 -1380 37275 -1260
rect 37330 -1380 37450 -1260
rect 37495 -1380 37615 -1260
rect 37660 -1380 37780 -1260
rect 37825 -1380 37945 -1260
rect 38000 -1380 38120 -1260
rect 38165 -1380 38285 -1260
rect 38330 -1380 38450 -1260
rect 38495 -1380 38615 -1260
rect 38670 -1380 38790 -1260
rect 38835 -1380 38955 -1260
rect 39000 -1380 39120 -1260
rect 39165 -1380 39285 -1260
rect 39340 -1380 39460 -1260
rect 39505 -1380 39625 -1260
rect 39670 -1380 39790 -1260
rect 39835 -1380 39955 -1260
rect 40010 -1380 40130 -1260
rect 40175 -1380 40295 -1260
rect 40340 -1380 40460 -1260
rect 40505 -1380 40625 -1260
rect 40680 -1380 40800 -1260
rect 40845 -1380 40965 -1260
rect 41010 -1380 41130 -1260
rect 41175 -1380 41295 -1260
rect 41350 -1380 41470 -1260
rect 41515 -1380 41635 -1260
rect 41680 -1380 41800 -1260
rect 41845 -1380 41965 -1260
rect 36485 -1545 36605 -1425
rect 36660 -1545 36780 -1425
rect 36825 -1545 36945 -1425
rect 36990 -1545 37110 -1425
rect 37155 -1545 37275 -1425
rect 37330 -1545 37450 -1425
rect 37495 -1545 37615 -1425
rect 37660 -1545 37780 -1425
rect 37825 -1545 37945 -1425
rect 38000 -1545 38120 -1425
rect 38165 -1545 38285 -1425
rect 38330 -1545 38450 -1425
rect 38495 -1545 38615 -1425
rect 38670 -1545 38790 -1425
rect 38835 -1545 38955 -1425
rect 39000 -1545 39120 -1425
rect 39165 -1545 39285 -1425
rect 39340 -1545 39460 -1425
rect 39505 -1545 39625 -1425
rect 39670 -1545 39790 -1425
rect 39835 -1545 39955 -1425
rect 40010 -1545 40130 -1425
rect 40175 -1545 40295 -1425
rect 40340 -1545 40460 -1425
rect 40505 -1545 40625 -1425
rect 40680 -1545 40800 -1425
rect 40845 -1545 40965 -1425
rect 41010 -1545 41130 -1425
rect 41175 -1545 41295 -1425
rect 41350 -1545 41470 -1425
rect 41515 -1545 41635 -1425
rect 41680 -1545 41800 -1425
rect 41845 -1545 41965 -1425
rect 36485 -1710 36605 -1590
rect 36660 -1710 36780 -1590
rect 36825 -1710 36945 -1590
rect 36990 -1710 37110 -1590
rect 37155 -1710 37275 -1590
rect 37330 -1710 37450 -1590
rect 37495 -1710 37615 -1590
rect 37660 -1710 37780 -1590
rect 37825 -1710 37945 -1590
rect 38000 -1710 38120 -1590
rect 38165 -1710 38285 -1590
rect 38330 -1710 38450 -1590
rect 38495 -1710 38615 -1590
rect 38670 -1710 38790 -1590
rect 38835 -1710 38955 -1590
rect 39000 -1710 39120 -1590
rect 39165 -1710 39285 -1590
rect 39340 -1710 39460 -1590
rect 39505 -1710 39625 -1590
rect 39670 -1710 39790 -1590
rect 39835 -1710 39955 -1590
rect 40010 -1710 40130 -1590
rect 40175 -1710 40295 -1590
rect 40340 -1710 40460 -1590
rect 40505 -1710 40625 -1590
rect 40680 -1710 40800 -1590
rect 40845 -1710 40965 -1590
rect 41010 -1710 41130 -1590
rect 41175 -1710 41295 -1590
rect 41350 -1710 41470 -1590
rect 41515 -1710 41635 -1590
rect 41680 -1710 41800 -1590
rect 41845 -1710 41965 -1590
rect 36485 -1875 36605 -1755
rect 36660 -1875 36780 -1755
rect 36825 -1875 36945 -1755
rect 36990 -1875 37110 -1755
rect 37155 -1875 37275 -1755
rect 37330 -1875 37450 -1755
rect 37495 -1875 37615 -1755
rect 37660 -1875 37780 -1755
rect 37825 -1875 37945 -1755
rect 38000 -1875 38120 -1755
rect 38165 -1875 38285 -1755
rect 38330 -1875 38450 -1755
rect 38495 -1875 38615 -1755
rect 38670 -1875 38790 -1755
rect 38835 -1875 38955 -1755
rect 39000 -1875 39120 -1755
rect 39165 -1875 39285 -1755
rect 39340 -1875 39460 -1755
rect 39505 -1875 39625 -1755
rect 39670 -1875 39790 -1755
rect 39835 -1875 39955 -1755
rect 40010 -1875 40130 -1755
rect 40175 -1875 40295 -1755
rect 40340 -1875 40460 -1755
rect 40505 -1875 40625 -1755
rect 40680 -1875 40800 -1755
rect 40845 -1875 40965 -1755
rect 41010 -1875 41130 -1755
rect 41175 -1875 41295 -1755
rect 41350 -1875 41470 -1755
rect 41515 -1875 41635 -1755
rect 41680 -1875 41800 -1755
rect 41845 -1875 41965 -1755
rect 36485 -2050 36605 -1930
rect 36660 -2050 36780 -1930
rect 36825 -2050 36945 -1930
rect 36990 -2050 37110 -1930
rect 37155 -2050 37275 -1930
rect 37330 -2050 37450 -1930
rect 37495 -2050 37615 -1930
rect 37660 -2050 37780 -1930
rect 37825 -2050 37945 -1930
rect 38000 -2050 38120 -1930
rect 38165 -2050 38285 -1930
rect 38330 -2050 38450 -1930
rect 38495 -2050 38615 -1930
rect 38670 -2050 38790 -1930
rect 38835 -2050 38955 -1930
rect 39000 -2050 39120 -1930
rect 39165 -2050 39285 -1930
rect 39340 -2050 39460 -1930
rect 39505 -2050 39625 -1930
rect 39670 -2050 39790 -1930
rect 39835 -2050 39955 -1930
rect 40010 -2050 40130 -1930
rect 40175 -2050 40295 -1930
rect 40340 -2050 40460 -1930
rect 40505 -2050 40625 -1930
rect 40680 -2050 40800 -1930
rect 40845 -2050 40965 -1930
rect 41010 -2050 41130 -1930
rect 41175 -2050 41295 -1930
rect 41350 -2050 41470 -1930
rect 41515 -2050 41635 -1930
rect 41680 -2050 41800 -1930
rect 41845 -2050 41965 -1930
rect 36485 -2215 36605 -2095
rect 36660 -2215 36780 -2095
rect 36825 -2215 36945 -2095
rect 36990 -2215 37110 -2095
rect 37155 -2215 37275 -2095
rect 37330 -2215 37450 -2095
rect 37495 -2215 37615 -2095
rect 37660 -2215 37780 -2095
rect 37825 -2215 37945 -2095
rect 38000 -2215 38120 -2095
rect 38165 -2215 38285 -2095
rect 38330 -2215 38450 -2095
rect 38495 -2215 38615 -2095
rect 38670 -2215 38790 -2095
rect 38835 -2215 38955 -2095
rect 39000 -2215 39120 -2095
rect 39165 -2215 39285 -2095
rect 39340 -2215 39460 -2095
rect 39505 -2215 39625 -2095
rect 39670 -2215 39790 -2095
rect 39835 -2215 39955 -2095
rect 40010 -2215 40130 -2095
rect 40175 -2215 40295 -2095
rect 40340 -2215 40460 -2095
rect 40505 -2215 40625 -2095
rect 40680 -2215 40800 -2095
rect 40845 -2215 40965 -2095
rect 41010 -2215 41130 -2095
rect 41175 -2215 41295 -2095
rect 41350 -2215 41470 -2095
rect 41515 -2215 41635 -2095
rect 41680 -2215 41800 -2095
rect 41845 -2215 41965 -2095
rect 36485 -2380 36605 -2260
rect 36660 -2380 36780 -2260
rect 36825 -2380 36945 -2260
rect 36990 -2380 37110 -2260
rect 37155 -2380 37275 -2260
rect 37330 -2380 37450 -2260
rect 37495 -2380 37615 -2260
rect 37660 -2380 37780 -2260
rect 37825 -2380 37945 -2260
rect 38000 -2380 38120 -2260
rect 38165 -2380 38285 -2260
rect 38330 -2380 38450 -2260
rect 38495 -2380 38615 -2260
rect 38670 -2380 38790 -2260
rect 38835 -2380 38955 -2260
rect 39000 -2380 39120 -2260
rect 39165 -2380 39285 -2260
rect 39340 -2380 39460 -2260
rect 39505 -2380 39625 -2260
rect 39670 -2380 39790 -2260
rect 39835 -2380 39955 -2260
rect 40010 -2380 40130 -2260
rect 40175 -2380 40295 -2260
rect 40340 -2380 40460 -2260
rect 40505 -2380 40625 -2260
rect 40680 -2380 40800 -2260
rect 40845 -2380 40965 -2260
rect 41010 -2380 41130 -2260
rect 41175 -2380 41295 -2260
rect 41350 -2380 41470 -2260
rect 41515 -2380 41635 -2260
rect 41680 -2380 41800 -2260
rect 41845 -2380 41965 -2260
rect 36485 -2545 36605 -2425
rect 36660 -2545 36780 -2425
rect 36825 -2545 36945 -2425
rect 36990 -2545 37110 -2425
rect 37155 -2545 37275 -2425
rect 37330 -2545 37450 -2425
rect 37495 -2545 37615 -2425
rect 37660 -2545 37780 -2425
rect 37825 -2545 37945 -2425
rect 38000 -2545 38120 -2425
rect 38165 -2545 38285 -2425
rect 38330 -2545 38450 -2425
rect 38495 -2545 38615 -2425
rect 38670 -2545 38790 -2425
rect 38835 -2545 38955 -2425
rect 39000 -2545 39120 -2425
rect 39165 -2545 39285 -2425
rect 39340 -2545 39460 -2425
rect 39505 -2545 39625 -2425
rect 39670 -2545 39790 -2425
rect 39835 -2545 39955 -2425
rect 40010 -2545 40130 -2425
rect 40175 -2545 40295 -2425
rect 40340 -2545 40460 -2425
rect 40505 -2545 40625 -2425
rect 40680 -2545 40800 -2425
rect 40845 -2545 40965 -2425
rect 41010 -2545 41130 -2425
rect 41175 -2545 41295 -2425
rect 41350 -2545 41470 -2425
rect 41515 -2545 41635 -2425
rect 41680 -2545 41800 -2425
rect 41845 -2545 41965 -2425
rect 36485 -2720 36605 -2600
rect 36660 -2720 36780 -2600
rect 36825 -2720 36945 -2600
rect 36990 -2720 37110 -2600
rect 37155 -2720 37275 -2600
rect 37330 -2720 37450 -2600
rect 37495 -2720 37615 -2600
rect 37660 -2720 37780 -2600
rect 37825 -2720 37945 -2600
rect 38000 -2720 38120 -2600
rect 38165 -2720 38285 -2600
rect 38330 -2720 38450 -2600
rect 38495 -2720 38615 -2600
rect 38670 -2720 38790 -2600
rect 38835 -2720 38955 -2600
rect 39000 -2720 39120 -2600
rect 39165 -2720 39285 -2600
rect 39340 -2720 39460 -2600
rect 39505 -2720 39625 -2600
rect 39670 -2720 39790 -2600
rect 39835 -2720 39955 -2600
rect 40010 -2720 40130 -2600
rect 40175 -2720 40295 -2600
rect 40340 -2720 40460 -2600
rect 40505 -2720 40625 -2600
rect 40680 -2720 40800 -2600
rect 40845 -2720 40965 -2600
rect 41010 -2720 41130 -2600
rect 41175 -2720 41295 -2600
rect 41350 -2720 41470 -2600
rect 41515 -2720 41635 -2600
rect 41680 -2720 41800 -2600
rect 41845 -2720 41965 -2600
rect 36485 -2885 36605 -2765
rect 36660 -2885 36780 -2765
rect 36825 -2885 36945 -2765
rect 36990 -2885 37110 -2765
rect 37155 -2885 37275 -2765
rect 37330 -2885 37450 -2765
rect 37495 -2885 37615 -2765
rect 37660 -2885 37780 -2765
rect 37825 -2885 37945 -2765
rect 38000 -2885 38120 -2765
rect 38165 -2885 38285 -2765
rect 38330 -2885 38450 -2765
rect 38495 -2885 38615 -2765
rect 38670 -2885 38790 -2765
rect 38835 -2885 38955 -2765
rect 39000 -2885 39120 -2765
rect 39165 -2885 39285 -2765
rect 39340 -2885 39460 -2765
rect 39505 -2885 39625 -2765
rect 39670 -2885 39790 -2765
rect 39835 -2885 39955 -2765
rect 40010 -2885 40130 -2765
rect 40175 -2885 40295 -2765
rect 40340 -2885 40460 -2765
rect 40505 -2885 40625 -2765
rect 40680 -2885 40800 -2765
rect 40845 -2885 40965 -2765
rect 41010 -2885 41130 -2765
rect 41175 -2885 41295 -2765
rect 41350 -2885 41470 -2765
rect 41515 -2885 41635 -2765
rect 41680 -2885 41800 -2765
rect 41845 -2885 41965 -2765
rect 36485 -3050 36605 -2930
rect 36660 -3050 36780 -2930
rect 36825 -3050 36945 -2930
rect 36990 -3050 37110 -2930
rect 37155 -3050 37275 -2930
rect 37330 -3050 37450 -2930
rect 37495 -3050 37615 -2930
rect 37660 -3050 37780 -2930
rect 37825 -3050 37945 -2930
rect 38000 -3050 38120 -2930
rect 38165 -3050 38285 -2930
rect 38330 -3050 38450 -2930
rect 38495 -3050 38615 -2930
rect 38670 -3050 38790 -2930
rect 38835 -3050 38955 -2930
rect 39000 -3050 39120 -2930
rect 39165 -3050 39285 -2930
rect 39340 -3050 39460 -2930
rect 39505 -3050 39625 -2930
rect 39670 -3050 39790 -2930
rect 39835 -3050 39955 -2930
rect 40010 -3050 40130 -2930
rect 40175 -3050 40295 -2930
rect 40340 -3050 40460 -2930
rect 40505 -3050 40625 -2930
rect 40680 -3050 40800 -2930
rect 40845 -3050 40965 -2930
rect 41010 -3050 41130 -2930
rect 41175 -3050 41295 -2930
rect 41350 -3050 41470 -2930
rect 41515 -3050 41635 -2930
rect 41680 -3050 41800 -2930
rect 41845 -3050 41965 -2930
rect 36485 -3215 36605 -3095
rect 36660 -3215 36780 -3095
rect 36825 -3215 36945 -3095
rect 36990 -3215 37110 -3095
rect 37155 -3215 37275 -3095
rect 37330 -3215 37450 -3095
rect 37495 -3215 37615 -3095
rect 37660 -3215 37780 -3095
rect 37825 -3215 37945 -3095
rect 38000 -3215 38120 -3095
rect 38165 -3215 38285 -3095
rect 38330 -3215 38450 -3095
rect 38495 -3215 38615 -3095
rect 38670 -3215 38790 -3095
rect 38835 -3215 38955 -3095
rect 39000 -3215 39120 -3095
rect 39165 -3215 39285 -3095
rect 39340 -3215 39460 -3095
rect 39505 -3215 39625 -3095
rect 39670 -3215 39790 -3095
rect 39835 -3215 39955 -3095
rect 40010 -3215 40130 -3095
rect 40175 -3215 40295 -3095
rect 40340 -3215 40460 -3095
rect 40505 -3215 40625 -3095
rect 40680 -3215 40800 -3095
rect 40845 -3215 40965 -3095
rect 41010 -3215 41130 -3095
rect 41175 -3215 41295 -3095
rect 41350 -3215 41470 -3095
rect 41515 -3215 41635 -3095
rect 41680 -3215 41800 -3095
rect 41845 -3215 41965 -3095
rect 36485 -3390 36605 -3270
rect 36660 -3390 36780 -3270
rect 36825 -3390 36945 -3270
rect 36990 -3390 37110 -3270
rect 37155 -3390 37275 -3270
rect 37330 -3390 37450 -3270
rect 37495 -3390 37615 -3270
rect 37660 -3390 37780 -3270
rect 37825 -3390 37945 -3270
rect 38000 -3390 38120 -3270
rect 38165 -3390 38285 -3270
rect 38330 -3390 38450 -3270
rect 38495 -3390 38615 -3270
rect 38670 -3390 38790 -3270
rect 38835 -3390 38955 -3270
rect 39000 -3390 39120 -3270
rect 39165 -3390 39285 -3270
rect 39340 -3390 39460 -3270
rect 39505 -3390 39625 -3270
rect 39670 -3390 39790 -3270
rect 39835 -3390 39955 -3270
rect 40010 -3390 40130 -3270
rect 40175 -3390 40295 -3270
rect 40340 -3390 40460 -3270
rect 40505 -3390 40625 -3270
rect 40680 -3390 40800 -3270
rect 40845 -3390 40965 -3270
rect 41010 -3390 41130 -3270
rect 41175 -3390 41295 -3270
rect 41350 -3390 41470 -3270
rect 41515 -3390 41635 -3270
rect 41680 -3390 41800 -3270
rect 41845 -3390 41965 -3270
rect 36485 -3555 36605 -3435
rect 36660 -3555 36780 -3435
rect 36825 -3555 36945 -3435
rect 36990 -3555 37110 -3435
rect 37155 -3555 37275 -3435
rect 37330 -3555 37450 -3435
rect 37495 -3555 37615 -3435
rect 37660 -3555 37780 -3435
rect 37825 -3555 37945 -3435
rect 38000 -3555 38120 -3435
rect 38165 -3555 38285 -3435
rect 38330 -3555 38450 -3435
rect 38495 -3555 38615 -3435
rect 38670 -3555 38790 -3435
rect 38835 -3555 38955 -3435
rect 39000 -3555 39120 -3435
rect 39165 -3555 39285 -3435
rect 39340 -3555 39460 -3435
rect 39505 -3555 39625 -3435
rect 39670 -3555 39790 -3435
rect 39835 -3555 39955 -3435
rect 40010 -3555 40130 -3435
rect 40175 -3555 40295 -3435
rect 40340 -3555 40460 -3435
rect 40505 -3555 40625 -3435
rect 40680 -3555 40800 -3435
rect 40845 -3555 40965 -3435
rect 41010 -3555 41130 -3435
rect 41175 -3555 41295 -3435
rect 41350 -3555 41470 -3435
rect 41515 -3555 41635 -3435
rect 41680 -3555 41800 -3435
rect 41845 -3555 41965 -3435
rect 36485 -3720 36605 -3600
rect 36660 -3720 36780 -3600
rect 36825 -3720 36945 -3600
rect 36990 -3720 37110 -3600
rect 37155 -3720 37275 -3600
rect 37330 -3720 37450 -3600
rect 37495 -3720 37615 -3600
rect 37660 -3720 37780 -3600
rect 37825 -3720 37945 -3600
rect 38000 -3720 38120 -3600
rect 38165 -3720 38285 -3600
rect 38330 -3720 38450 -3600
rect 38495 -3720 38615 -3600
rect 38670 -3720 38790 -3600
rect 38835 -3720 38955 -3600
rect 39000 -3720 39120 -3600
rect 39165 -3720 39285 -3600
rect 39340 -3720 39460 -3600
rect 39505 -3720 39625 -3600
rect 39670 -3720 39790 -3600
rect 39835 -3720 39955 -3600
rect 40010 -3720 40130 -3600
rect 40175 -3720 40295 -3600
rect 40340 -3720 40460 -3600
rect 40505 -3720 40625 -3600
rect 40680 -3720 40800 -3600
rect 40845 -3720 40965 -3600
rect 41010 -3720 41130 -3600
rect 41175 -3720 41295 -3600
rect 41350 -3720 41470 -3600
rect 41515 -3720 41635 -3600
rect 41680 -3720 41800 -3600
rect 41845 -3720 41965 -3600
rect 36485 -3885 36605 -3765
rect 36660 -3885 36780 -3765
rect 36825 -3885 36945 -3765
rect 36990 -3885 37110 -3765
rect 37155 -3885 37275 -3765
rect 37330 -3885 37450 -3765
rect 37495 -3885 37615 -3765
rect 37660 -3885 37780 -3765
rect 37825 -3885 37945 -3765
rect 38000 -3885 38120 -3765
rect 38165 -3885 38285 -3765
rect 38330 -3885 38450 -3765
rect 38495 -3885 38615 -3765
rect 38670 -3885 38790 -3765
rect 38835 -3885 38955 -3765
rect 39000 -3885 39120 -3765
rect 39165 -3885 39285 -3765
rect 39340 -3885 39460 -3765
rect 39505 -3885 39625 -3765
rect 39670 -3885 39790 -3765
rect 39835 -3885 39955 -3765
rect 40010 -3885 40130 -3765
rect 40175 -3885 40295 -3765
rect 40340 -3885 40460 -3765
rect 40505 -3885 40625 -3765
rect 40680 -3885 40800 -3765
rect 40845 -3885 40965 -3765
rect 41010 -3885 41130 -3765
rect 41175 -3885 41295 -3765
rect 41350 -3885 41470 -3765
rect 41515 -3885 41635 -3765
rect 41680 -3885 41800 -3765
rect 41845 -3885 41965 -3765
rect 36485 -4060 36605 -3940
rect 36660 -4060 36780 -3940
rect 36825 -4060 36945 -3940
rect 36990 -4060 37110 -3940
rect 37155 -4060 37275 -3940
rect 37330 -4060 37450 -3940
rect 37495 -4060 37615 -3940
rect 37660 -4060 37780 -3940
rect 37825 -4060 37945 -3940
rect 38000 -4060 38120 -3940
rect 38165 -4060 38285 -3940
rect 38330 -4060 38450 -3940
rect 38495 -4060 38615 -3940
rect 38670 -4060 38790 -3940
rect 38835 -4060 38955 -3940
rect 39000 -4060 39120 -3940
rect 39165 -4060 39285 -3940
rect 39340 -4060 39460 -3940
rect 39505 -4060 39625 -3940
rect 39670 -4060 39790 -3940
rect 39835 -4060 39955 -3940
rect 40010 -4060 40130 -3940
rect 40175 -4060 40295 -3940
rect 40340 -4060 40460 -3940
rect 40505 -4060 40625 -3940
rect 40680 -4060 40800 -3940
rect 40845 -4060 40965 -3940
rect 41010 -4060 41130 -3940
rect 41175 -4060 41295 -3940
rect 41350 -4060 41470 -3940
rect 41515 -4060 41635 -3940
rect 41680 -4060 41800 -3940
rect 41845 -4060 41965 -3940
rect 42175 1300 42295 1420
rect 42350 1300 42470 1420
rect 42515 1300 42635 1420
rect 42680 1300 42800 1420
rect 42845 1300 42965 1420
rect 43020 1300 43140 1420
rect 43185 1300 43305 1420
rect 43350 1300 43470 1420
rect 43515 1300 43635 1420
rect 43690 1300 43810 1420
rect 43855 1300 43975 1420
rect 44020 1300 44140 1420
rect 44185 1300 44305 1420
rect 44360 1300 44480 1420
rect 44525 1300 44645 1420
rect 44690 1300 44810 1420
rect 44855 1300 44975 1420
rect 45030 1300 45150 1420
rect 45195 1300 45315 1420
rect 45360 1300 45480 1420
rect 45525 1300 45645 1420
rect 45700 1300 45820 1420
rect 45865 1300 45985 1420
rect 46030 1300 46150 1420
rect 46195 1300 46315 1420
rect 46370 1300 46490 1420
rect 46535 1300 46655 1420
rect 46700 1300 46820 1420
rect 46865 1300 46985 1420
rect 47040 1300 47160 1420
rect 47205 1300 47325 1420
rect 47370 1300 47490 1420
rect 47535 1300 47655 1420
rect 42175 1135 42295 1255
rect 42350 1135 42470 1255
rect 42515 1135 42635 1255
rect 42680 1135 42800 1255
rect 42845 1135 42965 1255
rect 43020 1135 43140 1255
rect 43185 1135 43305 1255
rect 43350 1135 43470 1255
rect 43515 1135 43635 1255
rect 43690 1135 43810 1255
rect 43855 1135 43975 1255
rect 44020 1135 44140 1255
rect 44185 1135 44305 1255
rect 44360 1135 44480 1255
rect 44525 1135 44645 1255
rect 44690 1135 44810 1255
rect 44855 1135 44975 1255
rect 45030 1135 45150 1255
rect 45195 1135 45315 1255
rect 45360 1135 45480 1255
rect 45525 1135 45645 1255
rect 45700 1135 45820 1255
rect 45865 1135 45985 1255
rect 46030 1135 46150 1255
rect 46195 1135 46315 1255
rect 46370 1135 46490 1255
rect 46535 1135 46655 1255
rect 46700 1135 46820 1255
rect 46865 1135 46985 1255
rect 47040 1135 47160 1255
rect 47205 1135 47325 1255
rect 47370 1135 47490 1255
rect 47535 1135 47655 1255
rect 42175 970 42295 1090
rect 42350 970 42470 1090
rect 42515 970 42635 1090
rect 42680 970 42800 1090
rect 42845 970 42965 1090
rect 43020 970 43140 1090
rect 43185 970 43305 1090
rect 43350 970 43470 1090
rect 43515 970 43635 1090
rect 43690 970 43810 1090
rect 43855 970 43975 1090
rect 44020 970 44140 1090
rect 44185 970 44305 1090
rect 44360 970 44480 1090
rect 44525 970 44645 1090
rect 44690 970 44810 1090
rect 44855 970 44975 1090
rect 45030 970 45150 1090
rect 45195 970 45315 1090
rect 45360 970 45480 1090
rect 45525 970 45645 1090
rect 45700 970 45820 1090
rect 45865 970 45985 1090
rect 46030 970 46150 1090
rect 46195 970 46315 1090
rect 46370 970 46490 1090
rect 46535 970 46655 1090
rect 46700 970 46820 1090
rect 46865 970 46985 1090
rect 47040 970 47160 1090
rect 47205 970 47325 1090
rect 47370 970 47490 1090
rect 47535 970 47655 1090
rect 42175 805 42295 925
rect 42350 805 42470 925
rect 42515 805 42635 925
rect 42680 805 42800 925
rect 42845 805 42965 925
rect 43020 805 43140 925
rect 43185 805 43305 925
rect 43350 805 43470 925
rect 43515 805 43635 925
rect 43690 805 43810 925
rect 43855 805 43975 925
rect 44020 805 44140 925
rect 44185 805 44305 925
rect 44360 805 44480 925
rect 44525 805 44645 925
rect 44690 805 44810 925
rect 44855 805 44975 925
rect 45030 805 45150 925
rect 45195 805 45315 925
rect 45360 805 45480 925
rect 45525 805 45645 925
rect 45700 805 45820 925
rect 45865 805 45985 925
rect 46030 805 46150 925
rect 46195 805 46315 925
rect 46370 805 46490 925
rect 46535 805 46655 925
rect 46700 805 46820 925
rect 46865 805 46985 925
rect 47040 805 47160 925
rect 47205 805 47325 925
rect 47370 805 47490 925
rect 47535 805 47655 925
rect 42175 630 42295 750
rect 42350 630 42470 750
rect 42515 630 42635 750
rect 42680 630 42800 750
rect 42845 630 42965 750
rect 43020 630 43140 750
rect 43185 630 43305 750
rect 43350 630 43470 750
rect 43515 630 43635 750
rect 43690 630 43810 750
rect 43855 630 43975 750
rect 44020 630 44140 750
rect 44185 630 44305 750
rect 44360 630 44480 750
rect 44525 630 44645 750
rect 44690 630 44810 750
rect 44855 630 44975 750
rect 45030 630 45150 750
rect 45195 630 45315 750
rect 45360 630 45480 750
rect 45525 630 45645 750
rect 45700 630 45820 750
rect 45865 630 45985 750
rect 46030 630 46150 750
rect 46195 630 46315 750
rect 46370 630 46490 750
rect 46535 630 46655 750
rect 46700 630 46820 750
rect 46865 630 46985 750
rect 47040 630 47160 750
rect 47205 630 47325 750
rect 47370 630 47490 750
rect 47535 630 47655 750
rect 42175 465 42295 585
rect 42350 465 42470 585
rect 42515 465 42635 585
rect 42680 465 42800 585
rect 42845 465 42965 585
rect 43020 465 43140 585
rect 43185 465 43305 585
rect 43350 465 43470 585
rect 43515 465 43635 585
rect 43690 465 43810 585
rect 43855 465 43975 585
rect 44020 465 44140 585
rect 44185 465 44305 585
rect 44360 465 44480 585
rect 44525 465 44645 585
rect 44690 465 44810 585
rect 44855 465 44975 585
rect 45030 465 45150 585
rect 45195 465 45315 585
rect 45360 465 45480 585
rect 45525 465 45645 585
rect 45700 465 45820 585
rect 45865 465 45985 585
rect 46030 465 46150 585
rect 46195 465 46315 585
rect 46370 465 46490 585
rect 46535 465 46655 585
rect 46700 465 46820 585
rect 46865 465 46985 585
rect 47040 465 47160 585
rect 47205 465 47325 585
rect 47370 465 47490 585
rect 47535 465 47655 585
rect 42175 300 42295 420
rect 42350 300 42470 420
rect 42515 300 42635 420
rect 42680 300 42800 420
rect 42845 300 42965 420
rect 43020 300 43140 420
rect 43185 300 43305 420
rect 43350 300 43470 420
rect 43515 300 43635 420
rect 43690 300 43810 420
rect 43855 300 43975 420
rect 44020 300 44140 420
rect 44185 300 44305 420
rect 44360 300 44480 420
rect 44525 300 44645 420
rect 44690 300 44810 420
rect 44855 300 44975 420
rect 45030 300 45150 420
rect 45195 300 45315 420
rect 45360 300 45480 420
rect 45525 300 45645 420
rect 45700 300 45820 420
rect 45865 300 45985 420
rect 46030 300 46150 420
rect 46195 300 46315 420
rect 46370 300 46490 420
rect 46535 300 46655 420
rect 46700 300 46820 420
rect 46865 300 46985 420
rect 47040 300 47160 420
rect 47205 300 47325 420
rect 47370 300 47490 420
rect 47535 300 47655 420
rect 42175 135 42295 255
rect 42350 135 42470 255
rect 42515 135 42635 255
rect 42680 135 42800 255
rect 42845 135 42965 255
rect 43020 135 43140 255
rect 43185 135 43305 255
rect 43350 135 43470 255
rect 43515 135 43635 255
rect 43690 135 43810 255
rect 43855 135 43975 255
rect 44020 135 44140 255
rect 44185 135 44305 255
rect 44360 135 44480 255
rect 44525 135 44645 255
rect 44690 135 44810 255
rect 44855 135 44975 255
rect 45030 135 45150 255
rect 45195 135 45315 255
rect 45360 135 45480 255
rect 45525 135 45645 255
rect 45700 135 45820 255
rect 45865 135 45985 255
rect 46030 135 46150 255
rect 46195 135 46315 255
rect 46370 135 46490 255
rect 46535 135 46655 255
rect 46700 135 46820 255
rect 46865 135 46985 255
rect 47040 135 47160 255
rect 47205 135 47325 255
rect 47370 135 47490 255
rect 47535 135 47655 255
rect 42175 -40 42295 80
rect 42350 -40 42470 80
rect 42515 -40 42635 80
rect 42680 -40 42800 80
rect 42845 -40 42965 80
rect 43020 -40 43140 80
rect 43185 -40 43305 80
rect 43350 -40 43470 80
rect 43515 -40 43635 80
rect 43690 -40 43810 80
rect 43855 -40 43975 80
rect 44020 -40 44140 80
rect 44185 -40 44305 80
rect 44360 -40 44480 80
rect 44525 -40 44645 80
rect 44690 -40 44810 80
rect 44855 -40 44975 80
rect 45030 -40 45150 80
rect 45195 -40 45315 80
rect 45360 -40 45480 80
rect 45525 -40 45645 80
rect 45700 -40 45820 80
rect 45865 -40 45985 80
rect 46030 -40 46150 80
rect 46195 -40 46315 80
rect 46370 -40 46490 80
rect 46535 -40 46655 80
rect 46700 -40 46820 80
rect 46865 -40 46985 80
rect 47040 -40 47160 80
rect 47205 -40 47325 80
rect 47370 -40 47490 80
rect 47535 -40 47655 80
rect 42175 -205 42295 -85
rect 42350 -205 42470 -85
rect 42515 -205 42635 -85
rect 42680 -205 42800 -85
rect 42845 -205 42965 -85
rect 43020 -205 43140 -85
rect 43185 -205 43305 -85
rect 43350 -205 43470 -85
rect 43515 -205 43635 -85
rect 43690 -205 43810 -85
rect 43855 -205 43975 -85
rect 44020 -205 44140 -85
rect 44185 -205 44305 -85
rect 44360 -205 44480 -85
rect 44525 -205 44645 -85
rect 44690 -205 44810 -85
rect 44855 -205 44975 -85
rect 45030 -205 45150 -85
rect 45195 -205 45315 -85
rect 45360 -205 45480 -85
rect 45525 -205 45645 -85
rect 45700 -205 45820 -85
rect 45865 -205 45985 -85
rect 46030 -205 46150 -85
rect 46195 -205 46315 -85
rect 46370 -205 46490 -85
rect 46535 -205 46655 -85
rect 46700 -205 46820 -85
rect 46865 -205 46985 -85
rect 47040 -205 47160 -85
rect 47205 -205 47325 -85
rect 47370 -205 47490 -85
rect 47535 -205 47655 -85
rect 42175 -370 42295 -250
rect 42350 -370 42470 -250
rect 42515 -370 42635 -250
rect 42680 -370 42800 -250
rect 42845 -370 42965 -250
rect 43020 -370 43140 -250
rect 43185 -370 43305 -250
rect 43350 -370 43470 -250
rect 43515 -370 43635 -250
rect 43690 -370 43810 -250
rect 43855 -370 43975 -250
rect 44020 -370 44140 -250
rect 44185 -370 44305 -250
rect 44360 -370 44480 -250
rect 44525 -370 44645 -250
rect 44690 -370 44810 -250
rect 44855 -370 44975 -250
rect 45030 -370 45150 -250
rect 45195 -370 45315 -250
rect 45360 -370 45480 -250
rect 45525 -370 45645 -250
rect 45700 -370 45820 -250
rect 45865 -370 45985 -250
rect 46030 -370 46150 -250
rect 46195 -370 46315 -250
rect 46370 -370 46490 -250
rect 46535 -370 46655 -250
rect 46700 -370 46820 -250
rect 46865 -370 46985 -250
rect 47040 -370 47160 -250
rect 47205 -370 47325 -250
rect 47370 -370 47490 -250
rect 47535 -370 47655 -250
rect 42175 -535 42295 -415
rect 42350 -535 42470 -415
rect 42515 -535 42635 -415
rect 42680 -535 42800 -415
rect 42845 -535 42965 -415
rect 43020 -535 43140 -415
rect 43185 -535 43305 -415
rect 43350 -535 43470 -415
rect 43515 -535 43635 -415
rect 43690 -535 43810 -415
rect 43855 -535 43975 -415
rect 44020 -535 44140 -415
rect 44185 -535 44305 -415
rect 44360 -535 44480 -415
rect 44525 -535 44645 -415
rect 44690 -535 44810 -415
rect 44855 -535 44975 -415
rect 45030 -535 45150 -415
rect 45195 -535 45315 -415
rect 45360 -535 45480 -415
rect 45525 -535 45645 -415
rect 45700 -535 45820 -415
rect 45865 -535 45985 -415
rect 46030 -535 46150 -415
rect 46195 -535 46315 -415
rect 46370 -535 46490 -415
rect 46535 -535 46655 -415
rect 46700 -535 46820 -415
rect 46865 -535 46985 -415
rect 47040 -535 47160 -415
rect 47205 -535 47325 -415
rect 47370 -535 47490 -415
rect 47535 -535 47655 -415
rect 42175 -710 42295 -590
rect 42350 -710 42470 -590
rect 42515 -710 42635 -590
rect 42680 -710 42800 -590
rect 42845 -710 42965 -590
rect 43020 -710 43140 -590
rect 43185 -710 43305 -590
rect 43350 -710 43470 -590
rect 43515 -710 43635 -590
rect 43690 -710 43810 -590
rect 43855 -710 43975 -590
rect 44020 -710 44140 -590
rect 44185 -710 44305 -590
rect 44360 -710 44480 -590
rect 44525 -710 44645 -590
rect 44690 -710 44810 -590
rect 44855 -710 44975 -590
rect 45030 -710 45150 -590
rect 45195 -710 45315 -590
rect 45360 -710 45480 -590
rect 45525 -710 45645 -590
rect 45700 -710 45820 -590
rect 45865 -710 45985 -590
rect 46030 -710 46150 -590
rect 46195 -710 46315 -590
rect 46370 -710 46490 -590
rect 46535 -710 46655 -590
rect 46700 -710 46820 -590
rect 46865 -710 46985 -590
rect 47040 -710 47160 -590
rect 47205 -710 47325 -590
rect 47370 -710 47490 -590
rect 47535 -710 47655 -590
rect 42175 -875 42295 -755
rect 42350 -875 42470 -755
rect 42515 -875 42635 -755
rect 42680 -875 42800 -755
rect 42845 -875 42965 -755
rect 43020 -875 43140 -755
rect 43185 -875 43305 -755
rect 43350 -875 43470 -755
rect 43515 -875 43635 -755
rect 43690 -875 43810 -755
rect 43855 -875 43975 -755
rect 44020 -875 44140 -755
rect 44185 -875 44305 -755
rect 44360 -875 44480 -755
rect 44525 -875 44645 -755
rect 44690 -875 44810 -755
rect 44855 -875 44975 -755
rect 45030 -875 45150 -755
rect 45195 -875 45315 -755
rect 45360 -875 45480 -755
rect 45525 -875 45645 -755
rect 45700 -875 45820 -755
rect 45865 -875 45985 -755
rect 46030 -875 46150 -755
rect 46195 -875 46315 -755
rect 46370 -875 46490 -755
rect 46535 -875 46655 -755
rect 46700 -875 46820 -755
rect 46865 -875 46985 -755
rect 47040 -875 47160 -755
rect 47205 -875 47325 -755
rect 47370 -875 47490 -755
rect 47535 -875 47655 -755
rect 42175 -1040 42295 -920
rect 42350 -1040 42470 -920
rect 42515 -1040 42635 -920
rect 42680 -1040 42800 -920
rect 42845 -1040 42965 -920
rect 43020 -1040 43140 -920
rect 43185 -1040 43305 -920
rect 43350 -1040 43470 -920
rect 43515 -1040 43635 -920
rect 43690 -1040 43810 -920
rect 43855 -1040 43975 -920
rect 44020 -1040 44140 -920
rect 44185 -1040 44305 -920
rect 44360 -1040 44480 -920
rect 44525 -1040 44645 -920
rect 44690 -1040 44810 -920
rect 44855 -1040 44975 -920
rect 45030 -1040 45150 -920
rect 45195 -1040 45315 -920
rect 45360 -1040 45480 -920
rect 45525 -1040 45645 -920
rect 45700 -1040 45820 -920
rect 45865 -1040 45985 -920
rect 46030 -1040 46150 -920
rect 46195 -1040 46315 -920
rect 46370 -1040 46490 -920
rect 46535 -1040 46655 -920
rect 46700 -1040 46820 -920
rect 46865 -1040 46985 -920
rect 47040 -1040 47160 -920
rect 47205 -1040 47325 -920
rect 47370 -1040 47490 -920
rect 47535 -1040 47655 -920
rect 42175 -1205 42295 -1085
rect 42350 -1205 42470 -1085
rect 42515 -1205 42635 -1085
rect 42680 -1205 42800 -1085
rect 42845 -1205 42965 -1085
rect 43020 -1205 43140 -1085
rect 43185 -1205 43305 -1085
rect 43350 -1205 43470 -1085
rect 43515 -1205 43635 -1085
rect 43690 -1205 43810 -1085
rect 43855 -1205 43975 -1085
rect 44020 -1205 44140 -1085
rect 44185 -1205 44305 -1085
rect 44360 -1205 44480 -1085
rect 44525 -1205 44645 -1085
rect 44690 -1205 44810 -1085
rect 44855 -1205 44975 -1085
rect 45030 -1205 45150 -1085
rect 45195 -1205 45315 -1085
rect 45360 -1205 45480 -1085
rect 45525 -1205 45645 -1085
rect 45700 -1205 45820 -1085
rect 45865 -1205 45985 -1085
rect 46030 -1205 46150 -1085
rect 46195 -1205 46315 -1085
rect 46370 -1205 46490 -1085
rect 46535 -1205 46655 -1085
rect 46700 -1205 46820 -1085
rect 46865 -1205 46985 -1085
rect 47040 -1205 47160 -1085
rect 47205 -1205 47325 -1085
rect 47370 -1205 47490 -1085
rect 47535 -1205 47655 -1085
rect 42175 -1380 42295 -1260
rect 42350 -1380 42470 -1260
rect 42515 -1380 42635 -1260
rect 42680 -1380 42800 -1260
rect 42845 -1380 42965 -1260
rect 43020 -1380 43140 -1260
rect 43185 -1380 43305 -1260
rect 43350 -1380 43470 -1260
rect 43515 -1380 43635 -1260
rect 43690 -1380 43810 -1260
rect 43855 -1380 43975 -1260
rect 44020 -1380 44140 -1260
rect 44185 -1380 44305 -1260
rect 44360 -1380 44480 -1260
rect 44525 -1380 44645 -1260
rect 44690 -1380 44810 -1260
rect 44855 -1380 44975 -1260
rect 45030 -1380 45150 -1260
rect 45195 -1380 45315 -1260
rect 45360 -1380 45480 -1260
rect 45525 -1380 45645 -1260
rect 45700 -1380 45820 -1260
rect 45865 -1380 45985 -1260
rect 46030 -1380 46150 -1260
rect 46195 -1380 46315 -1260
rect 46370 -1380 46490 -1260
rect 46535 -1380 46655 -1260
rect 46700 -1380 46820 -1260
rect 46865 -1380 46985 -1260
rect 47040 -1380 47160 -1260
rect 47205 -1380 47325 -1260
rect 47370 -1380 47490 -1260
rect 47535 -1380 47655 -1260
rect 42175 -1545 42295 -1425
rect 42350 -1545 42470 -1425
rect 42515 -1545 42635 -1425
rect 42680 -1545 42800 -1425
rect 42845 -1545 42965 -1425
rect 43020 -1545 43140 -1425
rect 43185 -1545 43305 -1425
rect 43350 -1545 43470 -1425
rect 43515 -1545 43635 -1425
rect 43690 -1545 43810 -1425
rect 43855 -1545 43975 -1425
rect 44020 -1545 44140 -1425
rect 44185 -1545 44305 -1425
rect 44360 -1545 44480 -1425
rect 44525 -1545 44645 -1425
rect 44690 -1545 44810 -1425
rect 44855 -1545 44975 -1425
rect 45030 -1545 45150 -1425
rect 45195 -1545 45315 -1425
rect 45360 -1545 45480 -1425
rect 45525 -1545 45645 -1425
rect 45700 -1545 45820 -1425
rect 45865 -1545 45985 -1425
rect 46030 -1545 46150 -1425
rect 46195 -1545 46315 -1425
rect 46370 -1545 46490 -1425
rect 46535 -1545 46655 -1425
rect 46700 -1545 46820 -1425
rect 46865 -1545 46985 -1425
rect 47040 -1545 47160 -1425
rect 47205 -1545 47325 -1425
rect 47370 -1545 47490 -1425
rect 47535 -1545 47655 -1425
rect 42175 -1710 42295 -1590
rect 42350 -1710 42470 -1590
rect 42515 -1710 42635 -1590
rect 42680 -1710 42800 -1590
rect 42845 -1710 42965 -1590
rect 43020 -1710 43140 -1590
rect 43185 -1710 43305 -1590
rect 43350 -1710 43470 -1590
rect 43515 -1710 43635 -1590
rect 43690 -1710 43810 -1590
rect 43855 -1710 43975 -1590
rect 44020 -1710 44140 -1590
rect 44185 -1710 44305 -1590
rect 44360 -1710 44480 -1590
rect 44525 -1710 44645 -1590
rect 44690 -1710 44810 -1590
rect 44855 -1710 44975 -1590
rect 45030 -1710 45150 -1590
rect 45195 -1710 45315 -1590
rect 45360 -1710 45480 -1590
rect 45525 -1710 45645 -1590
rect 45700 -1710 45820 -1590
rect 45865 -1710 45985 -1590
rect 46030 -1710 46150 -1590
rect 46195 -1710 46315 -1590
rect 46370 -1710 46490 -1590
rect 46535 -1710 46655 -1590
rect 46700 -1710 46820 -1590
rect 46865 -1710 46985 -1590
rect 47040 -1710 47160 -1590
rect 47205 -1710 47325 -1590
rect 47370 -1710 47490 -1590
rect 47535 -1710 47655 -1590
rect 42175 -1875 42295 -1755
rect 42350 -1875 42470 -1755
rect 42515 -1875 42635 -1755
rect 42680 -1875 42800 -1755
rect 42845 -1875 42965 -1755
rect 43020 -1875 43140 -1755
rect 43185 -1875 43305 -1755
rect 43350 -1875 43470 -1755
rect 43515 -1875 43635 -1755
rect 43690 -1875 43810 -1755
rect 43855 -1875 43975 -1755
rect 44020 -1875 44140 -1755
rect 44185 -1875 44305 -1755
rect 44360 -1875 44480 -1755
rect 44525 -1875 44645 -1755
rect 44690 -1875 44810 -1755
rect 44855 -1875 44975 -1755
rect 45030 -1875 45150 -1755
rect 45195 -1875 45315 -1755
rect 45360 -1875 45480 -1755
rect 45525 -1875 45645 -1755
rect 45700 -1875 45820 -1755
rect 45865 -1875 45985 -1755
rect 46030 -1875 46150 -1755
rect 46195 -1875 46315 -1755
rect 46370 -1875 46490 -1755
rect 46535 -1875 46655 -1755
rect 46700 -1875 46820 -1755
rect 46865 -1875 46985 -1755
rect 47040 -1875 47160 -1755
rect 47205 -1875 47325 -1755
rect 47370 -1875 47490 -1755
rect 47535 -1875 47655 -1755
rect 42175 -2050 42295 -1930
rect 42350 -2050 42470 -1930
rect 42515 -2050 42635 -1930
rect 42680 -2050 42800 -1930
rect 42845 -2050 42965 -1930
rect 43020 -2050 43140 -1930
rect 43185 -2050 43305 -1930
rect 43350 -2050 43470 -1930
rect 43515 -2050 43635 -1930
rect 43690 -2050 43810 -1930
rect 43855 -2050 43975 -1930
rect 44020 -2050 44140 -1930
rect 44185 -2050 44305 -1930
rect 44360 -2050 44480 -1930
rect 44525 -2050 44645 -1930
rect 44690 -2050 44810 -1930
rect 44855 -2050 44975 -1930
rect 45030 -2050 45150 -1930
rect 45195 -2050 45315 -1930
rect 45360 -2050 45480 -1930
rect 45525 -2050 45645 -1930
rect 45700 -2050 45820 -1930
rect 45865 -2050 45985 -1930
rect 46030 -2050 46150 -1930
rect 46195 -2050 46315 -1930
rect 46370 -2050 46490 -1930
rect 46535 -2050 46655 -1930
rect 46700 -2050 46820 -1930
rect 46865 -2050 46985 -1930
rect 47040 -2050 47160 -1930
rect 47205 -2050 47325 -1930
rect 47370 -2050 47490 -1930
rect 47535 -2050 47655 -1930
rect 42175 -2215 42295 -2095
rect 42350 -2215 42470 -2095
rect 42515 -2215 42635 -2095
rect 42680 -2215 42800 -2095
rect 42845 -2215 42965 -2095
rect 43020 -2215 43140 -2095
rect 43185 -2215 43305 -2095
rect 43350 -2215 43470 -2095
rect 43515 -2215 43635 -2095
rect 43690 -2215 43810 -2095
rect 43855 -2215 43975 -2095
rect 44020 -2215 44140 -2095
rect 44185 -2215 44305 -2095
rect 44360 -2215 44480 -2095
rect 44525 -2215 44645 -2095
rect 44690 -2215 44810 -2095
rect 44855 -2215 44975 -2095
rect 45030 -2215 45150 -2095
rect 45195 -2215 45315 -2095
rect 45360 -2215 45480 -2095
rect 45525 -2215 45645 -2095
rect 45700 -2215 45820 -2095
rect 45865 -2215 45985 -2095
rect 46030 -2215 46150 -2095
rect 46195 -2215 46315 -2095
rect 46370 -2215 46490 -2095
rect 46535 -2215 46655 -2095
rect 46700 -2215 46820 -2095
rect 46865 -2215 46985 -2095
rect 47040 -2215 47160 -2095
rect 47205 -2215 47325 -2095
rect 47370 -2215 47490 -2095
rect 47535 -2215 47655 -2095
rect 42175 -2380 42295 -2260
rect 42350 -2380 42470 -2260
rect 42515 -2380 42635 -2260
rect 42680 -2380 42800 -2260
rect 42845 -2380 42965 -2260
rect 43020 -2380 43140 -2260
rect 43185 -2380 43305 -2260
rect 43350 -2380 43470 -2260
rect 43515 -2380 43635 -2260
rect 43690 -2380 43810 -2260
rect 43855 -2380 43975 -2260
rect 44020 -2380 44140 -2260
rect 44185 -2380 44305 -2260
rect 44360 -2380 44480 -2260
rect 44525 -2380 44645 -2260
rect 44690 -2380 44810 -2260
rect 44855 -2380 44975 -2260
rect 45030 -2380 45150 -2260
rect 45195 -2380 45315 -2260
rect 45360 -2380 45480 -2260
rect 45525 -2380 45645 -2260
rect 45700 -2380 45820 -2260
rect 45865 -2380 45985 -2260
rect 46030 -2380 46150 -2260
rect 46195 -2380 46315 -2260
rect 46370 -2380 46490 -2260
rect 46535 -2380 46655 -2260
rect 46700 -2380 46820 -2260
rect 46865 -2380 46985 -2260
rect 47040 -2380 47160 -2260
rect 47205 -2380 47325 -2260
rect 47370 -2380 47490 -2260
rect 47535 -2380 47655 -2260
rect 42175 -2545 42295 -2425
rect 42350 -2545 42470 -2425
rect 42515 -2545 42635 -2425
rect 42680 -2545 42800 -2425
rect 42845 -2545 42965 -2425
rect 43020 -2545 43140 -2425
rect 43185 -2545 43305 -2425
rect 43350 -2545 43470 -2425
rect 43515 -2545 43635 -2425
rect 43690 -2545 43810 -2425
rect 43855 -2545 43975 -2425
rect 44020 -2545 44140 -2425
rect 44185 -2545 44305 -2425
rect 44360 -2545 44480 -2425
rect 44525 -2545 44645 -2425
rect 44690 -2545 44810 -2425
rect 44855 -2545 44975 -2425
rect 45030 -2545 45150 -2425
rect 45195 -2545 45315 -2425
rect 45360 -2545 45480 -2425
rect 45525 -2545 45645 -2425
rect 45700 -2545 45820 -2425
rect 45865 -2545 45985 -2425
rect 46030 -2545 46150 -2425
rect 46195 -2545 46315 -2425
rect 46370 -2545 46490 -2425
rect 46535 -2545 46655 -2425
rect 46700 -2545 46820 -2425
rect 46865 -2545 46985 -2425
rect 47040 -2545 47160 -2425
rect 47205 -2545 47325 -2425
rect 47370 -2545 47490 -2425
rect 47535 -2545 47655 -2425
rect 42175 -2720 42295 -2600
rect 42350 -2720 42470 -2600
rect 42515 -2720 42635 -2600
rect 42680 -2720 42800 -2600
rect 42845 -2720 42965 -2600
rect 43020 -2720 43140 -2600
rect 43185 -2720 43305 -2600
rect 43350 -2720 43470 -2600
rect 43515 -2720 43635 -2600
rect 43690 -2720 43810 -2600
rect 43855 -2720 43975 -2600
rect 44020 -2720 44140 -2600
rect 44185 -2720 44305 -2600
rect 44360 -2720 44480 -2600
rect 44525 -2720 44645 -2600
rect 44690 -2720 44810 -2600
rect 44855 -2720 44975 -2600
rect 45030 -2720 45150 -2600
rect 45195 -2720 45315 -2600
rect 45360 -2720 45480 -2600
rect 45525 -2720 45645 -2600
rect 45700 -2720 45820 -2600
rect 45865 -2720 45985 -2600
rect 46030 -2720 46150 -2600
rect 46195 -2720 46315 -2600
rect 46370 -2720 46490 -2600
rect 46535 -2720 46655 -2600
rect 46700 -2720 46820 -2600
rect 46865 -2720 46985 -2600
rect 47040 -2720 47160 -2600
rect 47205 -2720 47325 -2600
rect 47370 -2720 47490 -2600
rect 47535 -2720 47655 -2600
rect 42175 -2885 42295 -2765
rect 42350 -2885 42470 -2765
rect 42515 -2885 42635 -2765
rect 42680 -2885 42800 -2765
rect 42845 -2885 42965 -2765
rect 43020 -2885 43140 -2765
rect 43185 -2885 43305 -2765
rect 43350 -2885 43470 -2765
rect 43515 -2885 43635 -2765
rect 43690 -2885 43810 -2765
rect 43855 -2885 43975 -2765
rect 44020 -2885 44140 -2765
rect 44185 -2885 44305 -2765
rect 44360 -2885 44480 -2765
rect 44525 -2885 44645 -2765
rect 44690 -2885 44810 -2765
rect 44855 -2885 44975 -2765
rect 45030 -2885 45150 -2765
rect 45195 -2885 45315 -2765
rect 45360 -2885 45480 -2765
rect 45525 -2885 45645 -2765
rect 45700 -2885 45820 -2765
rect 45865 -2885 45985 -2765
rect 46030 -2885 46150 -2765
rect 46195 -2885 46315 -2765
rect 46370 -2885 46490 -2765
rect 46535 -2885 46655 -2765
rect 46700 -2885 46820 -2765
rect 46865 -2885 46985 -2765
rect 47040 -2885 47160 -2765
rect 47205 -2885 47325 -2765
rect 47370 -2885 47490 -2765
rect 47535 -2885 47655 -2765
rect 42175 -3050 42295 -2930
rect 42350 -3050 42470 -2930
rect 42515 -3050 42635 -2930
rect 42680 -3050 42800 -2930
rect 42845 -3050 42965 -2930
rect 43020 -3050 43140 -2930
rect 43185 -3050 43305 -2930
rect 43350 -3050 43470 -2930
rect 43515 -3050 43635 -2930
rect 43690 -3050 43810 -2930
rect 43855 -3050 43975 -2930
rect 44020 -3050 44140 -2930
rect 44185 -3050 44305 -2930
rect 44360 -3050 44480 -2930
rect 44525 -3050 44645 -2930
rect 44690 -3050 44810 -2930
rect 44855 -3050 44975 -2930
rect 45030 -3050 45150 -2930
rect 45195 -3050 45315 -2930
rect 45360 -3050 45480 -2930
rect 45525 -3050 45645 -2930
rect 45700 -3050 45820 -2930
rect 45865 -3050 45985 -2930
rect 46030 -3050 46150 -2930
rect 46195 -3050 46315 -2930
rect 46370 -3050 46490 -2930
rect 46535 -3050 46655 -2930
rect 46700 -3050 46820 -2930
rect 46865 -3050 46985 -2930
rect 47040 -3050 47160 -2930
rect 47205 -3050 47325 -2930
rect 47370 -3050 47490 -2930
rect 47535 -3050 47655 -2930
rect 42175 -3215 42295 -3095
rect 42350 -3215 42470 -3095
rect 42515 -3215 42635 -3095
rect 42680 -3215 42800 -3095
rect 42845 -3215 42965 -3095
rect 43020 -3215 43140 -3095
rect 43185 -3215 43305 -3095
rect 43350 -3215 43470 -3095
rect 43515 -3215 43635 -3095
rect 43690 -3215 43810 -3095
rect 43855 -3215 43975 -3095
rect 44020 -3215 44140 -3095
rect 44185 -3215 44305 -3095
rect 44360 -3215 44480 -3095
rect 44525 -3215 44645 -3095
rect 44690 -3215 44810 -3095
rect 44855 -3215 44975 -3095
rect 45030 -3215 45150 -3095
rect 45195 -3215 45315 -3095
rect 45360 -3215 45480 -3095
rect 45525 -3215 45645 -3095
rect 45700 -3215 45820 -3095
rect 45865 -3215 45985 -3095
rect 46030 -3215 46150 -3095
rect 46195 -3215 46315 -3095
rect 46370 -3215 46490 -3095
rect 46535 -3215 46655 -3095
rect 46700 -3215 46820 -3095
rect 46865 -3215 46985 -3095
rect 47040 -3215 47160 -3095
rect 47205 -3215 47325 -3095
rect 47370 -3215 47490 -3095
rect 47535 -3215 47655 -3095
rect 42175 -3390 42295 -3270
rect 42350 -3390 42470 -3270
rect 42515 -3390 42635 -3270
rect 42680 -3390 42800 -3270
rect 42845 -3390 42965 -3270
rect 43020 -3390 43140 -3270
rect 43185 -3390 43305 -3270
rect 43350 -3390 43470 -3270
rect 43515 -3390 43635 -3270
rect 43690 -3390 43810 -3270
rect 43855 -3390 43975 -3270
rect 44020 -3390 44140 -3270
rect 44185 -3390 44305 -3270
rect 44360 -3390 44480 -3270
rect 44525 -3390 44645 -3270
rect 44690 -3390 44810 -3270
rect 44855 -3390 44975 -3270
rect 45030 -3390 45150 -3270
rect 45195 -3390 45315 -3270
rect 45360 -3390 45480 -3270
rect 45525 -3390 45645 -3270
rect 45700 -3390 45820 -3270
rect 45865 -3390 45985 -3270
rect 46030 -3390 46150 -3270
rect 46195 -3390 46315 -3270
rect 46370 -3390 46490 -3270
rect 46535 -3390 46655 -3270
rect 46700 -3390 46820 -3270
rect 46865 -3390 46985 -3270
rect 47040 -3390 47160 -3270
rect 47205 -3390 47325 -3270
rect 47370 -3390 47490 -3270
rect 47535 -3390 47655 -3270
rect 42175 -3555 42295 -3435
rect 42350 -3555 42470 -3435
rect 42515 -3555 42635 -3435
rect 42680 -3555 42800 -3435
rect 42845 -3555 42965 -3435
rect 43020 -3555 43140 -3435
rect 43185 -3555 43305 -3435
rect 43350 -3555 43470 -3435
rect 43515 -3555 43635 -3435
rect 43690 -3555 43810 -3435
rect 43855 -3555 43975 -3435
rect 44020 -3555 44140 -3435
rect 44185 -3555 44305 -3435
rect 44360 -3555 44480 -3435
rect 44525 -3555 44645 -3435
rect 44690 -3555 44810 -3435
rect 44855 -3555 44975 -3435
rect 45030 -3555 45150 -3435
rect 45195 -3555 45315 -3435
rect 45360 -3555 45480 -3435
rect 45525 -3555 45645 -3435
rect 45700 -3555 45820 -3435
rect 45865 -3555 45985 -3435
rect 46030 -3555 46150 -3435
rect 46195 -3555 46315 -3435
rect 46370 -3555 46490 -3435
rect 46535 -3555 46655 -3435
rect 46700 -3555 46820 -3435
rect 46865 -3555 46985 -3435
rect 47040 -3555 47160 -3435
rect 47205 -3555 47325 -3435
rect 47370 -3555 47490 -3435
rect 47535 -3555 47655 -3435
rect 42175 -3720 42295 -3600
rect 42350 -3720 42470 -3600
rect 42515 -3720 42635 -3600
rect 42680 -3720 42800 -3600
rect 42845 -3720 42965 -3600
rect 43020 -3720 43140 -3600
rect 43185 -3720 43305 -3600
rect 43350 -3720 43470 -3600
rect 43515 -3720 43635 -3600
rect 43690 -3720 43810 -3600
rect 43855 -3720 43975 -3600
rect 44020 -3720 44140 -3600
rect 44185 -3720 44305 -3600
rect 44360 -3720 44480 -3600
rect 44525 -3720 44645 -3600
rect 44690 -3720 44810 -3600
rect 44855 -3720 44975 -3600
rect 45030 -3720 45150 -3600
rect 45195 -3720 45315 -3600
rect 45360 -3720 45480 -3600
rect 45525 -3720 45645 -3600
rect 45700 -3720 45820 -3600
rect 45865 -3720 45985 -3600
rect 46030 -3720 46150 -3600
rect 46195 -3720 46315 -3600
rect 46370 -3720 46490 -3600
rect 46535 -3720 46655 -3600
rect 46700 -3720 46820 -3600
rect 46865 -3720 46985 -3600
rect 47040 -3720 47160 -3600
rect 47205 -3720 47325 -3600
rect 47370 -3720 47490 -3600
rect 47535 -3720 47655 -3600
rect 42175 -3885 42295 -3765
rect 42350 -3885 42470 -3765
rect 42515 -3885 42635 -3765
rect 42680 -3885 42800 -3765
rect 42845 -3885 42965 -3765
rect 43020 -3885 43140 -3765
rect 43185 -3885 43305 -3765
rect 43350 -3885 43470 -3765
rect 43515 -3885 43635 -3765
rect 43690 -3885 43810 -3765
rect 43855 -3885 43975 -3765
rect 44020 -3885 44140 -3765
rect 44185 -3885 44305 -3765
rect 44360 -3885 44480 -3765
rect 44525 -3885 44645 -3765
rect 44690 -3885 44810 -3765
rect 44855 -3885 44975 -3765
rect 45030 -3885 45150 -3765
rect 45195 -3885 45315 -3765
rect 45360 -3885 45480 -3765
rect 45525 -3885 45645 -3765
rect 45700 -3885 45820 -3765
rect 45865 -3885 45985 -3765
rect 46030 -3885 46150 -3765
rect 46195 -3885 46315 -3765
rect 46370 -3885 46490 -3765
rect 46535 -3885 46655 -3765
rect 46700 -3885 46820 -3765
rect 46865 -3885 46985 -3765
rect 47040 -3885 47160 -3765
rect 47205 -3885 47325 -3765
rect 47370 -3885 47490 -3765
rect 47535 -3885 47655 -3765
rect 42175 -4060 42295 -3940
rect 42350 -4060 42470 -3940
rect 42515 -4060 42635 -3940
rect 42680 -4060 42800 -3940
rect 42845 -4060 42965 -3940
rect 43020 -4060 43140 -3940
rect 43185 -4060 43305 -3940
rect 43350 -4060 43470 -3940
rect 43515 -4060 43635 -3940
rect 43690 -4060 43810 -3940
rect 43855 -4060 43975 -3940
rect 44020 -4060 44140 -3940
rect 44185 -4060 44305 -3940
rect 44360 -4060 44480 -3940
rect 44525 -4060 44645 -3940
rect 44690 -4060 44810 -3940
rect 44855 -4060 44975 -3940
rect 45030 -4060 45150 -3940
rect 45195 -4060 45315 -3940
rect 45360 -4060 45480 -3940
rect 45525 -4060 45645 -3940
rect 45700 -4060 45820 -3940
rect 45865 -4060 45985 -3940
rect 46030 -4060 46150 -3940
rect 46195 -4060 46315 -3940
rect 46370 -4060 46490 -3940
rect 46535 -4060 46655 -3940
rect 46700 -4060 46820 -3940
rect 46865 -4060 46985 -3940
rect 47040 -4060 47160 -3940
rect 47205 -4060 47325 -3940
rect 47370 -4060 47490 -3940
rect 47535 -4060 47655 -3940
rect 47865 1300 47985 1420
rect 48040 1300 48160 1420
rect 48205 1300 48325 1420
rect 48370 1300 48490 1420
rect 48535 1300 48655 1420
rect 48710 1300 48830 1420
rect 48875 1300 48995 1420
rect 49040 1300 49160 1420
rect 49205 1300 49325 1420
rect 49380 1300 49500 1420
rect 49545 1300 49665 1420
rect 49710 1300 49830 1420
rect 49875 1300 49995 1420
rect 50050 1300 50170 1420
rect 50215 1300 50335 1420
rect 50380 1300 50500 1420
rect 50545 1300 50665 1420
rect 50720 1300 50840 1420
rect 50885 1300 51005 1420
rect 51050 1300 51170 1420
rect 51215 1300 51335 1420
rect 51390 1300 51510 1420
rect 51555 1300 51675 1420
rect 51720 1300 51840 1420
rect 51885 1300 52005 1420
rect 52060 1300 52180 1420
rect 52225 1300 52345 1420
rect 52390 1300 52510 1420
rect 52555 1300 52675 1420
rect 52730 1300 52850 1420
rect 52895 1300 53015 1420
rect 53060 1300 53180 1420
rect 53225 1300 53345 1420
rect 47865 1135 47985 1255
rect 48040 1135 48160 1255
rect 48205 1135 48325 1255
rect 48370 1135 48490 1255
rect 48535 1135 48655 1255
rect 48710 1135 48830 1255
rect 48875 1135 48995 1255
rect 49040 1135 49160 1255
rect 49205 1135 49325 1255
rect 49380 1135 49500 1255
rect 49545 1135 49665 1255
rect 49710 1135 49830 1255
rect 49875 1135 49995 1255
rect 50050 1135 50170 1255
rect 50215 1135 50335 1255
rect 50380 1135 50500 1255
rect 50545 1135 50665 1255
rect 50720 1135 50840 1255
rect 50885 1135 51005 1255
rect 51050 1135 51170 1255
rect 51215 1135 51335 1255
rect 51390 1135 51510 1255
rect 51555 1135 51675 1255
rect 51720 1135 51840 1255
rect 51885 1135 52005 1255
rect 52060 1135 52180 1255
rect 52225 1135 52345 1255
rect 52390 1135 52510 1255
rect 52555 1135 52675 1255
rect 52730 1135 52850 1255
rect 52895 1135 53015 1255
rect 53060 1135 53180 1255
rect 53225 1135 53345 1255
rect 47865 970 47985 1090
rect 48040 970 48160 1090
rect 48205 970 48325 1090
rect 48370 970 48490 1090
rect 48535 970 48655 1090
rect 48710 970 48830 1090
rect 48875 970 48995 1090
rect 49040 970 49160 1090
rect 49205 970 49325 1090
rect 49380 970 49500 1090
rect 49545 970 49665 1090
rect 49710 970 49830 1090
rect 49875 970 49995 1090
rect 50050 970 50170 1090
rect 50215 970 50335 1090
rect 50380 970 50500 1090
rect 50545 970 50665 1090
rect 50720 970 50840 1090
rect 50885 970 51005 1090
rect 51050 970 51170 1090
rect 51215 970 51335 1090
rect 51390 970 51510 1090
rect 51555 970 51675 1090
rect 51720 970 51840 1090
rect 51885 970 52005 1090
rect 52060 970 52180 1090
rect 52225 970 52345 1090
rect 52390 970 52510 1090
rect 52555 970 52675 1090
rect 52730 970 52850 1090
rect 52895 970 53015 1090
rect 53060 970 53180 1090
rect 53225 970 53345 1090
rect 47865 805 47985 925
rect 48040 805 48160 925
rect 48205 805 48325 925
rect 48370 805 48490 925
rect 48535 805 48655 925
rect 48710 805 48830 925
rect 48875 805 48995 925
rect 49040 805 49160 925
rect 49205 805 49325 925
rect 49380 805 49500 925
rect 49545 805 49665 925
rect 49710 805 49830 925
rect 49875 805 49995 925
rect 50050 805 50170 925
rect 50215 805 50335 925
rect 50380 805 50500 925
rect 50545 805 50665 925
rect 50720 805 50840 925
rect 50885 805 51005 925
rect 51050 805 51170 925
rect 51215 805 51335 925
rect 51390 805 51510 925
rect 51555 805 51675 925
rect 51720 805 51840 925
rect 51885 805 52005 925
rect 52060 805 52180 925
rect 52225 805 52345 925
rect 52390 805 52510 925
rect 52555 805 52675 925
rect 52730 805 52850 925
rect 52895 805 53015 925
rect 53060 805 53180 925
rect 53225 805 53345 925
rect 47865 630 47985 750
rect 48040 630 48160 750
rect 48205 630 48325 750
rect 48370 630 48490 750
rect 48535 630 48655 750
rect 48710 630 48830 750
rect 48875 630 48995 750
rect 49040 630 49160 750
rect 49205 630 49325 750
rect 49380 630 49500 750
rect 49545 630 49665 750
rect 49710 630 49830 750
rect 49875 630 49995 750
rect 50050 630 50170 750
rect 50215 630 50335 750
rect 50380 630 50500 750
rect 50545 630 50665 750
rect 50720 630 50840 750
rect 50885 630 51005 750
rect 51050 630 51170 750
rect 51215 630 51335 750
rect 51390 630 51510 750
rect 51555 630 51675 750
rect 51720 630 51840 750
rect 51885 630 52005 750
rect 52060 630 52180 750
rect 52225 630 52345 750
rect 52390 630 52510 750
rect 52555 630 52675 750
rect 52730 630 52850 750
rect 52895 630 53015 750
rect 53060 630 53180 750
rect 53225 630 53345 750
rect 47865 465 47985 585
rect 48040 465 48160 585
rect 48205 465 48325 585
rect 48370 465 48490 585
rect 48535 465 48655 585
rect 48710 465 48830 585
rect 48875 465 48995 585
rect 49040 465 49160 585
rect 49205 465 49325 585
rect 49380 465 49500 585
rect 49545 465 49665 585
rect 49710 465 49830 585
rect 49875 465 49995 585
rect 50050 465 50170 585
rect 50215 465 50335 585
rect 50380 465 50500 585
rect 50545 465 50665 585
rect 50720 465 50840 585
rect 50885 465 51005 585
rect 51050 465 51170 585
rect 51215 465 51335 585
rect 51390 465 51510 585
rect 51555 465 51675 585
rect 51720 465 51840 585
rect 51885 465 52005 585
rect 52060 465 52180 585
rect 52225 465 52345 585
rect 52390 465 52510 585
rect 52555 465 52675 585
rect 52730 465 52850 585
rect 52895 465 53015 585
rect 53060 465 53180 585
rect 53225 465 53345 585
rect 47865 300 47985 420
rect 48040 300 48160 420
rect 48205 300 48325 420
rect 48370 300 48490 420
rect 48535 300 48655 420
rect 48710 300 48830 420
rect 48875 300 48995 420
rect 49040 300 49160 420
rect 49205 300 49325 420
rect 49380 300 49500 420
rect 49545 300 49665 420
rect 49710 300 49830 420
rect 49875 300 49995 420
rect 50050 300 50170 420
rect 50215 300 50335 420
rect 50380 300 50500 420
rect 50545 300 50665 420
rect 50720 300 50840 420
rect 50885 300 51005 420
rect 51050 300 51170 420
rect 51215 300 51335 420
rect 51390 300 51510 420
rect 51555 300 51675 420
rect 51720 300 51840 420
rect 51885 300 52005 420
rect 52060 300 52180 420
rect 52225 300 52345 420
rect 52390 300 52510 420
rect 52555 300 52675 420
rect 52730 300 52850 420
rect 52895 300 53015 420
rect 53060 300 53180 420
rect 53225 300 53345 420
rect 47865 135 47985 255
rect 48040 135 48160 255
rect 48205 135 48325 255
rect 48370 135 48490 255
rect 48535 135 48655 255
rect 48710 135 48830 255
rect 48875 135 48995 255
rect 49040 135 49160 255
rect 49205 135 49325 255
rect 49380 135 49500 255
rect 49545 135 49665 255
rect 49710 135 49830 255
rect 49875 135 49995 255
rect 50050 135 50170 255
rect 50215 135 50335 255
rect 50380 135 50500 255
rect 50545 135 50665 255
rect 50720 135 50840 255
rect 50885 135 51005 255
rect 51050 135 51170 255
rect 51215 135 51335 255
rect 51390 135 51510 255
rect 51555 135 51675 255
rect 51720 135 51840 255
rect 51885 135 52005 255
rect 52060 135 52180 255
rect 52225 135 52345 255
rect 52390 135 52510 255
rect 52555 135 52675 255
rect 52730 135 52850 255
rect 52895 135 53015 255
rect 53060 135 53180 255
rect 53225 135 53345 255
rect 47865 -40 47985 80
rect 48040 -40 48160 80
rect 48205 -40 48325 80
rect 48370 -40 48490 80
rect 48535 -40 48655 80
rect 48710 -40 48830 80
rect 48875 -40 48995 80
rect 49040 -40 49160 80
rect 49205 -40 49325 80
rect 49380 -40 49500 80
rect 49545 -40 49665 80
rect 49710 -40 49830 80
rect 49875 -40 49995 80
rect 50050 -40 50170 80
rect 50215 -40 50335 80
rect 50380 -40 50500 80
rect 50545 -40 50665 80
rect 50720 -40 50840 80
rect 50885 -40 51005 80
rect 51050 -40 51170 80
rect 51215 -40 51335 80
rect 51390 -40 51510 80
rect 51555 -40 51675 80
rect 51720 -40 51840 80
rect 51885 -40 52005 80
rect 52060 -40 52180 80
rect 52225 -40 52345 80
rect 52390 -40 52510 80
rect 52555 -40 52675 80
rect 52730 -40 52850 80
rect 52895 -40 53015 80
rect 53060 -40 53180 80
rect 53225 -40 53345 80
rect 47865 -205 47985 -85
rect 48040 -205 48160 -85
rect 48205 -205 48325 -85
rect 48370 -205 48490 -85
rect 48535 -205 48655 -85
rect 48710 -205 48830 -85
rect 48875 -205 48995 -85
rect 49040 -205 49160 -85
rect 49205 -205 49325 -85
rect 49380 -205 49500 -85
rect 49545 -205 49665 -85
rect 49710 -205 49830 -85
rect 49875 -205 49995 -85
rect 50050 -205 50170 -85
rect 50215 -205 50335 -85
rect 50380 -205 50500 -85
rect 50545 -205 50665 -85
rect 50720 -205 50840 -85
rect 50885 -205 51005 -85
rect 51050 -205 51170 -85
rect 51215 -205 51335 -85
rect 51390 -205 51510 -85
rect 51555 -205 51675 -85
rect 51720 -205 51840 -85
rect 51885 -205 52005 -85
rect 52060 -205 52180 -85
rect 52225 -205 52345 -85
rect 52390 -205 52510 -85
rect 52555 -205 52675 -85
rect 52730 -205 52850 -85
rect 52895 -205 53015 -85
rect 53060 -205 53180 -85
rect 53225 -205 53345 -85
rect 47865 -370 47985 -250
rect 48040 -370 48160 -250
rect 48205 -370 48325 -250
rect 48370 -370 48490 -250
rect 48535 -370 48655 -250
rect 48710 -370 48830 -250
rect 48875 -370 48995 -250
rect 49040 -370 49160 -250
rect 49205 -370 49325 -250
rect 49380 -370 49500 -250
rect 49545 -370 49665 -250
rect 49710 -370 49830 -250
rect 49875 -370 49995 -250
rect 50050 -370 50170 -250
rect 50215 -370 50335 -250
rect 50380 -370 50500 -250
rect 50545 -370 50665 -250
rect 50720 -370 50840 -250
rect 50885 -370 51005 -250
rect 51050 -370 51170 -250
rect 51215 -370 51335 -250
rect 51390 -370 51510 -250
rect 51555 -370 51675 -250
rect 51720 -370 51840 -250
rect 51885 -370 52005 -250
rect 52060 -370 52180 -250
rect 52225 -370 52345 -250
rect 52390 -370 52510 -250
rect 52555 -370 52675 -250
rect 52730 -370 52850 -250
rect 52895 -370 53015 -250
rect 53060 -370 53180 -250
rect 53225 -370 53345 -250
rect 47865 -535 47985 -415
rect 48040 -535 48160 -415
rect 48205 -535 48325 -415
rect 48370 -535 48490 -415
rect 48535 -535 48655 -415
rect 48710 -535 48830 -415
rect 48875 -535 48995 -415
rect 49040 -535 49160 -415
rect 49205 -535 49325 -415
rect 49380 -535 49500 -415
rect 49545 -535 49665 -415
rect 49710 -535 49830 -415
rect 49875 -535 49995 -415
rect 50050 -535 50170 -415
rect 50215 -535 50335 -415
rect 50380 -535 50500 -415
rect 50545 -535 50665 -415
rect 50720 -535 50840 -415
rect 50885 -535 51005 -415
rect 51050 -535 51170 -415
rect 51215 -535 51335 -415
rect 51390 -535 51510 -415
rect 51555 -535 51675 -415
rect 51720 -535 51840 -415
rect 51885 -535 52005 -415
rect 52060 -535 52180 -415
rect 52225 -535 52345 -415
rect 52390 -535 52510 -415
rect 52555 -535 52675 -415
rect 52730 -535 52850 -415
rect 52895 -535 53015 -415
rect 53060 -535 53180 -415
rect 53225 -535 53345 -415
rect 47865 -710 47985 -590
rect 48040 -710 48160 -590
rect 48205 -710 48325 -590
rect 48370 -710 48490 -590
rect 48535 -710 48655 -590
rect 48710 -710 48830 -590
rect 48875 -710 48995 -590
rect 49040 -710 49160 -590
rect 49205 -710 49325 -590
rect 49380 -710 49500 -590
rect 49545 -710 49665 -590
rect 49710 -710 49830 -590
rect 49875 -710 49995 -590
rect 50050 -710 50170 -590
rect 50215 -710 50335 -590
rect 50380 -710 50500 -590
rect 50545 -710 50665 -590
rect 50720 -710 50840 -590
rect 50885 -710 51005 -590
rect 51050 -710 51170 -590
rect 51215 -710 51335 -590
rect 51390 -710 51510 -590
rect 51555 -710 51675 -590
rect 51720 -710 51840 -590
rect 51885 -710 52005 -590
rect 52060 -710 52180 -590
rect 52225 -710 52345 -590
rect 52390 -710 52510 -590
rect 52555 -710 52675 -590
rect 52730 -710 52850 -590
rect 52895 -710 53015 -590
rect 53060 -710 53180 -590
rect 53225 -710 53345 -590
rect 47865 -875 47985 -755
rect 48040 -875 48160 -755
rect 48205 -875 48325 -755
rect 48370 -875 48490 -755
rect 48535 -875 48655 -755
rect 48710 -875 48830 -755
rect 48875 -875 48995 -755
rect 49040 -875 49160 -755
rect 49205 -875 49325 -755
rect 49380 -875 49500 -755
rect 49545 -875 49665 -755
rect 49710 -875 49830 -755
rect 49875 -875 49995 -755
rect 50050 -875 50170 -755
rect 50215 -875 50335 -755
rect 50380 -875 50500 -755
rect 50545 -875 50665 -755
rect 50720 -875 50840 -755
rect 50885 -875 51005 -755
rect 51050 -875 51170 -755
rect 51215 -875 51335 -755
rect 51390 -875 51510 -755
rect 51555 -875 51675 -755
rect 51720 -875 51840 -755
rect 51885 -875 52005 -755
rect 52060 -875 52180 -755
rect 52225 -875 52345 -755
rect 52390 -875 52510 -755
rect 52555 -875 52675 -755
rect 52730 -875 52850 -755
rect 52895 -875 53015 -755
rect 53060 -875 53180 -755
rect 53225 -875 53345 -755
rect 47865 -1040 47985 -920
rect 48040 -1040 48160 -920
rect 48205 -1040 48325 -920
rect 48370 -1040 48490 -920
rect 48535 -1040 48655 -920
rect 48710 -1040 48830 -920
rect 48875 -1040 48995 -920
rect 49040 -1040 49160 -920
rect 49205 -1040 49325 -920
rect 49380 -1040 49500 -920
rect 49545 -1040 49665 -920
rect 49710 -1040 49830 -920
rect 49875 -1040 49995 -920
rect 50050 -1040 50170 -920
rect 50215 -1040 50335 -920
rect 50380 -1040 50500 -920
rect 50545 -1040 50665 -920
rect 50720 -1040 50840 -920
rect 50885 -1040 51005 -920
rect 51050 -1040 51170 -920
rect 51215 -1040 51335 -920
rect 51390 -1040 51510 -920
rect 51555 -1040 51675 -920
rect 51720 -1040 51840 -920
rect 51885 -1040 52005 -920
rect 52060 -1040 52180 -920
rect 52225 -1040 52345 -920
rect 52390 -1040 52510 -920
rect 52555 -1040 52675 -920
rect 52730 -1040 52850 -920
rect 52895 -1040 53015 -920
rect 53060 -1040 53180 -920
rect 53225 -1040 53345 -920
rect 47865 -1205 47985 -1085
rect 48040 -1205 48160 -1085
rect 48205 -1205 48325 -1085
rect 48370 -1205 48490 -1085
rect 48535 -1205 48655 -1085
rect 48710 -1205 48830 -1085
rect 48875 -1205 48995 -1085
rect 49040 -1205 49160 -1085
rect 49205 -1205 49325 -1085
rect 49380 -1205 49500 -1085
rect 49545 -1205 49665 -1085
rect 49710 -1205 49830 -1085
rect 49875 -1205 49995 -1085
rect 50050 -1205 50170 -1085
rect 50215 -1205 50335 -1085
rect 50380 -1205 50500 -1085
rect 50545 -1205 50665 -1085
rect 50720 -1205 50840 -1085
rect 50885 -1205 51005 -1085
rect 51050 -1205 51170 -1085
rect 51215 -1205 51335 -1085
rect 51390 -1205 51510 -1085
rect 51555 -1205 51675 -1085
rect 51720 -1205 51840 -1085
rect 51885 -1205 52005 -1085
rect 52060 -1205 52180 -1085
rect 52225 -1205 52345 -1085
rect 52390 -1205 52510 -1085
rect 52555 -1205 52675 -1085
rect 52730 -1205 52850 -1085
rect 52895 -1205 53015 -1085
rect 53060 -1205 53180 -1085
rect 53225 -1205 53345 -1085
rect 47865 -1380 47985 -1260
rect 48040 -1380 48160 -1260
rect 48205 -1380 48325 -1260
rect 48370 -1380 48490 -1260
rect 48535 -1380 48655 -1260
rect 48710 -1380 48830 -1260
rect 48875 -1380 48995 -1260
rect 49040 -1380 49160 -1260
rect 49205 -1380 49325 -1260
rect 49380 -1380 49500 -1260
rect 49545 -1380 49665 -1260
rect 49710 -1380 49830 -1260
rect 49875 -1380 49995 -1260
rect 50050 -1380 50170 -1260
rect 50215 -1380 50335 -1260
rect 50380 -1380 50500 -1260
rect 50545 -1380 50665 -1260
rect 50720 -1380 50840 -1260
rect 50885 -1380 51005 -1260
rect 51050 -1380 51170 -1260
rect 51215 -1380 51335 -1260
rect 51390 -1380 51510 -1260
rect 51555 -1380 51675 -1260
rect 51720 -1380 51840 -1260
rect 51885 -1380 52005 -1260
rect 52060 -1380 52180 -1260
rect 52225 -1380 52345 -1260
rect 52390 -1380 52510 -1260
rect 52555 -1380 52675 -1260
rect 52730 -1380 52850 -1260
rect 52895 -1380 53015 -1260
rect 53060 -1380 53180 -1260
rect 53225 -1380 53345 -1260
rect 47865 -1545 47985 -1425
rect 48040 -1545 48160 -1425
rect 48205 -1545 48325 -1425
rect 48370 -1545 48490 -1425
rect 48535 -1545 48655 -1425
rect 48710 -1545 48830 -1425
rect 48875 -1545 48995 -1425
rect 49040 -1545 49160 -1425
rect 49205 -1545 49325 -1425
rect 49380 -1545 49500 -1425
rect 49545 -1545 49665 -1425
rect 49710 -1545 49830 -1425
rect 49875 -1545 49995 -1425
rect 50050 -1545 50170 -1425
rect 50215 -1545 50335 -1425
rect 50380 -1545 50500 -1425
rect 50545 -1545 50665 -1425
rect 50720 -1545 50840 -1425
rect 50885 -1545 51005 -1425
rect 51050 -1545 51170 -1425
rect 51215 -1545 51335 -1425
rect 51390 -1545 51510 -1425
rect 51555 -1545 51675 -1425
rect 51720 -1545 51840 -1425
rect 51885 -1545 52005 -1425
rect 52060 -1545 52180 -1425
rect 52225 -1545 52345 -1425
rect 52390 -1545 52510 -1425
rect 52555 -1545 52675 -1425
rect 52730 -1545 52850 -1425
rect 52895 -1545 53015 -1425
rect 53060 -1545 53180 -1425
rect 53225 -1545 53345 -1425
rect 47865 -1710 47985 -1590
rect 48040 -1710 48160 -1590
rect 48205 -1710 48325 -1590
rect 48370 -1710 48490 -1590
rect 48535 -1710 48655 -1590
rect 48710 -1710 48830 -1590
rect 48875 -1710 48995 -1590
rect 49040 -1710 49160 -1590
rect 49205 -1710 49325 -1590
rect 49380 -1710 49500 -1590
rect 49545 -1710 49665 -1590
rect 49710 -1710 49830 -1590
rect 49875 -1710 49995 -1590
rect 50050 -1710 50170 -1590
rect 50215 -1710 50335 -1590
rect 50380 -1710 50500 -1590
rect 50545 -1710 50665 -1590
rect 50720 -1710 50840 -1590
rect 50885 -1710 51005 -1590
rect 51050 -1710 51170 -1590
rect 51215 -1710 51335 -1590
rect 51390 -1710 51510 -1590
rect 51555 -1710 51675 -1590
rect 51720 -1710 51840 -1590
rect 51885 -1710 52005 -1590
rect 52060 -1710 52180 -1590
rect 52225 -1710 52345 -1590
rect 52390 -1710 52510 -1590
rect 52555 -1710 52675 -1590
rect 52730 -1710 52850 -1590
rect 52895 -1710 53015 -1590
rect 53060 -1710 53180 -1590
rect 53225 -1710 53345 -1590
rect 47865 -1875 47985 -1755
rect 48040 -1875 48160 -1755
rect 48205 -1875 48325 -1755
rect 48370 -1875 48490 -1755
rect 48535 -1875 48655 -1755
rect 48710 -1875 48830 -1755
rect 48875 -1875 48995 -1755
rect 49040 -1875 49160 -1755
rect 49205 -1875 49325 -1755
rect 49380 -1875 49500 -1755
rect 49545 -1875 49665 -1755
rect 49710 -1875 49830 -1755
rect 49875 -1875 49995 -1755
rect 50050 -1875 50170 -1755
rect 50215 -1875 50335 -1755
rect 50380 -1875 50500 -1755
rect 50545 -1875 50665 -1755
rect 50720 -1875 50840 -1755
rect 50885 -1875 51005 -1755
rect 51050 -1875 51170 -1755
rect 51215 -1875 51335 -1755
rect 51390 -1875 51510 -1755
rect 51555 -1875 51675 -1755
rect 51720 -1875 51840 -1755
rect 51885 -1875 52005 -1755
rect 52060 -1875 52180 -1755
rect 52225 -1875 52345 -1755
rect 52390 -1875 52510 -1755
rect 52555 -1875 52675 -1755
rect 52730 -1875 52850 -1755
rect 52895 -1875 53015 -1755
rect 53060 -1875 53180 -1755
rect 53225 -1875 53345 -1755
rect 47865 -2050 47985 -1930
rect 48040 -2050 48160 -1930
rect 48205 -2050 48325 -1930
rect 48370 -2050 48490 -1930
rect 48535 -2050 48655 -1930
rect 48710 -2050 48830 -1930
rect 48875 -2050 48995 -1930
rect 49040 -2050 49160 -1930
rect 49205 -2050 49325 -1930
rect 49380 -2050 49500 -1930
rect 49545 -2050 49665 -1930
rect 49710 -2050 49830 -1930
rect 49875 -2050 49995 -1930
rect 50050 -2050 50170 -1930
rect 50215 -2050 50335 -1930
rect 50380 -2050 50500 -1930
rect 50545 -2050 50665 -1930
rect 50720 -2050 50840 -1930
rect 50885 -2050 51005 -1930
rect 51050 -2050 51170 -1930
rect 51215 -2050 51335 -1930
rect 51390 -2050 51510 -1930
rect 51555 -2050 51675 -1930
rect 51720 -2050 51840 -1930
rect 51885 -2050 52005 -1930
rect 52060 -2050 52180 -1930
rect 52225 -2050 52345 -1930
rect 52390 -2050 52510 -1930
rect 52555 -2050 52675 -1930
rect 52730 -2050 52850 -1930
rect 52895 -2050 53015 -1930
rect 53060 -2050 53180 -1930
rect 53225 -2050 53345 -1930
rect 47865 -2215 47985 -2095
rect 48040 -2215 48160 -2095
rect 48205 -2215 48325 -2095
rect 48370 -2215 48490 -2095
rect 48535 -2215 48655 -2095
rect 48710 -2215 48830 -2095
rect 48875 -2215 48995 -2095
rect 49040 -2215 49160 -2095
rect 49205 -2215 49325 -2095
rect 49380 -2215 49500 -2095
rect 49545 -2215 49665 -2095
rect 49710 -2215 49830 -2095
rect 49875 -2215 49995 -2095
rect 50050 -2215 50170 -2095
rect 50215 -2215 50335 -2095
rect 50380 -2215 50500 -2095
rect 50545 -2215 50665 -2095
rect 50720 -2215 50840 -2095
rect 50885 -2215 51005 -2095
rect 51050 -2215 51170 -2095
rect 51215 -2215 51335 -2095
rect 51390 -2215 51510 -2095
rect 51555 -2215 51675 -2095
rect 51720 -2215 51840 -2095
rect 51885 -2215 52005 -2095
rect 52060 -2215 52180 -2095
rect 52225 -2215 52345 -2095
rect 52390 -2215 52510 -2095
rect 52555 -2215 52675 -2095
rect 52730 -2215 52850 -2095
rect 52895 -2215 53015 -2095
rect 53060 -2215 53180 -2095
rect 53225 -2215 53345 -2095
rect 47865 -2380 47985 -2260
rect 48040 -2380 48160 -2260
rect 48205 -2380 48325 -2260
rect 48370 -2380 48490 -2260
rect 48535 -2380 48655 -2260
rect 48710 -2380 48830 -2260
rect 48875 -2380 48995 -2260
rect 49040 -2380 49160 -2260
rect 49205 -2380 49325 -2260
rect 49380 -2380 49500 -2260
rect 49545 -2380 49665 -2260
rect 49710 -2380 49830 -2260
rect 49875 -2380 49995 -2260
rect 50050 -2380 50170 -2260
rect 50215 -2380 50335 -2260
rect 50380 -2380 50500 -2260
rect 50545 -2380 50665 -2260
rect 50720 -2380 50840 -2260
rect 50885 -2380 51005 -2260
rect 51050 -2380 51170 -2260
rect 51215 -2380 51335 -2260
rect 51390 -2380 51510 -2260
rect 51555 -2380 51675 -2260
rect 51720 -2380 51840 -2260
rect 51885 -2380 52005 -2260
rect 52060 -2380 52180 -2260
rect 52225 -2380 52345 -2260
rect 52390 -2380 52510 -2260
rect 52555 -2380 52675 -2260
rect 52730 -2380 52850 -2260
rect 52895 -2380 53015 -2260
rect 53060 -2380 53180 -2260
rect 53225 -2380 53345 -2260
rect 47865 -2545 47985 -2425
rect 48040 -2545 48160 -2425
rect 48205 -2545 48325 -2425
rect 48370 -2545 48490 -2425
rect 48535 -2545 48655 -2425
rect 48710 -2545 48830 -2425
rect 48875 -2545 48995 -2425
rect 49040 -2545 49160 -2425
rect 49205 -2545 49325 -2425
rect 49380 -2545 49500 -2425
rect 49545 -2545 49665 -2425
rect 49710 -2545 49830 -2425
rect 49875 -2545 49995 -2425
rect 50050 -2545 50170 -2425
rect 50215 -2545 50335 -2425
rect 50380 -2545 50500 -2425
rect 50545 -2545 50665 -2425
rect 50720 -2545 50840 -2425
rect 50885 -2545 51005 -2425
rect 51050 -2545 51170 -2425
rect 51215 -2545 51335 -2425
rect 51390 -2545 51510 -2425
rect 51555 -2545 51675 -2425
rect 51720 -2545 51840 -2425
rect 51885 -2545 52005 -2425
rect 52060 -2545 52180 -2425
rect 52225 -2545 52345 -2425
rect 52390 -2545 52510 -2425
rect 52555 -2545 52675 -2425
rect 52730 -2545 52850 -2425
rect 52895 -2545 53015 -2425
rect 53060 -2545 53180 -2425
rect 53225 -2545 53345 -2425
rect 47865 -2720 47985 -2600
rect 48040 -2720 48160 -2600
rect 48205 -2720 48325 -2600
rect 48370 -2720 48490 -2600
rect 48535 -2720 48655 -2600
rect 48710 -2720 48830 -2600
rect 48875 -2720 48995 -2600
rect 49040 -2720 49160 -2600
rect 49205 -2720 49325 -2600
rect 49380 -2720 49500 -2600
rect 49545 -2720 49665 -2600
rect 49710 -2720 49830 -2600
rect 49875 -2720 49995 -2600
rect 50050 -2720 50170 -2600
rect 50215 -2720 50335 -2600
rect 50380 -2720 50500 -2600
rect 50545 -2720 50665 -2600
rect 50720 -2720 50840 -2600
rect 50885 -2720 51005 -2600
rect 51050 -2720 51170 -2600
rect 51215 -2720 51335 -2600
rect 51390 -2720 51510 -2600
rect 51555 -2720 51675 -2600
rect 51720 -2720 51840 -2600
rect 51885 -2720 52005 -2600
rect 52060 -2720 52180 -2600
rect 52225 -2720 52345 -2600
rect 52390 -2720 52510 -2600
rect 52555 -2720 52675 -2600
rect 52730 -2720 52850 -2600
rect 52895 -2720 53015 -2600
rect 53060 -2720 53180 -2600
rect 53225 -2720 53345 -2600
rect 47865 -2885 47985 -2765
rect 48040 -2885 48160 -2765
rect 48205 -2885 48325 -2765
rect 48370 -2885 48490 -2765
rect 48535 -2885 48655 -2765
rect 48710 -2885 48830 -2765
rect 48875 -2885 48995 -2765
rect 49040 -2885 49160 -2765
rect 49205 -2885 49325 -2765
rect 49380 -2885 49500 -2765
rect 49545 -2885 49665 -2765
rect 49710 -2885 49830 -2765
rect 49875 -2885 49995 -2765
rect 50050 -2885 50170 -2765
rect 50215 -2885 50335 -2765
rect 50380 -2885 50500 -2765
rect 50545 -2885 50665 -2765
rect 50720 -2885 50840 -2765
rect 50885 -2885 51005 -2765
rect 51050 -2885 51170 -2765
rect 51215 -2885 51335 -2765
rect 51390 -2885 51510 -2765
rect 51555 -2885 51675 -2765
rect 51720 -2885 51840 -2765
rect 51885 -2885 52005 -2765
rect 52060 -2885 52180 -2765
rect 52225 -2885 52345 -2765
rect 52390 -2885 52510 -2765
rect 52555 -2885 52675 -2765
rect 52730 -2885 52850 -2765
rect 52895 -2885 53015 -2765
rect 53060 -2885 53180 -2765
rect 53225 -2885 53345 -2765
rect 47865 -3050 47985 -2930
rect 48040 -3050 48160 -2930
rect 48205 -3050 48325 -2930
rect 48370 -3050 48490 -2930
rect 48535 -3050 48655 -2930
rect 48710 -3050 48830 -2930
rect 48875 -3050 48995 -2930
rect 49040 -3050 49160 -2930
rect 49205 -3050 49325 -2930
rect 49380 -3050 49500 -2930
rect 49545 -3050 49665 -2930
rect 49710 -3050 49830 -2930
rect 49875 -3050 49995 -2930
rect 50050 -3050 50170 -2930
rect 50215 -3050 50335 -2930
rect 50380 -3050 50500 -2930
rect 50545 -3050 50665 -2930
rect 50720 -3050 50840 -2930
rect 50885 -3050 51005 -2930
rect 51050 -3050 51170 -2930
rect 51215 -3050 51335 -2930
rect 51390 -3050 51510 -2930
rect 51555 -3050 51675 -2930
rect 51720 -3050 51840 -2930
rect 51885 -3050 52005 -2930
rect 52060 -3050 52180 -2930
rect 52225 -3050 52345 -2930
rect 52390 -3050 52510 -2930
rect 52555 -3050 52675 -2930
rect 52730 -3050 52850 -2930
rect 52895 -3050 53015 -2930
rect 53060 -3050 53180 -2930
rect 53225 -3050 53345 -2930
rect 47865 -3215 47985 -3095
rect 48040 -3215 48160 -3095
rect 48205 -3215 48325 -3095
rect 48370 -3215 48490 -3095
rect 48535 -3215 48655 -3095
rect 48710 -3215 48830 -3095
rect 48875 -3215 48995 -3095
rect 49040 -3215 49160 -3095
rect 49205 -3215 49325 -3095
rect 49380 -3215 49500 -3095
rect 49545 -3215 49665 -3095
rect 49710 -3215 49830 -3095
rect 49875 -3215 49995 -3095
rect 50050 -3215 50170 -3095
rect 50215 -3215 50335 -3095
rect 50380 -3215 50500 -3095
rect 50545 -3215 50665 -3095
rect 50720 -3215 50840 -3095
rect 50885 -3215 51005 -3095
rect 51050 -3215 51170 -3095
rect 51215 -3215 51335 -3095
rect 51390 -3215 51510 -3095
rect 51555 -3215 51675 -3095
rect 51720 -3215 51840 -3095
rect 51885 -3215 52005 -3095
rect 52060 -3215 52180 -3095
rect 52225 -3215 52345 -3095
rect 52390 -3215 52510 -3095
rect 52555 -3215 52675 -3095
rect 52730 -3215 52850 -3095
rect 52895 -3215 53015 -3095
rect 53060 -3215 53180 -3095
rect 53225 -3215 53345 -3095
rect 47865 -3390 47985 -3270
rect 48040 -3390 48160 -3270
rect 48205 -3390 48325 -3270
rect 48370 -3390 48490 -3270
rect 48535 -3390 48655 -3270
rect 48710 -3390 48830 -3270
rect 48875 -3390 48995 -3270
rect 49040 -3390 49160 -3270
rect 49205 -3390 49325 -3270
rect 49380 -3390 49500 -3270
rect 49545 -3390 49665 -3270
rect 49710 -3390 49830 -3270
rect 49875 -3390 49995 -3270
rect 50050 -3390 50170 -3270
rect 50215 -3390 50335 -3270
rect 50380 -3390 50500 -3270
rect 50545 -3390 50665 -3270
rect 50720 -3390 50840 -3270
rect 50885 -3390 51005 -3270
rect 51050 -3390 51170 -3270
rect 51215 -3390 51335 -3270
rect 51390 -3390 51510 -3270
rect 51555 -3390 51675 -3270
rect 51720 -3390 51840 -3270
rect 51885 -3390 52005 -3270
rect 52060 -3390 52180 -3270
rect 52225 -3390 52345 -3270
rect 52390 -3390 52510 -3270
rect 52555 -3390 52675 -3270
rect 52730 -3390 52850 -3270
rect 52895 -3390 53015 -3270
rect 53060 -3390 53180 -3270
rect 53225 -3390 53345 -3270
rect 47865 -3555 47985 -3435
rect 48040 -3555 48160 -3435
rect 48205 -3555 48325 -3435
rect 48370 -3555 48490 -3435
rect 48535 -3555 48655 -3435
rect 48710 -3555 48830 -3435
rect 48875 -3555 48995 -3435
rect 49040 -3555 49160 -3435
rect 49205 -3555 49325 -3435
rect 49380 -3555 49500 -3435
rect 49545 -3555 49665 -3435
rect 49710 -3555 49830 -3435
rect 49875 -3555 49995 -3435
rect 50050 -3555 50170 -3435
rect 50215 -3555 50335 -3435
rect 50380 -3555 50500 -3435
rect 50545 -3555 50665 -3435
rect 50720 -3555 50840 -3435
rect 50885 -3555 51005 -3435
rect 51050 -3555 51170 -3435
rect 51215 -3555 51335 -3435
rect 51390 -3555 51510 -3435
rect 51555 -3555 51675 -3435
rect 51720 -3555 51840 -3435
rect 51885 -3555 52005 -3435
rect 52060 -3555 52180 -3435
rect 52225 -3555 52345 -3435
rect 52390 -3555 52510 -3435
rect 52555 -3555 52675 -3435
rect 52730 -3555 52850 -3435
rect 52895 -3555 53015 -3435
rect 53060 -3555 53180 -3435
rect 53225 -3555 53345 -3435
rect 47865 -3720 47985 -3600
rect 48040 -3720 48160 -3600
rect 48205 -3720 48325 -3600
rect 48370 -3720 48490 -3600
rect 48535 -3720 48655 -3600
rect 48710 -3720 48830 -3600
rect 48875 -3720 48995 -3600
rect 49040 -3720 49160 -3600
rect 49205 -3720 49325 -3600
rect 49380 -3720 49500 -3600
rect 49545 -3720 49665 -3600
rect 49710 -3720 49830 -3600
rect 49875 -3720 49995 -3600
rect 50050 -3720 50170 -3600
rect 50215 -3720 50335 -3600
rect 50380 -3720 50500 -3600
rect 50545 -3720 50665 -3600
rect 50720 -3720 50840 -3600
rect 50885 -3720 51005 -3600
rect 51050 -3720 51170 -3600
rect 51215 -3720 51335 -3600
rect 51390 -3720 51510 -3600
rect 51555 -3720 51675 -3600
rect 51720 -3720 51840 -3600
rect 51885 -3720 52005 -3600
rect 52060 -3720 52180 -3600
rect 52225 -3720 52345 -3600
rect 52390 -3720 52510 -3600
rect 52555 -3720 52675 -3600
rect 52730 -3720 52850 -3600
rect 52895 -3720 53015 -3600
rect 53060 -3720 53180 -3600
rect 53225 -3720 53345 -3600
rect 47865 -3885 47985 -3765
rect 48040 -3885 48160 -3765
rect 48205 -3885 48325 -3765
rect 48370 -3885 48490 -3765
rect 48535 -3885 48655 -3765
rect 48710 -3885 48830 -3765
rect 48875 -3885 48995 -3765
rect 49040 -3885 49160 -3765
rect 49205 -3885 49325 -3765
rect 49380 -3885 49500 -3765
rect 49545 -3885 49665 -3765
rect 49710 -3885 49830 -3765
rect 49875 -3885 49995 -3765
rect 50050 -3885 50170 -3765
rect 50215 -3885 50335 -3765
rect 50380 -3885 50500 -3765
rect 50545 -3885 50665 -3765
rect 50720 -3885 50840 -3765
rect 50885 -3885 51005 -3765
rect 51050 -3885 51170 -3765
rect 51215 -3885 51335 -3765
rect 51390 -3885 51510 -3765
rect 51555 -3885 51675 -3765
rect 51720 -3885 51840 -3765
rect 51885 -3885 52005 -3765
rect 52060 -3885 52180 -3765
rect 52225 -3885 52345 -3765
rect 52390 -3885 52510 -3765
rect 52555 -3885 52675 -3765
rect 52730 -3885 52850 -3765
rect 52895 -3885 53015 -3765
rect 53060 -3885 53180 -3765
rect 53225 -3885 53345 -3765
rect 47865 -4060 47985 -3940
rect 48040 -4060 48160 -3940
rect 48205 -4060 48325 -3940
rect 48370 -4060 48490 -3940
rect 48535 -4060 48655 -3940
rect 48710 -4060 48830 -3940
rect 48875 -4060 48995 -3940
rect 49040 -4060 49160 -3940
rect 49205 -4060 49325 -3940
rect 49380 -4060 49500 -3940
rect 49545 -4060 49665 -3940
rect 49710 -4060 49830 -3940
rect 49875 -4060 49995 -3940
rect 50050 -4060 50170 -3940
rect 50215 -4060 50335 -3940
rect 50380 -4060 50500 -3940
rect 50545 -4060 50665 -3940
rect 50720 -4060 50840 -3940
rect 50885 -4060 51005 -3940
rect 51050 -4060 51170 -3940
rect 51215 -4060 51335 -3940
rect 51390 -4060 51510 -3940
rect 51555 -4060 51675 -3940
rect 51720 -4060 51840 -3940
rect 51885 -4060 52005 -3940
rect 52060 -4060 52180 -3940
rect 52225 -4060 52345 -3940
rect 52390 -4060 52510 -3940
rect 52555 -4060 52675 -3940
rect 52730 -4060 52850 -3940
rect 52895 -4060 53015 -3940
rect 53060 -4060 53180 -3940
rect 53225 -4060 53345 -3940
rect 30795 -4390 30915 -4270
rect 30960 -4390 31080 -4270
rect 31125 -4390 31245 -4270
rect 31290 -4390 31410 -4270
rect 31465 -4390 31585 -4270
rect 31630 -4390 31750 -4270
rect 31795 -4390 31915 -4270
rect 31960 -4390 32080 -4270
rect 32135 -4390 32255 -4270
rect 32300 -4390 32420 -4270
rect 32465 -4390 32585 -4270
rect 32630 -4390 32750 -4270
rect 32805 -4390 32925 -4270
rect 32970 -4390 33090 -4270
rect 33135 -4390 33255 -4270
rect 33300 -4390 33420 -4270
rect 33475 -4390 33595 -4270
rect 33640 -4390 33760 -4270
rect 33805 -4390 33925 -4270
rect 33970 -4390 34090 -4270
rect 34145 -4390 34265 -4270
rect 34310 -4390 34430 -4270
rect 34475 -4390 34595 -4270
rect 34640 -4390 34760 -4270
rect 34815 -4390 34935 -4270
rect 34980 -4390 35100 -4270
rect 35145 -4390 35265 -4270
rect 35310 -4390 35430 -4270
rect 35485 -4390 35605 -4270
rect 35650 -4390 35770 -4270
rect 35815 -4390 35935 -4270
rect 35980 -4390 36100 -4270
rect 36155 -4390 36275 -4270
rect 30795 -4565 30915 -4445
rect 30960 -4565 31080 -4445
rect 31125 -4565 31245 -4445
rect 31290 -4565 31410 -4445
rect 31465 -4565 31585 -4445
rect 31630 -4565 31750 -4445
rect 31795 -4565 31915 -4445
rect 31960 -4565 32080 -4445
rect 32135 -4565 32255 -4445
rect 32300 -4565 32420 -4445
rect 32465 -4565 32585 -4445
rect 32630 -4565 32750 -4445
rect 32805 -4565 32925 -4445
rect 32970 -4565 33090 -4445
rect 33135 -4565 33255 -4445
rect 33300 -4565 33420 -4445
rect 33475 -4565 33595 -4445
rect 33640 -4565 33760 -4445
rect 33805 -4565 33925 -4445
rect 33970 -4565 34090 -4445
rect 34145 -4565 34265 -4445
rect 34310 -4565 34430 -4445
rect 34475 -4565 34595 -4445
rect 34640 -4565 34760 -4445
rect 34815 -4565 34935 -4445
rect 34980 -4565 35100 -4445
rect 35145 -4565 35265 -4445
rect 35310 -4565 35430 -4445
rect 35485 -4565 35605 -4445
rect 35650 -4565 35770 -4445
rect 35815 -4565 35935 -4445
rect 35980 -4565 36100 -4445
rect 36155 -4565 36275 -4445
rect 30795 -4730 30915 -4610
rect 30960 -4730 31080 -4610
rect 31125 -4730 31245 -4610
rect 31290 -4730 31410 -4610
rect 31465 -4730 31585 -4610
rect 31630 -4730 31750 -4610
rect 31795 -4730 31915 -4610
rect 31960 -4730 32080 -4610
rect 32135 -4730 32255 -4610
rect 32300 -4730 32420 -4610
rect 32465 -4730 32585 -4610
rect 32630 -4730 32750 -4610
rect 32805 -4730 32925 -4610
rect 32970 -4730 33090 -4610
rect 33135 -4730 33255 -4610
rect 33300 -4730 33420 -4610
rect 33475 -4730 33595 -4610
rect 33640 -4730 33760 -4610
rect 33805 -4730 33925 -4610
rect 33970 -4730 34090 -4610
rect 34145 -4730 34265 -4610
rect 34310 -4730 34430 -4610
rect 34475 -4730 34595 -4610
rect 34640 -4730 34760 -4610
rect 34815 -4730 34935 -4610
rect 34980 -4730 35100 -4610
rect 35145 -4730 35265 -4610
rect 35310 -4730 35430 -4610
rect 35485 -4730 35605 -4610
rect 35650 -4730 35770 -4610
rect 35815 -4730 35935 -4610
rect 35980 -4730 36100 -4610
rect 36155 -4730 36275 -4610
rect 30795 -4895 30915 -4775
rect 30960 -4895 31080 -4775
rect 31125 -4895 31245 -4775
rect 31290 -4895 31410 -4775
rect 31465 -4895 31585 -4775
rect 31630 -4895 31750 -4775
rect 31795 -4895 31915 -4775
rect 31960 -4895 32080 -4775
rect 32135 -4895 32255 -4775
rect 32300 -4895 32420 -4775
rect 32465 -4895 32585 -4775
rect 32630 -4895 32750 -4775
rect 32805 -4895 32925 -4775
rect 32970 -4895 33090 -4775
rect 33135 -4895 33255 -4775
rect 33300 -4895 33420 -4775
rect 33475 -4895 33595 -4775
rect 33640 -4895 33760 -4775
rect 33805 -4895 33925 -4775
rect 33970 -4895 34090 -4775
rect 34145 -4895 34265 -4775
rect 34310 -4895 34430 -4775
rect 34475 -4895 34595 -4775
rect 34640 -4895 34760 -4775
rect 34815 -4895 34935 -4775
rect 34980 -4895 35100 -4775
rect 35145 -4895 35265 -4775
rect 35310 -4895 35430 -4775
rect 35485 -4895 35605 -4775
rect 35650 -4895 35770 -4775
rect 35815 -4895 35935 -4775
rect 35980 -4895 36100 -4775
rect 36155 -4895 36275 -4775
rect 30795 -5060 30915 -4940
rect 30960 -5060 31080 -4940
rect 31125 -5060 31245 -4940
rect 31290 -5060 31410 -4940
rect 31465 -5060 31585 -4940
rect 31630 -5060 31750 -4940
rect 31795 -5060 31915 -4940
rect 31960 -5060 32080 -4940
rect 32135 -5060 32255 -4940
rect 32300 -5060 32420 -4940
rect 32465 -5060 32585 -4940
rect 32630 -5060 32750 -4940
rect 32805 -5060 32925 -4940
rect 32970 -5060 33090 -4940
rect 33135 -5060 33255 -4940
rect 33300 -5060 33420 -4940
rect 33475 -5060 33595 -4940
rect 33640 -5060 33760 -4940
rect 33805 -5060 33925 -4940
rect 33970 -5060 34090 -4940
rect 34145 -5060 34265 -4940
rect 34310 -5060 34430 -4940
rect 34475 -5060 34595 -4940
rect 34640 -5060 34760 -4940
rect 34815 -5060 34935 -4940
rect 34980 -5060 35100 -4940
rect 35145 -5060 35265 -4940
rect 35310 -5060 35430 -4940
rect 35485 -5060 35605 -4940
rect 35650 -5060 35770 -4940
rect 35815 -5060 35935 -4940
rect 35980 -5060 36100 -4940
rect 36155 -5060 36275 -4940
rect 30795 -5235 30915 -5115
rect 30960 -5235 31080 -5115
rect 31125 -5235 31245 -5115
rect 31290 -5235 31410 -5115
rect 31465 -5235 31585 -5115
rect 31630 -5235 31750 -5115
rect 31795 -5235 31915 -5115
rect 31960 -5235 32080 -5115
rect 32135 -5235 32255 -5115
rect 32300 -5235 32420 -5115
rect 32465 -5235 32585 -5115
rect 32630 -5235 32750 -5115
rect 32805 -5235 32925 -5115
rect 32970 -5235 33090 -5115
rect 33135 -5235 33255 -5115
rect 33300 -5235 33420 -5115
rect 33475 -5235 33595 -5115
rect 33640 -5235 33760 -5115
rect 33805 -5235 33925 -5115
rect 33970 -5235 34090 -5115
rect 34145 -5235 34265 -5115
rect 34310 -5235 34430 -5115
rect 34475 -5235 34595 -5115
rect 34640 -5235 34760 -5115
rect 34815 -5235 34935 -5115
rect 34980 -5235 35100 -5115
rect 35145 -5235 35265 -5115
rect 35310 -5235 35430 -5115
rect 35485 -5235 35605 -5115
rect 35650 -5235 35770 -5115
rect 35815 -5235 35935 -5115
rect 35980 -5235 36100 -5115
rect 36155 -5235 36275 -5115
rect 30795 -5400 30915 -5280
rect 30960 -5400 31080 -5280
rect 31125 -5400 31245 -5280
rect 31290 -5400 31410 -5280
rect 31465 -5400 31585 -5280
rect 31630 -5400 31750 -5280
rect 31795 -5400 31915 -5280
rect 31960 -5400 32080 -5280
rect 32135 -5400 32255 -5280
rect 32300 -5400 32420 -5280
rect 32465 -5400 32585 -5280
rect 32630 -5400 32750 -5280
rect 32805 -5400 32925 -5280
rect 32970 -5400 33090 -5280
rect 33135 -5400 33255 -5280
rect 33300 -5400 33420 -5280
rect 33475 -5400 33595 -5280
rect 33640 -5400 33760 -5280
rect 33805 -5400 33925 -5280
rect 33970 -5400 34090 -5280
rect 34145 -5400 34265 -5280
rect 34310 -5400 34430 -5280
rect 34475 -5400 34595 -5280
rect 34640 -5400 34760 -5280
rect 34815 -5400 34935 -5280
rect 34980 -5400 35100 -5280
rect 35145 -5400 35265 -5280
rect 35310 -5400 35430 -5280
rect 35485 -5400 35605 -5280
rect 35650 -5400 35770 -5280
rect 35815 -5400 35935 -5280
rect 35980 -5400 36100 -5280
rect 36155 -5400 36275 -5280
rect 30795 -5565 30915 -5445
rect 30960 -5565 31080 -5445
rect 31125 -5565 31245 -5445
rect 31290 -5565 31410 -5445
rect 31465 -5565 31585 -5445
rect 31630 -5565 31750 -5445
rect 31795 -5565 31915 -5445
rect 31960 -5565 32080 -5445
rect 32135 -5565 32255 -5445
rect 32300 -5565 32420 -5445
rect 32465 -5565 32585 -5445
rect 32630 -5565 32750 -5445
rect 32805 -5565 32925 -5445
rect 32970 -5565 33090 -5445
rect 33135 -5565 33255 -5445
rect 33300 -5565 33420 -5445
rect 33475 -5565 33595 -5445
rect 33640 -5565 33760 -5445
rect 33805 -5565 33925 -5445
rect 33970 -5565 34090 -5445
rect 34145 -5565 34265 -5445
rect 34310 -5565 34430 -5445
rect 34475 -5565 34595 -5445
rect 34640 -5565 34760 -5445
rect 34815 -5565 34935 -5445
rect 34980 -5565 35100 -5445
rect 35145 -5565 35265 -5445
rect 35310 -5565 35430 -5445
rect 35485 -5565 35605 -5445
rect 35650 -5565 35770 -5445
rect 35815 -5565 35935 -5445
rect 35980 -5565 36100 -5445
rect 36155 -5565 36275 -5445
rect 30795 -5730 30915 -5610
rect 30960 -5730 31080 -5610
rect 31125 -5730 31245 -5610
rect 31290 -5730 31410 -5610
rect 31465 -5730 31585 -5610
rect 31630 -5730 31750 -5610
rect 31795 -5730 31915 -5610
rect 31960 -5730 32080 -5610
rect 32135 -5730 32255 -5610
rect 32300 -5730 32420 -5610
rect 32465 -5730 32585 -5610
rect 32630 -5730 32750 -5610
rect 32805 -5730 32925 -5610
rect 32970 -5730 33090 -5610
rect 33135 -5730 33255 -5610
rect 33300 -5730 33420 -5610
rect 33475 -5730 33595 -5610
rect 33640 -5730 33760 -5610
rect 33805 -5730 33925 -5610
rect 33970 -5730 34090 -5610
rect 34145 -5730 34265 -5610
rect 34310 -5730 34430 -5610
rect 34475 -5730 34595 -5610
rect 34640 -5730 34760 -5610
rect 34815 -5730 34935 -5610
rect 34980 -5730 35100 -5610
rect 35145 -5730 35265 -5610
rect 35310 -5730 35430 -5610
rect 35485 -5730 35605 -5610
rect 35650 -5730 35770 -5610
rect 35815 -5730 35935 -5610
rect 35980 -5730 36100 -5610
rect 36155 -5730 36275 -5610
rect 30795 -5905 30915 -5785
rect 30960 -5905 31080 -5785
rect 31125 -5905 31245 -5785
rect 31290 -5905 31410 -5785
rect 31465 -5905 31585 -5785
rect 31630 -5905 31750 -5785
rect 31795 -5905 31915 -5785
rect 31960 -5905 32080 -5785
rect 32135 -5905 32255 -5785
rect 32300 -5905 32420 -5785
rect 32465 -5905 32585 -5785
rect 32630 -5905 32750 -5785
rect 32805 -5905 32925 -5785
rect 32970 -5905 33090 -5785
rect 33135 -5905 33255 -5785
rect 33300 -5905 33420 -5785
rect 33475 -5905 33595 -5785
rect 33640 -5905 33760 -5785
rect 33805 -5905 33925 -5785
rect 33970 -5905 34090 -5785
rect 34145 -5905 34265 -5785
rect 34310 -5905 34430 -5785
rect 34475 -5905 34595 -5785
rect 34640 -5905 34760 -5785
rect 34815 -5905 34935 -5785
rect 34980 -5905 35100 -5785
rect 35145 -5905 35265 -5785
rect 35310 -5905 35430 -5785
rect 35485 -5905 35605 -5785
rect 35650 -5905 35770 -5785
rect 35815 -5905 35935 -5785
rect 35980 -5905 36100 -5785
rect 36155 -5905 36275 -5785
rect 30795 -6070 30915 -5950
rect 30960 -6070 31080 -5950
rect 31125 -6070 31245 -5950
rect 31290 -6070 31410 -5950
rect 31465 -6070 31585 -5950
rect 31630 -6070 31750 -5950
rect 31795 -6070 31915 -5950
rect 31960 -6070 32080 -5950
rect 32135 -6070 32255 -5950
rect 32300 -6070 32420 -5950
rect 32465 -6070 32585 -5950
rect 32630 -6070 32750 -5950
rect 32805 -6070 32925 -5950
rect 32970 -6070 33090 -5950
rect 33135 -6070 33255 -5950
rect 33300 -6070 33420 -5950
rect 33475 -6070 33595 -5950
rect 33640 -6070 33760 -5950
rect 33805 -6070 33925 -5950
rect 33970 -6070 34090 -5950
rect 34145 -6070 34265 -5950
rect 34310 -6070 34430 -5950
rect 34475 -6070 34595 -5950
rect 34640 -6070 34760 -5950
rect 34815 -6070 34935 -5950
rect 34980 -6070 35100 -5950
rect 35145 -6070 35265 -5950
rect 35310 -6070 35430 -5950
rect 35485 -6070 35605 -5950
rect 35650 -6070 35770 -5950
rect 35815 -6070 35935 -5950
rect 35980 -6070 36100 -5950
rect 36155 -6070 36275 -5950
rect 30795 -6235 30915 -6115
rect 30960 -6235 31080 -6115
rect 31125 -6235 31245 -6115
rect 31290 -6235 31410 -6115
rect 31465 -6235 31585 -6115
rect 31630 -6235 31750 -6115
rect 31795 -6235 31915 -6115
rect 31960 -6235 32080 -6115
rect 32135 -6235 32255 -6115
rect 32300 -6235 32420 -6115
rect 32465 -6235 32585 -6115
rect 32630 -6235 32750 -6115
rect 32805 -6235 32925 -6115
rect 32970 -6235 33090 -6115
rect 33135 -6235 33255 -6115
rect 33300 -6235 33420 -6115
rect 33475 -6235 33595 -6115
rect 33640 -6235 33760 -6115
rect 33805 -6235 33925 -6115
rect 33970 -6235 34090 -6115
rect 34145 -6235 34265 -6115
rect 34310 -6235 34430 -6115
rect 34475 -6235 34595 -6115
rect 34640 -6235 34760 -6115
rect 34815 -6235 34935 -6115
rect 34980 -6235 35100 -6115
rect 35145 -6235 35265 -6115
rect 35310 -6235 35430 -6115
rect 35485 -6235 35605 -6115
rect 35650 -6235 35770 -6115
rect 35815 -6235 35935 -6115
rect 35980 -6235 36100 -6115
rect 36155 -6235 36275 -6115
rect 30795 -6400 30915 -6280
rect 30960 -6400 31080 -6280
rect 31125 -6400 31245 -6280
rect 31290 -6400 31410 -6280
rect 31465 -6400 31585 -6280
rect 31630 -6400 31750 -6280
rect 31795 -6400 31915 -6280
rect 31960 -6400 32080 -6280
rect 32135 -6400 32255 -6280
rect 32300 -6400 32420 -6280
rect 32465 -6400 32585 -6280
rect 32630 -6400 32750 -6280
rect 32805 -6400 32925 -6280
rect 32970 -6400 33090 -6280
rect 33135 -6400 33255 -6280
rect 33300 -6400 33420 -6280
rect 33475 -6400 33595 -6280
rect 33640 -6400 33760 -6280
rect 33805 -6400 33925 -6280
rect 33970 -6400 34090 -6280
rect 34145 -6400 34265 -6280
rect 34310 -6400 34430 -6280
rect 34475 -6400 34595 -6280
rect 34640 -6400 34760 -6280
rect 34815 -6400 34935 -6280
rect 34980 -6400 35100 -6280
rect 35145 -6400 35265 -6280
rect 35310 -6400 35430 -6280
rect 35485 -6400 35605 -6280
rect 35650 -6400 35770 -6280
rect 35815 -6400 35935 -6280
rect 35980 -6400 36100 -6280
rect 36155 -6400 36275 -6280
rect 30795 -6575 30915 -6455
rect 30960 -6575 31080 -6455
rect 31125 -6575 31245 -6455
rect 31290 -6575 31410 -6455
rect 31465 -6575 31585 -6455
rect 31630 -6575 31750 -6455
rect 31795 -6575 31915 -6455
rect 31960 -6575 32080 -6455
rect 32135 -6575 32255 -6455
rect 32300 -6575 32420 -6455
rect 32465 -6575 32585 -6455
rect 32630 -6575 32750 -6455
rect 32805 -6575 32925 -6455
rect 32970 -6575 33090 -6455
rect 33135 -6575 33255 -6455
rect 33300 -6575 33420 -6455
rect 33475 -6575 33595 -6455
rect 33640 -6575 33760 -6455
rect 33805 -6575 33925 -6455
rect 33970 -6575 34090 -6455
rect 34145 -6575 34265 -6455
rect 34310 -6575 34430 -6455
rect 34475 -6575 34595 -6455
rect 34640 -6575 34760 -6455
rect 34815 -6575 34935 -6455
rect 34980 -6575 35100 -6455
rect 35145 -6575 35265 -6455
rect 35310 -6575 35430 -6455
rect 35485 -6575 35605 -6455
rect 35650 -6575 35770 -6455
rect 35815 -6575 35935 -6455
rect 35980 -6575 36100 -6455
rect 36155 -6575 36275 -6455
rect 30795 -6740 30915 -6620
rect 30960 -6740 31080 -6620
rect 31125 -6740 31245 -6620
rect 31290 -6740 31410 -6620
rect 31465 -6740 31585 -6620
rect 31630 -6740 31750 -6620
rect 31795 -6740 31915 -6620
rect 31960 -6740 32080 -6620
rect 32135 -6740 32255 -6620
rect 32300 -6740 32420 -6620
rect 32465 -6740 32585 -6620
rect 32630 -6740 32750 -6620
rect 32805 -6740 32925 -6620
rect 32970 -6740 33090 -6620
rect 33135 -6740 33255 -6620
rect 33300 -6740 33420 -6620
rect 33475 -6740 33595 -6620
rect 33640 -6740 33760 -6620
rect 33805 -6740 33925 -6620
rect 33970 -6740 34090 -6620
rect 34145 -6740 34265 -6620
rect 34310 -6740 34430 -6620
rect 34475 -6740 34595 -6620
rect 34640 -6740 34760 -6620
rect 34815 -6740 34935 -6620
rect 34980 -6740 35100 -6620
rect 35145 -6740 35265 -6620
rect 35310 -6740 35430 -6620
rect 35485 -6740 35605 -6620
rect 35650 -6740 35770 -6620
rect 35815 -6740 35935 -6620
rect 35980 -6740 36100 -6620
rect 36155 -6740 36275 -6620
rect 30795 -6905 30915 -6785
rect 30960 -6905 31080 -6785
rect 31125 -6905 31245 -6785
rect 31290 -6905 31410 -6785
rect 31465 -6905 31585 -6785
rect 31630 -6905 31750 -6785
rect 31795 -6905 31915 -6785
rect 31960 -6905 32080 -6785
rect 32135 -6905 32255 -6785
rect 32300 -6905 32420 -6785
rect 32465 -6905 32585 -6785
rect 32630 -6905 32750 -6785
rect 32805 -6905 32925 -6785
rect 32970 -6905 33090 -6785
rect 33135 -6905 33255 -6785
rect 33300 -6905 33420 -6785
rect 33475 -6905 33595 -6785
rect 33640 -6905 33760 -6785
rect 33805 -6905 33925 -6785
rect 33970 -6905 34090 -6785
rect 34145 -6905 34265 -6785
rect 34310 -6905 34430 -6785
rect 34475 -6905 34595 -6785
rect 34640 -6905 34760 -6785
rect 34815 -6905 34935 -6785
rect 34980 -6905 35100 -6785
rect 35145 -6905 35265 -6785
rect 35310 -6905 35430 -6785
rect 35485 -6905 35605 -6785
rect 35650 -6905 35770 -6785
rect 35815 -6905 35935 -6785
rect 35980 -6905 36100 -6785
rect 36155 -6905 36275 -6785
rect 30795 -7070 30915 -6950
rect 30960 -7070 31080 -6950
rect 31125 -7070 31245 -6950
rect 31290 -7070 31410 -6950
rect 31465 -7070 31585 -6950
rect 31630 -7070 31750 -6950
rect 31795 -7070 31915 -6950
rect 31960 -7070 32080 -6950
rect 32135 -7070 32255 -6950
rect 32300 -7070 32420 -6950
rect 32465 -7070 32585 -6950
rect 32630 -7070 32750 -6950
rect 32805 -7070 32925 -6950
rect 32970 -7070 33090 -6950
rect 33135 -7070 33255 -6950
rect 33300 -7070 33420 -6950
rect 33475 -7070 33595 -6950
rect 33640 -7070 33760 -6950
rect 33805 -7070 33925 -6950
rect 33970 -7070 34090 -6950
rect 34145 -7070 34265 -6950
rect 34310 -7070 34430 -6950
rect 34475 -7070 34595 -6950
rect 34640 -7070 34760 -6950
rect 34815 -7070 34935 -6950
rect 34980 -7070 35100 -6950
rect 35145 -7070 35265 -6950
rect 35310 -7070 35430 -6950
rect 35485 -7070 35605 -6950
rect 35650 -7070 35770 -6950
rect 35815 -7070 35935 -6950
rect 35980 -7070 36100 -6950
rect 36155 -7070 36275 -6950
rect 30795 -7245 30915 -7125
rect 30960 -7245 31080 -7125
rect 31125 -7245 31245 -7125
rect 31290 -7245 31410 -7125
rect 31465 -7245 31585 -7125
rect 31630 -7245 31750 -7125
rect 31795 -7245 31915 -7125
rect 31960 -7245 32080 -7125
rect 32135 -7245 32255 -7125
rect 32300 -7245 32420 -7125
rect 32465 -7245 32585 -7125
rect 32630 -7245 32750 -7125
rect 32805 -7245 32925 -7125
rect 32970 -7245 33090 -7125
rect 33135 -7245 33255 -7125
rect 33300 -7245 33420 -7125
rect 33475 -7245 33595 -7125
rect 33640 -7245 33760 -7125
rect 33805 -7245 33925 -7125
rect 33970 -7245 34090 -7125
rect 34145 -7245 34265 -7125
rect 34310 -7245 34430 -7125
rect 34475 -7245 34595 -7125
rect 34640 -7245 34760 -7125
rect 34815 -7245 34935 -7125
rect 34980 -7245 35100 -7125
rect 35145 -7245 35265 -7125
rect 35310 -7245 35430 -7125
rect 35485 -7245 35605 -7125
rect 35650 -7245 35770 -7125
rect 35815 -7245 35935 -7125
rect 35980 -7245 36100 -7125
rect 36155 -7245 36275 -7125
rect 30795 -7410 30915 -7290
rect 30960 -7410 31080 -7290
rect 31125 -7410 31245 -7290
rect 31290 -7410 31410 -7290
rect 31465 -7410 31585 -7290
rect 31630 -7410 31750 -7290
rect 31795 -7410 31915 -7290
rect 31960 -7410 32080 -7290
rect 32135 -7410 32255 -7290
rect 32300 -7410 32420 -7290
rect 32465 -7410 32585 -7290
rect 32630 -7410 32750 -7290
rect 32805 -7410 32925 -7290
rect 32970 -7410 33090 -7290
rect 33135 -7410 33255 -7290
rect 33300 -7410 33420 -7290
rect 33475 -7410 33595 -7290
rect 33640 -7410 33760 -7290
rect 33805 -7410 33925 -7290
rect 33970 -7410 34090 -7290
rect 34145 -7410 34265 -7290
rect 34310 -7410 34430 -7290
rect 34475 -7410 34595 -7290
rect 34640 -7410 34760 -7290
rect 34815 -7410 34935 -7290
rect 34980 -7410 35100 -7290
rect 35145 -7410 35265 -7290
rect 35310 -7410 35430 -7290
rect 35485 -7410 35605 -7290
rect 35650 -7410 35770 -7290
rect 35815 -7410 35935 -7290
rect 35980 -7410 36100 -7290
rect 36155 -7410 36275 -7290
rect 30795 -7575 30915 -7455
rect 30960 -7575 31080 -7455
rect 31125 -7575 31245 -7455
rect 31290 -7575 31410 -7455
rect 31465 -7575 31585 -7455
rect 31630 -7575 31750 -7455
rect 31795 -7575 31915 -7455
rect 31960 -7575 32080 -7455
rect 32135 -7575 32255 -7455
rect 32300 -7575 32420 -7455
rect 32465 -7575 32585 -7455
rect 32630 -7575 32750 -7455
rect 32805 -7575 32925 -7455
rect 32970 -7575 33090 -7455
rect 33135 -7575 33255 -7455
rect 33300 -7575 33420 -7455
rect 33475 -7575 33595 -7455
rect 33640 -7575 33760 -7455
rect 33805 -7575 33925 -7455
rect 33970 -7575 34090 -7455
rect 34145 -7575 34265 -7455
rect 34310 -7575 34430 -7455
rect 34475 -7575 34595 -7455
rect 34640 -7575 34760 -7455
rect 34815 -7575 34935 -7455
rect 34980 -7575 35100 -7455
rect 35145 -7575 35265 -7455
rect 35310 -7575 35430 -7455
rect 35485 -7575 35605 -7455
rect 35650 -7575 35770 -7455
rect 35815 -7575 35935 -7455
rect 35980 -7575 36100 -7455
rect 36155 -7575 36275 -7455
rect 30795 -7740 30915 -7620
rect 30960 -7740 31080 -7620
rect 31125 -7740 31245 -7620
rect 31290 -7740 31410 -7620
rect 31465 -7740 31585 -7620
rect 31630 -7740 31750 -7620
rect 31795 -7740 31915 -7620
rect 31960 -7740 32080 -7620
rect 32135 -7740 32255 -7620
rect 32300 -7740 32420 -7620
rect 32465 -7740 32585 -7620
rect 32630 -7740 32750 -7620
rect 32805 -7740 32925 -7620
rect 32970 -7740 33090 -7620
rect 33135 -7740 33255 -7620
rect 33300 -7740 33420 -7620
rect 33475 -7740 33595 -7620
rect 33640 -7740 33760 -7620
rect 33805 -7740 33925 -7620
rect 33970 -7740 34090 -7620
rect 34145 -7740 34265 -7620
rect 34310 -7740 34430 -7620
rect 34475 -7740 34595 -7620
rect 34640 -7740 34760 -7620
rect 34815 -7740 34935 -7620
rect 34980 -7740 35100 -7620
rect 35145 -7740 35265 -7620
rect 35310 -7740 35430 -7620
rect 35485 -7740 35605 -7620
rect 35650 -7740 35770 -7620
rect 35815 -7740 35935 -7620
rect 35980 -7740 36100 -7620
rect 36155 -7740 36275 -7620
rect 30795 -7915 30915 -7795
rect 30960 -7915 31080 -7795
rect 31125 -7915 31245 -7795
rect 31290 -7915 31410 -7795
rect 31465 -7915 31585 -7795
rect 31630 -7915 31750 -7795
rect 31795 -7915 31915 -7795
rect 31960 -7915 32080 -7795
rect 32135 -7915 32255 -7795
rect 32300 -7915 32420 -7795
rect 32465 -7915 32585 -7795
rect 32630 -7915 32750 -7795
rect 32805 -7915 32925 -7795
rect 32970 -7915 33090 -7795
rect 33135 -7915 33255 -7795
rect 33300 -7915 33420 -7795
rect 33475 -7915 33595 -7795
rect 33640 -7915 33760 -7795
rect 33805 -7915 33925 -7795
rect 33970 -7915 34090 -7795
rect 34145 -7915 34265 -7795
rect 34310 -7915 34430 -7795
rect 34475 -7915 34595 -7795
rect 34640 -7915 34760 -7795
rect 34815 -7915 34935 -7795
rect 34980 -7915 35100 -7795
rect 35145 -7915 35265 -7795
rect 35310 -7915 35430 -7795
rect 35485 -7915 35605 -7795
rect 35650 -7915 35770 -7795
rect 35815 -7915 35935 -7795
rect 35980 -7915 36100 -7795
rect 36155 -7915 36275 -7795
rect 30795 -8080 30915 -7960
rect 30960 -8080 31080 -7960
rect 31125 -8080 31245 -7960
rect 31290 -8080 31410 -7960
rect 31465 -8080 31585 -7960
rect 31630 -8080 31750 -7960
rect 31795 -8080 31915 -7960
rect 31960 -8080 32080 -7960
rect 32135 -8080 32255 -7960
rect 32300 -8080 32420 -7960
rect 32465 -8080 32585 -7960
rect 32630 -8080 32750 -7960
rect 32805 -8080 32925 -7960
rect 32970 -8080 33090 -7960
rect 33135 -8080 33255 -7960
rect 33300 -8080 33420 -7960
rect 33475 -8080 33595 -7960
rect 33640 -8080 33760 -7960
rect 33805 -8080 33925 -7960
rect 33970 -8080 34090 -7960
rect 34145 -8080 34265 -7960
rect 34310 -8080 34430 -7960
rect 34475 -8080 34595 -7960
rect 34640 -8080 34760 -7960
rect 34815 -8080 34935 -7960
rect 34980 -8080 35100 -7960
rect 35145 -8080 35265 -7960
rect 35310 -8080 35430 -7960
rect 35485 -8080 35605 -7960
rect 35650 -8080 35770 -7960
rect 35815 -8080 35935 -7960
rect 35980 -8080 36100 -7960
rect 36155 -8080 36275 -7960
rect 30795 -8245 30915 -8125
rect 30960 -8245 31080 -8125
rect 31125 -8245 31245 -8125
rect 31290 -8245 31410 -8125
rect 31465 -8245 31585 -8125
rect 31630 -8245 31750 -8125
rect 31795 -8245 31915 -8125
rect 31960 -8245 32080 -8125
rect 32135 -8245 32255 -8125
rect 32300 -8245 32420 -8125
rect 32465 -8245 32585 -8125
rect 32630 -8245 32750 -8125
rect 32805 -8245 32925 -8125
rect 32970 -8245 33090 -8125
rect 33135 -8245 33255 -8125
rect 33300 -8245 33420 -8125
rect 33475 -8245 33595 -8125
rect 33640 -8245 33760 -8125
rect 33805 -8245 33925 -8125
rect 33970 -8245 34090 -8125
rect 34145 -8245 34265 -8125
rect 34310 -8245 34430 -8125
rect 34475 -8245 34595 -8125
rect 34640 -8245 34760 -8125
rect 34815 -8245 34935 -8125
rect 34980 -8245 35100 -8125
rect 35145 -8245 35265 -8125
rect 35310 -8245 35430 -8125
rect 35485 -8245 35605 -8125
rect 35650 -8245 35770 -8125
rect 35815 -8245 35935 -8125
rect 35980 -8245 36100 -8125
rect 36155 -8245 36275 -8125
rect 30795 -8410 30915 -8290
rect 30960 -8410 31080 -8290
rect 31125 -8410 31245 -8290
rect 31290 -8410 31410 -8290
rect 31465 -8410 31585 -8290
rect 31630 -8410 31750 -8290
rect 31795 -8410 31915 -8290
rect 31960 -8410 32080 -8290
rect 32135 -8410 32255 -8290
rect 32300 -8410 32420 -8290
rect 32465 -8410 32585 -8290
rect 32630 -8410 32750 -8290
rect 32805 -8410 32925 -8290
rect 32970 -8410 33090 -8290
rect 33135 -8410 33255 -8290
rect 33300 -8410 33420 -8290
rect 33475 -8410 33595 -8290
rect 33640 -8410 33760 -8290
rect 33805 -8410 33925 -8290
rect 33970 -8410 34090 -8290
rect 34145 -8410 34265 -8290
rect 34310 -8410 34430 -8290
rect 34475 -8410 34595 -8290
rect 34640 -8410 34760 -8290
rect 34815 -8410 34935 -8290
rect 34980 -8410 35100 -8290
rect 35145 -8410 35265 -8290
rect 35310 -8410 35430 -8290
rect 35485 -8410 35605 -8290
rect 35650 -8410 35770 -8290
rect 35815 -8410 35935 -8290
rect 35980 -8410 36100 -8290
rect 36155 -8410 36275 -8290
rect 30795 -8585 30915 -8465
rect 30960 -8585 31080 -8465
rect 31125 -8585 31245 -8465
rect 31290 -8585 31410 -8465
rect 31465 -8585 31585 -8465
rect 31630 -8585 31750 -8465
rect 31795 -8585 31915 -8465
rect 31960 -8585 32080 -8465
rect 32135 -8585 32255 -8465
rect 32300 -8585 32420 -8465
rect 32465 -8585 32585 -8465
rect 32630 -8585 32750 -8465
rect 32805 -8585 32925 -8465
rect 32970 -8585 33090 -8465
rect 33135 -8585 33255 -8465
rect 33300 -8585 33420 -8465
rect 33475 -8585 33595 -8465
rect 33640 -8585 33760 -8465
rect 33805 -8585 33925 -8465
rect 33970 -8585 34090 -8465
rect 34145 -8585 34265 -8465
rect 34310 -8585 34430 -8465
rect 34475 -8585 34595 -8465
rect 34640 -8585 34760 -8465
rect 34815 -8585 34935 -8465
rect 34980 -8585 35100 -8465
rect 35145 -8585 35265 -8465
rect 35310 -8585 35430 -8465
rect 35485 -8585 35605 -8465
rect 35650 -8585 35770 -8465
rect 35815 -8585 35935 -8465
rect 35980 -8585 36100 -8465
rect 36155 -8585 36275 -8465
rect 30795 -8750 30915 -8630
rect 30960 -8750 31080 -8630
rect 31125 -8750 31245 -8630
rect 31290 -8750 31410 -8630
rect 31465 -8750 31585 -8630
rect 31630 -8750 31750 -8630
rect 31795 -8750 31915 -8630
rect 31960 -8750 32080 -8630
rect 32135 -8750 32255 -8630
rect 32300 -8750 32420 -8630
rect 32465 -8750 32585 -8630
rect 32630 -8750 32750 -8630
rect 32805 -8750 32925 -8630
rect 32970 -8750 33090 -8630
rect 33135 -8750 33255 -8630
rect 33300 -8750 33420 -8630
rect 33475 -8750 33595 -8630
rect 33640 -8750 33760 -8630
rect 33805 -8750 33925 -8630
rect 33970 -8750 34090 -8630
rect 34145 -8750 34265 -8630
rect 34310 -8750 34430 -8630
rect 34475 -8750 34595 -8630
rect 34640 -8750 34760 -8630
rect 34815 -8750 34935 -8630
rect 34980 -8750 35100 -8630
rect 35145 -8750 35265 -8630
rect 35310 -8750 35430 -8630
rect 35485 -8750 35605 -8630
rect 35650 -8750 35770 -8630
rect 35815 -8750 35935 -8630
rect 35980 -8750 36100 -8630
rect 36155 -8750 36275 -8630
rect 30795 -8915 30915 -8795
rect 30960 -8915 31080 -8795
rect 31125 -8915 31245 -8795
rect 31290 -8915 31410 -8795
rect 31465 -8915 31585 -8795
rect 31630 -8915 31750 -8795
rect 31795 -8915 31915 -8795
rect 31960 -8915 32080 -8795
rect 32135 -8915 32255 -8795
rect 32300 -8915 32420 -8795
rect 32465 -8915 32585 -8795
rect 32630 -8915 32750 -8795
rect 32805 -8915 32925 -8795
rect 32970 -8915 33090 -8795
rect 33135 -8915 33255 -8795
rect 33300 -8915 33420 -8795
rect 33475 -8915 33595 -8795
rect 33640 -8915 33760 -8795
rect 33805 -8915 33925 -8795
rect 33970 -8915 34090 -8795
rect 34145 -8915 34265 -8795
rect 34310 -8915 34430 -8795
rect 34475 -8915 34595 -8795
rect 34640 -8915 34760 -8795
rect 34815 -8915 34935 -8795
rect 34980 -8915 35100 -8795
rect 35145 -8915 35265 -8795
rect 35310 -8915 35430 -8795
rect 35485 -8915 35605 -8795
rect 35650 -8915 35770 -8795
rect 35815 -8915 35935 -8795
rect 35980 -8915 36100 -8795
rect 36155 -8915 36275 -8795
rect 30795 -9080 30915 -8960
rect 30960 -9080 31080 -8960
rect 31125 -9080 31245 -8960
rect 31290 -9080 31410 -8960
rect 31465 -9080 31585 -8960
rect 31630 -9080 31750 -8960
rect 31795 -9080 31915 -8960
rect 31960 -9080 32080 -8960
rect 32135 -9080 32255 -8960
rect 32300 -9080 32420 -8960
rect 32465 -9080 32585 -8960
rect 32630 -9080 32750 -8960
rect 32805 -9080 32925 -8960
rect 32970 -9080 33090 -8960
rect 33135 -9080 33255 -8960
rect 33300 -9080 33420 -8960
rect 33475 -9080 33595 -8960
rect 33640 -9080 33760 -8960
rect 33805 -9080 33925 -8960
rect 33970 -9080 34090 -8960
rect 34145 -9080 34265 -8960
rect 34310 -9080 34430 -8960
rect 34475 -9080 34595 -8960
rect 34640 -9080 34760 -8960
rect 34815 -9080 34935 -8960
rect 34980 -9080 35100 -8960
rect 35145 -9080 35265 -8960
rect 35310 -9080 35430 -8960
rect 35485 -9080 35605 -8960
rect 35650 -9080 35770 -8960
rect 35815 -9080 35935 -8960
rect 35980 -9080 36100 -8960
rect 36155 -9080 36275 -8960
rect 30795 -9255 30915 -9135
rect 30960 -9255 31080 -9135
rect 31125 -9255 31245 -9135
rect 31290 -9255 31410 -9135
rect 31465 -9255 31585 -9135
rect 31630 -9255 31750 -9135
rect 31795 -9255 31915 -9135
rect 31960 -9255 32080 -9135
rect 32135 -9255 32255 -9135
rect 32300 -9255 32420 -9135
rect 32465 -9255 32585 -9135
rect 32630 -9255 32750 -9135
rect 32805 -9255 32925 -9135
rect 32970 -9255 33090 -9135
rect 33135 -9255 33255 -9135
rect 33300 -9255 33420 -9135
rect 33475 -9255 33595 -9135
rect 33640 -9255 33760 -9135
rect 33805 -9255 33925 -9135
rect 33970 -9255 34090 -9135
rect 34145 -9255 34265 -9135
rect 34310 -9255 34430 -9135
rect 34475 -9255 34595 -9135
rect 34640 -9255 34760 -9135
rect 34815 -9255 34935 -9135
rect 34980 -9255 35100 -9135
rect 35145 -9255 35265 -9135
rect 35310 -9255 35430 -9135
rect 35485 -9255 35605 -9135
rect 35650 -9255 35770 -9135
rect 35815 -9255 35935 -9135
rect 35980 -9255 36100 -9135
rect 36155 -9255 36275 -9135
rect 30795 -9420 30915 -9300
rect 30960 -9420 31080 -9300
rect 31125 -9420 31245 -9300
rect 31290 -9420 31410 -9300
rect 31465 -9420 31585 -9300
rect 31630 -9420 31750 -9300
rect 31795 -9420 31915 -9300
rect 31960 -9420 32080 -9300
rect 32135 -9420 32255 -9300
rect 32300 -9420 32420 -9300
rect 32465 -9420 32585 -9300
rect 32630 -9420 32750 -9300
rect 32805 -9420 32925 -9300
rect 32970 -9420 33090 -9300
rect 33135 -9420 33255 -9300
rect 33300 -9420 33420 -9300
rect 33475 -9420 33595 -9300
rect 33640 -9420 33760 -9300
rect 33805 -9420 33925 -9300
rect 33970 -9420 34090 -9300
rect 34145 -9420 34265 -9300
rect 34310 -9420 34430 -9300
rect 34475 -9420 34595 -9300
rect 34640 -9420 34760 -9300
rect 34815 -9420 34935 -9300
rect 34980 -9420 35100 -9300
rect 35145 -9420 35265 -9300
rect 35310 -9420 35430 -9300
rect 35485 -9420 35605 -9300
rect 35650 -9420 35770 -9300
rect 35815 -9420 35935 -9300
rect 35980 -9420 36100 -9300
rect 36155 -9420 36275 -9300
rect 30795 -9585 30915 -9465
rect 30960 -9585 31080 -9465
rect 31125 -9585 31245 -9465
rect 31290 -9585 31410 -9465
rect 31465 -9585 31585 -9465
rect 31630 -9585 31750 -9465
rect 31795 -9585 31915 -9465
rect 31960 -9585 32080 -9465
rect 32135 -9585 32255 -9465
rect 32300 -9585 32420 -9465
rect 32465 -9585 32585 -9465
rect 32630 -9585 32750 -9465
rect 32805 -9585 32925 -9465
rect 32970 -9585 33090 -9465
rect 33135 -9585 33255 -9465
rect 33300 -9585 33420 -9465
rect 33475 -9585 33595 -9465
rect 33640 -9585 33760 -9465
rect 33805 -9585 33925 -9465
rect 33970 -9585 34090 -9465
rect 34145 -9585 34265 -9465
rect 34310 -9585 34430 -9465
rect 34475 -9585 34595 -9465
rect 34640 -9585 34760 -9465
rect 34815 -9585 34935 -9465
rect 34980 -9585 35100 -9465
rect 35145 -9585 35265 -9465
rect 35310 -9585 35430 -9465
rect 35485 -9585 35605 -9465
rect 35650 -9585 35770 -9465
rect 35815 -9585 35935 -9465
rect 35980 -9585 36100 -9465
rect 36155 -9585 36275 -9465
rect 30795 -9750 30915 -9630
rect 30960 -9750 31080 -9630
rect 31125 -9750 31245 -9630
rect 31290 -9750 31410 -9630
rect 31465 -9750 31585 -9630
rect 31630 -9750 31750 -9630
rect 31795 -9750 31915 -9630
rect 31960 -9750 32080 -9630
rect 32135 -9750 32255 -9630
rect 32300 -9750 32420 -9630
rect 32465 -9750 32585 -9630
rect 32630 -9750 32750 -9630
rect 32805 -9750 32925 -9630
rect 32970 -9750 33090 -9630
rect 33135 -9750 33255 -9630
rect 33300 -9750 33420 -9630
rect 33475 -9750 33595 -9630
rect 33640 -9750 33760 -9630
rect 33805 -9750 33925 -9630
rect 33970 -9750 34090 -9630
rect 34145 -9750 34265 -9630
rect 34310 -9750 34430 -9630
rect 34475 -9750 34595 -9630
rect 34640 -9750 34760 -9630
rect 34815 -9750 34935 -9630
rect 34980 -9750 35100 -9630
rect 35145 -9750 35265 -9630
rect 35310 -9750 35430 -9630
rect 35485 -9750 35605 -9630
rect 35650 -9750 35770 -9630
rect 35815 -9750 35935 -9630
rect 35980 -9750 36100 -9630
rect 36155 -9750 36275 -9630
rect 36485 -4390 36605 -4270
rect 36650 -4390 36770 -4270
rect 36815 -4390 36935 -4270
rect 36980 -4390 37100 -4270
rect 37155 -4390 37275 -4270
rect 37320 -4390 37440 -4270
rect 37485 -4390 37605 -4270
rect 37650 -4390 37770 -4270
rect 37825 -4390 37945 -4270
rect 37990 -4390 38110 -4270
rect 38155 -4390 38275 -4270
rect 38320 -4390 38440 -4270
rect 38495 -4390 38615 -4270
rect 38660 -4390 38780 -4270
rect 38825 -4390 38945 -4270
rect 38990 -4390 39110 -4270
rect 39165 -4390 39285 -4270
rect 39330 -4390 39450 -4270
rect 39495 -4390 39615 -4270
rect 39660 -4390 39780 -4270
rect 39835 -4390 39955 -4270
rect 40000 -4390 40120 -4270
rect 40165 -4390 40285 -4270
rect 40330 -4390 40450 -4270
rect 40505 -4390 40625 -4270
rect 40670 -4390 40790 -4270
rect 40835 -4390 40955 -4270
rect 41000 -4390 41120 -4270
rect 41175 -4390 41295 -4270
rect 41340 -4390 41460 -4270
rect 41505 -4390 41625 -4270
rect 41670 -4390 41790 -4270
rect 41845 -4390 41965 -4270
rect 36485 -4565 36605 -4445
rect 36650 -4565 36770 -4445
rect 36815 -4565 36935 -4445
rect 36980 -4565 37100 -4445
rect 37155 -4565 37275 -4445
rect 37320 -4565 37440 -4445
rect 37485 -4565 37605 -4445
rect 37650 -4565 37770 -4445
rect 37825 -4565 37945 -4445
rect 37990 -4565 38110 -4445
rect 38155 -4565 38275 -4445
rect 38320 -4565 38440 -4445
rect 38495 -4565 38615 -4445
rect 38660 -4565 38780 -4445
rect 38825 -4565 38945 -4445
rect 38990 -4565 39110 -4445
rect 39165 -4565 39285 -4445
rect 39330 -4565 39450 -4445
rect 39495 -4565 39615 -4445
rect 39660 -4565 39780 -4445
rect 39835 -4565 39955 -4445
rect 40000 -4565 40120 -4445
rect 40165 -4565 40285 -4445
rect 40330 -4565 40450 -4445
rect 40505 -4565 40625 -4445
rect 40670 -4565 40790 -4445
rect 40835 -4565 40955 -4445
rect 41000 -4565 41120 -4445
rect 41175 -4565 41295 -4445
rect 41340 -4565 41460 -4445
rect 41505 -4565 41625 -4445
rect 41670 -4565 41790 -4445
rect 41845 -4565 41965 -4445
rect 36485 -4730 36605 -4610
rect 36650 -4730 36770 -4610
rect 36815 -4730 36935 -4610
rect 36980 -4730 37100 -4610
rect 37155 -4730 37275 -4610
rect 37320 -4730 37440 -4610
rect 37485 -4730 37605 -4610
rect 37650 -4730 37770 -4610
rect 37825 -4730 37945 -4610
rect 37990 -4730 38110 -4610
rect 38155 -4730 38275 -4610
rect 38320 -4730 38440 -4610
rect 38495 -4730 38615 -4610
rect 38660 -4730 38780 -4610
rect 38825 -4730 38945 -4610
rect 38990 -4730 39110 -4610
rect 39165 -4730 39285 -4610
rect 39330 -4730 39450 -4610
rect 39495 -4730 39615 -4610
rect 39660 -4730 39780 -4610
rect 39835 -4730 39955 -4610
rect 40000 -4730 40120 -4610
rect 40165 -4730 40285 -4610
rect 40330 -4730 40450 -4610
rect 40505 -4730 40625 -4610
rect 40670 -4730 40790 -4610
rect 40835 -4730 40955 -4610
rect 41000 -4730 41120 -4610
rect 41175 -4730 41295 -4610
rect 41340 -4730 41460 -4610
rect 41505 -4730 41625 -4610
rect 41670 -4730 41790 -4610
rect 41845 -4730 41965 -4610
rect 36485 -4895 36605 -4775
rect 36650 -4895 36770 -4775
rect 36815 -4895 36935 -4775
rect 36980 -4895 37100 -4775
rect 37155 -4895 37275 -4775
rect 37320 -4895 37440 -4775
rect 37485 -4895 37605 -4775
rect 37650 -4895 37770 -4775
rect 37825 -4895 37945 -4775
rect 37990 -4895 38110 -4775
rect 38155 -4895 38275 -4775
rect 38320 -4895 38440 -4775
rect 38495 -4895 38615 -4775
rect 38660 -4895 38780 -4775
rect 38825 -4895 38945 -4775
rect 38990 -4895 39110 -4775
rect 39165 -4895 39285 -4775
rect 39330 -4895 39450 -4775
rect 39495 -4895 39615 -4775
rect 39660 -4895 39780 -4775
rect 39835 -4895 39955 -4775
rect 40000 -4895 40120 -4775
rect 40165 -4895 40285 -4775
rect 40330 -4895 40450 -4775
rect 40505 -4895 40625 -4775
rect 40670 -4895 40790 -4775
rect 40835 -4895 40955 -4775
rect 41000 -4895 41120 -4775
rect 41175 -4895 41295 -4775
rect 41340 -4895 41460 -4775
rect 41505 -4895 41625 -4775
rect 41670 -4895 41790 -4775
rect 41845 -4895 41965 -4775
rect 36485 -5060 36605 -4940
rect 36650 -5060 36770 -4940
rect 36815 -5060 36935 -4940
rect 36980 -5060 37100 -4940
rect 37155 -5060 37275 -4940
rect 37320 -5060 37440 -4940
rect 37485 -5060 37605 -4940
rect 37650 -5060 37770 -4940
rect 37825 -5060 37945 -4940
rect 37990 -5060 38110 -4940
rect 38155 -5060 38275 -4940
rect 38320 -5060 38440 -4940
rect 38495 -5060 38615 -4940
rect 38660 -5060 38780 -4940
rect 38825 -5060 38945 -4940
rect 38990 -5060 39110 -4940
rect 39165 -5060 39285 -4940
rect 39330 -5060 39450 -4940
rect 39495 -5060 39615 -4940
rect 39660 -5060 39780 -4940
rect 39835 -5060 39955 -4940
rect 40000 -5060 40120 -4940
rect 40165 -5060 40285 -4940
rect 40330 -5060 40450 -4940
rect 40505 -5060 40625 -4940
rect 40670 -5060 40790 -4940
rect 40835 -5060 40955 -4940
rect 41000 -5060 41120 -4940
rect 41175 -5060 41295 -4940
rect 41340 -5060 41460 -4940
rect 41505 -5060 41625 -4940
rect 41670 -5060 41790 -4940
rect 41845 -5060 41965 -4940
rect 36485 -5235 36605 -5115
rect 36650 -5235 36770 -5115
rect 36815 -5235 36935 -5115
rect 36980 -5235 37100 -5115
rect 37155 -5235 37275 -5115
rect 37320 -5235 37440 -5115
rect 37485 -5235 37605 -5115
rect 37650 -5235 37770 -5115
rect 37825 -5235 37945 -5115
rect 37990 -5235 38110 -5115
rect 38155 -5235 38275 -5115
rect 38320 -5235 38440 -5115
rect 38495 -5235 38615 -5115
rect 38660 -5235 38780 -5115
rect 38825 -5235 38945 -5115
rect 38990 -5235 39110 -5115
rect 39165 -5235 39285 -5115
rect 39330 -5235 39450 -5115
rect 39495 -5235 39615 -5115
rect 39660 -5235 39780 -5115
rect 39835 -5235 39955 -5115
rect 40000 -5235 40120 -5115
rect 40165 -5235 40285 -5115
rect 40330 -5235 40450 -5115
rect 40505 -5235 40625 -5115
rect 40670 -5235 40790 -5115
rect 40835 -5235 40955 -5115
rect 41000 -5235 41120 -5115
rect 41175 -5235 41295 -5115
rect 41340 -5235 41460 -5115
rect 41505 -5235 41625 -5115
rect 41670 -5235 41790 -5115
rect 41845 -5235 41965 -5115
rect 36485 -5400 36605 -5280
rect 36650 -5400 36770 -5280
rect 36815 -5400 36935 -5280
rect 36980 -5400 37100 -5280
rect 37155 -5400 37275 -5280
rect 37320 -5400 37440 -5280
rect 37485 -5400 37605 -5280
rect 37650 -5400 37770 -5280
rect 37825 -5400 37945 -5280
rect 37990 -5400 38110 -5280
rect 38155 -5400 38275 -5280
rect 38320 -5400 38440 -5280
rect 38495 -5400 38615 -5280
rect 38660 -5400 38780 -5280
rect 38825 -5400 38945 -5280
rect 38990 -5400 39110 -5280
rect 39165 -5400 39285 -5280
rect 39330 -5400 39450 -5280
rect 39495 -5400 39615 -5280
rect 39660 -5400 39780 -5280
rect 39835 -5400 39955 -5280
rect 40000 -5400 40120 -5280
rect 40165 -5400 40285 -5280
rect 40330 -5400 40450 -5280
rect 40505 -5400 40625 -5280
rect 40670 -5400 40790 -5280
rect 40835 -5400 40955 -5280
rect 41000 -5400 41120 -5280
rect 41175 -5400 41295 -5280
rect 41340 -5400 41460 -5280
rect 41505 -5400 41625 -5280
rect 41670 -5400 41790 -5280
rect 41845 -5400 41965 -5280
rect 36485 -5565 36605 -5445
rect 36650 -5565 36770 -5445
rect 36815 -5565 36935 -5445
rect 36980 -5565 37100 -5445
rect 37155 -5565 37275 -5445
rect 37320 -5565 37440 -5445
rect 37485 -5565 37605 -5445
rect 37650 -5565 37770 -5445
rect 37825 -5565 37945 -5445
rect 37990 -5565 38110 -5445
rect 38155 -5565 38275 -5445
rect 38320 -5565 38440 -5445
rect 38495 -5565 38615 -5445
rect 38660 -5565 38780 -5445
rect 38825 -5565 38945 -5445
rect 38990 -5565 39110 -5445
rect 39165 -5565 39285 -5445
rect 39330 -5565 39450 -5445
rect 39495 -5565 39615 -5445
rect 39660 -5565 39780 -5445
rect 39835 -5565 39955 -5445
rect 40000 -5565 40120 -5445
rect 40165 -5565 40285 -5445
rect 40330 -5565 40450 -5445
rect 40505 -5565 40625 -5445
rect 40670 -5565 40790 -5445
rect 40835 -5565 40955 -5445
rect 41000 -5565 41120 -5445
rect 41175 -5565 41295 -5445
rect 41340 -5565 41460 -5445
rect 41505 -5565 41625 -5445
rect 41670 -5565 41790 -5445
rect 41845 -5565 41965 -5445
rect 36485 -5730 36605 -5610
rect 36650 -5730 36770 -5610
rect 36815 -5730 36935 -5610
rect 36980 -5730 37100 -5610
rect 37155 -5730 37275 -5610
rect 37320 -5730 37440 -5610
rect 37485 -5730 37605 -5610
rect 37650 -5730 37770 -5610
rect 37825 -5730 37945 -5610
rect 37990 -5730 38110 -5610
rect 38155 -5730 38275 -5610
rect 38320 -5730 38440 -5610
rect 38495 -5730 38615 -5610
rect 38660 -5730 38780 -5610
rect 38825 -5730 38945 -5610
rect 38990 -5730 39110 -5610
rect 39165 -5730 39285 -5610
rect 39330 -5730 39450 -5610
rect 39495 -5730 39615 -5610
rect 39660 -5730 39780 -5610
rect 39835 -5730 39955 -5610
rect 40000 -5730 40120 -5610
rect 40165 -5730 40285 -5610
rect 40330 -5730 40450 -5610
rect 40505 -5730 40625 -5610
rect 40670 -5730 40790 -5610
rect 40835 -5730 40955 -5610
rect 41000 -5730 41120 -5610
rect 41175 -5730 41295 -5610
rect 41340 -5730 41460 -5610
rect 41505 -5730 41625 -5610
rect 41670 -5730 41790 -5610
rect 41845 -5730 41965 -5610
rect 36485 -5905 36605 -5785
rect 36650 -5905 36770 -5785
rect 36815 -5905 36935 -5785
rect 36980 -5905 37100 -5785
rect 37155 -5905 37275 -5785
rect 37320 -5905 37440 -5785
rect 37485 -5905 37605 -5785
rect 37650 -5905 37770 -5785
rect 37825 -5905 37945 -5785
rect 37990 -5905 38110 -5785
rect 38155 -5905 38275 -5785
rect 38320 -5905 38440 -5785
rect 38495 -5905 38615 -5785
rect 38660 -5905 38780 -5785
rect 38825 -5905 38945 -5785
rect 38990 -5905 39110 -5785
rect 39165 -5905 39285 -5785
rect 39330 -5905 39450 -5785
rect 39495 -5905 39615 -5785
rect 39660 -5905 39780 -5785
rect 39835 -5905 39955 -5785
rect 40000 -5905 40120 -5785
rect 40165 -5905 40285 -5785
rect 40330 -5905 40450 -5785
rect 40505 -5905 40625 -5785
rect 40670 -5905 40790 -5785
rect 40835 -5905 40955 -5785
rect 41000 -5905 41120 -5785
rect 41175 -5905 41295 -5785
rect 41340 -5905 41460 -5785
rect 41505 -5905 41625 -5785
rect 41670 -5905 41790 -5785
rect 41845 -5905 41965 -5785
rect 36485 -6070 36605 -5950
rect 36650 -6070 36770 -5950
rect 36815 -6070 36935 -5950
rect 36980 -6070 37100 -5950
rect 37155 -6070 37275 -5950
rect 37320 -6070 37440 -5950
rect 37485 -6070 37605 -5950
rect 37650 -6070 37770 -5950
rect 37825 -6070 37945 -5950
rect 37990 -6070 38110 -5950
rect 38155 -6070 38275 -5950
rect 38320 -6070 38440 -5950
rect 38495 -6070 38615 -5950
rect 38660 -6070 38780 -5950
rect 38825 -6070 38945 -5950
rect 38990 -6070 39110 -5950
rect 39165 -6070 39285 -5950
rect 39330 -6070 39450 -5950
rect 39495 -6070 39615 -5950
rect 39660 -6070 39780 -5950
rect 39835 -6070 39955 -5950
rect 40000 -6070 40120 -5950
rect 40165 -6070 40285 -5950
rect 40330 -6070 40450 -5950
rect 40505 -6070 40625 -5950
rect 40670 -6070 40790 -5950
rect 40835 -6070 40955 -5950
rect 41000 -6070 41120 -5950
rect 41175 -6070 41295 -5950
rect 41340 -6070 41460 -5950
rect 41505 -6070 41625 -5950
rect 41670 -6070 41790 -5950
rect 41845 -6070 41965 -5950
rect 36485 -6235 36605 -6115
rect 36650 -6235 36770 -6115
rect 36815 -6235 36935 -6115
rect 36980 -6235 37100 -6115
rect 37155 -6235 37275 -6115
rect 37320 -6235 37440 -6115
rect 37485 -6235 37605 -6115
rect 37650 -6235 37770 -6115
rect 37825 -6235 37945 -6115
rect 37990 -6235 38110 -6115
rect 38155 -6235 38275 -6115
rect 38320 -6235 38440 -6115
rect 38495 -6235 38615 -6115
rect 38660 -6235 38780 -6115
rect 38825 -6235 38945 -6115
rect 38990 -6235 39110 -6115
rect 39165 -6235 39285 -6115
rect 39330 -6235 39450 -6115
rect 39495 -6235 39615 -6115
rect 39660 -6235 39780 -6115
rect 39835 -6235 39955 -6115
rect 40000 -6235 40120 -6115
rect 40165 -6235 40285 -6115
rect 40330 -6235 40450 -6115
rect 40505 -6235 40625 -6115
rect 40670 -6235 40790 -6115
rect 40835 -6235 40955 -6115
rect 41000 -6235 41120 -6115
rect 41175 -6235 41295 -6115
rect 41340 -6235 41460 -6115
rect 41505 -6235 41625 -6115
rect 41670 -6235 41790 -6115
rect 41845 -6235 41965 -6115
rect 36485 -6400 36605 -6280
rect 36650 -6400 36770 -6280
rect 36815 -6400 36935 -6280
rect 36980 -6400 37100 -6280
rect 37155 -6400 37275 -6280
rect 37320 -6400 37440 -6280
rect 37485 -6400 37605 -6280
rect 37650 -6400 37770 -6280
rect 37825 -6400 37945 -6280
rect 37990 -6400 38110 -6280
rect 38155 -6400 38275 -6280
rect 38320 -6400 38440 -6280
rect 38495 -6400 38615 -6280
rect 38660 -6400 38780 -6280
rect 38825 -6400 38945 -6280
rect 38990 -6400 39110 -6280
rect 39165 -6400 39285 -6280
rect 39330 -6400 39450 -6280
rect 39495 -6400 39615 -6280
rect 39660 -6400 39780 -6280
rect 39835 -6400 39955 -6280
rect 40000 -6400 40120 -6280
rect 40165 -6400 40285 -6280
rect 40330 -6400 40450 -6280
rect 40505 -6400 40625 -6280
rect 40670 -6400 40790 -6280
rect 40835 -6400 40955 -6280
rect 41000 -6400 41120 -6280
rect 41175 -6400 41295 -6280
rect 41340 -6400 41460 -6280
rect 41505 -6400 41625 -6280
rect 41670 -6400 41790 -6280
rect 41845 -6400 41965 -6280
rect 36485 -6575 36605 -6455
rect 36650 -6575 36770 -6455
rect 36815 -6575 36935 -6455
rect 36980 -6575 37100 -6455
rect 37155 -6575 37275 -6455
rect 37320 -6575 37440 -6455
rect 37485 -6575 37605 -6455
rect 37650 -6575 37770 -6455
rect 37825 -6575 37945 -6455
rect 37990 -6575 38110 -6455
rect 38155 -6575 38275 -6455
rect 38320 -6575 38440 -6455
rect 38495 -6575 38615 -6455
rect 38660 -6575 38780 -6455
rect 38825 -6575 38945 -6455
rect 38990 -6575 39110 -6455
rect 39165 -6575 39285 -6455
rect 39330 -6575 39450 -6455
rect 39495 -6575 39615 -6455
rect 39660 -6575 39780 -6455
rect 39835 -6575 39955 -6455
rect 40000 -6575 40120 -6455
rect 40165 -6575 40285 -6455
rect 40330 -6575 40450 -6455
rect 40505 -6575 40625 -6455
rect 40670 -6575 40790 -6455
rect 40835 -6575 40955 -6455
rect 41000 -6575 41120 -6455
rect 41175 -6575 41295 -6455
rect 41340 -6575 41460 -6455
rect 41505 -6575 41625 -6455
rect 41670 -6575 41790 -6455
rect 41845 -6575 41965 -6455
rect 36485 -6740 36605 -6620
rect 36650 -6740 36770 -6620
rect 36815 -6740 36935 -6620
rect 36980 -6740 37100 -6620
rect 37155 -6740 37275 -6620
rect 37320 -6740 37440 -6620
rect 37485 -6740 37605 -6620
rect 37650 -6740 37770 -6620
rect 37825 -6740 37945 -6620
rect 37990 -6740 38110 -6620
rect 38155 -6740 38275 -6620
rect 38320 -6740 38440 -6620
rect 38495 -6740 38615 -6620
rect 38660 -6740 38780 -6620
rect 38825 -6740 38945 -6620
rect 38990 -6740 39110 -6620
rect 39165 -6740 39285 -6620
rect 39330 -6740 39450 -6620
rect 39495 -6740 39615 -6620
rect 39660 -6740 39780 -6620
rect 39835 -6740 39955 -6620
rect 40000 -6740 40120 -6620
rect 40165 -6740 40285 -6620
rect 40330 -6740 40450 -6620
rect 40505 -6740 40625 -6620
rect 40670 -6740 40790 -6620
rect 40835 -6740 40955 -6620
rect 41000 -6740 41120 -6620
rect 41175 -6740 41295 -6620
rect 41340 -6740 41460 -6620
rect 41505 -6740 41625 -6620
rect 41670 -6740 41790 -6620
rect 41845 -6740 41965 -6620
rect 36485 -6905 36605 -6785
rect 36650 -6905 36770 -6785
rect 36815 -6905 36935 -6785
rect 36980 -6905 37100 -6785
rect 37155 -6905 37275 -6785
rect 37320 -6905 37440 -6785
rect 37485 -6905 37605 -6785
rect 37650 -6905 37770 -6785
rect 37825 -6905 37945 -6785
rect 37990 -6905 38110 -6785
rect 38155 -6905 38275 -6785
rect 38320 -6905 38440 -6785
rect 38495 -6905 38615 -6785
rect 38660 -6905 38780 -6785
rect 38825 -6905 38945 -6785
rect 38990 -6905 39110 -6785
rect 39165 -6905 39285 -6785
rect 39330 -6905 39450 -6785
rect 39495 -6905 39615 -6785
rect 39660 -6905 39780 -6785
rect 39835 -6905 39955 -6785
rect 40000 -6905 40120 -6785
rect 40165 -6905 40285 -6785
rect 40330 -6905 40450 -6785
rect 40505 -6905 40625 -6785
rect 40670 -6905 40790 -6785
rect 40835 -6905 40955 -6785
rect 41000 -6905 41120 -6785
rect 41175 -6905 41295 -6785
rect 41340 -6905 41460 -6785
rect 41505 -6905 41625 -6785
rect 41670 -6905 41790 -6785
rect 41845 -6905 41965 -6785
rect 36485 -7070 36605 -6950
rect 36650 -7070 36770 -6950
rect 36815 -7070 36935 -6950
rect 36980 -7070 37100 -6950
rect 37155 -7070 37275 -6950
rect 37320 -7070 37440 -6950
rect 37485 -7070 37605 -6950
rect 37650 -7070 37770 -6950
rect 37825 -7070 37945 -6950
rect 37990 -7070 38110 -6950
rect 38155 -7070 38275 -6950
rect 38320 -7070 38440 -6950
rect 38495 -7070 38615 -6950
rect 38660 -7070 38780 -6950
rect 38825 -7070 38945 -6950
rect 38990 -7070 39110 -6950
rect 39165 -7070 39285 -6950
rect 39330 -7070 39450 -6950
rect 39495 -7070 39615 -6950
rect 39660 -7070 39780 -6950
rect 39835 -7070 39955 -6950
rect 40000 -7070 40120 -6950
rect 40165 -7070 40285 -6950
rect 40330 -7070 40450 -6950
rect 40505 -7070 40625 -6950
rect 40670 -7070 40790 -6950
rect 40835 -7070 40955 -6950
rect 41000 -7070 41120 -6950
rect 41175 -7070 41295 -6950
rect 41340 -7070 41460 -6950
rect 41505 -7070 41625 -6950
rect 41670 -7070 41790 -6950
rect 41845 -7070 41965 -6950
rect 36485 -7245 36605 -7125
rect 36650 -7245 36770 -7125
rect 36815 -7245 36935 -7125
rect 36980 -7245 37100 -7125
rect 37155 -7245 37275 -7125
rect 37320 -7245 37440 -7125
rect 37485 -7245 37605 -7125
rect 37650 -7245 37770 -7125
rect 37825 -7245 37945 -7125
rect 37990 -7245 38110 -7125
rect 38155 -7245 38275 -7125
rect 38320 -7245 38440 -7125
rect 38495 -7245 38615 -7125
rect 38660 -7245 38780 -7125
rect 38825 -7245 38945 -7125
rect 38990 -7245 39110 -7125
rect 39165 -7245 39285 -7125
rect 39330 -7245 39450 -7125
rect 39495 -7245 39615 -7125
rect 39660 -7245 39780 -7125
rect 39835 -7245 39955 -7125
rect 40000 -7245 40120 -7125
rect 40165 -7245 40285 -7125
rect 40330 -7245 40450 -7125
rect 40505 -7245 40625 -7125
rect 40670 -7245 40790 -7125
rect 40835 -7245 40955 -7125
rect 41000 -7245 41120 -7125
rect 41175 -7245 41295 -7125
rect 41340 -7245 41460 -7125
rect 41505 -7245 41625 -7125
rect 41670 -7245 41790 -7125
rect 41845 -7245 41965 -7125
rect 36485 -7410 36605 -7290
rect 36650 -7410 36770 -7290
rect 36815 -7410 36935 -7290
rect 36980 -7410 37100 -7290
rect 37155 -7410 37275 -7290
rect 37320 -7410 37440 -7290
rect 37485 -7410 37605 -7290
rect 37650 -7410 37770 -7290
rect 37825 -7410 37945 -7290
rect 37990 -7410 38110 -7290
rect 38155 -7410 38275 -7290
rect 38320 -7410 38440 -7290
rect 38495 -7410 38615 -7290
rect 38660 -7410 38780 -7290
rect 38825 -7410 38945 -7290
rect 38990 -7410 39110 -7290
rect 39165 -7410 39285 -7290
rect 39330 -7410 39450 -7290
rect 39495 -7410 39615 -7290
rect 39660 -7410 39780 -7290
rect 39835 -7410 39955 -7290
rect 40000 -7410 40120 -7290
rect 40165 -7410 40285 -7290
rect 40330 -7410 40450 -7290
rect 40505 -7410 40625 -7290
rect 40670 -7410 40790 -7290
rect 40835 -7410 40955 -7290
rect 41000 -7410 41120 -7290
rect 41175 -7410 41295 -7290
rect 41340 -7410 41460 -7290
rect 41505 -7410 41625 -7290
rect 41670 -7410 41790 -7290
rect 41845 -7410 41965 -7290
rect 36485 -7575 36605 -7455
rect 36650 -7575 36770 -7455
rect 36815 -7575 36935 -7455
rect 36980 -7575 37100 -7455
rect 37155 -7575 37275 -7455
rect 37320 -7575 37440 -7455
rect 37485 -7575 37605 -7455
rect 37650 -7575 37770 -7455
rect 37825 -7575 37945 -7455
rect 37990 -7575 38110 -7455
rect 38155 -7575 38275 -7455
rect 38320 -7575 38440 -7455
rect 38495 -7575 38615 -7455
rect 38660 -7575 38780 -7455
rect 38825 -7575 38945 -7455
rect 38990 -7575 39110 -7455
rect 39165 -7575 39285 -7455
rect 39330 -7575 39450 -7455
rect 39495 -7575 39615 -7455
rect 39660 -7575 39780 -7455
rect 39835 -7575 39955 -7455
rect 40000 -7575 40120 -7455
rect 40165 -7575 40285 -7455
rect 40330 -7575 40450 -7455
rect 40505 -7575 40625 -7455
rect 40670 -7575 40790 -7455
rect 40835 -7575 40955 -7455
rect 41000 -7575 41120 -7455
rect 41175 -7575 41295 -7455
rect 41340 -7575 41460 -7455
rect 41505 -7575 41625 -7455
rect 41670 -7575 41790 -7455
rect 41845 -7575 41965 -7455
rect 36485 -7740 36605 -7620
rect 36650 -7740 36770 -7620
rect 36815 -7740 36935 -7620
rect 36980 -7740 37100 -7620
rect 37155 -7740 37275 -7620
rect 37320 -7740 37440 -7620
rect 37485 -7740 37605 -7620
rect 37650 -7740 37770 -7620
rect 37825 -7740 37945 -7620
rect 37990 -7740 38110 -7620
rect 38155 -7740 38275 -7620
rect 38320 -7740 38440 -7620
rect 38495 -7740 38615 -7620
rect 38660 -7740 38780 -7620
rect 38825 -7740 38945 -7620
rect 38990 -7740 39110 -7620
rect 39165 -7740 39285 -7620
rect 39330 -7740 39450 -7620
rect 39495 -7740 39615 -7620
rect 39660 -7740 39780 -7620
rect 39835 -7740 39955 -7620
rect 40000 -7740 40120 -7620
rect 40165 -7740 40285 -7620
rect 40330 -7740 40450 -7620
rect 40505 -7740 40625 -7620
rect 40670 -7740 40790 -7620
rect 40835 -7740 40955 -7620
rect 41000 -7740 41120 -7620
rect 41175 -7740 41295 -7620
rect 41340 -7740 41460 -7620
rect 41505 -7740 41625 -7620
rect 41670 -7740 41790 -7620
rect 41845 -7740 41965 -7620
rect 36485 -7915 36605 -7795
rect 36650 -7915 36770 -7795
rect 36815 -7915 36935 -7795
rect 36980 -7915 37100 -7795
rect 37155 -7915 37275 -7795
rect 37320 -7915 37440 -7795
rect 37485 -7915 37605 -7795
rect 37650 -7915 37770 -7795
rect 37825 -7915 37945 -7795
rect 37990 -7915 38110 -7795
rect 38155 -7915 38275 -7795
rect 38320 -7915 38440 -7795
rect 38495 -7915 38615 -7795
rect 38660 -7915 38780 -7795
rect 38825 -7915 38945 -7795
rect 38990 -7915 39110 -7795
rect 39165 -7915 39285 -7795
rect 39330 -7915 39450 -7795
rect 39495 -7915 39615 -7795
rect 39660 -7915 39780 -7795
rect 39835 -7915 39955 -7795
rect 40000 -7915 40120 -7795
rect 40165 -7915 40285 -7795
rect 40330 -7915 40450 -7795
rect 40505 -7915 40625 -7795
rect 40670 -7915 40790 -7795
rect 40835 -7915 40955 -7795
rect 41000 -7915 41120 -7795
rect 41175 -7915 41295 -7795
rect 41340 -7915 41460 -7795
rect 41505 -7915 41625 -7795
rect 41670 -7915 41790 -7795
rect 41845 -7915 41965 -7795
rect 36485 -8080 36605 -7960
rect 36650 -8080 36770 -7960
rect 36815 -8080 36935 -7960
rect 36980 -8080 37100 -7960
rect 37155 -8080 37275 -7960
rect 37320 -8080 37440 -7960
rect 37485 -8080 37605 -7960
rect 37650 -8080 37770 -7960
rect 37825 -8080 37945 -7960
rect 37990 -8080 38110 -7960
rect 38155 -8080 38275 -7960
rect 38320 -8080 38440 -7960
rect 38495 -8080 38615 -7960
rect 38660 -8080 38780 -7960
rect 38825 -8080 38945 -7960
rect 38990 -8080 39110 -7960
rect 39165 -8080 39285 -7960
rect 39330 -8080 39450 -7960
rect 39495 -8080 39615 -7960
rect 39660 -8080 39780 -7960
rect 39835 -8080 39955 -7960
rect 40000 -8080 40120 -7960
rect 40165 -8080 40285 -7960
rect 40330 -8080 40450 -7960
rect 40505 -8080 40625 -7960
rect 40670 -8080 40790 -7960
rect 40835 -8080 40955 -7960
rect 41000 -8080 41120 -7960
rect 41175 -8080 41295 -7960
rect 41340 -8080 41460 -7960
rect 41505 -8080 41625 -7960
rect 41670 -8080 41790 -7960
rect 41845 -8080 41965 -7960
rect 36485 -8245 36605 -8125
rect 36650 -8245 36770 -8125
rect 36815 -8245 36935 -8125
rect 36980 -8245 37100 -8125
rect 37155 -8245 37275 -8125
rect 37320 -8245 37440 -8125
rect 37485 -8245 37605 -8125
rect 37650 -8245 37770 -8125
rect 37825 -8245 37945 -8125
rect 37990 -8245 38110 -8125
rect 38155 -8245 38275 -8125
rect 38320 -8245 38440 -8125
rect 38495 -8245 38615 -8125
rect 38660 -8245 38780 -8125
rect 38825 -8245 38945 -8125
rect 38990 -8245 39110 -8125
rect 39165 -8245 39285 -8125
rect 39330 -8245 39450 -8125
rect 39495 -8245 39615 -8125
rect 39660 -8245 39780 -8125
rect 39835 -8245 39955 -8125
rect 40000 -8245 40120 -8125
rect 40165 -8245 40285 -8125
rect 40330 -8245 40450 -8125
rect 40505 -8245 40625 -8125
rect 40670 -8245 40790 -8125
rect 40835 -8245 40955 -8125
rect 41000 -8245 41120 -8125
rect 41175 -8245 41295 -8125
rect 41340 -8245 41460 -8125
rect 41505 -8245 41625 -8125
rect 41670 -8245 41790 -8125
rect 41845 -8245 41965 -8125
rect 36485 -8410 36605 -8290
rect 36650 -8410 36770 -8290
rect 36815 -8410 36935 -8290
rect 36980 -8410 37100 -8290
rect 37155 -8410 37275 -8290
rect 37320 -8410 37440 -8290
rect 37485 -8410 37605 -8290
rect 37650 -8410 37770 -8290
rect 37825 -8410 37945 -8290
rect 37990 -8410 38110 -8290
rect 38155 -8410 38275 -8290
rect 38320 -8410 38440 -8290
rect 38495 -8410 38615 -8290
rect 38660 -8410 38780 -8290
rect 38825 -8410 38945 -8290
rect 38990 -8410 39110 -8290
rect 39165 -8410 39285 -8290
rect 39330 -8410 39450 -8290
rect 39495 -8410 39615 -8290
rect 39660 -8410 39780 -8290
rect 39835 -8410 39955 -8290
rect 40000 -8410 40120 -8290
rect 40165 -8410 40285 -8290
rect 40330 -8410 40450 -8290
rect 40505 -8410 40625 -8290
rect 40670 -8410 40790 -8290
rect 40835 -8410 40955 -8290
rect 41000 -8410 41120 -8290
rect 41175 -8410 41295 -8290
rect 41340 -8410 41460 -8290
rect 41505 -8410 41625 -8290
rect 41670 -8410 41790 -8290
rect 41845 -8410 41965 -8290
rect 36485 -8585 36605 -8465
rect 36650 -8585 36770 -8465
rect 36815 -8585 36935 -8465
rect 36980 -8585 37100 -8465
rect 37155 -8585 37275 -8465
rect 37320 -8585 37440 -8465
rect 37485 -8585 37605 -8465
rect 37650 -8585 37770 -8465
rect 37825 -8585 37945 -8465
rect 37990 -8585 38110 -8465
rect 38155 -8585 38275 -8465
rect 38320 -8585 38440 -8465
rect 38495 -8585 38615 -8465
rect 38660 -8585 38780 -8465
rect 38825 -8585 38945 -8465
rect 38990 -8585 39110 -8465
rect 39165 -8585 39285 -8465
rect 39330 -8585 39450 -8465
rect 39495 -8585 39615 -8465
rect 39660 -8585 39780 -8465
rect 39835 -8585 39955 -8465
rect 40000 -8585 40120 -8465
rect 40165 -8585 40285 -8465
rect 40330 -8585 40450 -8465
rect 40505 -8585 40625 -8465
rect 40670 -8585 40790 -8465
rect 40835 -8585 40955 -8465
rect 41000 -8585 41120 -8465
rect 41175 -8585 41295 -8465
rect 41340 -8585 41460 -8465
rect 41505 -8585 41625 -8465
rect 41670 -8585 41790 -8465
rect 41845 -8585 41965 -8465
rect 36485 -8750 36605 -8630
rect 36650 -8750 36770 -8630
rect 36815 -8750 36935 -8630
rect 36980 -8750 37100 -8630
rect 37155 -8750 37275 -8630
rect 37320 -8750 37440 -8630
rect 37485 -8750 37605 -8630
rect 37650 -8750 37770 -8630
rect 37825 -8750 37945 -8630
rect 37990 -8750 38110 -8630
rect 38155 -8750 38275 -8630
rect 38320 -8750 38440 -8630
rect 38495 -8750 38615 -8630
rect 38660 -8750 38780 -8630
rect 38825 -8750 38945 -8630
rect 38990 -8750 39110 -8630
rect 39165 -8750 39285 -8630
rect 39330 -8750 39450 -8630
rect 39495 -8750 39615 -8630
rect 39660 -8750 39780 -8630
rect 39835 -8750 39955 -8630
rect 40000 -8750 40120 -8630
rect 40165 -8750 40285 -8630
rect 40330 -8750 40450 -8630
rect 40505 -8750 40625 -8630
rect 40670 -8750 40790 -8630
rect 40835 -8750 40955 -8630
rect 41000 -8750 41120 -8630
rect 41175 -8750 41295 -8630
rect 41340 -8750 41460 -8630
rect 41505 -8750 41625 -8630
rect 41670 -8750 41790 -8630
rect 41845 -8750 41965 -8630
rect 36485 -8915 36605 -8795
rect 36650 -8915 36770 -8795
rect 36815 -8915 36935 -8795
rect 36980 -8915 37100 -8795
rect 37155 -8915 37275 -8795
rect 37320 -8915 37440 -8795
rect 37485 -8915 37605 -8795
rect 37650 -8915 37770 -8795
rect 37825 -8915 37945 -8795
rect 37990 -8915 38110 -8795
rect 38155 -8915 38275 -8795
rect 38320 -8915 38440 -8795
rect 38495 -8915 38615 -8795
rect 38660 -8915 38780 -8795
rect 38825 -8915 38945 -8795
rect 38990 -8915 39110 -8795
rect 39165 -8915 39285 -8795
rect 39330 -8915 39450 -8795
rect 39495 -8915 39615 -8795
rect 39660 -8915 39780 -8795
rect 39835 -8915 39955 -8795
rect 40000 -8915 40120 -8795
rect 40165 -8915 40285 -8795
rect 40330 -8915 40450 -8795
rect 40505 -8915 40625 -8795
rect 40670 -8915 40790 -8795
rect 40835 -8915 40955 -8795
rect 41000 -8915 41120 -8795
rect 41175 -8915 41295 -8795
rect 41340 -8915 41460 -8795
rect 41505 -8915 41625 -8795
rect 41670 -8915 41790 -8795
rect 41845 -8915 41965 -8795
rect 36485 -9080 36605 -8960
rect 36650 -9080 36770 -8960
rect 36815 -9080 36935 -8960
rect 36980 -9080 37100 -8960
rect 37155 -9080 37275 -8960
rect 37320 -9080 37440 -8960
rect 37485 -9080 37605 -8960
rect 37650 -9080 37770 -8960
rect 37825 -9080 37945 -8960
rect 37990 -9080 38110 -8960
rect 38155 -9080 38275 -8960
rect 38320 -9080 38440 -8960
rect 38495 -9080 38615 -8960
rect 38660 -9080 38780 -8960
rect 38825 -9080 38945 -8960
rect 38990 -9080 39110 -8960
rect 39165 -9080 39285 -8960
rect 39330 -9080 39450 -8960
rect 39495 -9080 39615 -8960
rect 39660 -9080 39780 -8960
rect 39835 -9080 39955 -8960
rect 40000 -9080 40120 -8960
rect 40165 -9080 40285 -8960
rect 40330 -9080 40450 -8960
rect 40505 -9080 40625 -8960
rect 40670 -9080 40790 -8960
rect 40835 -9080 40955 -8960
rect 41000 -9080 41120 -8960
rect 41175 -9080 41295 -8960
rect 41340 -9080 41460 -8960
rect 41505 -9080 41625 -8960
rect 41670 -9080 41790 -8960
rect 41845 -9080 41965 -8960
rect 36485 -9255 36605 -9135
rect 36650 -9255 36770 -9135
rect 36815 -9255 36935 -9135
rect 36980 -9255 37100 -9135
rect 37155 -9255 37275 -9135
rect 37320 -9255 37440 -9135
rect 37485 -9255 37605 -9135
rect 37650 -9255 37770 -9135
rect 37825 -9255 37945 -9135
rect 37990 -9255 38110 -9135
rect 38155 -9255 38275 -9135
rect 38320 -9255 38440 -9135
rect 38495 -9255 38615 -9135
rect 38660 -9255 38780 -9135
rect 38825 -9255 38945 -9135
rect 38990 -9255 39110 -9135
rect 39165 -9255 39285 -9135
rect 39330 -9255 39450 -9135
rect 39495 -9255 39615 -9135
rect 39660 -9255 39780 -9135
rect 39835 -9255 39955 -9135
rect 40000 -9255 40120 -9135
rect 40165 -9255 40285 -9135
rect 40330 -9255 40450 -9135
rect 40505 -9255 40625 -9135
rect 40670 -9255 40790 -9135
rect 40835 -9255 40955 -9135
rect 41000 -9255 41120 -9135
rect 41175 -9255 41295 -9135
rect 41340 -9255 41460 -9135
rect 41505 -9255 41625 -9135
rect 41670 -9255 41790 -9135
rect 41845 -9255 41965 -9135
rect 36485 -9420 36605 -9300
rect 36650 -9420 36770 -9300
rect 36815 -9420 36935 -9300
rect 36980 -9420 37100 -9300
rect 37155 -9420 37275 -9300
rect 37320 -9420 37440 -9300
rect 37485 -9420 37605 -9300
rect 37650 -9420 37770 -9300
rect 37825 -9420 37945 -9300
rect 37990 -9420 38110 -9300
rect 38155 -9420 38275 -9300
rect 38320 -9420 38440 -9300
rect 38495 -9420 38615 -9300
rect 38660 -9420 38780 -9300
rect 38825 -9420 38945 -9300
rect 38990 -9420 39110 -9300
rect 39165 -9420 39285 -9300
rect 39330 -9420 39450 -9300
rect 39495 -9420 39615 -9300
rect 39660 -9420 39780 -9300
rect 39835 -9420 39955 -9300
rect 40000 -9420 40120 -9300
rect 40165 -9420 40285 -9300
rect 40330 -9420 40450 -9300
rect 40505 -9420 40625 -9300
rect 40670 -9420 40790 -9300
rect 40835 -9420 40955 -9300
rect 41000 -9420 41120 -9300
rect 41175 -9420 41295 -9300
rect 41340 -9420 41460 -9300
rect 41505 -9420 41625 -9300
rect 41670 -9420 41790 -9300
rect 41845 -9420 41965 -9300
rect 36485 -9585 36605 -9465
rect 36650 -9585 36770 -9465
rect 36815 -9585 36935 -9465
rect 36980 -9585 37100 -9465
rect 37155 -9585 37275 -9465
rect 37320 -9585 37440 -9465
rect 37485 -9585 37605 -9465
rect 37650 -9585 37770 -9465
rect 37825 -9585 37945 -9465
rect 37990 -9585 38110 -9465
rect 38155 -9585 38275 -9465
rect 38320 -9585 38440 -9465
rect 38495 -9585 38615 -9465
rect 38660 -9585 38780 -9465
rect 38825 -9585 38945 -9465
rect 38990 -9585 39110 -9465
rect 39165 -9585 39285 -9465
rect 39330 -9585 39450 -9465
rect 39495 -9585 39615 -9465
rect 39660 -9585 39780 -9465
rect 39835 -9585 39955 -9465
rect 40000 -9585 40120 -9465
rect 40165 -9585 40285 -9465
rect 40330 -9585 40450 -9465
rect 40505 -9585 40625 -9465
rect 40670 -9585 40790 -9465
rect 40835 -9585 40955 -9465
rect 41000 -9585 41120 -9465
rect 41175 -9585 41295 -9465
rect 41340 -9585 41460 -9465
rect 41505 -9585 41625 -9465
rect 41670 -9585 41790 -9465
rect 41845 -9585 41965 -9465
rect 36485 -9750 36605 -9630
rect 36650 -9750 36770 -9630
rect 36815 -9750 36935 -9630
rect 36980 -9750 37100 -9630
rect 37155 -9750 37275 -9630
rect 37320 -9750 37440 -9630
rect 37485 -9750 37605 -9630
rect 37650 -9750 37770 -9630
rect 37825 -9750 37945 -9630
rect 37990 -9750 38110 -9630
rect 38155 -9750 38275 -9630
rect 38320 -9750 38440 -9630
rect 38495 -9750 38615 -9630
rect 38660 -9750 38780 -9630
rect 38825 -9750 38945 -9630
rect 38990 -9750 39110 -9630
rect 39165 -9750 39285 -9630
rect 39330 -9750 39450 -9630
rect 39495 -9750 39615 -9630
rect 39660 -9750 39780 -9630
rect 39835 -9750 39955 -9630
rect 40000 -9750 40120 -9630
rect 40165 -9750 40285 -9630
rect 40330 -9750 40450 -9630
rect 40505 -9750 40625 -9630
rect 40670 -9750 40790 -9630
rect 40835 -9750 40955 -9630
rect 41000 -9750 41120 -9630
rect 41175 -9750 41295 -9630
rect 41340 -9750 41460 -9630
rect 41505 -9750 41625 -9630
rect 41670 -9750 41790 -9630
rect 41845 -9750 41965 -9630
rect 42175 -4390 42295 -4270
rect 42340 -4390 42460 -4270
rect 42505 -4390 42625 -4270
rect 42670 -4390 42790 -4270
rect 42845 -4390 42965 -4270
rect 43010 -4390 43130 -4270
rect 43175 -4390 43295 -4270
rect 43340 -4390 43460 -4270
rect 43515 -4390 43635 -4270
rect 43680 -4390 43800 -4270
rect 43845 -4390 43965 -4270
rect 44010 -4390 44130 -4270
rect 44185 -4390 44305 -4270
rect 44350 -4390 44470 -4270
rect 44515 -4390 44635 -4270
rect 44680 -4390 44800 -4270
rect 44855 -4390 44975 -4270
rect 45020 -4390 45140 -4270
rect 45185 -4390 45305 -4270
rect 45350 -4390 45470 -4270
rect 45525 -4390 45645 -4270
rect 45690 -4390 45810 -4270
rect 45855 -4390 45975 -4270
rect 46020 -4390 46140 -4270
rect 46195 -4390 46315 -4270
rect 46360 -4390 46480 -4270
rect 46525 -4390 46645 -4270
rect 46690 -4390 46810 -4270
rect 46865 -4390 46985 -4270
rect 47030 -4390 47150 -4270
rect 47195 -4390 47315 -4270
rect 47360 -4390 47480 -4270
rect 47535 -4390 47655 -4270
rect 42175 -4565 42295 -4445
rect 42340 -4565 42460 -4445
rect 42505 -4565 42625 -4445
rect 42670 -4565 42790 -4445
rect 42845 -4565 42965 -4445
rect 43010 -4565 43130 -4445
rect 43175 -4565 43295 -4445
rect 43340 -4565 43460 -4445
rect 43515 -4565 43635 -4445
rect 43680 -4565 43800 -4445
rect 43845 -4565 43965 -4445
rect 44010 -4565 44130 -4445
rect 44185 -4565 44305 -4445
rect 44350 -4565 44470 -4445
rect 44515 -4565 44635 -4445
rect 44680 -4565 44800 -4445
rect 44855 -4565 44975 -4445
rect 45020 -4565 45140 -4445
rect 45185 -4565 45305 -4445
rect 45350 -4565 45470 -4445
rect 45525 -4565 45645 -4445
rect 45690 -4565 45810 -4445
rect 45855 -4565 45975 -4445
rect 46020 -4565 46140 -4445
rect 46195 -4565 46315 -4445
rect 46360 -4565 46480 -4445
rect 46525 -4565 46645 -4445
rect 46690 -4565 46810 -4445
rect 46865 -4565 46985 -4445
rect 47030 -4565 47150 -4445
rect 47195 -4565 47315 -4445
rect 47360 -4565 47480 -4445
rect 47535 -4565 47655 -4445
rect 42175 -4730 42295 -4610
rect 42340 -4730 42460 -4610
rect 42505 -4730 42625 -4610
rect 42670 -4730 42790 -4610
rect 42845 -4730 42965 -4610
rect 43010 -4730 43130 -4610
rect 43175 -4730 43295 -4610
rect 43340 -4730 43460 -4610
rect 43515 -4730 43635 -4610
rect 43680 -4730 43800 -4610
rect 43845 -4730 43965 -4610
rect 44010 -4730 44130 -4610
rect 44185 -4730 44305 -4610
rect 44350 -4730 44470 -4610
rect 44515 -4730 44635 -4610
rect 44680 -4730 44800 -4610
rect 44855 -4730 44975 -4610
rect 45020 -4730 45140 -4610
rect 45185 -4730 45305 -4610
rect 45350 -4730 45470 -4610
rect 45525 -4730 45645 -4610
rect 45690 -4730 45810 -4610
rect 45855 -4730 45975 -4610
rect 46020 -4730 46140 -4610
rect 46195 -4730 46315 -4610
rect 46360 -4730 46480 -4610
rect 46525 -4730 46645 -4610
rect 46690 -4730 46810 -4610
rect 46865 -4730 46985 -4610
rect 47030 -4730 47150 -4610
rect 47195 -4730 47315 -4610
rect 47360 -4730 47480 -4610
rect 47535 -4730 47655 -4610
rect 42175 -4895 42295 -4775
rect 42340 -4895 42460 -4775
rect 42505 -4895 42625 -4775
rect 42670 -4895 42790 -4775
rect 42845 -4895 42965 -4775
rect 43010 -4895 43130 -4775
rect 43175 -4895 43295 -4775
rect 43340 -4895 43460 -4775
rect 43515 -4895 43635 -4775
rect 43680 -4895 43800 -4775
rect 43845 -4895 43965 -4775
rect 44010 -4895 44130 -4775
rect 44185 -4895 44305 -4775
rect 44350 -4895 44470 -4775
rect 44515 -4895 44635 -4775
rect 44680 -4895 44800 -4775
rect 44855 -4895 44975 -4775
rect 45020 -4895 45140 -4775
rect 45185 -4895 45305 -4775
rect 45350 -4895 45470 -4775
rect 45525 -4895 45645 -4775
rect 45690 -4895 45810 -4775
rect 45855 -4895 45975 -4775
rect 46020 -4895 46140 -4775
rect 46195 -4895 46315 -4775
rect 46360 -4895 46480 -4775
rect 46525 -4895 46645 -4775
rect 46690 -4895 46810 -4775
rect 46865 -4895 46985 -4775
rect 47030 -4895 47150 -4775
rect 47195 -4895 47315 -4775
rect 47360 -4895 47480 -4775
rect 47535 -4895 47655 -4775
rect 42175 -5060 42295 -4940
rect 42340 -5060 42460 -4940
rect 42505 -5060 42625 -4940
rect 42670 -5060 42790 -4940
rect 42845 -5060 42965 -4940
rect 43010 -5060 43130 -4940
rect 43175 -5060 43295 -4940
rect 43340 -5060 43460 -4940
rect 43515 -5060 43635 -4940
rect 43680 -5060 43800 -4940
rect 43845 -5060 43965 -4940
rect 44010 -5060 44130 -4940
rect 44185 -5060 44305 -4940
rect 44350 -5060 44470 -4940
rect 44515 -5060 44635 -4940
rect 44680 -5060 44800 -4940
rect 44855 -5060 44975 -4940
rect 45020 -5060 45140 -4940
rect 45185 -5060 45305 -4940
rect 45350 -5060 45470 -4940
rect 45525 -5060 45645 -4940
rect 45690 -5060 45810 -4940
rect 45855 -5060 45975 -4940
rect 46020 -5060 46140 -4940
rect 46195 -5060 46315 -4940
rect 46360 -5060 46480 -4940
rect 46525 -5060 46645 -4940
rect 46690 -5060 46810 -4940
rect 46865 -5060 46985 -4940
rect 47030 -5060 47150 -4940
rect 47195 -5060 47315 -4940
rect 47360 -5060 47480 -4940
rect 47535 -5060 47655 -4940
rect 42175 -5235 42295 -5115
rect 42340 -5235 42460 -5115
rect 42505 -5235 42625 -5115
rect 42670 -5235 42790 -5115
rect 42845 -5235 42965 -5115
rect 43010 -5235 43130 -5115
rect 43175 -5235 43295 -5115
rect 43340 -5235 43460 -5115
rect 43515 -5235 43635 -5115
rect 43680 -5235 43800 -5115
rect 43845 -5235 43965 -5115
rect 44010 -5235 44130 -5115
rect 44185 -5235 44305 -5115
rect 44350 -5235 44470 -5115
rect 44515 -5235 44635 -5115
rect 44680 -5235 44800 -5115
rect 44855 -5235 44975 -5115
rect 45020 -5235 45140 -5115
rect 45185 -5235 45305 -5115
rect 45350 -5235 45470 -5115
rect 45525 -5235 45645 -5115
rect 45690 -5235 45810 -5115
rect 45855 -5235 45975 -5115
rect 46020 -5235 46140 -5115
rect 46195 -5235 46315 -5115
rect 46360 -5235 46480 -5115
rect 46525 -5235 46645 -5115
rect 46690 -5235 46810 -5115
rect 46865 -5235 46985 -5115
rect 47030 -5235 47150 -5115
rect 47195 -5235 47315 -5115
rect 47360 -5235 47480 -5115
rect 47535 -5235 47655 -5115
rect 42175 -5400 42295 -5280
rect 42340 -5400 42460 -5280
rect 42505 -5400 42625 -5280
rect 42670 -5400 42790 -5280
rect 42845 -5400 42965 -5280
rect 43010 -5400 43130 -5280
rect 43175 -5400 43295 -5280
rect 43340 -5400 43460 -5280
rect 43515 -5400 43635 -5280
rect 43680 -5400 43800 -5280
rect 43845 -5400 43965 -5280
rect 44010 -5400 44130 -5280
rect 44185 -5400 44305 -5280
rect 44350 -5400 44470 -5280
rect 44515 -5400 44635 -5280
rect 44680 -5400 44800 -5280
rect 44855 -5400 44975 -5280
rect 45020 -5400 45140 -5280
rect 45185 -5400 45305 -5280
rect 45350 -5400 45470 -5280
rect 45525 -5400 45645 -5280
rect 45690 -5400 45810 -5280
rect 45855 -5400 45975 -5280
rect 46020 -5400 46140 -5280
rect 46195 -5400 46315 -5280
rect 46360 -5400 46480 -5280
rect 46525 -5400 46645 -5280
rect 46690 -5400 46810 -5280
rect 46865 -5400 46985 -5280
rect 47030 -5400 47150 -5280
rect 47195 -5400 47315 -5280
rect 47360 -5400 47480 -5280
rect 47535 -5400 47655 -5280
rect 42175 -5565 42295 -5445
rect 42340 -5565 42460 -5445
rect 42505 -5565 42625 -5445
rect 42670 -5565 42790 -5445
rect 42845 -5565 42965 -5445
rect 43010 -5565 43130 -5445
rect 43175 -5565 43295 -5445
rect 43340 -5565 43460 -5445
rect 43515 -5565 43635 -5445
rect 43680 -5565 43800 -5445
rect 43845 -5565 43965 -5445
rect 44010 -5565 44130 -5445
rect 44185 -5565 44305 -5445
rect 44350 -5565 44470 -5445
rect 44515 -5565 44635 -5445
rect 44680 -5565 44800 -5445
rect 44855 -5565 44975 -5445
rect 45020 -5565 45140 -5445
rect 45185 -5565 45305 -5445
rect 45350 -5565 45470 -5445
rect 45525 -5565 45645 -5445
rect 45690 -5565 45810 -5445
rect 45855 -5565 45975 -5445
rect 46020 -5565 46140 -5445
rect 46195 -5565 46315 -5445
rect 46360 -5565 46480 -5445
rect 46525 -5565 46645 -5445
rect 46690 -5565 46810 -5445
rect 46865 -5565 46985 -5445
rect 47030 -5565 47150 -5445
rect 47195 -5565 47315 -5445
rect 47360 -5565 47480 -5445
rect 47535 -5565 47655 -5445
rect 42175 -5730 42295 -5610
rect 42340 -5730 42460 -5610
rect 42505 -5730 42625 -5610
rect 42670 -5730 42790 -5610
rect 42845 -5730 42965 -5610
rect 43010 -5730 43130 -5610
rect 43175 -5730 43295 -5610
rect 43340 -5730 43460 -5610
rect 43515 -5730 43635 -5610
rect 43680 -5730 43800 -5610
rect 43845 -5730 43965 -5610
rect 44010 -5730 44130 -5610
rect 44185 -5730 44305 -5610
rect 44350 -5730 44470 -5610
rect 44515 -5730 44635 -5610
rect 44680 -5730 44800 -5610
rect 44855 -5730 44975 -5610
rect 45020 -5730 45140 -5610
rect 45185 -5730 45305 -5610
rect 45350 -5730 45470 -5610
rect 45525 -5730 45645 -5610
rect 45690 -5730 45810 -5610
rect 45855 -5730 45975 -5610
rect 46020 -5730 46140 -5610
rect 46195 -5730 46315 -5610
rect 46360 -5730 46480 -5610
rect 46525 -5730 46645 -5610
rect 46690 -5730 46810 -5610
rect 46865 -5730 46985 -5610
rect 47030 -5730 47150 -5610
rect 47195 -5730 47315 -5610
rect 47360 -5730 47480 -5610
rect 47535 -5730 47655 -5610
rect 42175 -5905 42295 -5785
rect 42340 -5905 42460 -5785
rect 42505 -5905 42625 -5785
rect 42670 -5905 42790 -5785
rect 42845 -5905 42965 -5785
rect 43010 -5905 43130 -5785
rect 43175 -5905 43295 -5785
rect 43340 -5905 43460 -5785
rect 43515 -5905 43635 -5785
rect 43680 -5905 43800 -5785
rect 43845 -5905 43965 -5785
rect 44010 -5905 44130 -5785
rect 44185 -5905 44305 -5785
rect 44350 -5905 44470 -5785
rect 44515 -5905 44635 -5785
rect 44680 -5905 44800 -5785
rect 44855 -5905 44975 -5785
rect 45020 -5905 45140 -5785
rect 45185 -5905 45305 -5785
rect 45350 -5905 45470 -5785
rect 45525 -5905 45645 -5785
rect 45690 -5905 45810 -5785
rect 45855 -5905 45975 -5785
rect 46020 -5905 46140 -5785
rect 46195 -5905 46315 -5785
rect 46360 -5905 46480 -5785
rect 46525 -5905 46645 -5785
rect 46690 -5905 46810 -5785
rect 46865 -5905 46985 -5785
rect 47030 -5905 47150 -5785
rect 47195 -5905 47315 -5785
rect 47360 -5905 47480 -5785
rect 47535 -5905 47655 -5785
rect 42175 -6070 42295 -5950
rect 42340 -6070 42460 -5950
rect 42505 -6070 42625 -5950
rect 42670 -6070 42790 -5950
rect 42845 -6070 42965 -5950
rect 43010 -6070 43130 -5950
rect 43175 -6070 43295 -5950
rect 43340 -6070 43460 -5950
rect 43515 -6070 43635 -5950
rect 43680 -6070 43800 -5950
rect 43845 -6070 43965 -5950
rect 44010 -6070 44130 -5950
rect 44185 -6070 44305 -5950
rect 44350 -6070 44470 -5950
rect 44515 -6070 44635 -5950
rect 44680 -6070 44800 -5950
rect 44855 -6070 44975 -5950
rect 45020 -6070 45140 -5950
rect 45185 -6070 45305 -5950
rect 45350 -6070 45470 -5950
rect 45525 -6070 45645 -5950
rect 45690 -6070 45810 -5950
rect 45855 -6070 45975 -5950
rect 46020 -6070 46140 -5950
rect 46195 -6070 46315 -5950
rect 46360 -6070 46480 -5950
rect 46525 -6070 46645 -5950
rect 46690 -6070 46810 -5950
rect 46865 -6070 46985 -5950
rect 47030 -6070 47150 -5950
rect 47195 -6070 47315 -5950
rect 47360 -6070 47480 -5950
rect 47535 -6070 47655 -5950
rect 42175 -6235 42295 -6115
rect 42340 -6235 42460 -6115
rect 42505 -6235 42625 -6115
rect 42670 -6235 42790 -6115
rect 42845 -6235 42965 -6115
rect 43010 -6235 43130 -6115
rect 43175 -6235 43295 -6115
rect 43340 -6235 43460 -6115
rect 43515 -6235 43635 -6115
rect 43680 -6235 43800 -6115
rect 43845 -6235 43965 -6115
rect 44010 -6235 44130 -6115
rect 44185 -6235 44305 -6115
rect 44350 -6235 44470 -6115
rect 44515 -6235 44635 -6115
rect 44680 -6235 44800 -6115
rect 44855 -6235 44975 -6115
rect 45020 -6235 45140 -6115
rect 45185 -6235 45305 -6115
rect 45350 -6235 45470 -6115
rect 45525 -6235 45645 -6115
rect 45690 -6235 45810 -6115
rect 45855 -6235 45975 -6115
rect 46020 -6235 46140 -6115
rect 46195 -6235 46315 -6115
rect 46360 -6235 46480 -6115
rect 46525 -6235 46645 -6115
rect 46690 -6235 46810 -6115
rect 46865 -6235 46985 -6115
rect 47030 -6235 47150 -6115
rect 47195 -6235 47315 -6115
rect 47360 -6235 47480 -6115
rect 47535 -6235 47655 -6115
rect 42175 -6400 42295 -6280
rect 42340 -6400 42460 -6280
rect 42505 -6400 42625 -6280
rect 42670 -6400 42790 -6280
rect 42845 -6400 42965 -6280
rect 43010 -6400 43130 -6280
rect 43175 -6400 43295 -6280
rect 43340 -6400 43460 -6280
rect 43515 -6400 43635 -6280
rect 43680 -6400 43800 -6280
rect 43845 -6400 43965 -6280
rect 44010 -6400 44130 -6280
rect 44185 -6400 44305 -6280
rect 44350 -6400 44470 -6280
rect 44515 -6400 44635 -6280
rect 44680 -6400 44800 -6280
rect 44855 -6400 44975 -6280
rect 45020 -6400 45140 -6280
rect 45185 -6400 45305 -6280
rect 45350 -6400 45470 -6280
rect 45525 -6400 45645 -6280
rect 45690 -6400 45810 -6280
rect 45855 -6400 45975 -6280
rect 46020 -6400 46140 -6280
rect 46195 -6400 46315 -6280
rect 46360 -6400 46480 -6280
rect 46525 -6400 46645 -6280
rect 46690 -6400 46810 -6280
rect 46865 -6400 46985 -6280
rect 47030 -6400 47150 -6280
rect 47195 -6400 47315 -6280
rect 47360 -6400 47480 -6280
rect 47535 -6400 47655 -6280
rect 42175 -6575 42295 -6455
rect 42340 -6575 42460 -6455
rect 42505 -6575 42625 -6455
rect 42670 -6575 42790 -6455
rect 42845 -6575 42965 -6455
rect 43010 -6575 43130 -6455
rect 43175 -6575 43295 -6455
rect 43340 -6575 43460 -6455
rect 43515 -6575 43635 -6455
rect 43680 -6575 43800 -6455
rect 43845 -6575 43965 -6455
rect 44010 -6575 44130 -6455
rect 44185 -6575 44305 -6455
rect 44350 -6575 44470 -6455
rect 44515 -6575 44635 -6455
rect 44680 -6575 44800 -6455
rect 44855 -6575 44975 -6455
rect 45020 -6575 45140 -6455
rect 45185 -6575 45305 -6455
rect 45350 -6575 45470 -6455
rect 45525 -6575 45645 -6455
rect 45690 -6575 45810 -6455
rect 45855 -6575 45975 -6455
rect 46020 -6575 46140 -6455
rect 46195 -6575 46315 -6455
rect 46360 -6575 46480 -6455
rect 46525 -6575 46645 -6455
rect 46690 -6575 46810 -6455
rect 46865 -6575 46985 -6455
rect 47030 -6575 47150 -6455
rect 47195 -6575 47315 -6455
rect 47360 -6575 47480 -6455
rect 47535 -6575 47655 -6455
rect 42175 -6740 42295 -6620
rect 42340 -6740 42460 -6620
rect 42505 -6740 42625 -6620
rect 42670 -6740 42790 -6620
rect 42845 -6740 42965 -6620
rect 43010 -6740 43130 -6620
rect 43175 -6740 43295 -6620
rect 43340 -6740 43460 -6620
rect 43515 -6740 43635 -6620
rect 43680 -6740 43800 -6620
rect 43845 -6740 43965 -6620
rect 44010 -6740 44130 -6620
rect 44185 -6740 44305 -6620
rect 44350 -6740 44470 -6620
rect 44515 -6740 44635 -6620
rect 44680 -6740 44800 -6620
rect 44855 -6740 44975 -6620
rect 45020 -6740 45140 -6620
rect 45185 -6740 45305 -6620
rect 45350 -6740 45470 -6620
rect 45525 -6740 45645 -6620
rect 45690 -6740 45810 -6620
rect 45855 -6740 45975 -6620
rect 46020 -6740 46140 -6620
rect 46195 -6740 46315 -6620
rect 46360 -6740 46480 -6620
rect 46525 -6740 46645 -6620
rect 46690 -6740 46810 -6620
rect 46865 -6740 46985 -6620
rect 47030 -6740 47150 -6620
rect 47195 -6740 47315 -6620
rect 47360 -6740 47480 -6620
rect 47535 -6740 47655 -6620
rect 42175 -6905 42295 -6785
rect 42340 -6905 42460 -6785
rect 42505 -6905 42625 -6785
rect 42670 -6905 42790 -6785
rect 42845 -6905 42965 -6785
rect 43010 -6905 43130 -6785
rect 43175 -6905 43295 -6785
rect 43340 -6905 43460 -6785
rect 43515 -6905 43635 -6785
rect 43680 -6905 43800 -6785
rect 43845 -6905 43965 -6785
rect 44010 -6905 44130 -6785
rect 44185 -6905 44305 -6785
rect 44350 -6905 44470 -6785
rect 44515 -6905 44635 -6785
rect 44680 -6905 44800 -6785
rect 44855 -6905 44975 -6785
rect 45020 -6905 45140 -6785
rect 45185 -6905 45305 -6785
rect 45350 -6905 45470 -6785
rect 45525 -6905 45645 -6785
rect 45690 -6905 45810 -6785
rect 45855 -6905 45975 -6785
rect 46020 -6905 46140 -6785
rect 46195 -6905 46315 -6785
rect 46360 -6905 46480 -6785
rect 46525 -6905 46645 -6785
rect 46690 -6905 46810 -6785
rect 46865 -6905 46985 -6785
rect 47030 -6905 47150 -6785
rect 47195 -6905 47315 -6785
rect 47360 -6905 47480 -6785
rect 47535 -6905 47655 -6785
rect 42175 -7070 42295 -6950
rect 42340 -7070 42460 -6950
rect 42505 -7070 42625 -6950
rect 42670 -7070 42790 -6950
rect 42845 -7070 42965 -6950
rect 43010 -7070 43130 -6950
rect 43175 -7070 43295 -6950
rect 43340 -7070 43460 -6950
rect 43515 -7070 43635 -6950
rect 43680 -7070 43800 -6950
rect 43845 -7070 43965 -6950
rect 44010 -7070 44130 -6950
rect 44185 -7070 44305 -6950
rect 44350 -7070 44470 -6950
rect 44515 -7070 44635 -6950
rect 44680 -7070 44800 -6950
rect 44855 -7070 44975 -6950
rect 45020 -7070 45140 -6950
rect 45185 -7070 45305 -6950
rect 45350 -7070 45470 -6950
rect 45525 -7070 45645 -6950
rect 45690 -7070 45810 -6950
rect 45855 -7070 45975 -6950
rect 46020 -7070 46140 -6950
rect 46195 -7070 46315 -6950
rect 46360 -7070 46480 -6950
rect 46525 -7070 46645 -6950
rect 46690 -7070 46810 -6950
rect 46865 -7070 46985 -6950
rect 47030 -7070 47150 -6950
rect 47195 -7070 47315 -6950
rect 47360 -7070 47480 -6950
rect 47535 -7070 47655 -6950
rect 42175 -7245 42295 -7125
rect 42340 -7245 42460 -7125
rect 42505 -7245 42625 -7125
rect 42670 -7245 42790 -7125
rect 42845 -7245 42965 -7125
rect 43010 -7245 43130 -7125
rect 43175 -7245 43295 -7125
rect 43340 -7245 43460 -7125
rect 43515 -7245 43635 -7125
rect 43680 -7245 43800 -7125
rect 43845 -7245 43965 -7125
rect 44010 -7245 44130 -7125
rect 44185 -7245 44305 -7125
rect 44350 -7245 44470 -7125
rect 44515 -7245 44635 -7125
rect 44680 -7245 44800 -7125
rect 44855 -7245 44975 -7125
rect 45020 -7245 45140 -7125
rect 45185 -7245 45305 -7125
rect 45350 -7245 45470 -7125
rect 45525 -7245 45645 -7125
rect 45690 -7245 45810 -7125
rect 45855 -7245 45975 -7125
rect 46020 -7245 46140 -7125
rect 46195 -7245 46315 -7125
rect 46360 -7245 46480 -7125
rect 46525 -7245 46645 -7125
rect 46690 -7245 46810 -7125
rect 46865 -7245 46985 -7125
rect 47030 -7245 47150 -7125
rect 47195 -7245 47315 -7125
rect 47360 -7245 47480 -7125
rect 47535 -7245 47655 -7125
rect 42175 -7410 42295 -7290
rect 42340 -7410 42460 -7290
rect 42505 -7410 42625 -7290
rect 42670 -7410 42790 -7290
rect 42845 -7410 42965 -7290
rect 43010 -7410 43130 -7290
rect 43175 -7410 43295 -7290
rect 43340 -7410 43460 -7290
rect 43515 -7410 43635 -7290
rect 43680 -7410 43800 -7290
rect 43845 -7410 43965 -7290
rect 44010 -7410 44130 -7290
rect 44185 -7410 44305 -7290
rect 44350 -7410 44470 -7290
rect 44515 -7410 44635 -7290
rect 44680 -7410 44800 -7290
rect 44855 -7410 44975 -7290
rect 45020 -7410 45140 -7290
rect 45185 -7410 45305 -7290
rect 45350 -7410 45470 -7290
rect 45525 -7410 45645 -7290
rect 45690 -7410 45810 -7290
rect 45855 -7410 45975 -7290
rect 46020 -7410 46140 -7290
rect 46195 -7410 46315 -7290
rect 46360 -7410 46480 -7290
rect 46525 -7410 46645 -7290
rect 46690 -7410 46810 -7290
rect 46865 -7410 46985 -7290
rect 47030 -7410 47150 -7290
rect 47195 -7410 47315 -7290
rect 47360 -7410 47480 -7290
rect 47535 -7410 47655 -7290
rect 42175 -7575 42295 -7455
rect 42340 -7575 42460 -7455
rect 42505 -7575 42625 -7455
rect 42670 -7575 42790 -7455
rect 42845 -7575 42965 -7455
rect 43010 -7575 43130 -7455
rect 43175 -7575 43295 -7455
rect 43340 -7575 43460 -7455
rect 43515 -7575 43635 -7455
rect 43680 -7575 43800 -7455
rect 43845 -7575 43965 -7455
rect 44010 -7575 44130 -7455
rect 44185 -7575 44305 -7455
rect 44350 -7575 44470 -7455
rect 44515 -7575 44635 -7455
rect 44680 -7575 44800 -7455
rect 44855 -7575 44975 -7455
rect 45020 -7575 45140 -7455
rect 45185 -7575 45305 -7455
rect 45350 -7575 45470 -7455
rect 45525 -7575 45645 -7455
rect 45690 -7575 45810 -7455
rect 45855 -7575 45975 -7455
rect 46020 -7575 46140 -7455
rect 46195 -7575 46315 -7455
rect 46360 -7575 46480 -7455
rect 46525 -7575 46645 -7455
rect 46690 -7575 46810 -7455
rect 46865 -7575 46985 -7455
rect 47030 -7575 47150 -7455
rect 47195 -7575 47315 -7455
rect 47360 -7575 47480 -7455
rect 47535 -7575 47655 -7455
rect 42175 -7740 42295 -7620
rect 42340 -7740 42460 -7620
rect 42505 -7740 42625 -7620
rect 42670 -7740 42790 -7620
rect 42845 -7740 42965 -7620
rect 43010 -7740 43130 -7620
rect 43175 -7740 43295 -7620
rect 43340 -7740 43460 -7620
rect 43515 -7740 43635 -7620
rect 43680 -7740 43800 -7620
rect 43845 -7740 43965 -7620
rect 44010 -7740 44130 -7620
rect 44185 -7740 44305 -7620
rect 44350 -7740 44470 -7620
rect 44515 -7740 44635 -7620
rect 44680 -7740 44800 -7620
rect 44855 -7740 44975 -7620
rect 45020 -7740 45140 -7620
rect 45185 -7740 45305 -7620
rect 45350 -7740 45470 -7620
rect 45525 -7740 45645 -7620
rect 45690 -7740 45810 -7620
rect 45855 -7740 45975 -7620
rect 46020 -7740 46140 -7620
rect 46195 -7740 46315 -7620
rect 46360 -7740 46480 -7620
rect 46525 -7740 46645 -7620
rect 46690 -7740 46810 -7620
rect 46865 -7740 46985 -7620
rect 47030 -7740 47150 -7620
rect 47195 -7740 47315 -7620
rect 47360 -7740 47480 -7620
rect 47535 -7740 47655 -7620
rect 42175 -7915 42295 -7795
rect 42340 -7915 42460 -7795
rect 42505 -7915 42625 -7795
rect 42670 -7915 42790 -7795
rect 42845 -7915 42965 -7795
rect 43010 -7915 43130 -7795
rect 43175 -7915 43295 -7795
rect 43340 -7915 43460 -7795
rect 43515 -7915 43635 -7795
rect 43680 -7915 43800 -7795
rect 43845 -7915 43965 -7795
rect 44010 -7915 44130 -7795
rect 44185 -7915 44305 -7795
rect 44350 -7915 44470 -7795
rect 44515 -7915 44635 -7795
rect 44680 -7915 44800 -7795
rect 44855 -7915 44975 -7795
rect 45020 -7915 45140 -7795
rect 45185 -7915 45305 -7795
rect 45350 -7915 45470 -7795
rect 45525 -7915 45645 -7795
rect 45690 -7915 45810 -7795
rect 45855 -7915 45975 -7795
rect 46020 -7915 46140 -7795
rect 46195 -7915 46315 -7795
rect 46360 -7915 46480 -7795
rect 46525 -7915 46645 -7795
rect 46690 -7915 46810 -7795
rect 46865 -7915 46985 -7795
rect 47030 -7915 47150 -7795
rect 47195 -7915 47315 -7795
rect 47360 -7915 47480 -7795
rect 47535 -7915 47655 -7795
rect 42175 -8080 42295 -7960
rect 42340 -8080 42460 -7960
rect 42505 -8080 42625 -7960
rect 42670 -8080 42790 -7960
rect 42845 -8080 42965 -7960
rect 43010 -8080 43130 -7960
rect 43175 -8080 43295 -7960
rect 43340 -8080 43460 -7960
rect 43515 -8080 43635 -7960
rect 43680 -8080 43800 -7960
rect 43845 -8080 43965 -7960
rect 44010 -8080 44130 -7960
rect 44185 -8080 44305 -7960
rect 44350 -8080 44470 -7960
rect 44515 -8080 44635 -7960
rect 44680 -8080 44800 -7960
rect 44855 -8080 44975 -7960
rect 45020 -8080 45140 -7960
rect 45185 -8080 45305 -7960
rect 45350 -8080 45470 -7960
rect 45525 -8080 45645 -7960
rect 45690 -8080 45810 -7960
rect 45855 -8080 45975 -7960
rect 46020 -8080 46140 -7960
rect 46195 -8080 46315 -7960
rect 46360 -8080 46480 -7960
rect 46525 -8080 46645 -7960
rect 46690 -8080 46810 -7960
rect 46865 -8080 46985 -7960
rect 47030 -8080 47150 -7960
rect 47195 -8080 47315 -7960
rect 47360 -8080 47480 -7960
rect 47535 -8080 47655 -7960
rect 42175 -8245 42295 -8125
rect 42340 -8245 42460 -8125
rect 42505 -8245 42625 -8125
rect 42670 -8245 42790 -8125
rect 42845 -8245 42965 -8125
rect 43010 -8245 43130 -8125
rect 43175 -8245 43295 -8125
rect 43340 -8245 43460 -8125
rect 43515 -8245 43635 -8125
rect 43680 -8245 43800 -8125
rect 43845 -8245 43965 -8125
rect 44010 -8245 44130 -8125
rect 44185 -8245 44305 -8125
rect 44350 -8245 44470 -8125
rect 44515 -8245 44635 -8125
rect 44680 -8245 44800 -8125
rect 44855 -8245 44975 -8125
rect 45020 -8245 45140 -8125
rect 45185 -8245 45305 -8125
rect 45350 -8245 45470 -8125
rect 45525 -8245 45645 -8125
rect 45690 -8245 45810 -8125
rect 45855 -8245 45975 -8125
rect 46020 -8245 46140 -8125
rect 46195 -8245 46315 -8125
rect 46360 -8245 46480 -8125
rect 46525 -8245 46645 -8125
rect 46690 -8245 46810 -8125
rect 46865 -8245 46985 -8125
rect 47030 -8245 47150 -8125
rect 47195 -8245 47315 -8125
rect 47360 -8245 47480 -8125
rect 47535 -8245 47655 -8125
rect 42175 -8410 42295 -8290
rect 42340 -8410 42460 -8290
rect 42505 -8410 42625 -8290
rect 42670 -8410 42790 -8290
rect 42845 -8410 42965 -8290
rect 43010 -8410 43130 -8290
rect 43175 -8410 43295 -8290
rect 43340 -8410 43460 -8290
rect 43515 -8410 43635 -8290
rect 43680 -8410 43800 -8290
rect 43845 -8410 43965 -8290
rect 44010 -8410 44130 -8290
rect 44185 -8410 44305 -8290
rect 44350 -8410 44470 -8290
rect 44515 -8410 44635 -8290
rect 44680 -8410 44800 -8290
rect 44855 -8410 44975 -8290
rect 45020 -8410 45140 -8290
rect 45185 -8410 45305 -8290
rect 45350 -8410 45470 -8290
rect 45525 -8410 45645 -8290
rect 45690 -8410 45810 -8290
rect 45855 -8410 45975 -8290
rect 46020 -8410 46140 -8290
rect 46195 -8410 46315 -8290
rect 46360 -8410 46480 -8290
rect 46525 -8410 46645 -8290
rect 46690 -8410 46810 -8290
rect 46865 -8410 46985 -8290
rect 47030 -8410 47150 -8290
rect 47195 -8410 47315 -8290
rect 47360 -8410 47480 -8290
rect 47535 -8410 47655 -8290
rect 42175 -8585 42295 -8465
rect 42340 -8585 42460 -8465
rect 42505 -8585 42625 -8465
rect 42670 -8585 42790 -8465
rect 42845 -8585 42965 -8465
rect 43010 -8585 43130 -8465
rect 43175 -8585 43295 -8465
rect 43340 -8585 43460 -8465
rect 43515 -8585 43635 -8465
rect 43680 -8585 43800 -8465
rect 43845 -8585 43965 -8465
rect 44010 -8585 44130 -8465
rect 44185 -8585 44305 -8465
rect 44350 -8585 44470 -8465
rect 44515 -8585 44635 -8465
rect 44680 -8585 44800 -8465
rect 44855 -8585 44975 -8465
rect 45020 -8585 45140 -8465
rect 45185 -8585 45305 -8465
rect 45350 -8585 45470 -8465
rect 45525 -8585 45645 -8465
rect 45690 -8585 45810 -8465
rect 45855 -8585 45975 -8465
rect 46020 -8585 46140 -8465
rect 46195 -8585 46315 -8465
rect 46360 -8585 46480 -8465
rect 46525 -8585 46645 -8465
rect 46690 -8585 46810 -8465
rect 46865 -8585 46985 -8465
rect 47030 -8585 47150 -8465
rect 47195 -8585 47315 -8465
rect 47360 -8585 47480 -8465
rect 47535 -8585 47655 -8465
rect 42175 -8750 42295 -8630
rect 42340 -8750 42460 -8630
rect 42505 -8750 42625 -8630
rect 42670 -8750 42790 -8630
rect 42845 -8750 42965 -8630
rect 43010 -8750 43130 -8630
rect 43175 -8750 43295 -8630
rect 43340 -8750 43460 -8630
rect 43515 -8750 43635 -8630
rect 43680 -8750 43800 -8630
rect 43845 -8750 43965 -8630
rect 44010 -8750 44130 -8630
rect 44185 -8750 44305 -8630
rect 44350 -8750 44470 -8630
rect 44515 -8750 44635 -8630
rect 44680 -8750 44800 -8630
rect 44855 -8750 44975 -8630
rect 45020 -8750 45140 -8630
rect 45185 -8750 45305 -8630
rect 45350 -8750 45470 -8630
rect 45525 -8750 45645 -8630
rect 45690 -8750 45810 -8630
rect 45855 -8750 45975 -8630
rect 46020 -8750 46140 -8630
rect 46195 -8750 46315 -8630
rect 46360 -8750 46480 -8630
rect 46525 -8750 46645 -8630
rect 46690 -8750 46810 -8630
rect 46865 -8750 46985 -8630
rect 47030 -8750 47150 -8630
rect 47195 -8750 47315 -8630
rect 47360 -8750 47480 -8630
rect 47535 -8750 47655 -8630
rect 42175 -8915 42295 -8795
rect 42340 -8915 42460 -8795
rect 42505 -8915 42625 -8795
rect 42670 -8915 42790 -8795
rect 42845 -8915 42965 -8795
rect 43010 -8915 43130 -8795
rect 43175 -8915 43295 -8795
rect 43340 -8915 43460 -8795
rect 43515 -8915 43635 -8795
rect 43680 -8915 43800 -8795
rect 43845 -8915 43965 -8795
rect 44010 -8915 44130 -8795
rect 44185 -8915 44305 -8795
rect 44350 -8915 44470 -8795
rect 44515 -8915 44635 -8795
rect 44680 -8915 44800 -8795
rect 44855 -8915 44975 -8795
rect 45020 -8915 45140 -8795
rect 45185 -8915 45305 -8795
rect 45350 -8915 45470 -8795
rect 45525 -8915 45645 -8795
rect 45690 -8915 45810 -8795
rect 45855 -8915 45975 -8795
rect 46020 -8915 46140 -8795
rect 46195 -8915 46315 -8795
rect 46360 -8915 46480 -8795
rect 46525 -8915 46645 -8795
rect 46690 -8915 46810 -8795
rect 46865 -8915 46985 -8795
rect 47030 -8915 47150 -8795
rect 47195 -8915 47315 -8795
rect 47360 -8915 47480 -8795
rect 47535 -8915 47655 -8795
rect 42175 -9080 42295 -8960
rect 42340 -9080 42460 -8960
rect 42505 -9080 42625 -8960
rect 42670 -9080 42790 -8960
rect 42845 -9080 42965 -8960
rect 43010 -9080 43130 -8960
rect 43175 -9080 43295 -8960
rect 43340 -9080 43460 -8960
rect 43515 -9080 43635 -8960
rect 43680 -9080 43800 -8960
rect 43845 -9080 43965 -8960
rect 44010 -9080 44130 -8960
rect 44185 -9080 44305 -8960
rect 44350 -9080 44470 -8960
rect 44515 -9080 44635 -8960
rect 44680 -9080 44800 -8960
rect 44855 -9080 44975 -8960
rect 45020 -9080 45140 -8960
rect 45185 -9080 45305 -8960
rect 45350 -9080 45470 -8960
rect 45525 -9080 45645 -8960
rect 45690 -9080 45810 -8960
rect 45855 -9080 45975 -8960
rect 46020 -9080 46140 -8960
rect 46195 -9080 46315 -8960
rect 46360 -9080 46480 -8960
rect 46525 -9080 46645 -8960
rect 46690 -9080 46810 -8960
rect 46865 -9080 46985 -8960
rect 47030 -9080 47150 -8960
rect 47195 -9080 47315 -8960
rect 47360 -9080 47480 -8960
rect 47535 -9080 47655 -8960
rect 42175 -9255 42295 -9135
rect 42340 -9255 42460 -9135
rect 42505 -9255 42625 -9135
rect 42670 -9255 42790 -9135
rect 42845 -9255 42965 -9135
rect 43010 -9255 43130 -9135
rect 43175 -9255 43295 -9135
rect 43340 -9255 43460 -9135
rect 43515 -9255 43635 -9135
rect 43680 -9255 43800 -9135
rect 43845 -9255 43965 -9135
rect 44010 -9255 44130 -9135
rect 44185 -9255 44305 -9135
rect 44350 -9255 44470 -9135
rect 44515 -9255 44635 -9135
rect 44680 -9255 44800 -9135
rect 44855 -9255 44975 -9135
rect 45020 -9255 45140 -9135
rect 45185 -9255 45305 -9135
rect 45350 -9255 45470 -9135
rect 45525 -9255 45645 -9135
rect 45690 -9255 45810 -9135
rect 45855 -9255 45975 -9135
rect 46020 -9255 46140 -9135
rect 46195 -9255 46315 -9135
rect 46360 -9255 46480 -9135
rect 46525 -9255 46645 -9135
rect 46690 -9255 46810 -9135
rect 46865 -9255 46985 -9135
rect 47030 -9255 47150 -9135
rect 47195 -9255 47315 -9135
rect 47360 -9255 47480 -9135
rect 47535 -9255 47655 -9135
rect 42175 -9420 42295 -9300
rect 42340 -9420 42460 -9300
rect 42505 -9420 42625 -9300
rect 42670 -9420 42790 -9300
rect 42845 -9420 42965 -9300
rect 43010 -9420 43130 -9300
rect 43175 -9420 43295 -9300
rect 43340 -9420 43460 -9300
rect 43515 -9420 43635 -9300
rect 43680 -9420 43800 -9300
rect 43845 -9420 43965 -9300
rect 44010 -9420 44130 -9300
rect 44185 -9420 44305 -9300
rect 44350 -9420 44470 -9300
rect 44515 -9420 44635 -9300
rect 44680 -9420 44800 -9300
rect 44855 -9420 44975 -9300
rect 45020 -9420 45140 -9300
rect 45185 -9420 45305 -9300
rect 45350 -9420 45470 -9300
rect 45525 -9420 45645 -9300
rect 45690 -9420 45810 -9300
rect 45855 -9420 45975 -9300
rect 46020 -9420 46140 -9300
rect 46195 -9420 46315 -9300
rect 46360 -9420 46480 -9300
rect 46525 -9420 46645 -9300
rect 46690 -9420 46810 -9300
rect 46865 -9420 46985 -9300
rect 47030 -9420 47150 -9300
rect 47195 -9420 47315 -9300
rect 47360 -9420 47480 -9300
rect 47535 -9420 47655 -9300
rect 42175 -9585 42295 -9465
rect 42340 -9585 42460 -9465
rect 42505 -9585 42625 -9465
rect 42670 -9585 42790 -9465
rect 42845 -9585 42965 -9465
rect 43010 -9585 43130 -9465
rect 43175 -9585 43295 -9465
rect 43340 -9585 43460 -9465
rect 43515 -9585 43635 -9465
rect 43680 -9585 43800 -9465
rect 43845 -9585 43965 -9465
rect 44010 -9585 44130 -9465
rect 44185 -9585 44305 -9465
rect 44350 -9585 44470 -9465
rect 44515 -9585 44635 -9465
rect 44680 -9585 44800 -9465
rect 44855 -9585 44975 -9465
rect 45020 -9585 45140 -9465
rect 45185 -9585 45305 -9465
rect 45350 -9585 45470 -9465
rect 45525 -9585 45645 -9465
rect 45690 -9585 45810 -9465
rect 45855 -9585 45975 -9465
rect 46020 -9585 46140 -9465
rect 46195 -9585 46315 -9465
rect 46360 -9585 46480 -9465
rect 46525 -9585 46645 -9465
rect 46690 -9585 46810 -9465
rect 46865 -9585 46985 -9465
rect 47030 -9585 47150 -9465
rect 47195 -9585 47315 -9465
rect 47360 -9585 47480 -9465
rect 47535 -9585 47655 -9465
rect 42175 -9750 42295 -9630
rect 42340 -9750 42460 -9630
rect 42505 -9750 42625 -9630
rect 42670 -9750 42790 -9630
rect 42845 -9750 42965 -9630
rect 43010 -9750 43130 -9630
rect 43175 -9750 43295 -9630
rect 43340 -9750 43460 -9630
rect 43515 -9750 43635 -9630
rect 43680 -9750 43800 -9630
rect 43845 -9750 43965 -9630
rect 44010 -9750 44130 -9630
rect 44185 -9750 44305 -9630
rect 44350 -9750 44470 -9630
rect 44515 -9750 44635 -9630
rect 44680 -9750 44800 -9630
rect 44855 -9750 44975 -9630
rect 45020 -9750 45140 -9630
rect 45185 -9750 45305 -9630
rect 45350 -9750 45470 -9630
rect 45525 -9750 45645 -9630
rect 45690 -9750 45810 -9630
rect 45855 -9750 45975 -9630
rect 46020 -9750 46140 -9630
rect 46195 -9750 46315 -9630
rect 46360 -9750 46480 -9630
rect 46525 -9750 46645 -9630
rect 46690 -9750 46810 -9630
rect 46865 -9750 46985 -9630
rect 47030 -9750 47150 -9630
rect 47195 -9750 47315 -9630
rect 47360 -9750 47480 -9630
rect 47535 -9750 47655 -9630
rect 47865 -4390 47985 -4270
rect 48030 -4390 48150 -4270
rect 48195 -4390 48315 -4270
rect 48360 -4390 48480 -4270
rect 48535 -4390 48655 -4270
rect 48700 -4390 48820 -4270
rect 48865 -4390 48985 -4270
rect 49030 -4390 49150 -4270
rect 49205 -4390 49325 -4270
rect 49370 -4390 49490 -4270
rect 49535 -4390 49655 -4270
rect 49700 -4390 49820 -4270
rect 49875 -4390 49995 -4270
rect 50040 -4390 50160 -4270
rect 50205 -4390 50325 -4270
rect 50370 -4390 50490 -4270
rect 50545 -4390 50665 -4270
rect 50710 -4390 50830 -4270
rect 50875 -4390 50995 -4270
rect 51040 -4390 51160 -4270
rect 51215 -4390 51335 -4270
rect 51380 -4390 51500 -4270
rect 51545 -4390 51665 -4270
rect 51710 -4390 51830 -4270
rect 51885 -4390 52005 -4270
rect 52050 -4390 52170 -4270
rect 52215 -4390 52335 -4270
rect 52380 -4390 52500 -4270
rect 52555 -4390 52675 -4270
rect 52720 -4390 52840 -4270
rect 52885 -4390 53005 -4270
rect 53050 -4390 53170 -4270
rect 53225 -4390 53345 -4270
rect 47865 -4565 47985 -4445
rect 48030 -4565 48150 -4445
rect 48195 -4565 48315 -4445
rect 48360 -4565 48480 -4445
rect 48535 -4565 48655 -4445
rect 48700 -4565 48820 -4445
rect 48865 -4565 48985 -4445
rect 49030 -4565 49150 -4445
rect 49205 -4565 49325 -4445
rect 49370 -4565 49490 -4445
rect 49535 -4565 49655 -4445
rect 49700 -4565 49820 -4445
rect 49875 -4565 49995 -4445
rect 50040 -4565 50160 -4445
rect 50205 -4565 50325 -4445
rect 50370 -4565 50490 -4445
rect 50545 -4565 50665 -4445
rect 50710 -4565 50830 -4445
rect 50875 -4565 50995 -4445
rect 51040 -4565 51160 -4445
rect 51215 -4565 51335 -4445
rect 51380 -4565 51500 -4445
rect 51545 -4565 51665 -4445
rect 51710 -4565 51830 -4445
rect 51885 -4565 52005 -4445
rect 52050 -4565 52170 -4445
rect 52215 -4565 52335 -4445
rect 52380 -4565 52500 -4445
rect 52555 -4565 52675 -4445
rect 52720 -4565 52840 -4445
rect 52885 -4565 53005 -4445
rect 53050 -4565 53170 -4445
rect 53225 -4565 53345 -4445
rect 47865 -4730 47985 -4610
rect 48030 -4730 48150 -4610
rect 48195 -4730 48315 -4610
rect 48360 -4730 48480 -4610
rect 48535 -4730 48655 -4610
rect 48700 -4730 48820 -4610
rect 48865 -4730 48985 -4610
rect 49030 -4730 49150 -4610
rect 49205 -4730 49325 -4610
rect 49370 -4730 49490 -4610
rect 49535 -4730 49655 -4610
rect 49700 -4730 49820 -4610
rect 49875 -4730 49995 -4610
rect 50040 -4730 50160 -4610
rect 50205 -4730 50325 -4610
rect 50370 -4730 50490 -4610
rect 50545 -4730 50665 -4610
rect 50710 -4730 50830 -4610
rect 50875 -4730 50995 -4610
rect 51040 -4730 51160 -4610
rect 51215 -4730 51335 -4610
rect 51380 -4730 51500 -4610
rect 51545 -4730 51665 -4610
rect 51710 -4730 51830 -4610
rect 51885 -4730 52005 -4610
rect 52050 -4730 52170 -4610
rect 52215 -4730 52335 -4610
rect 52380 -4730 52500 -4610
rect 52555 -4730 52675 -4610
rect 52720 -4730 52840 -4610
rect 52885 -4730 53005 -4610
rect 53050 -4730 53170 -4610
rect 53225 -4730 53345 -4610
rect 47865 -4895 47985 -4775
rect 48030 -4895 48150 -4775
rect 48195 -4895 48315 -4775
rect 48360 -4895 48480 -4775
rect 48535 -4895 48655 -4775
rect 48700 -4895 48820 -4775
rect 48865 -4895 48985 -4775
rect 49030 -4895 49150 -4775
rect 49205 -4895 49325 -4775
rect 49370 -4895 49490 -4775
rect 49535 -4895 49655 -4775
rect 49700 -4895 49820 -4775
rect 49875 -4895 49995 -4775
rect 50040 -4895 50160 -4775
rect 50205 -4895 50325 -4775
rect 50370 -4895 50490 -4775
rect 50545 -4895 50665 -4775
rect 50710 -4895 50830 -4775
rect 50875 -4895 50995 -4775
rect 51040 -4895 51160 -4775
rect 51215 -4895 51335 -4775
rect 51380 -4895 51500 -4775
rect 51545 -4895 51665 -4775
rect 51710 -4895 51830 -4775
rect 51885 -4895 52005 -4775
rect 52050 -4895 52170 -4775
rect 52215 -4895 52335 -4775
rect 52380 -4895 52500 -4775
rect 52555 -4895 52675 -4775
rect 52720 -4895 52840 -4775
rect 52885 -4895 53005 -4775
rect 53050 -4895 53170 -4775
rect 53225 -4895 53345 -4775
rect 47865 -5060 47985 -4940
rect 48030 -5060 48150 -4940
rect 48195 -5060 48315 -4940
rect 48360 -5060 48480 -4940
rect 48535 -5060 48655 -4940
rect 48700 -5060 48820 -4940
rect 48865 -5060 48985 -4940
rect 49030 -5060 49150 -4940
rect 49205 -5060 49325 -4940
rect 49370 -5060 49490 -4940
rect 49535 -5060 49655 -4940
rect 49700 -5060 49820 -4940
rect 49875 -5060 49995 -4940
rect 50040 -5060 50160 -4940
rect 50205 -5060 50325 -4940
rect 50370 -5060 50490 -4940
rect 50545 -5060 50665 -4940
rect 50710 -5060 50830 -4940
rect 50875 -5060 50995 -4940
rect 51040 -5060 51160 -4940
rect 51215 -5060 51335 -4940
rect 51380 -5060 51500 -4940
rect 51545 -5060 51665 -4940
rect 51710 -5060 51830 -4940
rect 51885 -5060 52005 -4940
rect 52050 -5060 52170 -4940
rect 52215 -5060 52335 -4940
rect 52380 -5060 52500 -4940
rect 52555 -5060 52675 -4940
rect 52720 -5060 52840 -4940
rect 52885 -5060 53005 -4940
rect 53050 -5060 53170 -4940
rect 53225 -5060 53345 -4940
rect 47865 -5235 47985 -5115
rect 48030 -5235 48150 -5115
rect 48195 -5235 48315 -5115
rect 48360 -5235 48480 -5115
rect 48535 -5235 48655 -5115
rect 48700 -5235 48820 -5115
rect 48865 -5235 48985 -5115
rect 49030 -5235 49150 -5115
rect 49205 -5235 49325 -5115
rect 49370 -5235 49490 -5115
rect 49535 -5235 49655 -5115
rect 49700 -5235 49820 -5115
rect 49875 -5235 49995 -5115
rect 50040 -5235 50160 -5115
rect 50205 -5235 50325 -5115
rect 50370 -5235 50490 -5115
rect 50545 -5235 50665 -5115
rect 50710 -5235 50830 -5115
rect 50875 -5235 50995 -5115
rect 51040 -5235 51160 -5115
rect 51215 -5235 51335 -5115
rect 51380 -5235 51500 -5115
rect 51545 -5235 51665 -5115
rect 51710 -5235 51830 -5115
rect 51885 -5235 52005 -5115
rect 52050 -5235 52170 -5115
rect 52215 -5235 52335 -5115
rect 52380 -5235 52500 -5115
rect 52555 -5235 52675 -5115
rect 52720 -5235 52840 -5115
rect 52885 -5235 53005 -5115
rect 53050 -5235 53170 -5115
rect 53225 -5235 53345 -5115
rect 47865 -5400 47985 -5280
rect 48030 -5400 48150 -5280
rect 48195 -5400 48315 -5280
rect 48360 -5400 48480 -5280
rect 48535 -5400 48655 -5280
rect 48700 -5400 48820 -5280
rect 48865 -5400 48985 -5280
rect 49030 -5400 49150 -5280
rect 49205 -5400 49325 -5280
rect 49370 -5400 49490 -5280
rect 49535 -5400 49655 -5280
rect 49700 -5400 49820 -5280
rect 49875 -5400 49995 -5280
rect 50040 -5400 50160 -5280
rect 50205 -5400 50325 -5280
rect 50370 -5400 50490 -5280
rect 50545 -5400 50665 -5280
rect 50710 -5400 50830 -5280
rect 50875 -5400 50995 -5280
rect 51040 -5400 51160 -5280
rect 51215 -5400 51335 -5280
rect 51380 -5400 51500 -5280
rect 51545 -5400 51665 -5280
rect 51710 -5400 51830 -5280
rect 51885 -5400 52005 -5280
rect 52050 -5400 52170 -5280
rect 52215 -5400 52335 -5280
rect 52380 -5400 52500 -5280
rect 52555 -5400 52675 -5280
rect 52720 -5400 52840 -5280
rect 52885 -5400 53005 -5280
rect 53050 -5400 53170 -5280
rect 53225 -5400 53345 -5280
rect 47865 -5565 47985 -5445
rect 48030 -5565 48150 -5445
rect 48195 -5565 48315 -5445
rect 48360 -5565 48480 -5445
rect 48535 -5565 48655 -5445
rect 48700 -5565 48820 -5445
rect 48865 -5565 48985 -5445
rect 49030 -5565 49150 -5445
rect 49205 -5565 49325 -5445
rect 49370 -5565 49490 -5445
rect 49535 -5565 49655 -5445
rect 49700 -5565 49820 -5445
rect 49875 -5565 49995 -5445
rect 50040 -5565 50160 -5445
rect 50205 -5565 50325 -5445
rect 50370 -5565 50490 -5445
rect 50545 -5565 50665 -5445
rect 50710 -5565 50830 -5445
rect 50875 -5565 50995 -5445
rect 51040 -5565 51160 -5445
rect 51215 -5565 51335 -5445
rect 51380 -5565 51500 -5445
rect 51545 -5565 51665 -5445
rect 51710 -5565 51830 -5445
rect 51885 -5565 52005 -5445
rect 52050 -5565 52170 -5445
rect 52215 -5565 52335 -5445
rect 52380 -5565 52500 -5445
rect 52555 -5565 52675 -5445
rect 52720 -5565 52840 -5445
rect 52885 -5565 53005 -5445
rect 53050 -5565 53170 -5445
rect 53225 -5565 53345 -5445
rect 47865 -5730 47985 -5610
rect 48030 -5730 48150 -5610
rect 48195 -5730 48315 -5610
rect 48360 -5730 48480 -5610
rect 48535 -5730 48655 -5610
rect 48700 -5730 48820 -5610
rect 48865 -5730 48985 -5610
rect 49030 -5730 49150 -5610
rect 49205 -5730 49325 -5610
rect 49370 -5730 49490 -5610
rect 49535 -5730 49655 -5610
rect 49700 -5730 49820 -5610
rect 49875 -5730 49995 -5610
rect 50040 -5730 50160 -5610
rect 50205 -5730 50325 -5610
rect 50370 -5730 50490 -5610
rect 50545 -5730 50665 -5610
rect 50710 -5730 50830 -5610
rect 50875 -5730 50995 -5610
rect 51040 -5730 51160 -5610
rect 51215 -5730 51335 -5610
rect 51380 -5730 51500 -5610
rect 51545 -5730 51665 -5610
rect 51710 -5730 51830 -5610
rect 51885 -5730 52005 -5610
rect 52050 -5730 52170 -5610
rect 52215 -5730 52335 -5610
rect 52380 -5730 52500 -5610
rect 52555 -5730 52675 -5610
rect 52720 -5730 52840 -5610
rect 52885 -5730 53005 -5610
rect 53050 -5730 53170 -5610
rect 53225 -5730 53345 -5610
rect 47865 -5905 47985 -5785
rect 48030 -5905 48150 -5785
rect 48195 -5905 48315 -5785
rect 48360 -5905 48480 -5785
rect 48535 -5905 48655 -5785
rect 48700 -5905 48820 -5785
rect 48865 -5905 48985 -5785
rect 49030 -5905 49150 -5785
rect 49205 -5905 49325 -5785
rect 49370 -5905 49490 -5785
rect 49535 -5905 49655 -5785
rect 49700 -5905 49820 -5785
rect 49875 -5905 49995 -5785
rect 50040 -5905 50160 -5785
rect 50205 -5905 50325 -5785
rect 50370 -5905 50490 -5785
rect 50545 -5905 50665 -5785
rect 50710 -5905 50830 -5785
rect 50875 -5905 50995 -5785
rect 51040 -5905 51160 -5785
rect 51215 -5905 51335 -5785
rect 51380 -5905 51500 -5785
rect 51545 -5905 51665 -5785
rect 51710 -5905 51830 -5785
rect 51885 -5905 52005 -5785
rect 52050 -5905 52170 -5785
rect 52215 -5905 52335 -5785
rect 52380 -5905 52500 -5785
rect 52555 -5905 52675 -5785
rect 52720 -5905 52840 -5785
rect 52885 -5905 53005 -5785
rect 53050 -5905 53170 -5785
rect 53225 -5905 53345 -5785
rect 47865 -6070 47985 -5950
rect 48030 -6070 48150 -5950
rect 48195 -6070 48315 -5950
rect 48360 -6070 48480 -5950
rect 48535 -6070 48655 -5950
rect 48700 -6070 48820 -5950
rect 48865 -6070 48985 -5950
rect 49030 -6070 49150 -5950
rect 49205 -6070 49325 -5950
rect 49370 -6070 49490 -5950
rect 49535 -6070 49655 -5950
rect 49700 -6070 49820 -5950
rect 49875 -6070 49995 -5950
rect 50040 -6070 50160 -5950
rect 50205 -6070 50325 -5950
rect 50370 -6070 50490 -5950
rect 50545 -6070 50665 -5950
rect 50710 -6070 50830 -5950
rect 50875 -6070 50995 -5950
rect 51040 -6070 51160 -5950
rect 51215 -6070 51335 -5950
rect 51380 -6070 51500 -5950
rect 51545 -6070 51665 -5950
rect 51710 -6070 51830 -5950
rect 51885 -6070 52005 -5950
rect 52050 -6070 52170 -5950
rect 52215 -6070 52335 -5950
rect 52380 -6070 52500 -5950
rect 52555 -6070 52675 -5950
rect 52720 -6070 52840 -5950
rect 52885 -6070 53005 -5950
rect 53050 -6070 53170 -5950
rect 53225 -6070 53345 -5950
rect 47865 -6235 47985 -6115
rect 48030 -6235 48150 -6115
rect 48195 -6235 48315 -6115
rect 48360 -6235 48480 -6115
rect 48535 -6235 48655 -6115
rect 48700 -6235 48820 -6115
rect 48865 -6235 48985 -6115
rect 49030 -6235 49150 -6115
rect 49205 -6235 49325 -6115
rect 49370 -6235 49490 -6115
rect 49535 -6235 49655 -6115
rect 49700 -6235 49820 -6115
rect 49875 -6235 49995 -6115
rect 50040 -6235 50160 -6115
rect 50205 -6235 50325 -6115
rect 50370 -6235 50490 -6115
rect 50545 -6235 50665 -6115
rect 50710 -6235 50830 -6115
rect 50875 -6235 50995 -6115
rect 51040 -6235 51160 -6115
rect 51215 -6235 51335 -6115
rect 51380 -6235 51500 -6115
rect 51545 -6235 51665 -6115
rect 51710 -6235 51830 -6115
rect 51885 -6235 52005 -6115
rect 52050 -6235 52170 -6115
rect 52215 -6235 52335 -6115
rect 52380 -6235 52500 -6115
rect 52555 -6235 52675 -6115
rect 52720 -6235 52840 -6115
rect 52885 -6235 53005 -6115
rect 53050 -6235 53170 -6115
rect 53225 -6235 53345 -6115
rect 47865 -6400 47985 -6280
rect 48030 -6400 48150 -6280
rect 48195 -6400 48315 -6280
rect 48360 -6400 48480 -6280
rect 48535 -6400 48655 -6280
rect 48700 -6400 48820 -6280
rect 48865 -6400 48985 -6280
rect 49030 -6400 49150 -6280
rect 49205 -6400 49325 -6280
rect 49370 -6400 49490 -6280
rect 49535 -6400 49655 -6280
rect 49700 -6400 49820 -6280
rect 49875 -6400 49995 -6280
rect 50040 -6400 50160 -6280
rect 50205 -6400 50325 -6280
rect 50370 -6400 50490 -6280
rect 50545 -6400 50665 -6280
rect 50710 -6400 50830 -6280
rect 50875 -6400 50995 -6280
rect 51040 -6400 51160 -6280
rect 51215 -6400 51335 -6280
rect 51380 -6400 51500 -6280
rect 51545 -6400 51665 -6280
rect 51710 -6400 51830 -6280
rect 51885 -6400 52005 -6280
rect 52050 -6400 52170 -6280
rect 52215 -6400 52335 -6280
rect 52380 -6400 52500 -6280
rect 52555 -6400 52675 -6280
rect 52720 -6400 52840 -6280
rect 52885 -6400 53005 -6280
rect 53050 -6400 53170 -6280
rect 53225 -6400 53345 -6280
rect 47865 -6575 47985 -6455
rect 48030 -6575 48150 -6455
rect 48195 -6575 48315 -6455
rect 48360 -6575 48480 -6455
rect 48535 -6575 48655 -6455
rect 48700 -6575 48820 -6455
rect 48865 -6575 48985 -6455
rect 49030 -6575 49150 -6455
rect 49205 -6575 49325 -6455
rect 49370 -6575 49490 -6455
rect 49535 -6575 49655 -6455
rect 49700 -6575 49820 -6455
rect 49875 -6575 49995 -6455
rect 50040 -6575 50160 -6455
rect 50205 -6575 50325 -6455
rect 50370 -6575 50490 -6455
rect 50545 -6575 50665 -6455
rect 50710 -6575 50830 -6455
rect 50875 -6575 50995 -6455
rect 51040 -6575 51160 -6455
rect 51215 -6575 51335 -6455
rect 51380 -6575 51500 -6455
rect 51545 -6575 51665 -6455
rect 51710 -6575 51830 -6455
rect 51885 -6575 52005 -6455
rect 52050 -6575 52170 -6455
rect 52215 -6575 52335 -6455
rect 52380 -6575 52500 -6455
rect 52555 -6575 52675 -6455
rect 52720 -6575 52840 -6455
rect 52885 -6575 53005 -6455
rect 53050 -6575 53170 -6455
rect 53225 -6575 53345 -6455
rect 47865 -6740 47985 -6620
rect 48030 -6740 48150 -6620
rect 48195 -6740 48315 -6620
rect 48360 -6740 48480 -6620
rect 48535 -6740 48655 -6620
rect 48700 -6740 48820 -6620
rect 48865 -6740 48985 -6620
rect 49030 -6740 49150 -6620
rect 49205 -6740 49325 -6620
rect 49370 -6740 49490 -6620
rect 49535 -6740 49655 -6620
rect 49700 -6740 49820 -6620
rect 49875 -6740 49995 -6620
rect 50040 -6740 50160 -6620
rect 50205 -6740 50325 -6620
rect 50370 -6740 50490 -6620
rect 50545 -6740 50665 -6620
rect 50710 -6740 50830 -6620
rect 50875 -6740 50995 -6620
rect 51040 -6740 51160 -6620
rect 51215 -6740 51335 -6620
rect 51380 -6740 51500 -6620
rect 51545 -6740 51665 -6620
rect 51710 -6740 51830 -6620
rect 51885 -6740 52005 -6620
rect 52050 -6740 52170 -6620
rect 52215 -6740 52335 -6620
rect 52380 -6740 52500 -6620
rect 52555 -6740 52675 -6620
rect 52720 -6740 52840 -6620
rect 52885 -6740 53005 -6620
rect 53050 -6740 53170 -6620
rect 53225 -6740 53345 -6620
rect 47865 -6905 47985 -6785
rect 48030 -6905 48150 -6785
rect 48195 -6905 48315 -6785
rect 48360 -6905 48480 -6785
rect 48535 -6905 48655 -6785
rect 48700 -6905 48820 -6785
rect 48865 -6905 48985 -6785
rect 49030 -6905 49150 -6785
rect 49205 -6905 49325 -6785
rect 49370 -6905 49490 -6785
rect 49535 -6905 49655 -6785
rect 49700 -6905 49820 -6785
rect 49875 -6905 49995 -6785
rect 50040 -6905 50160 -6785
rect 50205 -6905 50325 -6785
rect 50370 -6905 50490 -6785
rect 50545 -6905 50665 -6785
rect 50710 -6905 50830 -6785
rect 50875 -6905 50995 -6785
rect 51040 -6905 51160 -6785
rect 51215 -6905 51335 -6785
rect 51380 -6905 51500 -6785
rect 51545 -6905 51665 -6785
rect 51710 -6905 51830 -6785
rect 51885 -6905 52005 -6785
rect 52050 -6905 52170 -6785
rect 52215 -6905 52335 -6785
rect 52380 -6905 52500 -6785
rect 52555 -6905 52675 -6785
rect 52720 -6905 52840 -6785
rect 52885 -6905 53005 -6785
rect 53050 -6905 53170 -6785
rect 53225 -6905 53345 -6785
rect 47865 -7070 47985 -6950
rect 48030 -7070 48150 -6950
rect 48195 -7070 48315 -6950
rect 48360 -7070 48480 -6950
rect 48535 -7070 48655 -6950
rect 48700 -7070 48820 -6950
rect 48865 -7070 48985 -6950
rect 49030 -7070 49150 -6950
rect 49205 -7070 49325 -6950
rect 49370 -7070 49490 -6950
rect 49535 -7070 49655 -6950
rect 49700 -7070 49820 -6950
rect 49875 -7070 49995 -6950
rect 50040 -7070 50160 -6950
rect 50205 -7070 50325 -6950
rect 50370 -7070 50490 -6950
rect 50545 -7070 50665 -6950
rect 50710 -7070 50830 -6950
rect 50875 -7070 50995 -6950
rect 51040 -7070 51160 -6950
rect 51215 -7070 51335 -6950
rect 51380 -7070 51500 -6950
rect 51545 -7070 51665 -6950
rect 51710 -7070 51830 -6950
rect 51885 -7070 52005 -6950
rect 52050 -7070 52170 -6950
rect 52215 -7070 52335 -6950
rect 52380 -7070 52500 -6950
rect 52555 -7070 52675 -6950
rect 52720 -7070 52840 -6950
rect 52885 -7070 53005 -6950
rect 53050 -7070 53170 -6950
rect 53225 -7070 53345 -6950
rect 47865 -7245 47985 -7125
rect 48030 -7245 48150 -7125
rect 48195 -7245 48315 -7125
rect 48360 -7245 48480 -7125
rect 48535 -7245 48655 -7125
rect 48700 -7245 48820 -7125
rect 48865 -7245 48985 -7125
rect 49030 -7245 49150 -7125
rect 49205 -7245 49325 -7125
rect 49370 -7245 49490 -7125
rect 49535 -7245 49655 -7125
rect 49700 -7245 49820 -7125
rect 49875 -7245 49995 -7125
rect 50040 -7245 50160 -7125
rect 50205 -7245 50325 -7125
rect 50370 -7245 50490 -7125
rect 50545 -7245 50665 -7125
rect 50710 -7245 50830 -7125
rect 50875 -7245 50995 -7125
rect 51040 -7245 51160 -7125
rect 51215 -7245 51335 -7125
rect 51380 -7245 51500 -7125
rect 51545 -7245 51665 -7125
rect 51710 -7245 51830 -7125
rect 51885 -7245 52005 -7125
rect 52050 -7245 52170 -7125
rect 52215 -7245 52335 -7125
rect 52380 -7245 52500 -7125
rect 52555 -7245 52675 -7125
rect 52720 -7245 52840 -7125
rect 52885 -7245 53005 -7125
rect 53050 -7245 53170 -7125
rect 53225 -7245 53345 -7125
rect 47865 -7410 47985 -7290
rect 48030 -7410 48150 -7290
rect 48195 -7410 48315 -7290
rect 48360 -7410 48480 -7290
rect 48535 -7410 48655 -7290
rect 48700 -7410 48820 -7290
rect 48865 -7410 48985 -7290
rect 49030 -7410 49150 -7290
rect 49205 -7410 49325 -7290
rect 49370 -7410 49490 -7290
rect 49535 -7410 49655 -7290
rect 49700 -7410 49820 -7290
rect 49875 -7410 49995 -7290
rect 50040 -7410 50160 -7290
rect 50205 -7410 50325 -7290
rect 50370 -7410 50490 -7290
rect 50545 -7410 50665 -7290
rect 50710 -7410 50830 -7290
rect 50875 -7410 50995 -7290
rect 51040 -7410 51160 -7290
rect 51215 -7410 51335 -7290
rect 51380 -7410 51500 -7290
rect 51545 -7410 51665 -7290
rect 51710 -7410 51830 -7290
rect 51885 -7410 52005 -7290
rect 52050 -7410 52170 -7290
rect 52215 -7410 52335 -7290
rect 52380 -7410 52500 -7290
rect 52555 -7410 52675 -7290
rect 52720 -7410 52840 -7290
rect 52885 -7410 53005 -7290
rect 53050 -7410 53170 -7290
rect 53225 -7410 53345 -7290
rect 47865 -7575 47985 -7455
rect 48030 -7575 48150 -7455
rect 48195 -7575 48315 -7455
rect 48360 -7575 48480 -7455
rect 48535 -7575 48655 -7455
rect 48700 -7575 48820 -7455
rect 48865 -7575 48985 -7455
rect 49030 -7575 49150 -7455
rect 49205 -7575 49325 -7455
rect 49370 -7575 49490 -7455
rect 49535 -7575 49655 -7455
rect 49700 -7575 49820 -7455
rect 49875 -7575 49995 -7455
rect 50040 -7575 50160 -7455
rect 50205 -7575 50325 -7455
rect 50370 -7575 50490 -7455
rect 50545 -7575 50665 -7455
rect 50710 -7575 50830 -7455
rect 50875 -7575 50995 -7455
rect 51040 -7575 51160 -7455
rect 51215 -7575 51335 -7455
rect 51380 -7575 51500 -7455
rect 51545 -7575 51665 -7455
rect 51710 -7575 51830 -7455
rect 51885 -7575 52005 -7455
rect 52050 -7575 52170 -7455
rect 52215 -7575 52335 -7455
rect 52380 -7575 52500 -7455
rect 52555 -7575 52675 -7455
rect 52720 -7575 52840 -7455
rect 52885 -7575 53005 -7455
rect 53050 -7575 53170 -7455
rect 53225 -7575 53345 -7455
rect 47865 -7740 47985 -7620
rect 48030 -7740 48150 -7620
rect 48195 -7740 48315 -7620
rect 48360 -7740 48480 -7620
rect 48535 -7740 48655 -7620
rect 48700 -7740 48820 -7620
rect 48865 -7740 48985 -7620
rect 49030 -7740 49150 -7620
rect 49205 -7740 49325 -7620
rect 49370 -7740 49490 -7620
rect 49535 -7740 49655 -7620
rect 49700 -7740 49820 -7620
rect 49875 -7740 49995 -7620
rect 50040 -7740 50160 -7620
rect 50205 -7740 50325 -7620
rect 50370 -7740 50490 -7620
rect 50545 -7740 50665 -7620
rect 50710 -7740 50830 -7620
rect 50875 -7740 50995 -7620
rect 51040 -7740 51160 -7620
rect 51215 -7740 51335 -7620
rect 51380 -7740 51500 -7620
rect 51545 -7740 51665 -7620
rect 51710 -7740 51830 -7620
rect 51885 -7740 52005 -7620
rect 52050 -7740 52170 -7620
rect 52215 -7740 52335 -7620
rect 52380 -7740 52500 -7620
rect 52555 -7740 52675 -7620
rect 52720 -7740 52840 -7620
rect 52885 -7740 53005 -7620
rect 53050 -7740 53170 -7620
rect 53225 -7740 53345 -7620
rect 47865 -7915 47985 -7795
rect 48030 -7915 48150 -7795
rect 48195 -7915 48315 -7795
rect 48360 -7915 48480 -7795
rect 48535 -7915 48655 -7795
rect 48700 -7915 48820 -7795
rect 48865 -7915 48985 -7795
rect 49030 -7915 49150 -7795
rect 49205 -7915 49325 -7795
rect 49370 -7915 49490 -7795
rect 49535 -7915 49655 -7795
rect 49700 -7915 49820 -7795
rect 49875 -7915 49995 -7795
rect 50040 -7915 50160 -7795
rect 50205 -7915 50325 -7795
rect 50370 -7915 50490 -7795
rect 50545 -7915 50665 -7795
rect 50710 -7915 50830 -7795
rect 50875 -7915 50995 -7795
rect 51040 -7915 51160 -7795
rect 51215 -7915 51335 -7795
rect 51380 -7915 51500 -7795
rect 51545 -7915 51665 -7795
rect 51710 -7915 51830 -7795
rect 51885 -7915 52005 -7795
rect 52050 -7915 52170 -7795
rect 52215 -7915 52335 -7795
rect 52380 -7915 52500 -7795
rect 52555 -7915 52675 -7795
rect 52720 -7915 52840 -7795
rect 52885 -7915 53005 -7795
rect 53050 -7915 53170 -7795
rect 53225 -7915 53345 -7795
rect 47865 -8080 47985 -7960
rect 48030 -8080 48150 -7960
rect 48195 -8080 48315 -7960
rect 48360 -8080 48480 -7960
rect 48535 -8080 48655 -7960
rect 48700 -8080 48820 -7960
rect 48865 -8080 48985 -7960
rect 49030 -8080 49150 -7960
rect 49205 -8080 49325 -7960
rect 49370 -8080 49490 -7960
rect 49535 -8080 49655 -7960
rect 49700 -8080 49820 -7960
rect 49875 -8080 49995 -7960
rect 50040 -8080 50160 -7960
rect 50205 -8080 50325 -7960
rect 50370 -8080 50490 -7960
rect 50545 -8080 50665 -7960
rect 50710 -8080 50830 -7960
rect 50875 -8080 50995 -7960
rect 51040 -8080 51160 -7960
rect 51215 -8080 51335 -7960
rect 51380 -8080 51500 -7960
rect 51545 -8080 51665 -7960
rect 51710 -8080 51830 -7960
rect 51885 -8080 52005 -7960
rect 52050 -8080 52170 -7960
rect 52215 -8080 52335 -7960
rect 52380 -8080 52500 -7960
rect 52555 -8080 52675 -7960
rect 52720 -8080 52840 -7960
rect 52885 -8080 53005 -7960
rect 53050 -8080 53170 -7960
rect 53225 -8080 53345 -7960
rect 47865 -8245 47985 -8125
rect 48030 -8245 48150 -8125
rect 48195 -8245 48315 -8125
rect 48360 -8245 48480 -8125
rect 48535 -8245 48655 -8125
rect 48700 -8245 48820 -8125
rect 48865 -8245 48985 -8125
rect 49030 -8245 49150 -8125
rect 49205 -8245 49325 -8125
rect 49370 -8245 49490 -8125
rect 49535 -8245 49655 -8125
rect 49700 -8245 49820 -8125
rect 49875 -8245 49995 -8125
rect 50040 -8245 50160 -8125
rect 50205 -8245 50325 -8125
rect 50370 -8245 50490 -8125
rect 50545 -8245 50665 -8125
rect 50710 -8245 50830 -8125
rect 50875 -8245 50995 -8125
rect 51040 -8245 51160 -8125
rect 51215 -8245 51335 -8125
rect 51380 -8245 51500 -8125
rect 51545 -8245 51665 -8125
rect 51710 -8245 51830 -8125
rect 51885 -8245 52005 -8125
rect 52050 -8245 52170 -8125
rect 52215 -8245 52335 -8125
rect 52380 -8245 52500 -8125
rect 52555 -8245 52675 -8125
rect 52720 -8245 52840 -8125
rect 52885 -8245 53005 -8125
rect 53050 -8245 53170 -8125
rect 53225 -8245 53345 -8125
rect 47865 -8410 47985 -8290
rect 48030 -8410 48150 -8290
rect 48195 -8410 48315 -8290
rect 48360 -8410 48480 -8290
rect 48535 -8410 48655 -8290
rect 48700 -8410 48820 -8290
rect 48865 -8410 48985 -8290
rect 49030 -8410 49150 -8290
rect 49205 -8410 49325 -8290
rect 49370 -8410 49490 -8290
rect 49535 -8410 49655 -8290
rect 49700 -8410 49820 -8290
rect 49875 -8410 49995 -8290
rect 50040 -8410 50160 -8290
rect 50205 -8410 50325 -8290
rect 50370 -8410 50490 -8290
rect 50545 -8410 50665 -8290
rect 50710 -8410 50830 -8290
rect 50875 -8410 50995 -8290
rect 51040 -8410 51160 -8290
rect 51215 -8410 51335 -8290
rect 51380 -8410 51500 -8290
rect 51545 -8410 51665 -8290
rect 51710 -8410 51830 -8290
rect 51885 -8410 52005 -8290
rect 52050 -8410 52170 -8290
rect 52215 -8410 52335 -8290
rect 52380 -8410 52500 -8290
rect 52555 -8410 52675 -8290
rect 52720 -8410 52840 -8290
rect 52885 -8410 53005 -8290
rect 53050 -8410 53170 -8290
rect 53225 -8410 53345 -8290
rect 47865 -8585 47985 -8465
rect 48030 -8585 48150 -8465
rect 48195 -8585 48315 -8465
rect 48360 -8585 48480 -8465
rect 48535 -8585 48655 -8465
rect 48700 -8585 48820 -8465
rect 48865 -8585 48985 -8465
rect 49030 -8585 49150 -8465
rect 49205 -8585 49325 -8465
rect 49370 -8585 49490 -8465
rect 49535 -8585 49655 -8465
rect 49700 -8585 49820 -8465
rect 49875 -8585 49995 -8465
rect 50040 -8585 50160 -8465
rect 50205 -8585 50325 -8465
rect 50370 -8585 50490 -8465
rect 50545 -8585 50665 -8465
rect 50710 -8585 50830 -8465
rect 50875 -8585 50995 -8465
rect 51040 -8585 51160 -8465
rect 51215 -8585 51335 -8465
rect 51380 -8585 51500 -8465
rect 51545 -8585 51665 -8465
rect 51710 -8585 51830 -8465
rect 51885 -8585 52005 -8465
rect 52050 -8585 52170 -8465
rect 52215 -8585 52335 -8465
rect 52380 -8585 52500 -8465
rect 52555 -8585 52675 -8465
rect 52720 -8585 52840 -8465
rect 52885 -8585 53005 -8465
rect 53050 -8585 53170 -8465
rect 53225 -8585 53345 -8465
rect 47865 -8750 47985 -8630
rect 48030 -8750 48150 -8630
rect 48195 -8750 48315 -8630
rect 48360 -8750 48480 -8630
rect 48535 -8750 48655 -8630
rect 48700 -8750 48820 -8630
rect 48865 -8750 48985 -8630
rect 49030 -8750 49150 -8630
rect 49205 -8750 49325 -8630
rect 49370 -8750 49490 -8630
rect 49535 -8750 49655 -8630
rect 49700 -8750 49820 -8630
rect 49875 -8750 49995 -8630
rect 50040 -8750 50160 -8630
rect 50205 -8750 50325 -8630
rect 50370 -8750 50490 -8630
rect 50545 -8750 50665 -8630
rect 50710 -8750 50830 -8630
rect 50875 -8750 50995 -8630
rect 51040 -8750 51160 -8630
rect 51215 -8750 51335 -8630
rect 51380 -8750 51500 -8630
rect 51545 -8750 51665 -8630
rect 51710 -8750 51830 -8630
rect 51885 -8750 52005 -8630
rect 52050 -8750 52170 -8630
rect 52215 -8750 52335 -8630
rect 52380 -8750 52500 -8630
rect 52555 -8750 52675 -8630
rect 52720 -8750 52840 -8630
rect 52885 -8750 53005 -8630
rect 53050 -8750 53170 -8630
rect 53225 -8750 53345 -8630
rect 47865 -8915 47985 -8795
rect 48030 -8915 48150 -8795
rect 48195 -8915 48315 -8795
rect 48360 -8915 48480 -8795
rect 48535 -8915 48655 -8795
rect 48700 -8915 48820 -8795
rect 48865 -8915 48985 -8795
rect 49030 -8915 49150 -8795
rect 49205 -8915 49325 -8795
rect 49370 -8915 49490 -8795
rect 49535 -8915 49655 -8795
rect 49700 -8915 49820 -8795
rect 49875 -8915 49995 -8795
rect 50040 -8915 50160 -8795
rect 50205 -8915 50325 -8795
rect 50370 -8915 50490 -8795
rect 50545 -8915 50665 -8795
rect 50710 -8915 50830 -8795
rect 50875 -8915 50995 -8795
rect 51040 -8915 51160 -8795
rect 51215 -8915 51335 -8795
rect 51380 -8915 51500 -8795
rect 51545 -8915 51665 -8795
rect 51710 -8915 51830 -8795
rect 51885 -8915 52005 -8795
rect 52050 -8915 52170 -8795
rect 52215 -8915 52335 -8795
rect 52380 -8915 52500 -8795
rect 52555 -8915 52675 -8795
rect 52720 -8915 52840 -8795
rect 52885 -8915 53005 -8795
rect 53050 -8915 53170 -8795
rect 53225 -8915 53345 -8795
rect 47865 -9080 47985 -8960
rect 48030 -9080 48150 -8960
rect 48195 -9080 48315 -8960
rect 48360 -9080 48480 -8960
rect 48535 -9080 48655 -8960
rect 48700 -9080 48820 -8960
rect 48865 -9080 48985 -8960
rect 49030 -9080 49150 -8960
rect 49205 -9080 49325 -8960
rect 49370 -9080 49490 -8960
rect 49535 -9080 49655 -8960
rect 49700 -9080 49820 -8960
rect 49875 -9080 49995 -8960
rect 50040 -9080 50160 -8960
rect 50205 -9080 50325 -8960
rect 50370 -9080 50490 -8960
rect 50545 -9080 50665 -8960
rect 50710 -9080 50830 -8960
rect 50875 -9080 50995 -8960
rect 51040 -9080 51160 -8960
rect 51215 -9080 51335 -8960
rect 51380 -9080 51500 -8960
rect 51545 -9080 51665 -8960
rect 51710 -9080 51830 -8960
rect 51885 -9080 52005 -8960
rect 52050 -9080 52170 -8960
rect 52215 -9080 52335 -8960
rect 52380 -9080 52500 -8960
rect 52555 -9080 52675 -8960
rect 52720 -9080 52840 -8960
rect 52885 -9080 53005 -8960
rect 53050 -9080 53170 -8960
rect 53225 -9080 53345 -8960
rect 47865 -9255 47985 -9135
rect 48030 -9255 48150 -9135
rect 48195 -9255 48315 -9135
rect 48360 -9255 48480 -9135
rect 48535 -9255 48655 -9135
rect 48700 -9255 48820 -9135
rect 48865 -9255 48985 -9135
rect 49030 -9255 49150 -9135
rect 49205 -9255 49325 -9135
rect 49370 -9255 49490 -9135
rect 49535 -9255 49655 -9135
rect 49700 -9255 49820 -9135
rect 49875 -9255 49995 -9135
rect 50040 -9255 50160 -9135
rect 50205 -9255 50325 -9135
rect 50370 -9255 50490 -9135
rect 50545 -9255 50665 -9135
rect 50710 -9255 50830 -9135
rect 50875 -9255 50995 -9135
rect 51040 -9255 51160 -9135
rect 51215 -9255 51335 -9135
rect 51380 -9255 51500 -9135
rect 51545 -9255 51665 -9135
rect 51710 -9255 51830 -9135
rect 51885 -9255 52005 -9135
rect 52050 -9255 52170 -9135
rect 52215 -9255 52335 -9135
rect 52380 -9255 52500 -9135
rect 52555 -9255 52675 -9135
rect 52720 -9255 52840 -9135
rect 52885 -9255 53005 -9135
rect 53050 -9255 53170 -9135
rect 53225 -9255 53345 -9135
rect 47865 -9420 47985 -9300
rect 48030 -9420 48150 -9300
rect 48195 -9420 48315 -9300
rect 48360 -9420 48480 -9300
rect 48535 -9420 48655 -9300
rect 48700 -9420 48820 -9300
rect 48865 -9420 48985 -9300
rect 49030 -9420 49150 -9300
rect 49205 -9420 49325 -9300
rect 49370 -9420 49490 -9300
rect 49535 -9420 49655 -9300
rect 49700 -9420 49820 -9300
rect 49875 -9420 49995 -9300
rect 50040 -9420 50160 -9300
rect 50205 -9420 50325 -9300
rect 50370 -9420 50490 -9300
rect 50545 -9420 50665 -9300
rect 50710 -9420 50830 -9300
rect 50875 -9420 50995 -9300
rect 51040 -9420 51160 -9300
rect 51215 -9420 51335 -9300
rect 51380 -9420 51500 -9300
rect 51545 -9420 51665 -9300
rect 51710 -9420 51830 -9300
rect 51885 -9420 52005 -9300
rect 52050 -9420 52170 -9300
rect 52215 -9420 52335 -9300
rect 52380 -9420 52500 -9300
rect 52555 -9420 52675 -9300
rect 52720 -9420 52840 -9300
rect 52885 -9420 53005 -9300
rect 53050 -9420 53170 -9300
rect 53225 -9420 53345 -9300
rect 47865 -9585 47985 -9465
rect 48030 -9585 48150 -9465
rect 48195 -9585 48315 -9465
rect 48360 -9585 48480 -9465
rect 48535 -9585 48655 -9465
rect 48700 -9585 48820 -9465
rect 48865 -9585 48985 -9465
rect 49030 -9585 49150 -9465
rect 49205 -9585 49325 -9465
rect 49370 -9585 49490 -9465
rect 49535 -9585 49655 -9465
rect 49700 -9585 49820 -9465
rect 49875 -9585 49995 -9465
rect 50040 -9585 50160 -9465
rect 50205 -9585 50325 -9465
rect 50370 -9585 50490 -9465
rect 50545 -9585 50665 -9465
rect 50710 -9585 50830 -9465
rect 50875 -9585 50995 -9465
rect 51040 -9585 51160 -9465
rect 51215 -9585 51335 -9465
rect 51380 -9585 51500 -9465
rect 51545 -9585 51665 -9465
rect 51710 -9585 51830 -9465
rect 51885 -9585 52005 -9465
rect 52050 -9585 52170 -9465
rect 52215 -9585 52335 -9465
rect 52380 -9585 52500 -9465
rect 52555 -9585 52675 -9465
rect 52720 -9585 52840 -9465
rect 52885 -9585 53005 -9465
rect 53050 -9585 53170 -9465
rect 53225 -9585 53345 -9465
rect 47865 -9750 47985 -9630
rect 48030 -9750 48150 -9630
rect 48195 -9750 48315 -9630
rect 48360 -9750 48480 -9630
rect 48535 -9750 48655 -9630
rect 48700 -9750 48820 -9630
rect 48865 -9750 48985 -9630
rect 49030 -9750 49150 -9630
rect 49205 -9750 49325 -9630
rect 49370 -9750 49490 -9630
rect 49535 -9750 49655 -9630
rect 49700 -9750 49820 -9630
rect 49875 -9750 49995 -9630
rect 50040 -9750 50160 -9630
rect 50205 -9750 50325 -9630
rect 50370 -9750 50490 -9630
rect 50545 -9750 50665 -9630
rect 50710 -9750 50830 -9630
rect 50875 -9750 50995 -9630
rect 51040 -9750 51160 -9630
rect 51215 -9750 51335 -9630
rect 51380 -9750 51500 -9630
rect 51545 -9750 51665 -9630
rect 51710 -9750 51830 -9630
rect 51885 -9750 52005 -9630
rect 52050 -9750 52170 -9630
rect 52215 -9750 52335 -9630
rect 52380 -9750 52500 -9630
rect 52555 -9750 52675 -9630
rect 52720 -9750 52840 -9630
rect 52885 -9750 53005 -9630
rect 53050 -9750 53170 -9630
rect 53225 -9750 53345 -9630
rect 30795 -10170 30915 -10050
rect 30970 -10170 31090 -10050
rect 31135 -10170 31255 -10050
rect 31300 -10170 31420 -10050
rect 31465 -10170 31585 -10050
rect 31640 -10170 31760 -10050
rect 31805 -10170 31925 -10050
rect 31970 -10170 32090 -10050
rect 32135 -10170 32255 -10050
rect 32310 -10170 32430 -10050
rect 32475 -10170 32595 -10050
rect 32640 -10170 32760 -10050
rect 32805 -10170 32925 -10050
rect 32980 -10170 33100 -10050
rect 33145 -10170 33265 -10050
rect 33310 -10170 33430 -10050
rect 33475 -10170 33595 -10050
rect 33650 -10170 33770 -10050
rect 33815 -10170 33935 -10050
rect 33980 -10170 34100 -10050
rect 34145 -10170 34265 -10050
rect 34320 -10170 34440 -10050
rect 34485 -10170 34605 -10050
rect 34650 -10170 34770 -10050
rect 34815 -10170 34935 -10050
rect 34990 -10170 35110 -10050
rect 35155 -10170 35275 -10050
rect 35320 -10170 35440 -10050
rect 35485 -10170 35605 -10050
rect 35660 -10170 35780 -10050
rect 35825 -10170 35945 -10050
rect 35990 -10170 36110 -10050
rect 36155 -10170 36275 -10050
rect 30795 -10335 30915 -10215
rect 30970 -10335 31090 -10215
rect 31135 -10335 31255 -10215
rect 31300 -10335 31420 -10215
rect 31465 -10335 31585 -10215
rect 31640 -10335 31760 -10215
rect 31805 -10335 31925 -10215
rect 31970 -10335 32090 -10215
rect 32135 -10335 32255 -10215
rect 32310 -10335 32430 -10215
rect 32475 -10335 32595 -10215
rect 32640 -10335 32760 -10215
rect 32805 -10335 32925 -10215
rect 32980 -10335 33100 -10215
rect 33145 -10335 33265 -10215
rect 33310 -10335 33430 -10215
rect 33475 -10335 33595 -10215
rect 33650 -10335 33770 -10215
rect 33815 -10335 33935 -10215
rect 33980 -10335 34100 -10215
rect 34145 -10335 34265 -10215
rect 34320 -10335 34440 -10215
rect 34485 -10335 34605 -10215
rect 34650 -10335 34770 -10215
rect 34815 -10335 34935 -10215
rect 34990 -10335 35110 -10215
rect 35155 -10335 35275 -10215
rect 35320 -10335 35440 -10215
rect 35485 -10335 35605 -10215
rect 35660 -10335 35780 -10215
rect 35825 -10335 35945 -10215
rect 35990 -10335 36110 -10215
rect 36155 -10335 36275 -10215
rect 30795 -10500 30915 -10380
rect 30970 -10500 31090 -10380
rect 31135 -10500 31255 -10380
rect 31300 -10500 31420 -10380
rect 31465 -10500 31585 -10380
rect 31640 -10500 31760 -10380
rect 31805 -10500 31925 -10380
rect 31970 -10500 32090 -10380
rect 32135 -10500 32255 -10380
rect 32310 -10500 32430 -10380
rect 32475 -10500 32595 -10380
rect 32640 -10500 32760 -10380
rect 32805 -10500 32925 -10380
rect 32980 -10500 33100 -10380
rect 33145 -10500 33265 -10380
rect 33310 -10500 33430 -10380
rect 33475 -10500 33595 -10380
rect 33650 -10500 33770 -10380
rect 33815 -10500 33935 -10380
rect 33980 -10500 34100 -10380
rect 34145 -10500 34265 -10380
rect 34320 -10500 34440 -10380
rect 34485 -10500 34605 -10380
rect 34650 -10500 34770 -10380
rect 34815 -10500 34935 -10380
rect 34990 -10500 35110 -10380
rect 35155 -10500 35275 -10380
rect 35320 -10500 35440 -10380
rect 35485 -10500 35605 -10380
rect 35660 -10500 35780 -10380
rect 35825 -10500 35945 -10380
rect 35990 -10500 36110 -10380
rect 36155 -10500 36275 -10380
rect 30795 -10665 30915 -10545
rect 30970 -10665 31090 -10545
rect 31135 -10665 31255 -10545
rect 31300 -10665 31420 -10545
rect 31465 -10665 31585 -10545
rect 31640 -10665 31760 -10545
rect 31805 -10665 31925 -10545
rect 31970 -10665 32090 -10545
rect 32135 -10665 32255 -10545
rect 32310 -10665 32430 -10545
rect 32475 -10665 32595 -10545
rect 32640 -10665 32760 -10545
rect 32805 -10665 32925 -10545
rect 32980 -10665 33100 -10545
rect 33145 -10665 33265 -10545
rect 33310 -10665 33430 -10545
rect 33475 -10665 33595 -10545
rect 33650 -10665 33770 -10545
rect 33815 -10665 33935 -10545
rect 33980 -10665 34100 -10545
rect 34145 -10665 34265 -10545
rect 34320 -10665 34440 -10545
rect 34485 -10665 34605 -10545
rect 34650 -10665 34770 -10545
rect 34815 -10665 34935 -10545
rect 34990 -10665 35110 -10545
rect 35155 -10665 35275 -10545
rect 35320 -10665 35440 -10545
rect 35485 -10665 35605 -10545
rect 35660 -10665 35780 -10545
rect 35825 -10665 35945 -10545
rect 35990 -10665 36110 -10545
rect 36155 -10665 36275 -10545
rect 30795 -10840 30915 -10720
rect 30970 -10840 31090 -10720
rect 31135 -10840 31255 -10720
rect 31300 -10840 31420 -10720
rect 31465 -10840 31585 -10720
rect 31640 -10840 31760 -10720
rect 31805 -10840 31925 -10720
rect 31970 -10840 32090 -10720
rect 32135 -10840 32255 -10720
rect 32310 -10840 32430 -10720
rect 32475 -10840 32595 -10720
rect 32640 -10840 32760 -10720
rect 32805 -10840 32925 -10720
rect 32980 -10840 33100 -10720
rect 33145 -10840 33265 -10720
rect 33310 -10840 33430 -10720
rect 33475 -10840 33595 -10720
rect 33650 -10840 33770 -10720
rect 33815 -10840 33935 -10720
rect 33980 -10840 34100 -10720
rect 34145 -10840 34265 -10720
rect 34320 -10840 34440 -10720
rect 34485 -10840 34605 -10720
rect 34650 -10840 34770 -10720
rect 34815 -10840 34935 -10720
rect 34990 -10840 35110 -10720
rect 35155 -10840 35275 -10720
rect 35320 -10840 35440 -10720
rect 35485 -10840 35605 -10720
rect 35660 -10840 35780 -10720
rect 35825 -10840 35945 -10720
rect 35990 -10840 36110 -10720
rect 36155 -10840 36275 -10720
rect 30795 -11005 30915 -10885
rect 30970 -11005 31090 -10885
rect 31135 -11005 31255 -10885
rect 31300 -11005 31420 -10885
rect 31465 -11005 31585 -10885
rect 31640 -11005 31760 -10885
rect 31805 -11005 31925 -10885
rect 31970 -11005 32090 -10885
rect 32135 -11005 32255 -10885
rect 32310 -11005 32430 -10885
rect 32475 -11005 32595 -10885
rect 32640 -11005 32760 -10885
rect 32805 -11005 32925 -10885
rect 32980 -11005 33100 -10885
rect 33145 -11005 33265 -10885
rect 33310 -11005 33430 -10885
rect 33475 -11005 33595 -10885
rect 33650 -11005 33770 -10885
rect 33815 -11005 33935 -10885
rect 33980 -11005 34100 -10885
rect 34145 -11005 34265 -10885
rect 34320 -11005 34440 -10885
rect 34485 -11005 34605 -10885
rect 34650 -11005 34770 -10885
rect 34815 -11005 34935 -10885
rect 34990 -11005 35110 -10885
rect 35155 -11005 35275 -10885
rect 35320 -11005 35440 -10885
rect 35485 -11005 35605 -10885
rect 35660 -11005 35780 -10885
rect 35825 -11005 35945 -10885
rect 35990 -11005 36110 -10885
rect 36155 -11005 36275 -10885
rect 30795 -11170 30915 -11050
rect 30970 -11170 31090 -11050
rect 31135 -11170 31255 -11050
rect 31300 -11170 31420 -11050
rect 31465 -11170 31585 -11050
rect 31640 -11170 31760 -11050
rect 31805 -11170 31925 -11050
rect 31970 -11170 32090 -11050
rect 32135 -11170 32255 -11050
rect 32310 -11170 32430 -11050
rect 32475 -11170 32595 -11050
rect 32640 -11170 32760 -11050
rect 32805 -11170 32925 -11050
rect 32980 -11170 33100 -11050
rect 33145 -11170 33265 -11050
rect 33310 -11170 33430 -11050
rect 33475 -11170 33595 -11050
rect 33650 -11170 33770 -11050
rect 33815 -11170 33935 -11050
rect 33980 -11170 34100 -11050
rect 34145 -11170 34265 -11050
rect 34320 -11170 34440 -11050
rect 34485 -11170 34605 -11050
rect 34650 -11170 34770 -11050
rect 34815 -11170 34935 -11050
rect 34990 -11170 35110 -11050
rect 35155 -11170 35275 -11050
rect 35320 -11170 35440 -11050
rect 35485 -11170 35605 -11050
rect 35660 -11170 35780 -11050
rect 35825 -11170 35945 -11050
rect 35990 -11170 36110 -11050
rect 36155 -11170 36275 -11050
rect 30795 -11335 30915 -11215
rect 30970 -11335 31090 -11215
rect 31135 -11335 31255 -11215
rect 31300 -11335 31420 -11215
rect 31465 -11335 31585 -11215
rect 31640 -11335 31760 -11215
rect 31805 -11335 31925 -11215
rect 31970 -11335 32090 -11215
rect 32135 -11335 32255 -11215
rect 32310 -11335 32430 -11215
rect 32475 -11335 32595 -11215
rect 32640 -11335 32760 -11215
rect 32805 -11335 32925 -11215
rect 32980 -11335 33100 -11215
rect 33145 -11335 33265 -11215
rect 33310 -11335 33430 -11215
rect 33475 -11335 33595 -11215
rect 33650 -11335 33770 -11215
rect 33815 -11335 33935 -11215
rect 33980 -11335 34100 -11215
rect 34145 -11335 34265 -11215
rect 34320 -11335 34440 -11215
rect 34485 -11335 34605 -11215
rect 34650 -11335 34770 -11215
rect 34815 -11335 34935 -11215
rect 34990 -11335 35110 -11215
rect 35155 -11335 35275 -11215
rect 35320 -11335 35440 -11215
rect 35485 -11335 35605 -11215
rect 35660 -11335 35780 -11215
rect 35825 -11335 35945 -11215
rect 35990 -11335 36110 -11215
rect 36155 -11335 36275 -11215
rect 30795 -11510 30915 -11390
rect 30970 -11510 31090 -11390
rect 31135 -11510 31255 -11390
rect 31300 -11510 31420 -11390
rect 31465 -11510 31585 -11390
rect 31640 -11510 31760 -11390
rect 31805 -11510 31925 -11390
rect 31970 -11510 32090 -11390
rect 32135 -11510 32255 -11390
rect 32310 -11510 32430 -11390
rect 32475 -11510 32595 -11390
rect 32640 -11510 32760 -11390
rect 32805 -11510 32925 -11390
rect 32980 -11510 33100 -11390
rect 33145 -11510 33265 -11390
rect 33310 -11510 33430 -11390
rect 33475 -11510 33595 -11390
rect 33650 -11510 33770 -11390
rect 33815 -11510 33935 -11390
rect 33980 -11510 34100 -11390
rect 34145 -11510 34265 -11390
rect 34320 -11510 34440 -11390
rect 34485 -11510 34605 -11390
rect 34650 -11510 34770 -11390
rect 34815 -11510 34935 -11390
rect 34990 -11510 35110 -11390
rect 35155 -11510 35275 -11390
rect 35320 -11510 35440 -11390
rect 35485 -11510 35605 -11390
rect 35660 -11510 35780 -11390
rect 35825 -11510 35945 -11390
rect 35990 -11510 36110 -11390
rect 36155 -11510 36275 -11390
rect 30795 -11675 30915 -11555
rect 30970 -11675 31090 -11555
rect 31135 -11675 31255 -11555
rect 31300 -11675 31420 -11555
rect 31465 -11675 31585 -11555
rect 31640 -11675 31760 -11555
rect 31805 -11675 31925 -11555
rect 31970 -11675 32090 -11555
rect 32135 -11675 32255 -11555
rect 32310 -11675 32430 -11555
rect 32475 -11675 32595 -11555
rect 32640 -11675 32760 -11555
rect 32805 -11675 32925 -11555
rect 32980 -11675 33100 -11555
rect 33145 -11675 33265 -11555
rect 33310 -11675 33430 -11555
rect 33475 -11675 33595 -11555
rect 33650 -11675 33770 -11555
rect 33815 -11675 33935 -11555
rect 33980 -11675 34100 -11555
rect 34145 -11675 34265 -11555
rect 34320 -11675 34440 -11555
rect 34485 -11675 34605 -11555
rect 34650 -11675 34770 -11555
rect 34815 -11675 34935 -11555
rect 34990 -11675 35110 -11555
rect 35155 -11675 35275 -11555
rect 35320 -11675 35440 -11555
rect 35485 -11675 35605 -11555
rect 35660 -11675 35780 -11555
rect 35825 -11675 35945 -11555
rect 35990 -11675 36110 -11555
rect 36155 -11675 36275 -11555
rect 30795 -11840 30915 -11720
rect 30970 -11840 31090 -11720
rect 31135 -11840 31255 -11720
rect 31300 -11840 31420 -11720
rect 31465 -11840 31585 -11720
rect 31640 -11840 31760 -11720
rect 31805 -11840 31925 -11720
rect 31970 -11840 32090 -11720
rect 32135 -11840 32255 -11720
rect 32310 -11840 32430 -11720
rect 32475 -11840 32595 -11720
rect 32640 -11840 32760 -11720
rect 32805 -11840 32925 -11720
rect 32980 -11840 33100 -11720
rect 33145 -11840 33265 -11720
rect 33310 -11840 33430 -11720
rect 33475 -11840 33595 -11720
rect 33650 -11840 33770 -11720
rect 33815 -11840 33935 -11720
rect 33980 -11840 34100 -11720
rect 34145 -11840 34265 -11720
rect 34320 -11840 34440 -11720
rect 34485 -11840 34605 -11720
rect 34650 -11840 34770 -11720
rect 34815 -11840 34935 -11720
rect 34990 -11840 35110 -11720
rect 35155 -11840 35275 -11720
rect 35320 -11840 35440 -11720
rect 35485 -11840 35605 -11720
rect 35660 -11840 35780 -11720
rect 35825 -11840 35945 -11720
rect 35990 -11840 36110 -11720
rect 36155 -11840 36275 -11720
rect 30795 -12005 30915 -11885
rect 30970 -12005 31090 -11885
rect 31135 -12005 31255 -11885
rect 31300 -12005 31420 -11885
rect 31465 -12005 31585 -11885
rect 31640 -12005 31760 -11885
rect 31805 -12005 31925 -11885
rect 31970 -12005 32090 -11885
rect 32135 -12005 32255 -11885
rect 32310 -12005 32430 -11885
rect 32475 -12005 32595 -11885
rect 32640 -12005 32760 -11885
rect 32805 -12005 32925 -11885
rect 32980 -12005 33100 -11885
rect 33145 -12005 33265 -11885
rect 33310 -12005 33430 -11885
rect 33475 -12005 33595 -11885
rect 33650 -12005 33770 -11885
rect 33815 -12005 33935 -11885
rect 33980 -12005 34100 -11885
rect 34145 -12005 34265 -11885
rect 34320 -12005 34440 -11885
rect 34485 -12005 34605 -11885
rect 34650 -12005 34770 -11885
rect 34815 -12005 34935 -11885
rect 34990 -12005 35110 -11885
rect 35155 -12005 35275 -11885
rect 35320 -12005 35440 -11885
rect 35485 -12005 35605 -11885
rect 35660 -12005 35780 -11885
rect 35825 -12005 35945 -11885
rect 35990 -12005 36110 -11885
rect 36155 -12005 36275 -11885
rect 30795 -12180 30915 -12060
rect 30970 -12180 31090 -12060
rect 31135 -12180 31255 -12060
rect 31300 -12180 31420 -12060
rect 31465 -12180 31585 -12060
rect 31640 -12180 31760 -12060
rect 31805 -12180 31925 -12060
rect 31970 -12180 32090 -12060
rect 32135 -12180 32255 -12060
rect 32310 -12180 32430 -12060
rect 32475 -12180 32595 -12060
rect 32640 -12180 32760 -12060
rect 32805 -12180 32925 -12060
rect 32980 -12180 33100 -12060
rect 33145 -12180 33265 -12060
rect 33310 -12180 33430 -12060
rect 33475 -12180 33595 -12060
rect 33650 -12180 33770 -12060
rect 33815 -12180 33935 -12060
rect 33980 -12180 34100 -12060
rect 34145 -12180 34265 -12060
rect 34320 -12180 34440 -12060
rect 34485 -12180 34605 -12060
rect 34650 -12180 34770 -12060
rect 34815 -12180 34935 -12060
rect 34990 -12180 35110 -12060
rect 35155 -12180 35275 -12060
rect 35320 -12180 35440 -12060
rect 35485 -12180 35605 -12060
rect 35660 -12180 35780 -12060
rect 35825 -12180 35945 -12060
rect 35990 -12180 36110 -12060
rect 36155 -12180 36275 -12060
rect 30795 -12345 30915 -12225
rect 30970 -12345 31090 -12225
rect 31135 -12345 31255 -12225
rect 31300 -12345 31420 -12225
rect 31465 -12345 31585 -12225
rect 31640 -12345 31760 -12225
rect 31805 -12345 31925 -12225
rect 31970 -12345 32090 -12225
rect 32135 -12345 32255 -12225
rect 32310 -12345 32430 -12225
rect 32475 -12345 32595 -12225
rect 32640 -12345 32760 -12225
rect 32805 -12345 32925 -12225
rect 32980 -12345 33100 -12225
rect 33145 -12345 33265 -12225
rect 33310 -12345 33430 -12225
rect 33475 -12345 33595 -12225
rect 33650 -12345 33770 -12225
rect 33815 -12345 33935 -12225
rect 33980 -12345 34100 -12225
rect 34145 -12345 34265 -12225
rect 34320 -12345 34440 -12225
rect 34485 -12345 34605 -12225
rect 34650 -12345 34770 -12225
rect 34815 -12345 34935 -12225
rect 34990 -12345 35110 -12225
rect 35155 -12345 35275 -12225
rect 35320 -12345 35440 -12225
rect 35485 -12345 35605 -12225
rect 35660 -12345 35780 -12225
rect 35825 -12345 35945 -12225
rect 35990 -12345 36110 -12225
rect 36155 -12345 36275 -12225
rect 30795 -12510 30915 -12390
rect 30970 -12510 31090 -12390
rect 31135 -12510 31255 -12390
rect 31300 -12510 31420 -12390
rect 31465 -12510 31585 -12390
rect 31640 -12510 31760 -12390
rect 31805 -12510 31925 -12390
rect 31970 -12510 32090 -12390
rect 32135 -12510 32255 -12390
rect 32310 -12510 32430 -12390
rect 32475 -12510 32595 -12390
rect 32640 -12510 32760 -12390
rect 32805 -12510 32925 -12390
rect 32980 -12510 33100 -12390
rect 33145 -12510 33265 -12390
rect 33310 -12510 33430 -12390
rect 33475 -12510 33595 -12390
rect 33650 -12510 33770 -12390
rect 33815 -12510 33935 -12390
rect 33980 -12510 34100 -12390
rect 34145 -12510 34265 -12390
rect 34320 -12510 34440 -12390
rect 34485 -12510 34605 -12390
rect 34650 -12510 34770 -12390
rect 34815 -12510 34935 -12390
rect 34990 -12510 35110 -12390
rect 35155 -12510 35275 -12390
rect 35320 -12510 35440 -12390
rect 35485 -12510 35605 -12390
rect 35660 -12510 35780 -12390
rect 35825 -12510 35945 -12390
rect 35990 -12510 36110 -12390
rect 36155 -12510 36275 -12390
rect 30795 -12675 30915 -12555
rect 30970 -12675 31090 -12555
rect 31135 -12675 31255 -12555
rect 31300 -12675 31420 -12555
rect 31465 -12675 31585 -12555
rect 31640 -12675 31760 -12555
rect 31805 -12675 31925 -12555
rect 31970 -12675 32090 -12555
rect 32135 -12675 32255 -12555
rect 32310 -12675 32430 -12555
rect 32475 -12675 32595 -12555
rect 32640 -12675 32760 -12555
rect 32805 -12675 32925 -12555
rect 32980 -12675 33100 -12555
rect 33145 -12675 33265 -12555
rect 33310 -12675 33430 -12555
rect 33475 -12675 33595 -12555
rect 33650 -12675 33770 -12555
rect 33815 -12675 33935 -12555
rect 33980 -12675 34100 -12555
rect 34145 -12675 34265 -12555
rect 34320 -12675 34440 -12555
rect 34485 -12675 34605 -12555
rect 34650 -12675 34770 -12555
rect 34815 -12675 34935 -12555
rect 34990 -12675 35110 -12555
rect 35155 -12675 35275 -12555
rect 35320 -12675 35440 -12555
rect 35485 -12675 35605 -12555
rect 35660 -12675 35780 -12555
rect 35825 -12675 35945 -12555
rect 35990 -12675 36110 -12555
rect 36155 -12675 36275 -12555
rect 30795 -12850 30915 -12730
rect 30970 -12850 31090 -12730
rect 31135 -12850 31255 -12730
rect 31300 -12850 31420 -12730
rect 31465 -12850 31585 -12730
rect 31640 -12850 31760 -12730
rect 31805 -12850 31925 -12730
rect 31970 -12850 32090 -12730
rect 32135 -12850 32255 -12730
rect 32310 -12850 32430 -12730
rect 32475 -12850 32595 -12730
rect 32640 -12850 32760 -12730
rect 32805 -12850 32925 -12730
rect 32980 -12850 33100 -12730
rect 33145 -12850 33265 -12730
rect 33310 -12850 33430 -12730
rect 33475 -12850 33595 -12730
rect 33650 -12850 33770 -12730
rect 33815 -12850 33935 -12730
rect 33980 -12850 34100 -12730
rect 34145 -12850 34265 -12730
rect 34320 -12850 34440 -12730
rect 34485 -12850 34605 -12730
rect 34650 -12850 34770 -12730
rect 34815 -12850 34935 -12730
rect 34990 -12850 35110 -12730
rect 35155 -12850 35275 -12730
rect 35320 -12850 35440 -12730
rect 35485 -12850 35605 -12730
rect 35660 -12850 35780 -12730
rect 35825 -12850 35945 -12730
rect 35990 -12850 36110 -12730
rect 36155 -12850 36275 -12730
rect 30795 -13015 30915 -12895
rect 30970 -13015 31090 -12895
rect 31135 -13015 31255 -12895
rect 31300 -13015 31420 -12895
rect 31465 -13015 31585 -12895
rect 31640 -13015 31760 -12895
rect 31805 -13015 31925 -12895
rect 31970 -13015 32090 -12895
rect 32135 -13015 32255 -12895
rect 32310 -13015 32430 -12895
rect 32475 -13015 32595 -12895
rect 32640 -13015 32760 -12895
rect 32805 -13015 32925 -12895
rect 32980 -13015 33100 -12895
rect 33145 -13015 33265 -12895
rect 33310 -13015 33430 -12895
rect 33475 -13015 33595 -12895
rect 33650 -13015 33770 -12895
rect 33815 -13015 33935 -12895
rect 33980 -13015 34100 -12895
rect 34145 -13015 34265 -12895
rect 34320 -13015 34440 -12895
rect 34485 -13015 34605 -12895
rect 34650 -13015 34770 -12895
rect 34815 -13015 34935 -12895
rect 34990 -13015 35110 -12895
rect 35155 -13015 35275 -12895
rect 35320 -13015 35440 -12895
rect 35485 -13015 35605 -12895
rect 35660 -13015 35780 -12895
rect 35825 -13015 35945 -12895
rect 35990 -13015 36110 -12895
rect 36155 -13015 36275 -12895
rect 30795 -13180 30915 -13060
rect 30970 -13180 31090 -13060
rect 31135 -13180 31255 -13060
rect 31300 -13180 31420 -13060
rect 31465 -13180 31585 -13060
rect 31640 -13180 31760 -13060
rect 31805 -13180 31925 -13060
rect 31970 -13180 32090 -13060
rect 32135 -13180 32255 -13060
rect 32310 -13180 32430 -13060
rect 32475 -13180 32595 -13060
rect 32640 -13180 32760 -13060
rect 32805 -13180 32925 -13060
rect 32980 -13180 33100 -13060
rect 33145 -13180 33265 -13060
rect 33310 -13180 33430 -13060
rect 33475 -13180 33595 -13060
rect 33650 -13180 33770 -13060
rect 33815 -13180 33935 -13060
rect 33980 -13180 34100 -13060
rect 34145 -13180 34265 -13060
rect 34320 -13180 34440 -13060
rect 34485 -13180 34605 -13060
rect 34650 -13180 34770 -13060
rect 34815 -13180 34935 -13060
rect 34990 -13180 35110 -13060
rect 35155 -13180 35275 -13060
rect 35320 -13180 35440 -13060
rect 35485 -13180 35605 -13060
rect 35660 -13180 35780 -13060
rect 35825 -13180 35945 -13060
rect 35990 -13180 36110 -13060
rect 36155 -13180 36275 -13060
rect 30795 -13345 30915 -13225
rect 30970 -13345 31090 -13225
rect 31135 -13345 31255 -13225
rect 31300 -13345 31420 -13225
rect 31465 -13345 31585 -13225
rect 31640 -13345 31760 -13225
rect 31805 -13345 31925 -13225
rect 31970 -13345 32090 -13225
rect 32135 -13345 32255 -13225
rect 32310 -13345 32430 -13225
rect 32475 -13345 32595 -13225
rect 32640 -13345 32760 -13225
rect 32805 -13345 32925 -13225
rect 32980 -13345 33100 -13225
rect 33145 -13345 33265 -13225
rect 33310 -13345 33430 -13225
rect 33475 -13345 33595 -13225
rect 33650 -13345 33770 -13225
rect 33815 -13345 33935 -13225
rect 33980 -13345 34100 -13225
rect 34145 -13345 34265 -13225
rect 34320 -13345 34440 -13225
rect 34485 -13345 34605 -13225
rect 34650 -13345 34770 -13225
rect 34815 -13345 34935 -13225
rect 34990 -13345 35110 -13225
rect 35155 -13345 35275 -13225
rect 35320 -13345 35440 -13225
rect 35485 -13345 35605 -13225
rect 35660 -13345 35780 -13225
rect 35825 -13345 35945 -13225
rect 35990 -13345 36110 -13225
rect 36155 -13345 36275 -13225
rect 30795 -13520 30915 -13400
rect 30970 -13520 31090 -13400
rect 31135 -13520 31255 -13400
rect 31300 -13520 31420 -13400
rect 31465 -13520 31585 -13400
rect 31640 -13520 31760 -13400
rect 31805 -13520 31925 -13400
rect 31970 -13520 32090 -13400
rect 32135 -13520 32255 -13400
rect 32310 -13520 32430 -13400
rect 32475 -13520 32595 -13400
rect 32640 -13520 32760 -13400
rect 32805 -13520 32925 -13400
rect 32980 -13520 33100 -13400
rect 33145 -13520 33265 -13400
rect 33310 -13520 33430 -13400
rect 33475 -13520 33595 -13400
rect 33650 -13520 33770 -13400
rect 33815 -13520 33935 -13400
rect 33980 -13520 34100 -13400
rect 34145 -13520 34265 -13400
rect 34320 -13520 34440 -13400
rect 34485 -13520 34605 -13400
rect 34650 -13520 34770 -13400
rect 34815 -13520 34935 -13400
rect 34990 -13520 35110 -13400
rect 35155 -13520 35275 -13400
rect 35320 -13520 35440 -13400
rect 35485 -13520 35605 -13400
rect 35660 -13520 35780 -13400
rect 35825 -13520 35945 -13400
rect 35990 -13520 36110 -13400
rect 36155 -13520 36275 -13400
rect 30795 -13685 30915 -13565
rect 30970 -13685 31090 -13565
rect 31135 -13685 31255 -13565
rect 31300 -13685 31420 -13565
rect 31465 -13685 31585 -13565
rect 31640 -13685 31760 -13565
rect 31805 -13685 31925 -13565
rect 31970 -13685 32090 -13565
rect 32135 -13685 32255 -13565
rect 32310 -13685 32430 -13565
rect 32475 -13685 32595 -13565
rect 32640 -13685 32760 -13565
rect 32805 -13685 32925 -13565
rect 32980 -13685 33100 -13565
rect 33145 -13685 33265 -13565
rect 33310 -13685 33430 -13565
rect 33475 -13685 33595 -13565
rect 33650 -13685 33770 -13565
rect 33815 -13685 33935 -13565
rect 33980 -13685 34100 -13565
rect 34145 -13685 34265 -13565
rect 34320 -13685 34440 -13565
rect 34485 -13685 34605 -13565
rect 34650 -13685 34770 -13565
rect 34815 -13685 34935 -13565
rect 34990 -13685 35110 -13565
rect 35155 -13685 35275 -13565
rect 35320 -13685 35440 -13565
rect 35485 -13685 35605 -13565
rect 35660 -13685 35780 -13565
rect 35825 -13685 35945 -13565
rect 35990 -13685 36110 -13565
rect 36155 -13685 36275 -13565
rect 30795 -13850 30915 -13730
rect 30970 -13850 31090 -13730
rect 31135 -13850 31255 -13730
rect 31300 -13850 31420 -13730
rect 31465 -13850 31585 -13730
rect 31640 -13850 31760 -13730
rect 31805 -13850 31925 -13730
rect 31970 -13850 32090 -13730
rect 32135 -13850 32255 -13730
rect 32310 -13850 32430 -13730
rect 32475 -13850 32595 -13730
rect 32640 -13850 32760 -13730
rect 32805 -13850 32925 -13730
rect 32980 -13850 33100 -13730
rect 33145 -13850 33265 -13730
rect 33310 -13850 33430 -13730
rect 33475 -13850 33595 -13730
rect 33650 -13850 33770 -13730
rect 33815 -13850 33935 -13730
rect 33980 -13850 34100 -13730
rect 34145 -13850 34265 -13730
rect 34320 -13850 34440 -13730
rect 34485 -13850 34605 -13730
rect 34650 -13850 34770 -13730
rect 34815 -13850 34935 -13730
rect 34990 -13850 35110 -13730
rect 35155 -13850 35275 -13730
rect 35320 -13850 35440 -13730
rect 35485 -13850 35605 -13730
rect 35660 -13850 35780 -13730
rect 35825 -13850 35945 -13730
rect 35990 -13850 36110 -13730
rect 36155 -13850 36275 -13730
rect 30795 -14015 30915 -13895
rect 30970 -14015 31090 -13895
rect 31135 -14015 31255 -13895
rect 31300 -14015 31420 -13895
rect 31465 -14015 31585 -13895
rect 31640 -14015 31760 -13895
rect 31805 -14015 31925 -13895
rect 31970 -14015 32090 -13895
rect 32135 -14015 32255 -13895
rect 32310 -14015 32430 -13895
rect 32475 -14015 32595 -13895
rect 32640 -14015 32760 -13895
rect 32805 -14015 32925 -13895
rect 32980 -14015 33100 -13895
rect 33145 -14015 33265 -13895
rect 33310 -14015 33430 -13895
rect 33475 -14015 33595 -13895
rect 33650 -14015 33770 -13895
rect 33815 -14015 33935 -13895
rect 33980 -14015 34100 -13895
rect 34145 -14015 34265 -13895
rect 34320 -14015 34440 -13895
rect 34485 -14015 34605 -13895
rect 34650 -14015 34770 -13895
rect 34815 -14015 34935 -13895
rect 34990 -14015 35110 -13895
rect 35155 -14015 35275 -13895
rect 35320 -14015 35440 -13895
rect 35485 -14015 35605 -13895
rect 35660 -14015 35780 -13895
rect 35825 -14015 35945 -13895
rect 35990 -14015 36110 -13895
rect 36155 -14015 36275 -13895
rect 30795 -14190 30915 -14070
rect 30970 -14190 31090 -14070
rect 31135 -14190 31255 -14070
rect 31300 -14190 31420 -14070
rect 31465 -14190 31585 -14070
rect 31640 -14190 31760 -14070
rect 31805 -14190 31925 -14070
rect 31970 -14190 32090 -14070
rect 32135 -14190 32255 -14070
rect 32310 -14190 32430 -14070
rect 32475 -14190 32595 -14070
rect 32640 -14190 32760 -14070
rect 32805 -14190 32925 -14070
rect 32980 -14190 33100 -14070
rect 33145 -14190 33265 -14070
rect 33310 -14190 33430 -14070
rect 33475 -14190 33595 -14070
rect 33650 -14190 33770 -14070
rect 33815 -14190 33935 -14070
rect 33980 -14190 34100 -14070
rect 34145 -14190 34265 -14070
rect 34320 -14190 34440 -14070
rect 34485 -14190 34605 -14070
rect 34650 -14190 34770 -14070
rect 34815 -14190 34935 -14070
rect 34990 -14190 35110 -14070
rect 35155 -14190 35275 -14070
rect 35320 -14190 35440 -14070
rect 35485 -14190 35605 -14070
rect 35660 -14190 35780 -14070
rect 35825 -14190 35945 -14070
rect 35990 -14190 36110 -14070
rect 36155 -14190 36275 -14070
rect 30795 -14355 30915 -14235
rect 30970 -14355 31090 -14235
rect 31135 -14355 31255 -14235
rect 31300 -14355 31420 -14235
rect 31465 -14355 31585 -14235
rect 31640 -14355 31760 -14235
rect 31805 -14355 31925 -14235
rect 31970 -14355 32090 -14235
rect 32135 -14355 32255 -14235
rect 32310 -14355 32430 -14235
rect 32475 -14355 32595 -14235
rect 32640 -14355 32760 -14235
rect 32805 -14355 32925 -14235
rect 32980 -14355 33100 -14235
rect 33145 -14355 33265 -14235
rect 33310 -14355 33430 -14235
rect 33475 -14355 33595 -14235
rect 33650 -14355 33770 -14235
rect 33815 -14355 33935 -14235
rect 33980 -14355 34100 -14235
rect 34145 -14355 34265 -14235
rect 34320 -14355 34440 -14235
rect 34485 -14355 34605 -14235
rect 34650 -14355 34770 -14235
rect 34815 -14355 34935 -14235
rect 34990 -14355 35110 -14235
rect 35155 -14355 35275 -14235
rect 35320 -14355 35440 -14235
rect 35485 -14355 35605 -14235
rect 35660 -14355 35780 -14235
rect 35825 -14355 35945 -14235
rect 35990 -14355 36110 -14235
rect 36155 -14355 36275 -14235
rect 30795 -14520 30915 -14400
rect 30970 -14520 31090 -14400
rect 31135 -14520 31255 -14400
rect 31300 -14520 31420 -14400
rect 31465 -14520 31585 -14400
rect 31640 -14520 31760 -14400
rect 31805 -14520 31925 -14400
rect 31970 -14520 32090 -14400
rect 32135 -14520 32255 -14400
rect 32310 -14520 32430 -14400
rect 32475 -14520 32595 -14400
rect 32640 -14520 32760 -14400
rect 32805 -14520 32925 -14400
rect 32980 -14520 33100 -14400
rect 33145 -14520 33265 -14400
rect 33310 -14520 33430 -14400
rect 33475 -14520 33595 -14400
rect 33650 -14520 33770 -14400
rect 33815 -14520 33935 -14400
rect 33980 -14520 34100 -14400
rect 34145 -14520 34265 -14400
rect 34320 -14520 34440 -14400
rect 34485 -14520 34605 -14400
rect 34650 -14520 34770 -14400
rect 34815 -14520 34935 -14400
rect 34990 -14520 35110 -14400
rect 35155 -14520 35275 -14400
rect 35320 -14520 35440 -14400
rect 35485 -14520 35605 -14400
rect 35660 -14520 35780 -14400
rect 35825 -14520 35945 -14400
rect 35990 -14520 36110 -14400
rect 36155 -14520 36275 -14400
rect 30795 -14685 30915 -14565
rect 30970 -14685 31090 -14565
rect 31135 -14685 31255 -14565
rect 31300 -14685 31420 -14565
rect 31465 -14685 31585 -14565
rect 31640 -14685 31760 -14565
rect 31805 -14685 31925 -14565
rect 31970 -14685 32090 -14565
rect 32135 -14685 32255 -14565
rect 32310 -14685 32430 -14565
rect 32475 -14685 32595 -14565
rect 32640 -14685 32760 -14565
rect 32805 -14685 32925 -14565
rect 32980 -14685 33100 -14565
rect 33145 -14685 33265 -14565
rect 33310 -14685 33430 -14565
rect 33475 -14685 33595 -14565
rect 33650 -14685 33770 -14565
rect 33815 -14685 33935 -14565
rect 33980 -14685 34100 -14565
rect 34145 -14685 34265 -14565
rect 34320 -14685 34440 -14565
rect 34485 -14685 34605 -14565
rect 34650 -14685 34770 -14565
rect 34815 -14685 34935 -14565
rect 34990 -14685 35110 -14565
rect 35155 -14685 35275 -14565
rect 35320 -14685 35440 -14565
rect 35485 -14685 35605 -14565
rect 35660 -14685 35780 -14565
rect 35825 -14685 35945 -14565
rect 35990 -14685 36110 -14565
rect 36155 -14685 36275 -14565
rect 30795 -14860 30915 -14740
rect 30970 -14860 31090 -14740
rect 31135 -14860 31255 -14740
rect 31300 -14860 31420 -14740
rect 31465 -14860 31585 -14740
rect 31640 -14860 31760 -14740
rect 31805 -14860 31925 -14740
rect 31970 -14860 32090 -14740
rect 32135 -14860 32255 -14740
rect 32310 -14860 32430 -14740
rect 32475 -14860 32595 -14740
rect 32640 -14860 32760 -14740
rect 32805 -14860 32925 -14740
rect 32980 -14860 33100 -14740
rect 33145 -14860 33265 -14740
rect 33310 -14860 33430 -14740
rect 33475 -14860 33595 -14740
rect 33650 -14860 33770 -14740
rect 33815 -14860 33935 -14740
rect 33980 -14860 34100 -14740
rect 34145 -14860 34265 -14740
rect 34320 -14860 34440 -14740
rect 34485 -14860 34605 -14740
rect 34650 -14860 34770 -14740
rect 34815 -14860 34935 -14740
rect 34990 -14860 35110 -14740
rect 35155 -14860 35275 -14740
rect 35320 -14860 35440 -14740
rect 35485 -14860 35605 -14740
rect 35660 -14860 35780 -14740
rect 35825 -14860 35945 -14740
rect 35990 -14860 36110 -14740
rect 36155 -14860 36275 -14740
rect 30795 -15025 30915 -14905
rect 30970 -15025 31090 -14905
rect 31135 -15025 31255 -14905
rect 31300 -15025 31420 -14905
rect 31465 -15025 31585 -14905
rect 31640 -15025 31760 -14905
rect 31805 -15025 31925 -14905
rect 31970 -15025 32090 -14905
rect 32135 -15025 32255 -14905
rect 32310 -15025 32430 -14905
rect 32475 -15025 32595 -14905
rect 32640 -15025 32760 -14905
rect 32805 -15025 32925 -14905
rect 32980 -15025 33100 -14905
rect 33145 -15025 33265 -14905
rect 33310 -15025 33430 -14905
rect 33475 -15025 33595 -14905
rect 33650 -15025 33770 -14905
rect 33815 -15025 33935 -14905
rect 33980 -15025 34100 -14905
rect 34145 -15025 34265 -14905
rect 34320 -15025 34440 -14905
rect 34485 -15025 34605 -14905
rect 34650 -15025 34770 -14905
rect 34815 -15025 34935 -14905
rect 34990 -15025 35110 -14905
rect 35155 -15025 35275 -14905
rect 35320 -15025 35440 -14905
rect 35485 -15025 35605 -14905
rect 35660 -15025 35780 -14905
rect 35825 -15025 35945 -14905
rect 35990 -15025 36110 -14905
rect 36155 -15025 36275 -14905
rect 30795 -15190 30915 -15070
rect 30970 -15190 31090 -15070
rect 31135 -15190 31255 -15070
rect 31300 -15190 31420 -15070
rect 31465 -15190 31585 -15070
rect 31640 -15190 31760 -15070
rect 31805 -15190 31925 -15070
rect 31970 -15190 32090 -15070
rect 32135 -15190 32255 -15070
rect 32310 -15190 32430 -15070
rect 32475 -15190 32595 -15070
rect 32640 -15190 32760 -15070
rect 32805 -15190 32925 -15070
rect 32980 -15190 33100 -15070
rect 33145 -15190 33265 -15070
rect 33310 -15190 33430 -15070
rect 33475 -15190 33595 -15070
rect 33650 -15190 33770 -15070
rect 33815 -15190 33935 -15070
rect 33980 -15190 34100 -15070
rect 34145 -15190 34265 -15070
rect 34320 -15190 34440 -15070
rect 34485 -15190 34605 -15070
rect 34650 -15190 34770 -15070
rect 34815 -15190 34935 -15070
rect 34990 -15190 35110 -15070
rect 35155 -15190 35275 -15070
rect 35320 -15190 35440 -15070
rect 35485 -15190 35605 -15070
rect 35660 -15190 35780 -15070
rect 35825 -15190 35945 -15070
rect 35990 -15190 36110 -15070
rect 36155 -15190 36275 -15070
rect 30795 -15355 30915 -15235
rect 30970 -15355 31090 -15235
rect 31135 -15355 31255 -15235
rect 31300 -15355 31420 -15235
rect 31465 -15355 31585 -15235
rect 31640 -15355 31760 -15235
rect 31805 -15355 31925 -15235
rect 31970 -15355 32090 -15235
rect 32135 -15355 32255 -15235
rect 32310 -15355 32430 -15235
rect 32475 -15355 32595 -15235
rect 32640 -15355 32760 -15235
rect 32805 -15355 32925 -15235
rect 32980 -15355 33100 -15235
rect 33145 -15355 33265 -15235
rect 33310 -15355 33430 -15235
rect 33475 -15355 33595 -15235
rect 33650 -15355 33770 -15235
rect 33815 -15355 33935 -15235
rect 33980 -15355 34100 -15235
rect 34145 -15355 34265 -15235
rect 34320 -15355 34440 -15235
rect 34485 -15355 34605 -15235
rect 34650 -15355 34770 -15235
rect 34815 -15355 34935 -15235
rect 34990 -15355 35110 -15235
rect 35155 -15355 35275 -15235
rect 35320 -15355 35440 -15235
rect 35485 -15355 35605 -15235
rect 35660 -15355 35780 -15235
rect 35825 -15355 35945 -15235
rect 35990 -15355 36110 -15235
rect 36155 -15355 36275 -15235
rect 30795 -15530 30915 -15410
rect 30970 -15530 31090 -15410
rect 31135 -15530 31255 -15410
rect 31300 -15530 31420 -15410
rect 31465 -15530 31585 -15410
rect 31640 -15530 31760 -15410
rect 31805 -15530 31925 -15410
rect 31970 -15530 32090 -15410
rect 32135 -15530 32255 -15410
rect 32310 -15530 32430 -15410
rect 32475 -15530 32595 -15410
rect 32640 -15530 32760 -15410
rect 32805 -15530 32925 -15410
rect 32980 -15530 33100 -15410
rect 33145 -15530 33265 -15410
rect 33310 -15530 33430 -15410
rect 33475 -15530 33595 -15410
rect 33650 -15530 33770 -15410
rect 33815 -15530 33935 -15410
rect 33980 -15530 34100 -15410
rect 34145 -15530 34265 -15410
rect 34320 -15530 34440 -15410
rect 34485 -15530 34605 -15410
rect 34650 -15530 34770 -15410
rect 34815 -15530 34935 -15410
rect 34990 -15530 35110 -15410
rect 35155 -15530 35275 -15410
rect 35320 -15530 35440 -15410
rect 35485 -15530 35605 -15410
rect 35660 -15530 35780 -15410
rect 35825 -15530 35945 -15410
rect 35990 -15530 36110 -15410
rect 36155 -15530 36275 -15410
rect 36485 -10170 36605 -10050
rect 36660 -10170 36780 -10050
rect 36825 -10170 36945 -10050
rect 36990 -10170 37110 -10050
rect 37155 -10170 37275 -10050
rect 37330 -10170 37450 -10050
rect 37495 -10170 37615 -10050
rect 37660 -10170 37780 -10050
rect 37825 -10170 37945 -10050
rect 38000 -10170 38120 -10050
rect 38165 -10170 38285 -10050
rect 38330 -10170 38450 -10050
rect 38495 -10170 38615 -10050
rect 38670 -10170 38790 -10050
rect 38835 -10170 38955 -10050
rect 39000 -10170 39120 -10050
rect 39165 -10170 39285 -10050
rect 39340 -10170 39460 -10050
rect 39505 -10170 39625 -10050
rect 39670 -10170 39790 -10050
rect 39835 -10170 39955 -10050
rect 40010 -10170 40130 -10050
rect 40175 -10170 40295 -10050
rect 40340 -10170 40460 -10050
rect 40505 -10170 40625 -10050
rect 40680 -10170 40800 -10050
rect 40845 -10170 40965 -10050
rect 41010 -10170 41130 -10050
rect 41175 -10170 41295 -10050
rect 41350 -10170 41470 -10050
rect 41515 -10170 41635 -10050
rect 41680 -10170 41800 -10050
rect 41845 -10170 41965 -10050
rect 36485 -10335 36605 -10215
rect 36660 -10335 36780 -10215
rect 36825 -10335 36945 -10215
rect 36990 -10335 37110 -10215
rect 37155 -10335 37275 -10215
rect 37330 -10335 37450 -10215
rect 37495 -10335 37615 -10215
rect 37660 -10335 37780 -10215
rect 37825 -10335 37945 -10215
rect 38000 -10335 38120 -10215
rect 38165 -10335 38285 -10215
rect 38330 -10335 38450 -10215
rect 38495 -10335 38615 -10215
rect 38670 -10335 38790 -10215
rect 38835 -10335 38955 -10215
rect 39000 -10335 39120 -10215
rect 39165 -10335 39285 -10215
rect 39340 -10335 39460 -10215
rect 39505 -10335 39625 -10215
rect 39670 -10335 39790 -10215
rect 39835 -10335 39955 -10215
rect 40010 -10335 40130 -10215
rect 40175 -10335 40295 -10215
rect 40340 -10335 40460 -10215
rect 40505 -10335 40625 -10215
rect 40680 -10335 40800 -10215
rect 40845 -10335 40965 -10215
rect 41010 -10335 41130 -10215
rect 41175 -10335 41295 -10215
rect 41350 -10335 41470 -10215
rect 41515 -10335 41635 -10215
rect 41680 -10335 41800 -10215
rect 41845 -10335 41965 -10215
rect 36485 -10500 36605 -10380
rect 36660 -10500 36780 -10380
rect 36825 -10500 36945 -10380
rect 36990 -10500 37110 -10380
rect 37155 -10500 37275 -10380
rect 37330 -10500 37450 -10380
rect 37495 -10500 37615 -10380
rect 37660 -10500 37780 -10380
rect 37825 -10500 37945 -10380
rect 38000 -10500 38120 -10380
rect 38165 -10500 38285 -10380
rect 38330 -10500 38450 -10380
rect 38495 -10500 38615 -10380
rect 38670 -10500 38790 -10380
rect 38835 -10500 38955 -10380
rect 39000 -10500 39120 -10380
rect 39165 -10500 39285 -10380
rect 39340 -10500 39460 -10380
rect 39505 -10500 39625 -10380
rect 39670 -10500 39790 -10380
rect 39835 -10500 39955 -10380
rect 40010 -10500 40130 -10380
rect 40175 -10500 40295 -10380
rect 40340 -10500 40460 -10380
rect 40505 -10500 40625 -10380
rect 40680 -10500 40800 -10380
rect 40845 -10500 40965 -10380
rect 41010 -10500 41130 -10380
rect 41175 -10500 41295 -10380
rect 41350 -10500 41470 -10380
rect 41515 -10500 41635 -10380
rect 41680 -10500 41800 -10380
rect 41845 -10500 41965 -10380
rect 36485 -10665 36605 -10545
rect 36660 -10665 36780 -10545
rect 36825 -10665 36945 -10545
rect 36990 -10665 37110 -10545
rect 37155 -10665 37275 -10545
rect 37330 -10665 37450 -10545
rect 37495 -10665 37615 -10545
rect 37660 -10665 37780 -10545
rect 37825 -10665 37945 -10545
rect 38000 -10665 38120 -10545
rect 38165 -10665 38285 -10545
rect 38330 -10665 38450 -10545
rect 38495 -10665 38615 -10545
rect 38670 -10665 38790 -10545
rect 38835 -10665 38955 -10545
rect 39000 -10665 39120 -10545
rect 39165 -10665 39285 -10545
rect 39340 -10665 39460 -10545
rect 39505 -10665 39625 -10545
rect 39670 -10665 39790 -10545
rect 39835 -10665 39955 -10545
rect 40010 -10665 40130 -10545
rect 40175 -10665 40295 -10545
rect 40340 -10665 40460 -10545
rect 40505 -10665 40625 -10545
rect 40680 -10665 40800 -10545
rect 40845 -10665 40965 -10545
rect 41010 -10665 41130 -10545
rect 41175 -10665 41295 -10545
rect 41350 -10665 41470 -10545
rect 41515 -10665 41635 -10545
rect 41680 -10665 41800 -10545
rect 41845 -10665 41965 -10545
rect 36485 -10840 36605 -10720
rect 36660 -10840 36780 -10720
rect 36825 -10840 36945 -10720
rect 36990 -10840 37110 -10720
rect 37155 -10840 37275 -10720
rect 37330 -10840 37450 -10720
rect 37495 -10840 37615 -10720
rect 37660 -10840 37780 -10720
rect 37825 -10840 37945 -10720
rect 38000 -10840 38120 -10720
rect 38165 -10840 38285 -10720
rect 38330 -10840 38450 -10720
rect 38495 -10840 38615 -10720
rect 38670 -10840 38790 -10720
rect 38835 -10840 38955 -10720
rect 39000 -10840 39120 -10720
rect 39165 -10840 39285 -10720
rect 39340 -10840 39460 -10720
rect 39505 -10840 39625 -10720
rect 39670 -10840 39790 -10720
rect 39835 -10840 39955 -10720
rect 40010 -10840 40130 -10720
rect 40175 -10840 40295 -10720
rect 40340 -10840 40460 -10720
rect 40505 -10840 40625 -10720
rect 40680 -10840 40800 -10720
rect 40845 -10840 40965 -10720
rect 41010 -10840 41130 -10720
rect 41175 -10840 41295 -10720
rect 41350 -10840 41470 -10720
rect 41515 -10840 41635 -10720
rect 41680 -10840 41800 -10720
rect 41845 -10840 41965 -10720
rect 36485 -11005 36605 -10885
rect 36660 -11005 36780 -10885
rect 36825 -11005 36945 -10885
rect 36990 -11005 37110 -10885
rect 37155 -11005 37275 -10885
rect 37330 -11005 37450 -10885
rect 37495 -11005 37615 -10885
rect 37660 -11005 37780 -10885
rect 37825 -11005 37945 -10885
rect 38000 -11005 38120 -10885
rect 38165 -11005 38285 -10885
rect 38330 -11005 38450 -10885
rect 38495 -11005 38615 -10885
rect 38670 -11005 38790 -10885
rect 38835 -11005 38955 -10885
rect 39000 -11005 39120 -10885
rect 39165 -11005 39285 -10885
rect 39340 -11005 39460 -10885
rect 39505 -11005 39625 -10885
rect 39670 -11005 39790 -10885
rect 39835 -11005 39955 -10885
rect 40010 -11005 40130 -10885
rect 40175 -11005 40295 -10885
rect 40340 -11005 40460 -10885
rect 40505 -11005 40625 -10885
rect 40680 -11005 40800 -10885
rect 40845 -11005 40965 -10885
rect 41010 -11005 41130 -10885
rect 41175 -11005 41295 -10885
rect 41350 -11005 41470 -10885
rect 41515 -11005 41635 -10885
rect 41680 -11005 41800 -10885
rect 41845 -11005 41965 -10885
rect 36485 -11170 36605 -11050
rect 36660 -11170 36780 -11050
rect 36825 -11170 36945 -11050
rect 36990 -11170 37110 -11050
rect 37155 -11170 37275 -11050
rect 37330 -11170 37450 -11050
rect 37495 -11170 37615 -11050
rect 37660 -11170 37780 -11050
rect 37825 -11170 37945 -11050
rect 38000 -11170 38120 -11050
rect 38165 -11170 38285 -11050
rect 38330 -11170 38450 -11050
rect 38495 -11170 38615 -11050
rect 38670 -11170 38790 -11050
rect 38835 -11170 38955 -11050
rect 39000 -11170 39120 -11050
rect 39165 -11170 39285 -11050
rect 39340 -11170 39460 -11050
rect 39505 -11170 39625 -11050
rect 39670 -11170 39790 -11050
rect 39835 -11170 39955 -11050
rect 40010 -11170 40130 -11050
rect 40175 -11170 40295 -11050
rect 40340 -11170 40460 -11050
rect 40505 -11170 40625 -11050
rect 40680 -11170 40800 -11050
rect 40845 -11170 40965 -11050
rect 41010 -11170 41130 -11050
rect 41175 -11170 41295 -11050
rect 41350 -11170 41470 -11050
rect 41515 -11170 41635 -11050
rect 41680 -11170 41800 -11050
rect 41845 -11170 41965 -11050
rect 36485 -11335 36605 -11215
rect 36660 -11335 36780 -11215
rect 36825 -11335 36945 -11215
rect 36990 -11335 37110 -11215
rect 37155 -11335 37275 -11215
rect 37330 -11335 37450 -11215
rect 37495 -11335 37615 -11215
rect 37660 -11335 37780 -11215
rect 37825 -11335 37945 -11215
rect 38000 -11335 38120 -11215
rect 38165 -11335 38285 -11215
rect 38330 -11335 38450 -11215
rect 38495 -11335 38615 -11215
rect 38670 -11335 38790 -11215
rect 38835 -11335 38955 -11215
rect 39000 -11335 39120 -11215
rect 39165 -11335 39285 -11215
rect 39340 -11335 39460 -11215
rect 39505 -11335 39625 -11215
rect 39670 -11335 39790 -11215
rect 39835 -11335 39955 -11215
rect 40010 -11335 40130 -11215
rect 40175 -11335 40295 -11215
rect 40340 -11335 40460 -11215
rect 40505 -11335 40625 -11215
rect 40680 -11335 40800 -11215
rect 40845 -11335 40965 -11215
rect 41010 -11335 41130 -11215
rect 41175 -11335 41295 -11215
rect 41350 -11335 41470 -11215
rect 41515 -11335 41635 -11215
rect 41680 -11335 41800 -11215
rect 41845 -11335 41965 -11215
rect 36485 -11510 36605 -11390
rect 36660 -11510 36780 -11390
rect 36825 -11510 36945 -11390
rect 36990 -11510 37110 -11390
rect 37155 -11510 37275 -11390
rect 37330 -11510 37450 -11390
rect 37495 -11510 37615 -11390
rect 37660 -11510 37780 -11390
rect 37825 -11510 37945 -11390
rect 38000 -11510 38120 -11390
rect 38165 -11510 38285 -11390
rect 38330 -11510 38450 -11390
rect 38495 -11510 38615 -11390
rect 38670 -11510 38790 -11390
rect 38835 -11510 38955 -11390
rect 39000 -11510 39120 -11390
rect 39165 -11510 39285 -11390
rect 39340 -11510 39460 -11390
rect 39505 -11510 39625 -11390
rect 39670 -11510 39790 -11390
rect 39835 -11510 39955 -11390
rect 40010 -11510 40130 -11390
rect 40175 -11510 40295 -11390
rect 40340 -11510 40460 -11390
rect 40505 -11510 40625 -11390
rect 40680 -11510 40800 -11390
rect 40845 -11510 40965 -11390
rect 41010 -11510 41130 -11390
rect 41175 -11510 41295 -11390
rect 41350 -11510 41470 -11390
rect 41515 -11510 41635 -11390
rect 41680 -11510 41800 -11390
rect 41845 -11510 41965 -11390
rect 36485 -11675 36605 -11555
rect 36660 -11675 36780 -11555
rect 36825 -11675 36945 -11555
rect 36990 -11675 37110 -11555
rect 37155 -11675 37275 -11555
rect 37330 -11675 37450 -11555
rect 37495 -11675 37615 -11555
rect 37660 -11675 37780 -11555
rect 37825 -11675 37945 -11555
rect 38000 -11675 38120 -11555
rect 38165 -11675 38285 -11555
rect 38330 -11675 38450 -11555
rect 38495 -11675 38615 -11555
rect 38670 -11675 38790 -11555
rect 38835 -11675 38955 -11555
rect 39000 -11675 39120 -11555
rect 39165 -11675 39285 -11555
rect 39340 -11675 39460 -11555
rect 39505 -11675 39625 -11555
rect 39670 -11675 39790 -11555
rect 39835 -11675 39955 -11555
rect 40010 -11675 40130 -11555
rect 40175 -11675 40295 -11555
rect 40340 -11675 40460 -11555
rect 40505 -11675 40625 -11555
rect 40680 -11675 40800 -11555
rect 40845 -11675 40965 -11555
rect 41010 -11675 41130 -11555
rect 41175 -11675 41295 -11555
rect 41350 -11675 41470 -11555
rect 41515 -11675 41635 -11555
rect 41680 -11675 41800 -11555
rect 41845 -11675 41965 -11555
rect 36485 -11840 36605 -11720
rect 36660 -11840 36780 -11720
rect 36825 -11840 36945 -11720
rect 36990 -11840 37110 -11720
rect 37155 -11840 37275 -11720
rect 37330 -11840 37450 -11720
rect 37495 -11840 37615 -11720
rect 37660 -11840 37780 -11720
rect 37825 -11840 37945 -11720
rect 38000 -11840 38120 -11720
rect 38165 -11840 38285 -11720
rect 38330 -11840 38450 -11720
rect 38495 -11840 38615 -11720
rect 38670 -11840 38790 -11720
rect 38835 -11840 38955 -11720
rect 39000 -11840 39120 -11720
rect 39165 -11840 39285 -11720
rect 39340 -11840 39460 -11720
rect 39505 -11840 39625 -11720
rect 39670 -11840 39790 -11720
rect 39835 -11840 39955 -11720
rect 40010 -11840 40130 -11720
rect 40175 -11840 40295 -11720
rect 40340 -11840 40460 -11720
rect 40505 -11840 40625 -11720
rect 40680 -11840 40800 -11720
rect 40845 -11840 40965 -11720
rect 41010 -11840 41130 -11720
rect 41175 -11840 41295 -11720
rect 41350 -11840 41470 -11720
rect 41515 -11840 41635 -11720
rect 41680 -11840 41800 -11720
rect 41845 -11840 41965 -11720
rect 36485 -12005 36605 -11885
rect 36660 -12005 36780 -11885
rect 36825 -12005 36945 -11885
rect 36990 -12005 37110 -11885
rect 37155 -12005 37275 -11885
rect 37330 -12005 37450 -11885
rect 37495 -12005 37615 -11885
rect 37660 -12005 37780 -11885
rect 37825 -12005 37945 -11885
rect 38000 -12005 38120 -11885
rect 38165 -12005 38285 -11885
rect 38330 -12005 38450 -11885
rect 38495 -12005 38615 -11885
rect 38670 -12005 38790 -11885
rect 38835 -12005 38955 -11885
rect 39000 -12005 39120 -11885
rect 39165 -12005 39285 -11885
rect 39340 -12005 39460 -11885
rect 39505 -12005 39625 -11885
rect 39670 -12005 39790 -11885
rect 39835 -12005 39955 -11885
rect 40010 -12005 40130 -11885
rect 40175 -12005 40295 -11885
rect 40340 -12005 40460 -11885
rect 40505 -12005 40625 -11885
rect 40680 -12005 40800 -11885
rect 40845 -12005 40965 -11885
rect 41010 -12005 41130 -11885
rect 41175 -12005 41295 -11885
rect 41350 -12005 41470 -11885
rect 41515 -12005 41635 -11885
rect 41680 -12005 41800 -11885
rect 41845 -12005 41965 -11885
rect 36485 -12180 36605 -12060
rect 36660 -12180 36780 -12060
rect 36825 -12180 36945 -12060
rect 36990 -12180 37110 -12060
rect 37155 -12180 37275 -12060
rect 37330 -12180 37450 -12060
rect 37495 -12180 37615 -12060
rect 37660 -12180 37780 -12060
rect 37825 -12180 37945 -12060
rect 38000 -12180 38120 -12060
rect 38165 -12180 38285 -12060
rect 38330 -12180 38450 -12060
rect 38495 -12180 38615 -12060
rect 38670 -12180 38790 -12060
rect 38835 -12180 38955 -12060
rect 39000 -12180 39120 -12060
rect 39165 -12180 39285 -12060
rect 39340 -12180 39460 -12060
rect 39505 -12180 39625 -12060
rect 39670 -12180 39790 -12060
rect 39835 -12180 39955 -12060
rect 40010 -12180 40130 -12060
rect 40175 -12180 40295 -12060
rect 40340 -12180 40460 -12060
rect 40505 -12180 40625 -12060
rect 40680 -12180 40800 -12060
rect 40845 -12180 40965 -12060
rect 41010 -12180 41130 -12060
rect 41175 -12180 41295 -12060
rect 41350 -12180 41470 -12060
rect 41515 -12180 41635 -12060
rect 41680 -12180 41800 -12060
rect 41845 -12180 41965 -12060
rect 36485 -12345 36605 -12225
rect 36660 -12345 36780 -12225
rect 36825 -12345 36945 -12225
rect 36990 -12345 37110 -12225
rect 37155 -12345 37275 -12225
rect 37330 -12345 37450 -12225
rect 37495 -12345 37615 -12225
rect 37660 -12345 37780 -12225
rect 37825 -12345 37945 -12225
rect 38000 -12345 38120 -12225
rect 38165 -12345 38285 -12225
rect 38330 -12345 38450 -12225
rect 38495 -12345 38615 -12225
rect 38670 -12345 38790 -12225
rect 38835 -12345 38955 -12225
rect 39000 -12345 39120 -12225
rect 39165 -12345 39285 -12225
rect 39340 -12345 39460 -12225
rect 39505 -12345 39625 -12225
rect 39670 -12345 39790 -12225
rect 39835 -12345 39955 -12225
rect 40010 -12345 40130 -12225
rect 40175 -12345 40295 -12225
rect 40340 -12345 40460 -12225
rect 40505 -12345 40625 -12225
rect 40680 -12345 40800 -12225
rect 40845 -12345 40965 -12225
rect 41010 -12345 41130 -12225
rect 41175 -12345 41295 -12225
rect 41350 -12345 41470 -12225
rect 41515 -12345 41635 -12225
rect 41680 -12345 41800 -12225
rect 41845 -12345 41965 -12225
rect 36485 -12510 36605 -12390
rect 36660 -12510 36780 -12390
rect 36825 -12510 36945 -12390
rect 36990 -12510 37110 -12390
rect 37155 -12510 37275 -12390
rect 37330 -12510 37450 -12390
rect 37495 -12510 37615 -12390
rect 37660 -12510 37780 -12390
rect 37825 -12510 37945 -12390
rect 38000 -12510 38120 -12390
rect 38165 -12510 38285 -12390
rect 38330 -12510 38450 -12390
rect 38495 -12510 38615 -12390
rect 38670 -12510 38790 -12390
rect 38835 -12510 38955 -12390
rect 39000 -12510 39120 -12390
rect 39165 -12510 39285 -12390
rect 39340 -12510 39460 -12390
rect 39505 -12510 39625 -12390
rect 39670 -12510 39790 -12390
rect 39835 -12510 39955 -12390
rect 40010 -12510 40130 -12390
rect 40175 -12510 40295 -12390
rect 40340 -12510 40460 -12390
rect 40505 -12510 40625 -12390
rect 40680 -12510 40800 -12390
rect 40845 -12510 40965 -12390
rect 41010 -12510 41130 -12390
rect 41175 -12510 41295 -12390
rect 41350 -12510 41470 -12390
rect 41515 -12510 41635 -12390
rect 41680 -12510 41800 -12390
rect 41845 -12510 41965 -12390
rect 36485 -12675 36605 -12555
rect 36660 -12675 36780 -12555
rect 36825 -12675 36945 -12555
rect 36990 -12675 37110 -12555
rect 37155 -12675 37275 -12555
rect 37330 -12675 37450 -12555
rect 37495 -12675 37615 -12555
rect 37660 -12675 37780 -12555
rect 37825 -12675 37945 -12555
rect 38000 -12675 38120 -12555
rect 38165 -12675 38285 -12555
rect 38330 -12675 38450 -12555
rect 38495 -12675 38615 -12555
rect 38670 -12675 38790 -12555
rect 38835 -12675 38955 -12555
rect 39000 -12675 39120 -12555
rect 39165 -12675 39285 -12555
rect 39340 -12675 39460 -12555
rect 39505 -12675 39625 -12555
rect 39670 -12675 39790 -12555
rect 39835 -12675 39955 -12555
rect 40010 -12675 40130 -12555
rect 40175 -12675 40295 -12555
rect 40340 -12675 40460 -12555
rect 40505 -12675 40625 -12555
rect 40680 -12675 40800 -12555
rect 40845 -12675 40965 -12555
rect 41010 -12675 41130 -12555
rect 41175 -12675 41295 -12555
rect 41350 -12675 41470 -12555
rect 41515 -12675 41635 -12555
rect 41680 -12675 41800 -12555
rect 41845 -12675 41965 -12555
rect 36485 -12850 36605 -12730
rect 36660 -12850 36780 -12730
rect 36825 -12850 36945 -12730
rect 36990 -12850 37110 -12730
rect 37155 -12850 37275 -12730
rect 37330 -12850 37450 -12730
rect 37495 -12850 37615 -12730
rect 37660 -12850 37780 -12730
rect 37825 -12850 37945 -12730
rect 38000 -12850 38120 -12730
rect 38165 -12850 38285 -12730
rect 38330 -12850 38450 -12730
rect 38495 -12850 38615 -12730
rect 38670 -12850 38790 -12730
rect 38835 -12850 38955 -12730
rect 39000 -12850 39120 -12730
rect 39165 -12850 39285 -12730
rect 39340 -12850 39460 -12730
rect 39505 -12850 39625 -12730
rect 39670 -12850 39790 -12730
rect 39835 -12850 39955 -12730
rect 40010 -12850 40130 -12730
rect 40175 -12850 40295 -12730
rect 40340 -12850 40460 -12730
rect 40505 -12850 40625 -12730
rect 40680 -12850 40800 -12730
rect 40845 -12850 40965 -12730
rect 41010 -12850 41130 -12730
rect 41175 -12850 41295 -12730
rect 41350 -12850 41470 -12730
rect 41515 -12850 41635 -12730
rect 41680 -12850 41800 -12730
rect 41845 -12850 41965 -12730
rect 36485 -13015 36605 -12895
rect 36660 -13015 36780 -12895
rect 36825 -13015 36945 -12895
rect 36990 -13015 37110 -12895
rect 37155 -13015 37275 -12895
rect 37330 -13015 37450 -12895
rect 37495 -13015 37615 -12895
rect 37660 -13015 37780 -12895
rect 37825 -13015 37945 -12895
rect 38000 -13015 38120 -12895
rect 38165 -13015 38285 -12895
rect 38330 -13015 38450 -12895
rect 38495 -13015 38615 -12895
rect 38670 -13015 38790 -12895
rect 38835 -13015 38955 -12895
rect 39000 -13015 39120 -12895
rect 39165 -13015 39285 -12895
rect 39340 -13015 39460 -12895
rect 39505 -13015 39625 -12895
rect 39670 -13015 39790 -12895
rect 39835 -13015 39955 -12895
rect 40010 -13015 40130 -12895
rect 40175 -13015 40295 -12895
rect 40340 -13015 40460 -12895
rect 40505 -13015 40625 -12895
rect 40680 -13015 40800 -12895
rect 40845 -13015 40965 -12895
rect 41010 -13015 41130 -12895
rect 41175 -13015 41295 -12895
rect 41350 -13015 41470 -12895
rect 41515 -13015 41635 -12895
rect 41680 -13015 41800 -12895
rect 41845 -13015 41965 -12895
rect 36485 -13180 36605 -13060
rect 36660 -13180 36780 -13060
rect 36825 -13180 36945 -13060
rect 36990 -13180 37110 -13060
rect 37155 -13180 37275 -13060
rect 37330 -13180 37450 -13060
rect 37495 -13180 37615 -13060
rect 37660 -13180 37780 -13060
rect 37825 -13180 37945 -13060
rect 38000 -13180 38120 -13060
rect 38165 -13180 38285 -13060
rect 38330 -13180 38450 -13060
rect 38495 -13180 38615 -13060
rect 38670 -13180 38790 -13060
rect 38835 -13180 38955 -13060
rect 39000 -13180 39120 -13060
rect 39165 -13180 39285 -13060
rect 39340 -13180 39460 -13060
rect 39505 -13180 39625 -13060
rect 39670 -13180 39790 -13060
rect 39835 -13180 39955 -13060
rect 40010 -13180 40130 -13060
rect 40175 -13180 40295 -13060
rect 40340 -13180 40460 -13060
rect 40505 -13180 40625 -13060
rect 40680 -13180 40800 -13060
rect 40845 -13180 40965 -13060
rect 41010 -13180 41130 -13060
rect 41175 -13180 41295 -13060
rect 41350 -13180 41470 -13060
rect 41515 -13180 41635 -13060
rect 41680 -13180 41800 -13060
rect 41845 -13180 41965 -13060
rect 36485 -13345 36605 -13225
rect 36660 -13345 36780 -13225
rect 36825 -13345 36945 -13225
rect 36990 -13345 37110 -13225
rect 37155 -13345 37275 -13225
rect 37330 -13345 37450 -13225
rect 37495 -13345 37615 -13225
rect 37660 -13345 37780 -13225
rect 37825 -13345 37945 -13225
rect 38000 -13345 38120 -13225
rect 38165 -13345 38285 -13225
rect 38330 -13345 38450 -13225
rect 38495 -13345 38615 -13225
rect 38670 -13345 38790 -13225
rect 38835 -13345 38955 -13225
rect 39000 -13345 39120 -13225
rect 39165 -13345 39285 -13225
rect 39340 -13345 39460 -13225
rect 39505 -13345 39625 -13225
rect 39670 -13345 39790 -13225
rect 39835 -13345 39955 -13225
rect 40010 -13345 40130 -13225
rect 40175 -13345 40295 -13225
rect 40340 -13345 40460 -13225
rect 40505 -13345 40625 -13225
rect 40680 -13345 40800 -13225
rect 40845 -13345 40965 -13225
rect 41010 -13345 41130 -13225
rect 41175 -13345 41295 -13225
rect 41350 -13345 41470 -13225
rect 41515 -13345 41635 -13225
rect 41680 -13345 41800 -13225
rect 41845 -13345 41965 -13225
rect 36485 -13520 36605 -13400
rect 36660 -13520 36780 -13400
rect 36825 -13520 36945 -13400
rect 36990 -13520 37110 -13400
rect 37155 -13520 37275 -13400
rect 37330 -13520 37450 -13400
rect 37495 -13520 37615 -13400
rect 37660 -13520 37780 -13400
rect 37825 -13520 37945 -13400
rect 38000 -13520 38120 -13400
rect 38165 -13520 38285 -13400
rect 38330 -13520 38450 -13400
rect 38495 -13520 38615 -13400
rect 38670 -13520 38790 -13400
rect 38835 -13520 38955 -13400
rect 39000 -13520 39120 -13400
rect 39165 -13520 39285 -13400
rect 39340 -13520 39460 -13400
rect 39505 -13520 39625 -13400
rect 39670 -13520 39790 -13400
rect 39835 -13520 39955 -13400
rect 40010 -13520 40130 -13400
rect 40175 -13520 40295 -13400
rect 40340 -13520 40460 -13400
rect 40505 -13520 40625 -13400
rect 40680 -13520 40800 -13400
rect 40845 -13520 40965 -13400
rect 41010 -13520 41130 -13400
rect 41175 -13520 41295 -13400
rect 41350 -13520 41470 -13400
rect 41515 -13520 41635 -13400
rect 41680 -13520 41800 -13400
rect 41845 -13520 41965 -13400
rect 36485 -13685 36605 -13565
rect 36660 -13685 36780 -13565
rect 36825 -13685 36945 -13565
rect 36990 -13685 37110 -13565
rect 37155 -13685 37275 -13565
rect 37330 -13685 37450 -13565
rect 37495 -13685 37615 -13565
rect 37660 -13685 37780 -13565
rect 37825 -13685 37945 -13565
rect 38000 -13685 38120 -13565
rect 38165 -13685 38285 -13565
rect 38330 -13685 38450 -13565
rect 38495 -13685 38615 -13565
rect 38670 -13685 38790 -13565
rect 38835 -13685 38955 -13565
rect 39000 -13685 39120 -13565
rect 39165 -13685 39285 -13565
rect 39340 -13685 39460 -13565
rect 39505 -13685 39625 -13565
rect 39670 -13685 39790 -13565
rect 39835 -13685 39955 -13565
rect 40010 -13685 40130 -13565
rect 40175 -13685 40295 -13565
rect 40340 -13685 40460 -13565
rect 40505 -13685 40625 -13565
rect 40680 -13685 40800 -13565
rect 40845 -13685 40965 -13565
rect 41010 -13685 41130 -13565
rect 41175 -13685 41295 -13565
rect 41350 -13685 41470 -13565
rect 41515 -13685 41635 -13565
rect 41680 -13685 41800 -13565
rect 41845 -13685 41965 -13565
rect 36485 -13850 36605 -13730
rect 36660 -13850 36780 -13730
rect 36825 -13850 36945 -13730
rect 36990 -13850 37110 -13730
rect 37155 -13850 37275 -13730
rect 37330 -13850 37450 -13730
rect 37495 -13850 37615 -13730
rect 37660 -13850 37780 -13730
rect 37825 -13850 37945 -13730
rect 38000 -13850 38120 -13730
rect 38165 -13850 38285 -13730
rect 38330 -13850 38450 -13730
rect 38495 -13850 38615 -13730
rect 38670 -13850 38790 -13730
rect 38835 -13850 38955 -13730
rect 39000 -13850 39120 -13730
rect 39165 -13850 39285 -13730
rect 39340 -13850 39460 -13730
rect 39505 -13850 39625 -13730
rect 39670 -13850 39790 -13730
rect 39835 -13850 39955 -13730
rect 40010 -13850 40130 -13730
rect 40175 -13850 40295 -13730
rect 40340 -13850 40460 -13730
rect 40505 -13850 40625 -13730
rect 40680 -13850 40800 -13730
rect 40845 -13850 40965 -13730
rect 41010 -13850 41130 -13730
rect 41175 -13850 41295 -13730
rect 41350 -13850 41470 -13730
rect 41515 -13850 41635 -13730
rect 41680 -13850 41800 -13730
rect 41845 -13850 41965 -13730
rect 36485 -14015 36605 -13895
rect 36660 -14015 36780 -13895
rect 36825 -14015 36945 -13895
rect 36990 -14015 37110 -13895
rect 37155 -14015 37275 -13895
rect 37330 -14015 37450 -13895
rect 37495 -14015 37615 -13895
rect 37660 -14015 37780 -13895
rect 37825 -14015 37945 -13895
rect 38000 -14015 38120 -13895
rect 38165 -14015 38285 -13895
rect 38330 -14015 38450 -13895
rect 38495 -14015 38615 -13895
rect 38670 -14015 38790 -13895
rect 38835 -14015 38955 -13895
rect 39000 -14015 39120 -13895
rect 39165 -14015 39285 -13895
rect 39340 -14015 39460 -13895
rect 39505 -14015 39625 -13895
rect 39670 -14015 39790 -13895
rect 39835 -14015 39955 -13895
rect 40010 -14015 40130 -13895
rect 40175 -14015 40295 -13895
rect 40340 -14015 40460 -13895
rect 40505 -14015 40625 -13895
rect 40680 -14015 40800 -13895
rect 40845 -14015 40965 -13895
rect 41010 -14015 41130 -13895
rect 41175 -14015 41295 -13895
rect 41350 -14015 41470 -13895
rect 41515 -14015 41635 -13895
rect 41680 -14015 41800 -13895
rect 41845 -14015 41965 -13895
rect 36485 -14190 36605 -14070
rect 36660 -14190 36780 -14070
rect 36825 -14190 36945 -14070
rect 36990 -14190 37110 -14070
rect 37155 -14190 37275 -14070
rect 37330 -14190 37450 -14070
rect 37495 -14190 37615 -14070
rect 37660 -14190 37780 -14070
rect 37825 -14190 37945 -14070
rect 38000 -14190 38120 -14070
rect 38165 -14190 38285 -14070
rect 38330 -14190 38450 -14070
rect 38495 -14190 38615 -14070
rect 38670 -14190 38790 -14070
rect 38835 -14190 38955 -14070
rect 39000 -14190 39120 -14070
rect 39165 -14190 39285 -14070
rect 39340 -14190 39460 -14070
rect 39505 -14190 39625 -14070
rect 39670 -14190 39790 -14070
rect 39835 -14190 39955 -14070
rect 40010 -14190 40130 -14070
rect 40175 -14190 40295 -14070
rect 40340 -14190 40460 -14070
rect 40505 -14190 40625 -14070
rect 40680 -14190 40800 -14070
rect 40845 -14190 40965 -14070
rect 41010 -14190 41130 -14070
rect 41175 -14190 41295 -14070
rect 41350 -14190 41470 -14070
rect 41515 -14190 41635 -14070
rect 41680 -14190 41800 -14070
rect 41845 -14190 41965 -14070
rect 36485 -14355 36605 -14235
rect 36660 -14355 36780 -14235
rect 36825 -14355 36945 -14235
rect 36990 -14355 37110 -14235
rect 37155 -14355 37275 -14235
rect 37330 -14355 37450 -14235
rect 37495 -14355 37615 -14235
rect 37660 -14355 37780 -14235
rect 37825 -14355 37945 -14235
rect 38000 -14355 38120 -14235
rect 38165 -14355 38285 -14235
rect 38330 -14355 38450 -14235
rect 38495 -14355 38615 -14235
rect 38670 -14355 38790 -14235
rect 38835 -14355 38955 -14235
rect 39000 -14355 39120 -14235
rect 39165 -14355 39285 -14235
rect 39340 -14355 39460 -14235
rect 39505 -14355 39625 -14235
rect 39670 -14355 39790 -14235
rect 39835 -14355 39955 -14235
rect 40010 -14355 40130 -14235
rect 40175 -14355 40295 -14235
rect 40340 -14355 40460 -14235
rect 40505 -14355 40625 -14235
rect 40680 -14355 40800 -14235
rect 40845 -14355 40965 -14235
rect 41010 -14355 41130 -14235
rect 41175 -14355 41295 -14235
rect 41350 -14355 41470 -14235
rect 41515 -14355 41635 -14235
rect 41680 -14355 41800 -14235
rect 41845 -14355 41965 -14235
rect 36485 -14520 36605 -14400
rect 36660 -14520 36780 -14400
rect 36825 -14520 36945 -14400
rect 36990 -14520 37110 -14400
rect 37155 -14520 37275 -14400
rect 37330 -14520 37450 -14400
rect 37495 -14520 37615 -14400
rect 37660 -14520 37780 -14400
rect 37825 -14520 37945 -14400
rect 38000 -14520 38120 -14400
rect 38165 -14520 38285 -14400
rect 38330 -14520 38450 -14400
rect 38495 -14520 38615 -14400
rect 38670 -14520 38790 -14400
rect 38835 -14520 38955 -14400
rect 39000 -14520 39120 -14400
rect 39165 -14520 39285 -14400
rect 39340 -14520 39460 -14400
rect 39505 -14520 39625 -14400
rect 39670 -14520 39790 -14400
rect 39835 -14520 39955 -14400
rect 40010 -14520 40130 -14400
rect 40175 -14520 40295 -14400
rect 40340 -14520 40460 -14400
rect 40505 -14520 40625 -14400
rect 40680 -14520 40800 -14400
rect 40845 -14520 40965 -14400
rect 41010 -14520 41130 -14400
rect 41175 -14520 41295 -14400
rect 41350 -14520 41470 -14400
rect 41515 -14520 41635 -14400
rect 41680 -14520 41800 -14400
rect 41845 -14520 41965 -14400
rect 36485 -14685 36605 -14565
rect 36660 -14685 36780 -14565
rect 36825 -14685 36945 -14565
rect 36990 -14685 37110 -14565
rect 37155 -14685 37275 -14565
rect 37330 -14685 37450 -14565
rect 37495 -14685 37615 -14565
rect 37660 -14685 37780 -14565
rect 37825 -14685 37945 -14565
rect 38000 -14685 38120 -14565
rect 38165 -14685 38285 -14565
rect 38330 -14685 38450 -14565
rect 38495 -14685 38615 -14565
rect 38670 -14685 38790 -14565
rect 38835 -14685 38955 -14565
rect 39000 -14685 39120 -14565
rect 39165 -14685 39285 -14565
rect 39340 -14685 39460 -14565
rect 39505 -14685 39625 -14565
rect 39670 -14685 39790 -14565
rect 39835 -14685 39955 -14565
rect 40010 -14685 40130 -14565
rect 40175 -14685 40295 -14565
rect 40340 -14685 40460 -14565
rect 40505 -14685 40625 -14565
rect 40680 -14685 40800 -14565
rect 40845 -14685 40965 -14565
rect 41010 -14685 41130 -14565
rect 41175 -14685 41295 -14565
rect 41350 -14685 41470 -14565
rect 41515 -14685 41635 -14565
rect 41680 -14685 41800 -14565
rect 41845 -14685 41965 -14565
rect 36485 -14860 36605 -14740
rect 36660 -14860 36780 -14740
rect 36825 -14860 36945 -14740
rect 36990 -14860 37110 -14740
rect 37155 -14860 37275 -14740
rect 37330 -14860 37450 -14740
rect 37495 -14860 37615 -14740
rect 37660 -14860 37780 -14740
rect 37825 -14860 37945 -14740
rect 38000 -14860 38120 -14740
rect 38165 -14860 38285 -14740
rect 38330 -14860 38450 -14740
rect 38495 -14860 38615 -14740
rect 38670 -14860 38790 -14740
rect 38835 -14860 38955 -14740
rect 39000 -14860 39120 -14740
rect 39165 -14860 39285 -14740
rect 39340 -14860 39460 -14740
rect 39505 -14860 39625 -14740
rect 39670 -14860 39790 -14740
rect 39835 -14860 39955 -14740
rect 40010 -14860 40130 -14740
rect 40175 -14860 40295 -14740
rect 40340 -14860 40460 -14740
rect 40505 -14860 40625 -14740
rect 40680 -14860 40800 -14740
rect 40845 -14860 40965 -14740
rect 41010 -14860 41130 -14740
rect 41175 -14860 41295 -14740
rect 41350 -14860 41470 -14740
rect 41515 -14860 41635 -14740
rect 41680 -14860 41800 -14740
rect 41845 -14860 41965 -14740
rect 36485 -15025 36605 -14905
rect 36660 -15025 36780 -14905
rect 36825 -15025 36945 -14905
rect 36990 -15025 37110 -14905
rect 37155 -15025 37275 -14905
rect 37330 -15025 37450 -14905
rect 37495 -15025 37615 -14905
rect 37660 -15025 37780 -14905
rect 37825 -15025 37945 -14905
rect 38000 -15025 38120 -14905
rect 38165 -15025 38285 -14905
rect 38330 -15025 38450 -14905
rect 38495 -15025 38615 -14905
rect 38670 -15025 38790 -14905
rect 38835 -15025 38955 -14905
rect 39000 -15025 39120 -14905
rect 39165 -15025 39285 -14905
rect 39340 -15025 39460 -14905
rect 39505 -15025 39625 -14905
rect 39670 -15025 39790 -14905
rect 39835 -15025 39955 -14905
rect 40010 -15025 40130 -14905
rect 40175 -15025 40295 -14905
rect 40340 -15025 40460 -14905
rect 40505 -15025 40625 -14905
rect 40680 -15025 40800 -14905
rect 40845 -15025 40965 -14905
rect 41010 -15025 41130 -14905
rect 41175 -15025 41295 -14905
rect 41350 -15025 41470 -14905
rect 41515 -15025 41635 -14905
rect 41680 -15025 41800 -14905
rect 41845 -15025 41965 -14905
rect 36485 -15190 36605 -15070
rect 36660 -15190 36780 -15070
rect 36825 -15190 36945 -15070
rect 36990 -15190 37110 -15070
rect 37155 -15190 37275 -15070
rect 37330 -15190 37450 -15070
rect 37495 -15190 37615 -15070
rect 37660 -15190 37780 -15070
rect 37825 -15190 37945 -15070
rect 38000 -15190 38120 -15070
rect 38165 -15190 38285 -15070
rect 38330 -15190 38450 -15070
rect 38495 -15190 38615 -15070
rect 38670 -15190 38790 -15070
rect 38835 -15190 38955 -15070
rect 39000 -15190 39120 -15070
rect 39165 -15190 39285 -15070
rect 39340 -15190 39460 -15070
rect 39505 -15190 39625 -15070
rect 39670 -15190 39790 -15070
rect 39835 -15190 39955 -15070
rect 40010 -15190 40130 -15070
rect 40175 -15190 40295 -15070
rect 40340 -15190 40460 -15070
rect 40505 -15190 40625 -15070
rect 40680 -15190 40800 -15070
rect 40845 -15190 40965 -15070
rect 41010 -15190 41130 -15070
rect 41175 -15190 41295 -15070
rect 41350 -15190 41470 -15070
rect 41515 -15190 41635 -15070
rect 41680 -15190 41800 -15070
rect 41845 -15190 41965 -15070
rect 36485 -15355 36605 -15235
rect 36660 -15355 36780 -15235
rect 36825 -15355 36945 -15235
rect 36990 -15355 37110 -15235
rect 37155 -15355 37275 -15235
rect 37330 -15355 37450 -15235
rect 37495 -15355 37615 -15235
rect 37660 -15355 37780 -15235
rect 37825 -15355 37945 -15235
rect 38000 -15355 38120 -15235
rect 38165 -15355 38285 -15235
rect 38330 -15355 38450 -15235
rect 38495 -15355 38615 -15235
rect 38670 -15355 38790 -15235
rect 38835 -15355 38955 -15235
rect 39000 -15355 39120 -15235
rect 39165 -15355 39285 -15235
rect 39340 -15355 39460 -15235
rect 39505 -15355 39625 -15235
rect 39670 -15355 39790 -15235
rect 39835 -15355 39955 -15235
rect 40010 -15355 40130 -15235
rect 40175 -15355 40295 -15235
rect 40340 -15355 40460 -15235
rect 40505 -15355 40625 -15235
rect 40680 -15355 40800 -15235
rect 40845 -15355 40965 -15235
rect 41010 -15355 41130 -15235
rect 41175 -15355 41295 -15235
rect 41350 -15355 41470 -15235
rect 41515 -15355 41635 -15235
rect 41680 -15355 41800 -15235
rect 41845 -15355 41965 -15235
rect 36485 -15530 36605 -15410
rect 36660 -15530 36780 -15410
rect 36825 -15530 36945 -15410
rect 36990 -15530 37110 -15410
rect 37155 -15530 37275 -15410
rect 37330 -15530 37450 -15410
rect 37495 -15530 37615 -15410
rect 37660 -15530 37780 -15410
rect 37825 -15530 37945 -15410
rect 38000 -15530 38120 -15410
rect 38165 -15530 38285 -15410
rect 38330 -15530 38450 -15410
rect 38495 -15530 38615 -15410
rect 38670 -15530 38790 -15410
rect 38835 -15530 38955 -15410
rect 39000 -15530 39120 -15410
rect 39165 -15530 39285 -15410
rect 39340 -15530 39460 -15410
rect 39505 -15530 39625 -15410
rect 39670 -15530 39790 -15410
rect 39835 -15530 39955 -15410
rect 40010 -15530 40130 -15410
rect 40175 -15530 40295 -15410
rect 40340 -15530 40460 -15410
rect 40505 -15530 40625 -15410
rect 40680 -15530 40800 -15410
rect 40845 -15530 40965 -15410
rect 41010 -15530 41130 -15410
rect 41175 -15530 41295 -15410
rect 41350 -15530 41470 -15410
rect 41515 -15530 41635 -15410
rect 41680 -15530 41800 -15410
rect 41845 -15530 41965 -15410
rect 42175 -10170 42295 -10050
rect 42350 -10170 42470 -10050
rect 42515 -10170 42635 -10050
rect 42680 -10170 42800 -10050
rect 42845 -10170 42965 -10050
rect 43020 -10170 43140 -10050
rect 43185 -10170 43305 -10050
rect 43350 -10170 43470 -10050
rect 43515 -10170 43635 -10050
rect 43690 -10170 43810 -10050
rect 43855 -10170 43975 -10050
rect 44020 -10170 44140 -10050
rect 44185 -10170 44305 -10050
rect 44360 -10170 44480 -10050
rect 44525 -10170 44645 -10050
rect 44690 -10170 44810 -10050
rect 44855 -10170 44975 -10050
rect 45030 -10170 45150 -10050
rect 45195 -10170 45315 -10050
rect 45360 -10170 45480 -10050
rect 45525 -10170 45645 -10050
rect 45700 -10170 45820 -10050
rect 45865 -10170 45985 -10050
rect 46030 -10170 46150 -10050
rect 46195 -10170 46315 -10050
rect 46370 -10170 46490 -10050
rect 46535 -10170 46655 -10050
rect 46700 -10170 46820 -10050
rect 46865 -10170 46985 -10050
rect 47040 -10170 47160 -10050
rect 47205 -10170 47325 -10050
rect 47370 -10170 47490 -10050
rect 47535 -10170 47655 -10050
rect 42175 -10335 42295 -10215
rect 42350 -10335 42470 -10215
rect 42515 -10335 42635 -10215
rect 42680 -10335 42800 -10215
rect 42845 -10335 42965 -10215
rect 43020 -10335 43140 -10215
rect 43185 -10335 43305 -10215
rect 43350 -10335 43470 -10215
rect 43515 -10335 43635 -10215
rect 43690 -10335 43810 -10215
rect 43855 -10335 43975 -10215
rect 44020 -10335 44140 -10215
rect 44185 -10335 44305 -10215
rect 44360 -10335 44480 -10215
rect 44525 -10335 44645 -10215
rect 44690 -10335 44810 -10215
rect 44855 -10335 44975 -10215
rect 45030 -10335 45150 -10215
rect 45195 -10335 45315 -10215
rect 45360 -10335 45480 -10215
rect 45525 -10335 45645 -10215
rect 45700 -10335 45820 -10215
rect 45865 -10335 45985 -10215
rect 46030 -10335 46150 -10215
rect 46195 -10335 46315 -10215
rect 46370 -10335 46490 -10215
rect 46535 -10335 46655 -10215
rect 46700 -10335 46820 -10215
rect 46865 -10335 46985 -10215
rect 47040 -10335 47160 -10215
rect 47205 -10335 47325 -10215
rect 47370 -10335 47490 -10215
rect 47535 -10335 47655 -10215
rect 42175 -10500 42295 -10380
rect 42350 -10500 42470 -10380
rect 42515 -10500 42635 -10380
rect 42680 -10500 42800 -10380
rect 42845 -10500 42965 -10380
rect 43020 -10500 43140 -10380
rect 43185 -10500 43305 -10380
rect 43350 -10500 43470 -10380
rect 43515 -10500 43635 -10380
rect 43690 -10500 43810 -10380
rect 43855 -10500 43975 -10380
rect 44020 -10500 44140 -10380
rect 44185 -10500 44305 -10380
rect 44360 -10500 44480 -10380
rect 44525 -10500 44645 -10380
rect 44690 -10500 44810 -10380
rect 44855 -10500 44975 -10380
rect 45030 -10500 45150 -10380
rect 45195 -10500 45315 -10380
rect 45360 -10500 45480 -10380
rect 45525 -10500 45645 -10380
rect 45700 -10500 45820 -10380
rect 45865 -10500 45985 -10380
rect 46030 -10500 46150 -10380
rect 46195 -10500 46315 -10380
rect 46370 -10500 46490 -10380
rect 46535 -10500 46655 -10380
rect 46700 -10500 46820 -10380
rect 46865 -10500 46985 -10380
rect 47040 -10500 47160 -10380
rect 47205 -10500 47325 -10380
rect 47370 -10500 47490 -10380
rect 47535 -10500 47655 -10380
rect 42175 -10665 42295 -10545
rect 42350 -10665 42470 -10545
rect 42515 -10665 42635 -10545
rect 42680 -10665 42800 -10545
rect 42845 -10665 42965 -10545
rect 43020 -10665 43140 -10545
rect 43185 -10665 43305 -10545
rect 43350 -10665 43470 -10545
rect 43515 -10665 43635 -10545
rect 43690 -10665 43810 -10545
rect 43855 -10665 43975 -10545
rect 44020 -10665 44140 -10545
rect 44185 -10665 44305 -10545
rect 44360 -10665 44480 -10545
rect 44525 -10665 44645 -10545
rect 44690 -10665 44810 -10545
rect 44855 -10665 44975 -10545
rect 45030 -10665 45150 -10545
rect 45195 -10665 45315 -10545
rect 45360 -10665 45480 -10545
rect 45525 -10665 45645 -10545
rect 45700 -10665 45820 -10545
rect 45865 -10665 45985 -10545
rect 46030 -10665 46150 -10545
rect 46195 -10665 46315 -10545
rect 46370 -10665 46490 -10545
rect 46535 -10665 46655 -10545
rect 46700 -10665 46820 -10545
rect 46865 -10665 46985 -10545
rect 47040 -10665 47160 -10545
rect 47205 -10665 47325 -10545
rect 47370 -10665 47490 -10545
rect 47535 -10665 47655 -10545
rect 42175 -10840 42295 -10720
rect 42350 -10840 42470 -10720
rect 42515 -10840 42635 -10720
rect 42680 -10840 42800 -10720
rect 42845 -10840 42965 -10720
rect 43020 -10840 43140 -10720
rect 43185 -10840 43305 -10720
rect 43350 -10840 43470 -10720
rect 43515 -10840 43635 -10720
rect 43690 -10840 43810 -10720
rect 43855 -10840 43975 -10720
rect 44020 -10840 44140 -10720
rect 44185 -10840 44305 -10720
rect 44360 -10840 44480 -10720
rect 44525 -10840 44645 -10720
rect 44690 -10840 44810 -10720
rect 44855 -10840 44975 -10720
rect 45030 -10840 45150 -10720
rect 45195 -10840 45315 -10720
rect 45360 -10840 45480 -10720
rect 45525 -10840 45645 -10720
rect 45700 -10840 45820 -10720
rect 45865 -10840 45985 -10720
rect 46030 -10840 46150 -10720
rect 46195 -10840 46315 -10720
rect 46370 -10840 46490 -10720
rect 46535 -10840 46655 -10720
rect 46700 -10840 46820 -10720
rect 46865 -10840 46985 -10720
rect 47040 -10840 47160 -10720
rect 47205 -10840 47325 -10720
rect 47370 -10840 47490 -10720
rect 47535 -10840 47655 -10720
rect 42175 -11005 42295 -10885
rect 42350 -11005 42470 -10885
rect 42515 -11005 42635 -10885
rect 42680 -11005 42800 -10885
rect 42845 -11005 42965 -10885
rect 43020 -11005 43140 -10885
rect 43185 -11005 43305 -10885
rect 43350 -11005 43470 -10885
rect 43515 -11005 43635 -10885
rect 43690 -11005 43810 -10885
rect 43855 -11005 43975 -10885
rect 44020 -11005 44140 -10885
rect 44185 -11005 44305 -10885
rect 44360 -11005 44480 -10885
rect 44525 -11005 44645 -10885
rect 44690 -11005 44810 -10885
rect 44855 -11005 44975 -10885
rect 45030 -11005 45150 -10885
rect 45195 -11005 45315 -10885
rect 45360 -11005 45480 -10885
rect 45525 -11005 45645 -10885
rect 45700 -11005 45820 -10885
rect 45865 -11005 45985 -10885
rect 46030 -11005 46150 -10885
rect 46195 -11005 46315 -10885
rect 46370 -11005 46490 -10885
rect 46535 -11005 46655 -10885
rect 46700 -11005 46820 -10885
rect 46865 -11005 46985 -10885
rect 47040 -11005 47160 -10885
rect 47205 -11005 47325 -10885
rect 47370 -11005 47490 -10885
rect 47535 -11005 47655 -10885
rect 42175 -11170 42295 -11050
rect 42350 -11170 42470 -11050
rect 42515 -11170 42635 -11050
rect 42680 -11170 42800 -11050
rect 42845 -11170 42965 -11050
rect 43020 -11170 43140 -11050
rect 43185 -11170 43305 -11050
rect 43350 -11170 43470 -11050
rect 43515 -11170 43635 -11050
rect 43690 -11170 43810 -11050
rect 43855 -11170 43975 -11050
rect 44020 -11170 44140 -11050
rect 44185 -11170 44305 -11050
rect 44360 -11170 44480 -11050
rect 44525 -11170 44645 -11050
rect 44690 -11170 44810 -11050
rect 44855 -11170 44975 -11050
rect 45030 -11170 45150 -11050
rect 45195 -11170 45315 -11050
rect 45360 -11170 45480 -11050
rect 45525 -11170 45645 -11050
rect 45700 -11170 45820 -11050
rect 45865 -11170 45985 -11050
rect 46030 -11170 46150 -11050
rect 46195 -11170 46315 -11050
rect 46370 -11170 46490 -11050
rect 46535 -11170 46655 -11050
rect 46700 -11170 46820 -11050
rect 46865 -11170 46985 -11050
rect 47040 -11170 47160 -11050
rect 47205 -11170 47325 -11050
rect 47370 -11170 47490 -11050
rect 47535 -11170 47655 -11050
rect 42175 -11335 42295 -11215
rect 42350 -11335 42470 -11215
rect 42515 -11335 42635 -11215
rect 42680 -11335 42800 -11215
rect 42845 -11335 42965 -11215
rect 43020 -11335 43140 -11215
rect 43185 -11335 43305 -11215
rect 43350 -11335 43470 -11215
rect 43515 -11335 43635 -11215
rect 43690 -11335 43810 -11215
rect 43855 -11335 43975 -11215
rect 44020 -11335 44140 -11215
rect 44185 -11335 44305 -11215
rect 44360 -11335 44480 -11215
rect 44525 -11335 44645 -11215
rect 44690 -11335 44810 -11215
rect 44855 -11335 44975 -11215
rect 45030 -11335 45150 -11215
rect 45195 -11335 45315 -11215
rect 45360 -11335 45480 -11215
rect 45525 -11335 45645 -11215
rect 45700 -11335 45820 -11215
rect 45865 -11335 45985 -11215
rect 46030 -11335 46150 -11215
rect 46195 -11335 46315 -11215
rect 46370 -11335 46490 -11215
rect 46535 -11335 46655 -11215
rect 46700 -11335 46820 -11215
rect 46865 -11335 46985 -11215
rect 47040 -11335 47160 -11215
rect 47205 -11335 47325 -11215
rect 47370 -11335 47490 -11215
rect 47535 -11335 47655 -11215
rect 42175 -11510 42295 -11390
rect 42350 -11510 42470 -11390
rect 42515 -11510 42635 -11390
rect 42680 -11510 42800 -11390
rect 42845 -11510 42965 -11390
rect 43020 -11510 43140 -11390
rect 43185 -11510 43305 -11390
rect 43350 -11510 43470 -11390
rect 43515 -11510 43635 -11390
rect 43690 -11510 43810 -11390
rect 43855 -11510 43975 -11390
rect 44020 -11510 44140 -11390
rect 44185 -11510 44305 -11390
rect 44360 -11510 44480 -11390
rect 44525 -11510 44645 -11390
rect 44690 -11510 44810 -11390
rect 44855 -11510 44975 -11390
rect 45030 -11510 45150 -11390
rect 45195 -11510 45315 -11390
rect 45360 -11510 45480 -11390
rect 45525 -11510 45645 -11390
rect 45700 -11510 45820 -11390
rect 45865 -11510 45985 -11390
rect 46030 -11510 46150 -11390
rect 46195 -11510 46315 -11390
rect 46370 -11510 46490 -11390
rect 46535 -11510 46655 -11390
rect 46700 -11510 46820 -11390
rect 46865 -11510 46985 -11390
rect 47040 -11510 47160 -11390
rect 47205 -11510 47325 -11390
rect 47370 -11510 47490 -11390
rect 47535 -11510 47655 -11390
rect 42175 -11675 42295 -11555
rect 42350 -11675 42470 -11555
rect 42515 -11675 42635 -11555
rect 42680 -11675 42800 -11555
rect 42845 -11675 42965 -11555
rect 43020 -11675 43140 -11555
rect 43185 -11675 43305 -11555
rect 43350 -11675 43470 -11555
rect 43515 -11675 43635 -11555
rect 43690 -11675 43810 -11555
rect 43855 -11675 43975 -11555
rect 44020 -11675 44140 -11555
rect 44185 -11675 44305 -11555
rect 44360 -11675 44480 -11555
rect 44525 -11675 44645 -11555
rect 44690 -11675 44810 -11555
rect 44855 -11675 44975 -11555
rect 45030 -11675 45150 -11555
rect 45195 -11675 45315 -11555
rect 45360 -11675 45480 -11555
rect 45525 -11675 45645 -11555
rect 45700 -11675 45820 -11555
rect 45865 -11675 45985 -11555
rect 46030 -11675 46150 -11555
rect 46195 -11675 46315 -11555
rect 46370 -11675 46490 -11555
rect 46535 -11675 46655 -11555
rect 46700 -11675 46820 -11555
rect 46865 -11675 46985 -11555
rect 47040 -11675 47160 -11555
rect 47205 -11675 47325 -11555
rect 47370 -11675 47490 -11555
rect 47535 -11675 47655 -11555
rect 42175 -11840 42295 -11720
rect 42350 -11840 42470 -11720
rect 42515 -11840 42635 -11720
rect 42680 -11840 42800 -11720
rect 42845 -11840 42965 -11720
rect 43020 -11840 43140 -11720
rect 43185 -11840 43305 -11720
rect 43350 -11840 43470 -11720
rect 43515 -11840 43635 -11720
rect 43690 -11840 43810 -11720
rect 43855 -11840 43975 -11720
rect 44020 -11840 44140 -11720
rect 44185 -11840 44305 -11720
rect 44360 -11840 44480 -11720
rect 44525 -11840 44645 -11720
rect 44690 -11840 44810 -11720
rect 44855 -11840 44975 -11720
rect 45030 -11840 45150 -11720
rect 45195 -11840 45315 -11720
rect 45360 -11840 45480 -11720
rect 45525 -11840 45645 -11720
rect 45700 -11840 45820 -11720
rect 45865 -11840 45985 -11720
rect 46030 -11840 46150 -11720
rect 46195 -11840 46315 -11720
rect 46370 -11840 46490 -11720
rect 46535 -11840 46655 -11720
rect 46700 -11840 46820 -11720
rect 46865 -11840 46985 -11720
rect 47040 -11840 47160 -11720
rect 47205 -11840 47325 -11720
rect 47370 -11840 47490 -11720
rect 47535 -11840 47655 -11720
rect 42175 -12005 42295 -11885
rect 42350 -12005 42470 -11885
rect 42515 -12005 42635 -11885
rect 42680 -12005 42800 -11885
rect 42845 -12005 42965 -11885
rect 43020 -12005 43140 -11885
rect 43185 -12005 43305 -11885
rect 43350 -12005 43470 -11885
rect 43515 -12005 43635 -11885
rect 43690 -12005 43810 -11885
rect 43855 -12005 43975 -11885
rect 44020 -12005 44140 -11885
rect 44185 -12005 44305 -11885
rect 44360 -12005 44480 -11885
rect 44525 -12005 44645 -11885
rect 44690 -12005 44810 -11885
rect 44855 -12005 44975 -11885
rect 45030 -12005 45150 -11885
rect 45195 -12005 45315 -11885
rect 45360 -12005 45480 -11885
rect 45525 -12005 45645 -11885
rect 45700 -12005 45820 -11885
rect 45865 -12005 45985 -11885
rect 46030 -12005 46150 -11885
rect 46195 -12005 46315 -11885
rect 46370 -12005 46490 -11885
rect 46535 -12005 46655 -11885
rect 46700 -12005 46820 -11885
rect 46865 -12005 46985 -11885
rect 47040 -12005 47160 -11885
rect 47205 -12005 47325 -11885
rect 47370 -12005 47490 -11885
rect 47535 -12005 47655 -11885
rect 42175 -12180 42295 -12060
rect 42350 -12180 42470 -12060
rect 42515 -12180 42635 -12060
rect 42680 -12180 42800 -12060
rect 42845 -12180 42965 -12060
rect 43020 -12180 43140 -12060
rect 43185 -12180 43305 -12060
rect 43350 -12180 43470 -12060
rect 43515 -12180 43635 -12060
rect 43690 -12180 43810 -12060
rect 43855 -12180 43975 -12060
rect 44020 -12180 44140 -12060
rect 44185 -12180 44305 -12060
rect 44360 -12180 44480 -12060
rect 44525 -12180 44645 -12060
rect 44690 -12180 44810 -12060
rect 44855 -12180 44975 -12060
rect 45030 -12180 45150 -12060
rect 45195 -12180 45315 -12060
rect 45360 -12180 45480 -12060
rect 45525 -12180 45645 -12060
rect 45700 -12180 45820 -12060
rect 45865 -12180 45985 -12060
rect 46030 -12180 46150 -12060
rect 46195 -12180 46315 -12060
rect 46370 -12180 46490 -12060
rect 46535 -12180 46655 -12060
rect 46700 -12180 46820 -12060
rect 46865 -12180 46985 -12060
rect 47040 -12180 47160 -12060
rect 47205 -12180 47325 -12060
rect 47370 -12180 47490 -12060
rect 47535 -12180 47655 -12060
rect 42175 -12345 42295 -12225
rect 42350 -12345 42470 -12225
rect 42515 -12345 42635 -12225
rect 42680 -12345 42800 -12225
rect 42845 -12345 42965 -12225
rect 43020 -12345 43140 -12225
rect 43185 -12345 43305 -12225
rect 43350 -12345 43470 -12225
rect 43515 -12345 43635 -12225
rect 43690 -12345 43810 -12225
rect 43855 -12345 43975 -12225
rect 44020 -12345 44140 -12225
rect 44185 -12345 44305 -12225
rect 44360 -12345 44480 -12225
rect 44525 -12345 44645 -12225
rect 44690 -12345 44810 -12225
rect 44855 -12345 44975 -12225
rect 45030 -12345 45150 -12225
rect 45195 -12345 45315 -12225
rect 45360 -12345 45480 -12225
rect 45525 -12345 45645 -12225
rect 45700 -12345 45820 -12225
rect 45865 -12345 45985 -12225
rect 46030 -12345 46150 -12225
rect 46195 -12345 46315 -12225
rect 46370 -12345 46490 -12225
rect 46535 -12345 46655 -12225
rect 46700 -12345 46820 -12225
rect 46865 -12345 46985 -12225
rect 47040 -12345 47160 -12225
rect 47205 -12345 47325 -12225
rect 47370 -12345 47490 -12225
rect 47535 -12345 47655 -12225
rect 42175 -12510 42295 -12390
rect 42350 -12510 42470 -12390
rect 42515 -12510 42635 -12390
rect 42680 -12510 42800 -12390
rect 42845 -12510 42965 -12390
rect 43020 -12510 43140 -12390
rect 43185 -12510 43305 -12390
rect 43350 -12510 43470 -12390
rect 43515 -12510 43635 -12390
rect 43690 -12510 43810 -12390
rect 43855 -12510 43975 -12390
rect 44020 -12510 44140 -12390
rect 44185 -12510 44305 -12390
rect 44360 -12510 44480 -12390
rect 44525 -12510 44645 -12390
rect 44690 -12510 44810 -12390
rect 44855 -12510 44975 -12390
rect 45030 -12510 45150 -12390
rect 45195 -12510 45315 -12390
rect 45360 -12510 45480 -12390
rect 45525 -12510 45645 -12390
rect 45700 -12510 45820 -12390
rect 45865 -12510 45985 -12390
rect 46030 -12510 46150 -12390
rect 46195 -12510 46315 -12390
rect 46370 -12510 46490 -12390
rect 46535 -12510 46655 -12390
rect 46700 -12510 46820 -12390
rect 46865 -12510 46985 -12390
rect 47040 -12510 47160 -12390
rect 47205 -12510 47325 -12390
rect 47370 -12510 47490 -12390
rect 47535 -12510 47655 -12390
rect 42175 -12675 42295 -12555
rect 42350 -12675 42470 -12555
rect 42515 -12675 42635 -12555
rect 42680 -12675 42800 -12555
rect 42845 -12675 42965 -12555
rect 43020 -12675 43140 -12555
rect 43185 -12675 43305 -12555
rect 43350 -12675 43470 -12555
rect 43515 -12675 43635 -12555
rect 43690 -12675 43810 -12555
rect 43855 -12675 43975 -12555
rect 44020 -12675 44140 -12555
rect 44185 -12675 44305 -12555
rect 44360 -12675 44480 -12555
rect 44525 -12675 44645 -12555
rect 44690 -12675 44810 -12555
rect 44855 -12675 44975 -12555
rect 45030 -12675 45150 -12555
rect 45195 -12675 45315 -12555
rect 45360 -12675 45480 -12555
rect 45525 -12675 45645 -12555
rect 45700 -12675 45820 -12555
rect 45865 -12675 45985 -12555
rect 46030 -12675 46150 -12555
rect 46195 -12675 46315 -12555
rect 46370 -12675 46490 -12555
rect 46535 -12675 46655 -12555
rect 46700 -12675 46820 -12555
rect 46865 -12675 46985 -12555
rect 47040 -12675 47160 -12555
rect 47205 -12675 47325 -12555
rect 47370 -12675 47490 -12555
rect 47535 -12675 47655 -12555
rect 42175 -12850 42295 -12730
rect 42350 -12850 42470 -12730
rect 42515 -12850 42635 -12730
rect 42680 -12850 42800 -12730
rect 42845 -12850 42965 -12730
rect 43020 -12850 43140 -12730
rect 43185 -12850 43305 -12730
rect 43350 -12850 43470 -12730
rect 43515 -12850 43635 -12730
rect 43690 -12850 43810 -12730
rect 43855 -12850 43975 -12730
rect 44020 -12850 44140 -12730
rect 44185 -12850 44305 -12730
rect 44360 -12850 44480 -12730
rect 44525 -12850 44645 -12730
rect 44690 -12850 44810 -12730
rect 44855 -12850 44975 -12730
rect 45030 -12850 45150 -12730
rect 45195 -12850 45315 -12730
rect 45360 -12850 45480 -12730
rect 45525 -12850 45645 -12730
rect 45700 -12850 45820 -12730
rect 45865 -12850 45985 -12730
rect 46030 -12850 46150 -12730
rect 46195 -12850 46315 -12730
rect 46370 -12850 46490 -12730
rect 46535 -12850 46655 -12730
rect 46700 -12850 46820 -12730
rect 46865 -12850 46985 -12730
rect 47040 -12850 47160 -12730
rect 47205 -12850 47325 -12730
rect 47370 -12850 47490 -12730
rect 47535 -12850 47655 -12730
rect 42175 -13015 42295 -12895
rect 42350 -13015 42470 -12895
rect 42515 -13015 42635 -12895
rect 42680 -13015 42800 -12895
rect 42845 -13015 42965 -12895
rect 43020 -13015 43140 -12895
rect 43185 -13015 43305 -12895
rect 43350 -13015 43470 -12895
rect 43515 -13015 43635 -12895
rect 43690 -13015 43810 -12895
rect 43855 -13015 43975 -12895
rect 44020 -13015 44140 -12895
rect 44185 -13015 44305 -12895
rect 44360 -13015 44480 -12895
rect 44525 -13015 44645 -12895
rect 44690 -13015 44810 -12895
rect 44855 -13015 44975 -12895
rect 45030 -13015 45150 -12895
rect 45195 -13015 45315 -12895
rect 45360 -13015 45480 -12895
rect 45525 -13015 45645 -12895
rect 45700 -13015 45820 -12895
rect 45865 -13015 45985 -12895
rect 46030 -13015 46150 -12895
rect 46195 -13015 46315 -12895
rect 46370 -13015 46490 -12895
rect 46535 -13015 46655 -12895
rect 46700 -13015 46820 -12895
rect 46865 -13015 46985 -12895
rect 47040 -13015 47160 -12895
rect 47205 -13015 47325 -12895
rect 47370 -13015 47490 -12895
rect 47535 -13015 47655 -12895
rect 42175 -13180 42295 -13060
rect 42350 -13180 42470 -13060
rect 42515 -13180 42635 -13060
rect 42680 -13180 42800 -13060
rect 42845 -13180 42965 -13060
rect 43020 -13180 43140 -13060
rect 43185 -13180 43305 -13060
rect 43350 -13180 43470 -13060
rect 43515 -13180 43635 -13060
rect 43690 -13180 43810 -13060
rect 43855 -13180 43975 -13060
rect 44020 -13180 44140 -13060
rect 44185 -13180 44305 -13060
rect 44360 -13180 44480 -13060
rect 44525 -13180 44645 -13060
rect 44690 -13180 44810 -13060
rect 44855 -13180 44975 -13060
rect 45030 -13180 45150 -13060
rect 45195 -13180 45315 -13060
rect 45360 -13180 45480 -13060
rect 45525 -13180 45645 -13060
rect 45700 -13180 45820 -13060
rect 45865 -13180 45985 -13060
rect 46030 -13180 46150 -13060
rect 46195 -13180 46315 -13060
rect 46370 -13180 46490 -13060
rect 46535 -13180 46655 -13060
rect 46700 -13180 46820 -13060
rect 46865 -13180 46985 -13060
rect 47040 -13180 47160 -13060
rect 47205 -13180 47325 -13060
rect 47370 -13180 47490 -13060
rect 47535 -13180 47655 -13060
rect 42175 -13345 42295 -13225
rect 42350 -13345 42470 -13225
rect 42515 -13345 42635 -13225
rect 42680 -13345 42800 -13225
rect 42845 -13345 42965 -13225
rect 43020 -13345 43140 -13225
rect 43185 -13345 43305 -13225
rect 43350 -13345 43470 -13225
rect 43515 -13345 43635 -13225
rect 43690 -13345 43810 -13225
rect 43855 -13345 43975 -13225
rect 44020 -13345 44140 -13225
rect 44185 -13345 44305 -13225
rect 44360 -13345 44480 -13225
rect 44525 -13345 44645 -13225
rect 44690 -13345 44810 -13225
rect 44855 -13345 44975 -13225
rect 45030 -13345 45150 -13225
rect 45195 -13345 45315 -13225
rect 45360 -13345 45480 -13225
rect 45525 -13345 45645 -13225
rect 45700 -13345 45820 -13225
rect 45865 -13345 45985 -13225
rect 46030 -13345 46150 -13225
rect 46195 -13345 46315 -13225
rect 46370 -13345 46490 -13225
rect 46535 -13345 46655 -13225
rect 46700 -13345 46820 -13225
rect 46865 -13345 46985 -13225
rect 47040 -13345 47160 -13225
rect 47205 -13345 47325 -13225
rect 47370 -13345 47490 -13225
rect 47535 -13345 47655 -13225
rect 42175 -13520 42295 -13400
rect 42350 -13520 42470 -13400
rect 42515 -13520 42635 -13400
rect 42680 -13520 42800 -13400
rect 42845 -13520 42965 -13400
rect 43020 -13520 43140 -13400
rect 43185 -13520 43305 -13400
rect 43350 -13520 43470 -13400
rect 43515 -13520 43635 -13400
rect 43690 -13520 43810 -13400
rect 43855 -13520 43975 -13400
rect 44020 -13520 44140 -13400
rect 44185 -13520 44305 -13400
rect 44360 -13520 44480 -13400
rect 44525 -13520 44645 -13400
rect 44690 -13520 44810 -13400
rect 44855 -13520 44975 -13400
rect 45030 -13520 45150 -13400
rect 45195 -13520 45315 -13400
rect 45360 -13520 45480 -13400
rect 45525 -13520 45645 -13400
rect 45700 -13520 45820 -13400
rect 45865 -13520 45985 -13400
rect 46030 -13520 46150 -13400
rect 46195 -13520 46315 -13400
rect 46370 -13520 46490 -13400
rect 46535 -13520 46655 -13400
rect 46700 -13520 46820 -13400
rect 46865 -13520 46985 -13400
rect 47040 -13520 47160 -13400
rect 47205 -13520 47325 -13400
rect 47370 -13520 47490 -13400
rect 47535 -13520 47655 -13400
rect 42175 -13685 42295 -13565
rect 42350 -13685 42470 -13565
rect 42515 -13685 42635 -13565
rect 42680 -13685 42800 -13565
rect 42845 -13685 42965 -13565
rect 43020 -13685 43140 -13565
rect 43185 -13685 43305 -13565
rect 43350 -13685 43470 -13565
rect 43515 -13685 43635 -13565
rect 43690 -13685 43810 -13565
rect 43855 -13685 43975 -13565
rect 44020 -13685 44140 -13565
rect 44185 -13685 44305 -13565
rect 44360 -13685 44480 -13565
rect 44525 -13685 44645 -13565
rect 44690 -13685 44810 -13565
rect 44855 -13685 44975 -13565
rect 45030 -13685 45150 -13565
rect 45195 -13685 45315 -13565
rect 45360 -13685 45480 -13565
rect 45525 -13685 45645 -13565
rect 45700 -13685 45820 -13565
rect 45865 -13685 45985 -13565
rect 46030 -13685 46150 -13565
rect 46195 -13685 46315 -13565
rect 46370 -13685 46490 -13565
rect 46535 -13685 46655 -13565
rect 46700 -13685 46820 -13565
rect 46865 -13685 46985 -13565
rect 47040 -13685 47160 -13565
rect 47205 -13685 47325 -13565
rect 47370 -13685 47490 -13565
rect 47535 -13685 47655 -13565
rect 42175 -13850 42295 -13730
rect 42350 -13850 42470 -13730
rect 42515 -13850 42635 -13730
rect 42680 -13850 42800 -13730
rect 42845 -13850 42965 -13730
rect 43020 -13850 43140 -13730
rect 43185 -13850 43305 -13730
rect 43350 -13850 43470 -13730
rect 43515 -13850 43635 -13730
rect 43690 -13850 43810 -13730
rect 43855 -13850 43975 -13730
rect 44020 -13850 44140 -13730
rect 44185 -13850 44305 -13730
rect 44360 -13850 44480 -13730
rect 44525 -13850 44645 -13730
rect 44690 -13850 44810 -13730
rect 44855 -13850 44975 -13730
rect 45030 -13850 45150 -13730
rect 45195 -13850 45315 -13730
rect 45360 -13850 45480 -13730
rect 45525 -13850 45645 -13730
rect 45700 -13850 45820 -13730
rect 45865 -13850 45985 -13730
rect 46030 -13850 46150 -13730
rect 46195 -13850 46315 -13730
rect 46370 -13850 46490 -13730
rect 46535 -13850 46655 -13730
rect 46700 -13850 46820 -13730
rect 46865 -13850 46985 -13730
rect 47040 -13850 47160 -13730
rect 47205 -13850 47325 -13730
rect 47370 -13850 47490 -13730
rect 47535 -13850 47655 -13730
rect 42175 -14015 42295 -13895
rect 42350 -14015 42470 -13895
rect 42515 -14015 42635 -13895
rect 42680 -14015 42800 -13895
rect 42845 -14015 42965 -13895
rect 43020 -14015 43140 -13895
rect 43185 -14015 43305 -13895
rect 43350 -14015 43470 -13895
rect 43515 -14015 43635 -13895
rect 43690 -14015 43810 -13895
rect 43855 -14015 43975 -13895
rect 44020 -14015 44140 -13895
rect 44185 -14015 44305 -13895
rect 44360 -14015 44480 -13895
rect 44525 -14015 44645 -13895
rect 44690 -14015 44810 -13895
rect 44855 -14015 44975 -13895
rect 45030 -14015 45150 -13895
rect 45195 -14015 45315 -13895
rect 45360 -14015 45480 -13895
rect 45525 -14015 45645 -13895
rect 45700 -14015 45820 -13895
rect 45865 -14015 45985 -13895
rect 46030 -14015 46150 -13895
rect 46195 -14015 46315 -13895
rect 46370 -14015 46490 -13895
rect 46535 -14015 46655 -13895
rect 46700 -14015 46820 -13895
rect 46865 -14015 46985 -13895
rect 47040 -14015 47160 -13895
rect 47205 -14015 47325 -13895
rect 47370 -14015 47490 -13895
rect 47535 -14015 47655 -13895
rect 42175 -14190 42295 -14070
rect 42350 -14190 42470 -14070
rect 42515 -14190 42635 -14070
rect 42680 -14190 42800 -14070
rect 42845 -14190 42965 -14070
rect 43020 -14190 43140 -14070
rect 43185 -14190 43305 -14070
rect 43350 -14190 43470 -14070
rect 43515 -14190 43635 -14070
rect 43690 -14190 43810 -14070
rect 43855 -14190 43975 -14070
rect 44020 -14190 44140 -14070
rect 44185 -14190 44305 -14070
rect 44360 -14190 44480 -14070
rect 44525 -14190 44645 -14070
rect 44690 -14190 44810 -14070
rect 44855 -14190 44975 -14070
rect 45030 -14190 45150 -14070
rect 45195 -14190 45315 -14070
rect 45360 -14190 45480 -14070
rect 45525 -14190 45645 -14070
rect 45700 -14190 45820 -14070
rect 45865 -14190 45985 -14070
rect 46030 -14190 46150 -14070
rect 46195 -14190 46315 -14070
rect 46370 -14190 46490 -14070
rect 46535 -14190 46655 -14070
rect 46700 -14190 46820 -14070
rect 46865 -14190 46985 -14070
rect 47040 -14190 47160 -14070
rect 47205 -14190 47325 -14070
rect 47370 -14190 47490 -14070
rect 47535 -14190 47655 -14070
rect 42175 -14355 42295 -14235
rect 42350 -14355 42470 -14235
rect 42515 -14355 42635 -14235
rect 42680 -14355 42800 -14235
rect 42845 -14355 42965 -14235
rect 43020 -14355 43140 -14235
rect 43185 -14355 43305 -14235
rect 43350 -14355 43470 -14235
rect 43515 -14355 43635 -14235
rect 43690 -14355 43810 -14235
rect 43855 -14355 43975 -14235
rect 44020 -14355 44140 -14235
rect 44185 -14355 44305 -14235
rect 44360 -14355 44480 -14235
rect 44525 -14355 44645 -14235
rect 44690 -14355 44810 -14235
rect 44855 -14355 44975 -14235
rect 45030 -14355 45150 -14235
rect 45195 -14355 45315 -14235
rect 45360 -14355 45480 -14235
rect 45525 -14355 45645 -14235
rect 45700 -14355 45820 -14235
rect 45865 -14355 45985 -14235
rect 46030 -14355 46150 -14235
rect 46195 -14355 46315 -14235
rect 46370 -14355 46490 -14235
rect 46535 -14355 46655 -14235
rect 46700 -14355 46820 -14235
rect 46865 -14355 46985 -14235
rect 47040 -14355 47160 -14235
rect 47205 -14355 47325 -14235
rect 47370 -14355 47490 -14235
rect 47535 -14355 47655 -14235
rect 42175 -14520 42295 -14400
rect 42350 -14520 42470 -14400
rect 42515 -14520 42635 -14400
rect 42680 -14520 42800 -14400
rect 42845 -14520 42965 -14400
rect 43020 -14520 43140 -14400
rect 43185 -14520 43305 -14400
rect 43350 -14520 43470 -14400
rect 43515 -14520 43635 -14400
rect 43690 -14520 43810 -14400
rect 43855 -14520 43975 -14400
rect 44020 -14520 44140 -14400
rect 44185 -14520 44305 -14400
rect 44360 -14520 44480 -14400
rect 44525 -14520 44645 -14400
rect 44690 -14520 44810 -14400
rect 44855 -14520 44975 -14400
rect 45030 -14520 45150 -14400
rect 45195 -14520 45315 -14400
rect 45360 -14520 45480 -14400
rect 45525 -14520 45645 -14400
rect 45700 -14520 45820 -14400
rect 45865 -14520 45985 -14400
rect 46030 -14520 46150 -14400
rect 46195 -14520 46315 -14400
rect 46370 -14520 46490 -14400
rect 46535 -14520 46655 -14400
rect 46700 -14520 46820 -14400
rect 46865 -14520 46985 -14400
rect 47040 -14520 47160 -14400
rect 47205 -14520 47325 -14400
rect 47370 -14520 47490 -14400
rect 47535 -14520 47655 -14400
rect 42175 -14685 42295 -14565
rect 42350 -14685 42470 -14565
rect 42515 -14685 42635 -14565
rect 42680 -14685 42800 -14565
rect 42845 -14685 42965 -14565
rect 43020 -14685 43140 -14565
rect 43185 -14685 43305 -14565
rect 43350 -14685 43470 -14565
rect 43515 -14685 43635 -14565
rect 43690 -14685 43810 -14565
rect 43855 -14685 43975 -14565
rect 44020 -14685 44140 -14565
rect 44185 -14685 44305 -14565
rect 44360 -14685 44480 -14565
rect 44525 -14685 44645 -14565
rect 44690 -14685 44810 -14565
rect 44855 -14685 44975 -14565
rect 45030 -14685 45150 -14565
rect 45195 -14685 45315 -14565
rect 45360 -14685 45480 -14565
rect 45525 -14685 45645 -14565
rect 45700 -14685 45820 -14565
rect 45865 -14685 45985 -14565
rect 46030 -14685 46150 -14565
rect 46195 -14685 46315 -14565
rect 46370 -14685 46490 -14565
rect 46535 -14685 46655 -14565
rect 46700 -14685 46820 -14565
rect 46865 -14685 46985 -14565
rect 47040 -14685 47160 -14565
rect 47205 -14685 47325 -14565
rect 47370 -14685 47490 -14565
rect 47535 -14685 47655 -14565
rect 42175 -14860 42295 -14740
rect 42350 -14860 42470 -14740
rect 42515 -14860 42635 -14740
rect 42680 -14860 42800 -14740
rect 42845 -14860 42965 -14740
rect 43020 -14860 43140 -14740
rect 43185 -14860 43305 -14740
rect 43350 -14860 43470 -14740
rect 43515 -14860 43635 -14740
rect 43690 -14860 43810 -14740
rect 43855 -14860 43975 -14740
rect 44020 -14860 44140 -14740
rect 44185 -14860 44305 -14740
rect 44360 -14860 44480 -14740
rect 44525 -14860 44645 -14740
rect 44690 -14860 44810 -14740
rect 44855 -14860 44975 -14740
rect 45030 -14860 45150 -14740
rect 45195 -14860 45315 -14740
rect 45360 -14860 45480 -14740
rect 45525 -14860 45645 -14740
rect 45700 -14860 45820 -14740
rect 45865 -14860 45985 -14740
rect 46030 -14860 46150 -14740
rect 46195 -14860 46315 -14740
rect 46370 -14860 46490 -14740
rect 46535 -14860 46655 -14740
rect 46700 -14860 46820 -14740
rect 46865 -14860 46985 -14740
rect 47040 -14860 47160 -14740
rect 47205 -14860 47325 -14740
rect 47370 -14860 47490 -14740
rect 47535 -14860 47655 -14740
rect 42175 -15025 42295 -14905
rect 42350 -15025 42470 -14905
rect 42515 -15025 42635 -14905
rect 42680 -15025 42800 -14905
rect 42845 -15025 42965 -14905
rect 43020 -15025 43140 -14905
rect 43185 -15025 43305 -14905
rect 43350 -15025 43470 -14905
rect 43515 -15025 43635 -14905
rect 43690 -15025 43810 -14905
rect 43855 -15025 43975 -14905
rect 44020 -15025 44140 -14905
rect 44185 -15025 44305 -14905
rect 44360 -15025 44480 -14905
rect 44525 -15025 44645 -14905
rect 44690 -15025 44810 -14905
rect 44855 -15025 44975 -14905
rect 45030 -15025 45150 -14905
rect 45195 -15025 45315 -14905
rect 45360 -15025 45480 -14905
rect 45525 -15025 45645 -14905
rect 45700 -15025 45820 -14905
rect 45865 -15025 45985 -14905
rect 46030 -15025 46150 -14905
rect 46195 -15025 46315 -14905
rect 46370 -15025 46490 -14905
rect 46535 -15025 46655 -14905
rect 46700 -15025 46820 -14905
rect 46865 -15025 46985 -14905
rect 47040 -15025 47160 -14905
rect 47205 -15025 47325 -14905
rect 47370 -15025 47490 -14905
rect 47535 -15025 47655 -14905
rect 42175 -15190 42295 -15070
rect 42350 -15190 42470 -15070
rect 42515 -15190 42635 -15070
rect 42680 -15190 42800 -15070
rect 42845 -15190 42965 -15070
rect 43020 -15190 43140 -15070
rect 43185 -15190 43305 -15070
rect 43350 -15190 43470 -15070
rect 43515 -15190 43635 -15070
rect 43690 -15190 43810 -15070
rect 43855 -15190 43975 -15070
rect 44020 -15190 44140 -15070
rect 44185 -15190 44305 -15070
rect 44360 -15190 44480 -15070
rect 44525 -15190 44645 -15070
rect 44690 -15190 44810 -15070
rect 44855 -15190 44975 -15070
rect 45030 -15190 45150 -15070
rect 45195 -15190 45315 -15070
rect 45360 -15190 45480 -15070
rect 45525 -15190 45645 -15070
rect 45700 -15190 45820 -15070
rect 45865 -15190 45985 -15070
rect 46030 -15190 46150 -15070
rect 46195 -15190 46315 -15070
rect 46370 -15190 46490 -15070
rect 46535 -15190 46655 -15070
rect 46700 -15190 46820 -15070
rect 46865 -15190 46985 -15070
rect 47040 -15190 47160 -15070
rect 47205 -15190 47325 -15070
rect 47370 -15190 47490 -15070
rect 47535 -15190 47655 -15070
rect 42175 -15355 42295 -15235
rect 42350 -15355 42470 -15235
rect 42515 -15355 42635 -15235
rect 42680 -15355 42800 -15235
rect 42845 -15355 42965 -15235
rect 43020 -15355 43140 -15235
rect 43185 -15355 43305 -15235
rect 43350 -15355 43470 -15235
rect 43515 -15355 43635 -15235
rect 43690 -15355 43810 -15235
rect 43855 -15355 43975 -15235
rect 44020 -15355 44140 -15235
rect 44185 -15355 44305 -15235
rect 44360 -15355 44480 -15235
rect 44525 -15355 44645 -15235
rect 44690 -15355 44810 -15235
rect 44855 -15355 44975 -15235
rect 45030 -15355 45150 -15235
rect 45195 -15355 45315 -15235
rect 45360 -15355 45480 -15235
rect 45525 -15355 45645 -15235
rect 45700 -15355 45820 -15235
rect 45865 -15355 45985 -15235
rect 46030 -15355 46150 -15235
rect 46195 -15355 46315 -15235
rect 46370 -15355 46490 -15235
rect 46535 -15355 46655 -15235
rect 46700 -15355 46820 -15235
rect 46865 -15355 46985 -15235
rect 47040 -15355 47160 -15235
rect 47205 -15355 47325 -15235
rect 47370 -15355 47490 -15235
rect 47535 -15355 47655 -15235
rect 42175 -15530 42295 -15410
rect 42350 -15530 42470 -15410
rect 42515 -15530 42635 -15410
rect 42680 -15530 42800 -15410
rect 42845 -15530 42965 -15410
rect 43020 -15530 43140 -15410
rect 43185 -15530 43305 -15410
rect 43350 -15530 43470 -15410
rect 43515 -15530 43635 -15410
rect 43690 -15530 43810 -15410
rect 43855 -15530 43975 -15410
rect 44020 -15530 44140 -15410
rect 44185 -15530 44305 -15410
rect 44360 -15530 44480 -15410
rect 44525 -15530 44645 -15410
rect 44690 -15530 44810 -15410
rect 44855 -15530 44975 -15410
rect 45030 -15530 45150 -15410
rect 45195 -15530 45315 -15410
rect 45360 -15530 45480 -15410
rect 45525 -15530 45645 -15410
rect 45700 -15530 45820 -15410
rect 45865 -15530 45985 -15410
rect 46030 -15530 46150 -15410
rect 46195 -15530 46315 -15410
rect 46370 -15530 46490 -15410
rect 46535 -15530 46655 -15410
rect 46700 -15530 46820 -15410
rect 46865 -15530 46985 -15410
rect 47040 -15530 47160 -15410
rect 47205 -15530 47325 -15410
rect 47370 -15530 47490 -15410
rect 47535 -15530 47655 -15410
rect 47865 -10170 47985 -10050
rect 48040 -10170 48160 -10050
rect 48205 -10170 48325 -10050
rect 48370 -10170 48490 -10050
rect 48535 -10170 48655 -10050
rect 48710 -10170 48830 -10050
rect 48875 -10170 48995 -10050
rect 49040 -10170 49160 -10050
rect 49205 -10170 49325 -10050
rect 49380 -10170 49500 -10050
rect 49545 -10170 49665 -10050
rect 49710 -10170 49830 -10050
rect 49875 -10170 49995 -10050
rect 50050 -10170 50170 -10050
rect 50215 -10170 50335 -10050
rect 50380 -10170 50500 -10050
rect 50545 -10170 50665 -10050
rect 50720 -10170 50840 -10050
rect 50885 -10170 51005 -10050
rect 51050 -10170 51170 -10050
rect 51215 -10170 51335 -10050
rect 51390 -10170 51510 -10050
rect 51555 -10170 51675 -10050
rect 51720 -10170 51840 -10050
rect 51885 -10170 52005 -10050
rect 52060 -10170 52180 -10050
rect 52225 -10170 52345 -10050
rect 52390 -10170 52510 -10050
rect 52555 -10170 52675 -10050
rect 52730 -10170 52850 -10050
rect 52895 -10170 53015 -10050
rect 53060 -10170 53180 -10050
rect 53225 -10170 53345 -10050
rect 47865 -10335 47985 -10215
rect 48040 -10335 48160 -10215
rect 48205 -10335 48325 -10215
rect 48370 -10335 48490 -10215
rect 48535 -10335 48655 -10215
rect 48710 -10335 48830 -10215
rect 48875 -10335 48995 -10215
rect 49040 -10335 49160 -10215
rect 49205 -10335 49325 -10215
rect 49380 -10335 49500 -10215
rect 49545 -10335 49665 -10215
rect 49710 -10335 49830 -10215
rect 49875 -10335 49995 -10215
rect 50050 -10335 50170 -10215
rect 50215 -10335 50335 -10215
rect 50380 -10335 50500 -10215
rect 50545 -10335 50665 -10215
rect 50720 -10335 50840 -10215
rect 50885 -10335 51005 -10215
rect 51050 -10335 51170 -10215
rect 51215 -10335 51335 -10215
rect 51390 -10335 51510 -10215
rect 51555 -10335 51675 -10215
rect 51720 -10335 51840 -10215
rect 51885 -10335 52005 -10215
rect 52060 -10335 52180 -10215
rect 52225 -10335 52345 -10215
rect 52390 -10335 52510 -10215
rect 52555 -10335 52675 -10215
rect 52730 -10335 52850 -10215
rect 52895 -10335 53015 -10215
rect 53060 -10335 53180 -10215
rect 53225 -10335 53345 -10215
rect 47865 -10500 47985 -10380
rect 48040 -10500 48160 -10380
rect 48205 -10500 48325 -10380
rect 48370 -10500 48490 -10380
rect 48535 -10500 48655 -10380
rect 48710 -10500 48830 -10380
rect 48875 -10500 48995 -10380
rect 49040 -10500 49160 -10380
rect 49205 -10500 49325 -10380
rect 49380 -10500 49500 -10380
rect 49545 -10500 49665 -10380
rect 49710 -10500 49830 -10380
rect 49875 -10500 49995 -10380
rect 50050 -10500 50170 -10380
rect 50215 -10500 50335 -10380
rect 50380 -10500 50500 -10380
rect 50545 -10500 50665 -10380
rect 50720 -10500 50840 -10380
rect 50885 -10500 51005 -10380
rect 51050 -10500 51170 -10380
rect 51215 -10500 51335 -10380
rect 51390 -10500 51510 -10380
rect 51555 -10500 51675 -10380
rect 51720 -10500 51840 -10380
rect 51885 -10500 52005 -10380
rect 52060 -10500 52180 -10380
rect 52225 -10500 52345 -10380
rect 52390 -10500 52510 -10380
rect 52555 -10500 52675 -10380
rect 52730 -10500 52850 -10380
rect 52895 -10500 53015 -10380
rect 53060 -10500 53180 -10380
rect 53225 -10500 53345 -10380
rect 47865 -10665 47985 -10545
rect 48040 -10665 48160 -10545
rect 48205 -10665 48325 -10545
rect 48370 -10665 48490 -10545
rect 48535 -10665 48655 -10545
rect 48710 -10665 48830 -10545
rect 48875 -10665 48995 -10545
rect 49040 -10665 49160 -10545
rect 49205 -10665 49325 -10545
rect 49380 -10665 49500 -10545
rect 49545 -10665 49665 -10545
rect 49710 -10665 49830 -10545
rect 49875 -10665 49995 -10545
rect 50050 -10665 50170 -10545
rect 50215 -10665 50335 -10545
rect 50380 -10665 50500 -10545
rect 50545 -10665 50665 -10545
rect 50720 -10665 50840 -10545
rect 50885 -10665 51005 -10545
rect 51050 -10665 51170 -10545
rect 51215 -10665 51335 -10545
rect 51390 -10665 51510 -10545
rect 51555 -10665 51675 -10545
rect 51720 -10665 51840 -10545
rect 51885 -10665 52005 -10545
rect 52060 -10665 52180 -10545
rect 52225 -10665 52345 -10545
rect 52390 -10665 52510 -10545
rect 52555 -10665 52675 -10545
rect 52730 -10665 52850 -10545
rect 52895 -10665 53015 -10545
rect 53060 -10665 53180 -10545
rect 53225 -10665 53345 -10545
rect 47865 -10840 47985 -10720
rect 48040 -10840 48160 -10720
rect 48205 -10840 48325 -10720
rect 48370 -10840 48490 -10720
rect 48535 -10840 48655 -10720
rect 48710 -10840 48830 -10720
rect 48875 -10840 48995 -10720
rect 49040 -10840 49160 -10720
rect 49205 -10840 49325 -10720
rect 49380 -10840 49500 -10720
rect 49545 -10840 49665 -10720
rect 49710 -10840 49830 -10720
rect 49875 -10840 49995 -10720
rect 50050 -10840 50170 -10720
rect 50215 -10840 50335 -10720
rect 50380 -10840 50500 -10720
rect 50545 -10840 50665 -10720
rect 50720 -10840 50840 -10720
rect 50885 -10840 51005 -10720
rect 51050 -10840 51170 -10720
rect 51215 -10840 51335 -10720
rect 51390 -10840 51510 -10720
rect 51555 -10840 51675 -10720
rect 51720 -10840 51840 -10720
rect 51885 -10840 52005 -10720
rect 52060 -10840 52180 -10720
rect 52225 -10840 52345 -10720
rect 52390 -10840 52510 -10720
rect 52555 -10840 52675 -10720
rect 52730 -10840 52850 -10720
rect 52895 -10840 53015 -10720
rect 53060 -10840 53180 -10720
rect 53225 -10840 53345 -10720
rect 47865 -11005 47985 -10885
rect 48040 -11005 48160 -10885
rect 48205 -11005 48325 -10885
rect 48370 -11005 48490 -10885
rect 48535 -11005 48655 -10885
rect 48710 -11005 48830 -10885
rect 48875 -11005 48995 -10885
rect 49040 -11005 49160 -10885
rect 49205 -11005 49325 -10885
rect 49380 -11005 49500 -10885
rect 49545 -11005 49665 -10885
rect 49710 -11005 49830 -10885
rect 49875 -11005 49995 -10885
rect 50050 -11005 50170 -10885
rect 50215 -11005 50335 -10885
rect 50380 -11005 50500 -10885
rect 50545 -11005 50665 -10885
rect 50720 -11005 50840 -10885
rect 50885 -11005 51005 -10885
rect 51050 -11005 51170 -10885
rect 51215 -11005 51335 -10885
rect 51390 -11005 51510 -10885
rect 51555 -11005 51675 -10885
rect 51720 -11005 51840 -10885
rect 51885 -11005 52005 -10885
rect 52060 -11005 52180 -10885
rect 52225 -11005 52345 -10885
rect 52390 -11005 52510 -10885
rect 52555 -11005 52675 -10885
rect 52730 -11005 52850 -10885
rect 52895 -11005 53015 -10885
rect 53060 -11005 53180 -10885
rect 53225 -11005 53345 -10885
rect 47865 -11170 47985 -11050
rect 48040 -11170 48160 -11050
rect 48205 -11170 48325 -11050
rect 48370 -11170 48490 -11050
rect 48535 -11170 48655 -11050
rect 48710 -11170 48830 -11050
rect 48875 -11170 48995 -11050
rect 49040 -11170 49160 -11050
rect 49205 -11170 49325 -11050
rect 49380 -11170 49500 -11050
rect 49545 -11170 49665 -11050
rect 49710 -11170 49830 -11050
rect 49875 -11170 49995 -11050
rect 50050 -11170 50170 -11050
rect 50215 -11170 50335 -11050
rect 50380 -11170 50500 -11050
rect 50545 -11170 50665 -11050
rect 50720 -11170 50840 -11050
rect 50885 -11170 51005 -11050
rect 51050 -11170 51170 -11050
rect 51215 -11170 51335 -11050
rect 51390 -11170 51510 -11050
rect 51555 -11170 51675 -11050
rect 51720 -11170 51840 -11050
rect 51885 -11170 52005 -11050
rect 52060 -11170 52180 -11050
rect 52225 -11170 52345 -11050
rect 52390 -11170 52510 -11050
rect 52555 -11170 52675 -11050
rect 52730 -11170 52850 -11050
rect 52895 -11170 53015 -11050
rect 53060 -11170 53180 -11050
rect 53225 -11170 53345 -11050
rect 47865 -11335 47985 -11215
rect 48040 -11335 48160 -11215
rect 48205 -11335 48325 -11215
rect 48370 -11335 48490 -11215
rect 48535 -11335 48655 -11215
rect 48710 -11335 48830 -11215
rect 48875 -11335 48995 -11215
rect 49040 -11335 49160 -11215
rect 49205 -11335 49325 -11215
rect 49380 -11335 49500 -11215
rect 49545 -11335 49665 -11215
rect 49710 -11335 49830 -11215
rect 49875 -11335 49995 -11215
rect 50050 -11335 50170 -11215
rect 50215 -11335 50335 -11215
rect 50380 -11335 50500 -11215
rect 50545 -11335 50665 -11215
rect 50720 -11335 50840 -11215
rect 50885 -11335 51005 -11215
rect 51050 -11335 51170 -11215
rect 51215 -11335 51335 -11215
rect 51390 -11335 51510 -11215
rect 51555 -11335 51675 -11215
rect 51720 -11335 51840 -11215
rect 51885 -11335 52005 -11215
rect 52060 -11335 52180 -11215
rect 52225 -11335 52345 -11215
rect 52390 -11335 52510 -11215
rect 52555 -11335 52675 -11215
rect 52730 -11335 52850 -11215
rect 52895 -11335 53015 -11215
rect 53060 -11335 53180 -11215
rect 53225 -11335 53345 -11215
rect 47865 -11510 47985 -11390
rect 48040 -11510 48160 -11390
rect 48205 -11510 48325 -11390
rect 48370 -11510 48490 -11390
rect 48535 -11510 48655 -11390
rect 48710 -11510 48830 -11390
rect 48875 -11510 48995 -11390
rect 49040 -11510 49160 -11390
rect 49205 -11510 49325 -11390
rect 49380 -11510 49500 -11390
rect 49545 -11510 49665 -11390
rect 49710 -11510 49830 -11390
rect 49875 -11510 49995 -11390
rect 50050 -11510 50170 -11390
rect 50215 -11510 50335 -11390
rect 50380 -11510 50500 -11390
rect 50545 -11510 50665 -11390
rect 50720 -11510 50840 -11390
rect 50885 -11510 51005 -11390
rect 51050 -11510 51170 -11390
rect 51215 -11510 51335 -11390
rect 51390 -11510 51510 -11390
rect 51555 -11510 51675 -11390
rect 51720 -11510 51840 -11390
rect 51885 -11510 52005 -11390
rect 52060 -11510 52180 -11390
rect 52225 -11510 52345 -11390
rect 52390 -11510 52510 -11390
rect 52555 -11510 52675 -11390
rect 52730 -11510 52850 -11390
rect 52895 -11510 53015 -11390
rect 53060 -11510 53180 -11390
rect 53225 -11510 53345 -11390
rect 47865 -11675 47985 -11555
rect 48040 -11675 48160 -11555
rect 48205 -11675 48325 -11555
rect 48370 -11675 48490 -11555
rect 48535 -11675 48655 -11555
rect 48710 -11675 48830 -11555
rect 48875 -11675 48995 -11555
rect 49040 -11675 49160 -11555
rect 49205 -11675 49325 -11555
rect 49380 -11675 49500 -11555
rect 49545 -11675 49665 -11555
rect 49710 -11675 49830 -11555
rect 49875 -11675 49995 -11555
rect 50050 -11675 50170 -11555
rect 50215 -11675 50335 -11555
rect 50380 -11675 50500 -11555
rect 50545 -11675 50665 -11555
rect 50720 -11675 50840 -11555
rect 50885 -11675 51005 -11555
rect 51050 -11675 51170 -11555
rect 51215 -11675 51335 -11555
rect 51390 -11675 51510 -11555
rect 51555 -11675 51675 -11555
rect 51720 -11675 51840 -11555
rect 51885 -11675 52005 -11555
rect 52060 -11675 52180 -11555
rect 52225 -11675 52345 -11555
rect 52390 -11675 52510 -11555
rect 52555 -11675 52675 -11555
rect 52730 -11675 52850 -11555
rect 52895 -11675 53015 -11555
rect 53060 -11675 53180 -11555
rect 53225 -11675 53345 -11555
rect 47865 -11840 47985 -11720
rect 48040 -11840 48160 -11720
rect 48205 -11840 48325 -11720
rect 48370 -11840 48490 -11720
rect 48535 -11840 48655 -11720
rect 48710 -11840 48830 -11720
rect 48875 -11840 48995 -11720
rect 49040 -11840 49160 -11720
rect 49205 -11840 49325 -11720
rect 49380 -11840 49500 -11720
rect 49545 -11840 49665 -11720
rect 49710 -11840 49830 -11720
rect 49875 -11840 49995 -11720
rect 50050 -11840 50170 -11720
rect 50215 -11840 50335 -11720
rect 50380 -11840 50500 -11720
rect 50545 -11840 50665 -11720
rect 50720 -11840 50840 -11720
rect 50885 -11840 51005 -11720
rect 51050 -11840 51170 -11720
rect 51215 -11840 51335 -11720
rect 51390 -11840 51510 -11720
rect 51555 -11840 51675 -11720
rect 51720 -11840 51840 -11720
rect 51885 -11840 52005 -11720
rect 52060 -11840 52180 -11720
rect 52225 -11840 52345 -11720
rect 52390 -11840 52510 -11720
rect 52555 -11840 52675 -11720
rect 52730 -11840 52850 -11720
rect 52895 -11840 53015 -11720
rect 53060 -11840 53180 -11720
rect 53225 -11840 53345 -11720
rect 47865 -12005 47985 -11885
rect 48040 -12005 48160 -11885
rect 48205 -12005 48325 -11885
rect 48370 -12005 48490 -11885
rect 48535 -12005 48655 -11885
rect 48710 -12005 48830 -11885
rect 48875 -12005 48995 -11885
rect 49040 -12005 49160 -11885
rect 49205 -12005 49325 -11885
rect 49380 -12005 49500 -11885
rect 49545 -12005 49665 -11885
rect 49710 -12005 49830 -11885
rect 49875 -12005 49995 -11885
rect 50050 -12005 50170 -11885
rect 50215 -12005 50335 -11885
rect 50380 -12005 50500 -11885
rect 50545 -12005 50665 -11885
rect 50720 -12005 50840 -11885
rect 50885 -12005 51005 -11885
rect 51050 -12005 51170 -11885
rect 51215 -12005 51335 -11885
rect 51390 -12005 51510 -11885
rect 51555 -12005 51675 -11885
rect 51720 -12005 51840 -11885
rect 51885 -12005 52005 -11885
rect 52060 -12005 52180 -11885
rect 52225 -12005 52345 -11885
rect 52390 -12005 52510 -11885
rect 52555 -12005 52675 -11885
rect 52730 -12005 52850 -11885
rect 52895 -12005 53015 -11885
rect 53060 -12005 53180 -11885
rect 53225 -12005 53345 -11885
rect 47865 -12180 47985 -12060
rect 48040 -12180 48160 -12060
rect 48205 -12180 48325 -12060
rect 48370 -12180 48490 -12060
rect 48535 -12180 48655 -12060
rect 48710 -12180 48830 -12060
rect 48875 -12180 48995 -12060
rect 49040 -12180 49160 -12060
rect 49205 -12180 49325 -12060
rect 49380 -12180 49500 -12060
rect 49545 -12180 49665 -12060
rect 49710 -12180 49830 -12060
rect 49875 -12180 49995 -12060
rect 50050 -12180 50170 -12060
rect 50215 -12180 50335 -12060
rect 50380 -12180 50500 -12060
rect 50545 -12180 50665 -12060
rect 50720 -12180 50840 -12060
rect 50885 -12180 51005 -12060
rect 51050 -12180 51170 -12060
rect 51215 -12180 51335 -12060
rect 51390 -12180 51510 -12060
rect 51555 -12180 51675 -12060
rect 51720 -12180 51840 -12060
rect 51885 -12180 52005 -12060
rect 52060 -12180 52180 -12060
rect 52225 -12180 52345 -12060
rect 52390 -12180 52510 -12060
rect 52555 -12180 52675 -12060
rect 52730 -12180 52850 -12060
rect 52895 -12180 53015 -12060
rect 53060 -12180 53180 -12060
rect 53225 -12180 53345 -12060
rect 47865 -12345 47985 -12225
rect 48040 -12345 48160 -12225
rect 48205 -12345 48325 -12225
rect 48370 -12345 48490 -12225
rect 48535 -12345 48655 -12225
rect 48710 -12345 48830 -12225
rect 48875 -12345 48995 -12225
rect 49040 -12345 49160 -12225
rect 49205 -12345 49325 -12225
rect 49380 -12345 49500 -12225
rect 49545 -12345 49665 -12225
rect 49710 -12345 49830 -12225
rect 49875 -12345 49995 -12225
rect 50050 -12345 50170 -12225
rect 50215 -12345 50335 -12225
rect 50380 -12345 50500 -12225
rect 50545 -12345 50665 -12225
rect 50720 -12345 50840 -12225
rect 50885 -12345 51005 -12225
rect 51050 -12345 51170 -12225
rect 51215 -12345 51335 -12225
rect 51390 -12345 51510 -12225
rect 51555 -12345 51675 -12225
rect 51720 -12345 51840 -12225
rect 51885 -12345 52005 -12225
rect 52060 -12345 52180 -12225
rect 52225 -12345 52345 -12225
rect 52390 -12345 52510 -12225
rect 52555 -12345 52675 -12225
rect 52730 -12345 52850 -12225
rect 52895 -12345 53015 -12225
rect 53060 -12345 53180 -12225
rect 53225 -12345 53345 -12225
rect 47865 -12510 47985 -12390
rect 48040 -12510 48160 -12390
rect 48205 -12510 48325 -12390
rect 48370 -12510 48490 -12390
rect 48535 -12510 48655 -12390
rect 48710 -12510 48830 -12390
rect 48875 -12510 48995 -12390
rect 49040 -12510 49160 -12390
rect 49205 -12510 49325 -12390
rect 49380 -12510 49500 -12390
rect 49545 -12510 49665 -12390
rect 49710 -12510 49830 -12390
rect 49875 -12510 49995 -12390
rect 50050 -12510 50170 -12390
rect 50215 -12510 50335 -12390
rect 50380 -12510 50500 -12390
rect 50545 -12510 50665 -12390
rect 50720 -12510 50840 -12390
rect 50885 -12510 51005 -12390
rect 51050 -12510 51170 -12390
rect 51215 -12510 51335 -12390
rect 51390 -12510 51510 -12390
rect 51555 -12510 51675 -12390
rect 51720 -12510 51840 -12390
rect 51885 -12510 52005 -12390
rect 52060 -12510 52180 -12390
rect 52225 -12510 52345 -12390
rect 52390 -12510 52510 -12390
rect 52555 -12510 52675 -12390
rect 52730 -12510 52850 -12390
rect 52895 -12510 53015 -12390
rect 53060 -12510 53180 -12390
rect 53225 -12510 53345 -12390
rect 47865 -12675 47985 -12555
rect 48040 -12675 48160 -12555
rect 48205 -12675 48325 -12555
rect 48370 -12675 48490 -12555
rect 48535 -12675 48655 -12555
rect 48710 -12675 48830 -12555
rect 48875 -12675 48995 -12555
rect 49040 -12675 49160 -12555
rect 49205 -12675 49325 -12555
rect 49380 -12675 49500 -12555
rect 49545 -12675 49665 -12555
rect 49710 -12675 49830 -12555
rect 49875 -12675 49995 -12555
rect 50050 -12675 50170 -12555
rect 50215 -12675 50335 -12555
rect 50380 -12675 50500 -12555
rect 50545 -12675 50665 -12555
rect 50720 -12675 50840 -12555
rect 50885 -12675 51005 -12555
rect 51050 -12675 51170 -12555
rect 51215 -12675 51335 -12555
rect 51390 -12675 51510 -12555
rect 51555 -12675 51675 -12555
rect 51720 -12675 51840 -12555
rect 51885 -12675 52005 -12555
rect 52060 -12675 52180 -12555
rect 52225 -12675 52345 -12555
rect 52390 -12675 52510 -12555
rect 52555 -12675 52675 -12555
rect 52730 -12675 52850 -12555
rect 52895 -12675 53015 -12555
rect 53060 -12675 53180 -12555
rect 53225 -12675 53345 -12555
rect 47865 -12850 47985 -12730
rect 48040 -12850 48160 -12730
rect 48205 -12850 48325 -12730
rect 48370 -12850 48490 -12730
rect 48535 -12850 48655 -12730
rect 48710 -12850 48830 -12730
rect 48875 -12850 48995 -12730
rect 49040 -12850 49160 -12730
rect 49205 -12850 49325 -12730
rect 49380 -12850 49500 -12730
rect 49545 -12850 49665 -12730
rect 49710 -12850 49830 -12730
rect 49875 -12850 49995 -12730
rect 50050 -12850 50170 -12730
rect 50215 -12850 50335 -12730
rect 50380 -12850 50500 -12730
rect 50545 -12850 50665 -12730
rect 50720 -12850 50840 -12730
rect 50885 -12850 51005 -12730
rect 51050 -12850 51170 -12730
rect 51215 -12850 51335 -12730
rect 51390 -12850 51510 -12730
rect 51555 -12850 51675 -12730
rect 51720 -12850 51840 -12730
rect 51885 -12850 52005 -12730
rect 52060 -12850 52180 -12730
rect 52225 -12850 52345 -12730
rect 52390 -12850 52510 -12730
rect 52555 -12850 52675 -12730
rect 52730 -12850 52850 -12730
rect 52895 -12850 53015 -12730
rect 53060 -12850 53180 -12730
rect 53225 -12850 53345 -12730
rect 47865 -13015 47985 -12895
rect 48040 -13015 48160 -12895
rect 48205 -13015 48325 -12895
rect 48370 -13015 48490 -12895
rect 48535 -13015 48655 -12895
rect 48710 -13015 48830 -12895
rect 48875 -13015 48995 -12895
rect 49040 -13015 49160 -12895
rect 49205 -13015 49325 -12895
rect 49380 -13015 49500 -12895
rect 49545 -13015 49665 -12895
rect 49710 -13015 49830 -12895
rect 49875 -13015 49995 -12895
rect 50050 -13015 50170 -12895
rect 50215 -13015 50335 -12895
rect 50380 -13015 50500 -12895
rect 50545 -13015 50665 -12895
rect 50720 -13015 50840 -12895
rect 50885 -13015 51005 -12895
rect 51050 -13015 51170 -12895
rect 51215 -13015 51335 -12895
rect 51390 -13015 51510 -12895
rect 51555 -13015 51675 -12895
rect 51720 -13015 51840 -12895
rect 51885 -13015 52005 -12895
rect 52060 -13015 52180 -12895
rect 52225 -13015 52345 -12895
rect 52390 -13015 52510 -12895
rect 52555 -13015 52675 -12895
rect 52730 -13015 52850 -12895
rect 52895 -13015 53015 -12895
rect 53060 -13015 53180 -12895
rect 53225 -13015 53345 -12895
rect 47865 -13180 47985 -13060
rect 48040 -13180 48160 -13060
rect 48205 -13180 48325 -13060
rect 48370 -13180 48490 -13060
rect 48535 -13180 48655 -13060
rect 48710 -13180 48830 -13060
rect 48875 -13180 48995 -13060
rect 49040 -13180 49160 -13060
rect 49205 -13180 49325 -13060
rect 49380 -13180 49500 -13060
rect 49545 -13180 49665 -13060
rect 49710 -13180 49830 -13060
rect 49875 -13180 49995 -13060
rect 50050 -13180 50170 -13060
rect 50215 -13180 50335 -13060
rect 50380 -13180 50500 -13060
rect 50545 -13180 50665 -13060
rect 50720 -13180 50840 -13060
rect 50885 -13180 51005 -13060
rect 51050 -13180 51170 -13060
rect 51215 -13180 51335 -13060
rect 51390 -13180 51510 -13060
rect 51555 -13180 51675 -13060
rect 51720 -13180 51840 -13060
rect 51885 -13180 52005 -13060
rect 52060 -13180 52180 -13060
rect 52225 -13180 52345 -13060
rect 52390 -13180 52510 -13060
rect 52555 -13180 52675 -13060
rect 52730 -13180 52850 -13060
rect 52895 -13180 53015 -13060
rect 53060 -13180 53180 -13060
rect 53225 -13180 53345 -13060
rect 47865 -13345 47985 -13225
rect 48040 -13345 48160 -13225
rect 48205 -13345 48325 -13225
rect 48370 -13345 48490 -13225
rect 48535 -13345 48655 -13225
rect 48710 -13345 48830 -13225
rect 48875 -13345 48995 -13225
rect 49040 -13345 49160 -13225
rect 49205 -13345 49325 -13225
rect 49380 -13345 49500 -13225
rect 49545 -13345 49665 -13225
rect 49710 -13345 49830 -13225
rect 49875 -13345 49995 -13225
rect 50050 -13345 50170 -13225
rect 50215 -13345 50335 -13225
rect 50380 -13345 50500 -13225
rect 50545 -13345 50665 -13225
rect 50720 -13345 50840 -13225
rect 50885 -13345 51005 -13225
rect 51050 -13345 51170 -13225
rect 51215 -13345 51335 -13225
rect 51390 -13345 51510 -13225
rect 51555 -13345 51675 -13225
rect 51720 -13345 51840 -13225
rect 51885 -13345 52005 -13225
rect 52060 -13345 52180 -13225
rect 52225 -13345 52345 -13225
rect 52390 -13345 52510 -13225
rect 52555 -13345 52675 -13225
rect 52730 -13345 52850 -13225
rect 52895 -13345 53015 -13225
rect 53060 -13345 53180 -13225
rect 53225 -13345 53345 -13225
rect 47865 -13520 47985 -13400
rect 48040 -13520 48160 -13400
rect 48205 -13520 48325 -13400
rect 48370 -13520 48490 -13400
rect 48535 -13520 48655 -13400
rect 48710 -13520 48830 -13400
rect 48875 -13520 48995 -13400
rect 49040 -13520 49160 -13400
rect 49205 -13520 49325 -13400
rect 49380 -13520 49500 -13400
rect 49545 -13520 49665 -13400
rect 49710 -13520 49830 -13400
rect 49875 -13520 49995 -13400
rect 50050 -13520 50170 -13400
rect 50215 -13520 50335 -13400
rect 50380 -13520 50500 -13400
rect 50545 -13520 50665 -13400
rect 50720 -13520 50840 -13400
rect 50885 -13520 51005 -13400
rect 51050 -13520 51170 -13400
rect 51215 -13520 51335 -13400
rect 51390 -13520 51510 -13400
rect 51555 -13520 51675 -13400
rect 51720 -13520 51840 -13400
rect 51885 -13520 52005 -13400
rect 52060 -13520 52180 -13400
rect 52225 -13520 52345 -13400
rect 52390 -13520 52510 -13400
rect 52555 -13520 52675 -13400
rect 52730 -13520 52850 -13400
rect 52895 -13520 53015 -13400
rect 53060 -13520 53180 -13400
rect 53225 -13520 53345 -13400
rect 47865 -13685 47985 -13565
rect 48040 -13685 48160 -13565
rect 48205 -13685 48325 -13565
rect 48370 -13685 48490 -13565
rect 48535 -13685 48655 -13565
rect 48710 -13685 48830 -13565
rect 48875 -13685 48995 -13565
rect 49040 -13685 49160 -13565
rect 49205 -13685 49325 -13565
rect 49380 -13685 49500 -13565
rect 49545 -13685 49665 -13565
rect 49710 -13685 49830 -13565
rect 49875 -13685 49995 -13565
rect 50050 -13685 50170 -13565
rect 50215 -13685 50335 -13565
rect 50380 -13685 50500 -13565
rect 50545 -13685 50665 -13565
rect 50720 -13685 50840 -13565
rect 50885 -13685 51005 -13565
rect 51050 -13685 51170 -13565
rect 51215 -13685 51335 -13565
rect 51390 -13685 51510 -13565
rect 51555 -13685 51675 -13565
rect 51720 -13685 51840 -13565
rect 51885 -13685 52005 -13565
rect 52060 -13685 52180 -13565
rect 52225 -13685 52345 -13565
rect 52390 -13685 52510 -13565
rect 52555 -13685 52675 -13565
rect 52730 -13685 52850 -13565
rect 52895 -13685 53015 -13565
rect 53060 -13685 53180 -13565
rect 53225 -13685 53345 -13565
rect 47865 -13850 47985 -13730
rect 48040 -13850 48160 -13730
rect 48205 -13850 48325 -13730
rect 48370 -13850 48490 -13730
rect 48535 -13850 48655 -13730
rect 48710 -13850 48830 -13730
rect 48875 -13850 48995 -13730
rect 49040 -13850 49160 -13730
rect 49205 -13850 49325 -13730
rect 49380 -13850 49500 -13730
rect 49545 -13850 49665 -13730
rect 49710 -13850 49830 -13730
rect 49875 -13850 49995 -13730
rect 50050 -13850 50170 -13730
rect 50215 -13850 50335 -13730
rect 50380 -13850 50500 -13730
rect 50545 -13850 50665 -13730
rect 50720 -13850 50840 -13730
rect 50885 -13850 51005 -13730
rect 51050 -13850 51170 -13730
rect 51215 -13850 51335 -13730
rect 51390 -13850 51510 -13730
rect 51555 -13850 51675 -13730
rect 51720 -13850 51840 -13730
rect 51885 -13850 52005 -13730
rect 52060 -13850 52180 -13730
rect 52225 -13850 52345 -13730
rect 52390 -13850 52510 -13730
rect 52555 -13850 52675 -13730
rect 52730 -13850 52850 -13730
rect 52895 -13850 53015 -13730
rect 53060 -13850 53180 -13730
rect 53225 -13850 53345 -13730
rect 47865 -14015 47985 -13895
rect 48040 -14015 48160 -13895
rect 48205 -14015 48325 -13895
rect 48370 -14015 48490 -13895
rect 48535 -14015 48655 -13895
rect 48710 -14015 48830 -13895
rect 48875 -14015 48995 -13895
rect 49040 -14015 49160 -13895
rect 49205 -14015 49325 -13895
rect 49380 -14015 49500 -13895
rect 49545 -14015 49665 -13895
rect 49710 -14015 49830 -13895
rect 49875 -14015 49995 -13895
rect 50050 -14015 50170 -13895
rect 50215 -14015 50335 -13895
rect 50380 -14015 50500 -13895
rect 50545 -14015 50665 -13895
rect 50720 -14015 50840 -13895
rect 50885 -14015 51005 -13895
rect 51050 -14015 51170 -13895
rect 51215 -14015 51335 -13895
rect 51390 -14015 51510 -13895
rect 51555 -14015 51675 -13895
rect 51720 -14015 51840 -13895
rect 51885 -14015 52005 -13895
rect 52060 -14015 52180 -13895
rect 52225 -14015 52345 -13895
rect 52390 -14015 52510 -13895
rect 52555 -14015 52675 -13895
rect 52730 -14015 52850 -13895
rect 52895 -14015 53015 -13895
rect 53060 -14015 53180 -13895
rect 53225 -14015 53345 -13895
rect 47865 -14190 47985 -14070
rect 48040 -14190 48160 -14070
rect 48205 -14190 48325 -14070
rect 48370 -14190 48490 -14070
rect 48535 -14190 48655 -14070
rect 48710 -14190 48830 -14070
rect 48875 -14190 48995 -14070
rect 49040 -14190 49160 -14070
rect 49205 -14190 49325 -14070
rect 49380 -14190 49500 -14070
rect 49545 -14190 49665 -14070
rect 49710 -14190 49830 -14070
rect 49875 -14190 49995 -14070
rect 50050 -14190 50170 -14070
rect 50215 -14190 50335 -14070
rect 50380 -14190 50500 -14070
rect 50545 -14190 50665 -14070
rect 50720 -14190 50840 -14070
rect 50885 -14190 51005 -14070
rect 51050 -14190 51170 -14070
rect 51215 -14190 51335 -14070
rect 51390 -14190 51510 -14070
rect 51555 -14190 51675 -14070
rect 51720 -14190 51840 -14070
rect 51885 -14190 52005 -14070
rect 52060 -14190 52180 -14070
rect 52225 -14190 52345 -14070
rect 52390 -14190 52510 -14070
rect 52555 -14190 52675 -14070
rect 52730 -14190 52850 -14070
rect 52895 -14190 53015 -14070
rect 53060 -14190 53180 -14070
rect 53225 -14190 53345 -14070
rect 47865 -14355 47985 -14235
rect 48040 -14355 48160 -14235
rect 48205 -14355 48325 -14235
rect 48370 -14355 48490 -14235
rect 48535 -14355 48655 -14235
rect 48710 -14355 48830 -14235
rect 48875 -14355 48995 -14235
rect 49040 -14355 49160 -14235
rect 49205 -14355 49325 -14235
rect 49380 -14355 49500 -14235
rect 49545 -14355 49665 -14235
rect 49710 -14355 49830 -14235
rect 49875 -14355 49995 -14235
rect 50050 -14355 50170 -14235
rect 50215 -14355 50335 -14235
rect 50380 -14355 50500 -14235
rect 50545 -14355 50665 -14235
rect 50720 -14355 50840 -14235
rect 50885 -14355 51005 -14235
rect 51050 -14355 51170 -14235
rect 51215 -14355 51335 -14235
rect 51390 -14355 51510 -14235
rect 51555 -14355 51675 -14235
rect 51720 -14355 51840 -14235
rect 51885 -14355 52005 -14235
rect 52060 -14355 52180 -14235
rect 52225 -14355 52345 -14235
rect 52390 -14355 52510 -14235
rect 52555 -14355 52675 -14235
rect 52730 -14355 52850 -14235
rect 52895 -14355 53015 -14235
rect 53060 -14355 53180 -14235
rect 53225 -14355 53345 -14235
rect 47865 -14520 47985 -14400
rect 48040 -14520 48160 -14400
rect 48205 -14520 48325 -14400
rect 48370 -14520 48490 -14400
rect 48535 -14520 48655 -14400
rect 48710 -14520 48830 -14400
rect 48875 -14520 48995 -14400
rect 49040 -14520 49160 -14400
rect 49205 -14520 49325 -14400
rect 49380 -14520 49500 -14400
rect 49545 -14520 49665 -14400
rect 49710 -14520 49830 -14400
rect 49875 -14520 49995 -14400
rect 50050 -14520 50170 -14400
rect 50215 -14520 50335 -14400
rect 50380 -14520 50500 -14400
rect 50545 -14520 50665 -14400
rect 50720 -14520 50840 -14400
rect 50885 -14520 51005 -14400
rect 51050 -14520 51170 -14400
rect 51215 -14520 51335 -14400
rect 51390 -14520 51510 -14400
rect 51555 -14520 51675 -14400
rect 51720 -14520 51840 -14400
rect 51885 -14520 52005 -14400
rect 52060 -14520 52180 -14400
rect 52225 -14520 52345 -14400
rect 52390 -14520 52510 -14400
rect 52555 -14520 52675 -14400
rect 52730 -14520 52850 -14400
rect 52895 -14520 53015 -14400
rect 53060 -14520 53180 -14400
rect 53225 -14520 53345 -14400
rect 47865 -14685 47985 -14565
rect 48040 -14685 48160 -14565
rect 48205 -14685 48325 -14565
rect 48370 -14685 48490 -14565
rect 48535 -14685 48655 -14565
rect 48710 -14685 48830 -14565
rect 48875 -14685 48995 -14565
rect 49040 -14685 49160 -14565
rect 49205 -14685 49325 -14565
rect 49380 -14685 49500 -14565
rect 49545 -14685 49665 -14565
rect 49710 -14685 49830 -14565
rect 49875 -14685 49995 -14565
rect 50050 -14685 50170 -14565
rect 50215 -14685 50335 -14565
rect 50380 -14685 50500 -14565
rect 50545 -14685 50665 -14565
rect 50720 -14685 50840 -14565
rect 50885 -14685 51005 -14565
rect 51050 -14685 51170 -14565
rect 51215 -14685 51335 -14565
rect 51390 -14685 51510 -14565
rect 51555 -14685 51675 -14565
rect 51720 -14685 51840 -14565
rect 51885 -14685 52005 -14565
rect 52060 -14685 52180 -14565
rect 52225 -14685 52345 -14565
rect 52390 -14685 52510 -14565
rect 52555 -14685 52675 -14565
rect 52730 -14685 52850 -14565
rect 52895 -14685 53015 -14565
rect 53060 -14685 53180 -14565
rect 53225 -14685 53345 -14565
rect 47865 -14860 47985 -14740
rect 48040 -14860 48160 -14740
rect 48205 -14860 48325 -14740
rect 48370 -14860 48490 -14740
rect 48535 -14860 48655 -14740
rect 48710 -14860 48830 -14740
rect 48875 -14860 48995 -14740
rect 49040 -14860 49160 -14740
rect 49205 -14860 49325 -14740
rect 49380 -14860 49500 -14740
rect 49545 -14860 49665 -14740
rect 49710 -14860 49830 -14740
rect 49875 -14860 49995 -14740
rect 50050 -14860 50170 -14740
rect 50215 -14860 50335 -14740
rect 50380 -14860 50500 -14740
rect 50545 -14860 50665 -14740
rect 50720 -14860 50840 -14740
rect 50885 -14860 51005 -14740
rect 51050 -14860 51170 -14740
rect 51215 -14860 51335 -14740
rect 51390 -14860 51510 -14740
rect 51555 -14860 51675 -14740
rect 51720 -14860 51840 -14740
rect 51885 -14860 52005 -14740
rect 52060 -14860 52180 -14740
rect 52225 -14860 52345 -14740
rect 52390 -14860 52510 -14740
rect 52555 -14860 52675 -14740
rect 52730 -14860 52850 -14740
rect 52895 -14860 53015 -14740
rect 53060 -14860 53180 -14740
rect 53225 -14860 53345 -14740
rect 47865 -15025 47985 -14905
rect 48040 -15025 48160 -14905
rect 48205 -15025 48325 -14905
rect 48370 -15025 48490 -14905
rect 48535 -15025 48655 -14905
rect 48710 -15025 48830 -14905
rect 48875 -15025 48995 -14905
rect 49040 -15025 49160 -14905
rect 49205 -15025 49325 -14905
rect 49380 -15025 49500 -14905
rect 49545 -15025 49665 -14905
rect 49710 -15025 49830 -14905
rect 49875 -15025 49995 -14905
rect 50050 -15025 50170 -14905
rect 50215 -15025 50335 -14905
rect 50380 -15025 50500 -14905
rect 50545 -15025 50665 -14905
rect 50720 -15025 50840 -14905
rect 50885 -15025 51005 -14905
rect 51050 -15025 51170 -14905
rect 51215 -15025 51335 -14905
rect 51390 -15025 51510 -14905
rect 51555 -15025 51675 -14905
rect 51720 -15025 51840 -14905
rect 51885 -15025 52005 -14905
rect 52060 -15025 52180 -14905
rect 52225 -15025 52345 -14905
rect 52390 -15025 52510 -14905
rect 52555 -15025 52675 -14905
rect 52730 -15025 52850 -14905
rect 52895 -15025 53015 -14905
rect 53060 -15025 53180 -14905
rect 53225 -15025 53345 -14905
rect 47865 -15190 47985 -15070
rect 48040 -15190 48160 -15070
rect 48205 -15190 48325 -15070
rect 48370 -15190 48490 -15070
rect 48535 -15190 48655 -15070
rect 48710 -15190 48830 -15070
rect 48875 -15190 48995 -15070
rect 49040 -15190 49160 -15070
rect 49205 -15190 49325 -15070
rect 49380 -15190 49500 -15070
rect 49545 -15190 49665 -15070
rect 49710 -15190 49830 -15070
rect 49875 -15190 49995 -15070
rect 50050 -15190 50170 -15070
rect 50215 -15190 50335 -15070
rect 50380 -15190 50500 -15070
rect 50545 -15190 50665 -15070
rect 50720 -15190 50840 -15070
rect 50885 -15190 51005 -15070
rect 51050 -15190 51170 -15070
rect 51215 -15190 51335 -15070
rect 51390 -15190 51510 -15070
rect 51555 -15190 51675 -15070
rect 51720 -15190 51840 -15070
rect 51885 -15190 52005 -15070
rect 52060 -15190 52180 -15070
rect 52225 -15190 52345 -15070
rect 52390 -15190 52510 -15070
rect 52555 -15190 52675 -15070
rect 52730 -15190 52850 -15070
rect 52895 -15190 53015 -15070
rect 53060 -15190 53180 -15070
rect 53225 -15190 53345 -15070
rect 47865 -15355 47985 -15235
rect 48040 -15355 48160 -15235
rect 48205 -15355 48325 -15235
rect 48370 -15355 48490 -15235
rect 48535 -15355 48655 -15235
rect 48710 -15355 48830 -15235
rect 48875 -15355 48995 -15235
rect 49040 -15355 49160 -15235
rect 49205 -15355 49325 -15235
rect 49380 -15355 49500 -15235
rect 49545 -15355 49665 -15235
rect 49710 -15355 49830 -15235
rect 49875 -15355 49995 -15235
rect 50050 -15355 50170 -15235
rect 50215 -15355 50335 -15235
rect 50380 -15355 50500 -15235
rect 50545 -15355 50665 -15235
rect 50720 -15355 50840 -15235
rect 50885 -15355 51005 -15235
rect 51050 -15355 51170 -15235
rect 51215 -15355 51335 -15235
rect 51390 -15355 51510 -15235
rect 51555 -15355 51675 -15235
rect 51720 -15355 51840 -15235
rect 51885 -15355 52005 -15235
rect 52060 -15355 52180 -15235
rect 52225 -15355 52345 -15235
rect 52390 -15355 52510 -15235
rect 52555 -15355 52675 -15235
rect 52730 -15355 52850 -15235
rect 52895 -15355 53015 -15235
rect 53060 -15355 53180 -15235
rect 53225 -15355 53345 -15235
rect 47865 -15530 47985 -15410
rect 48040 -15530 48160 -15410
rect 48205 -15530 48325 -15410
rect 48370 -15530 48490 -15410
rect 48535 -15530 48655 -15410
rect 48710 -15530 48830 -15410
rect 48875 -15530 48995 -15410
rect 49040 -15530 49160 -15410
rect 49205 -15530 49325 -15410
rect 49380 -15530 49500 -15410
rect 49545 -15530 49665 -15410
rect 49710 -15530 49830 -15410
rect 49875 -15530 49995 -15410
rect 50050 -15530 50170 -15410
rect 50215 -15530 50335 -15410
rect 50380 -15530 50500 -15410
rect 50545 -15530 50665 -15410
rect 50720 -15530 50840 -15410
rect 50885 -15530 51005 -15410
rect 51050 -15530 51170 -15410
rect 51215 -15530 51335 -15410
rect 51390 -15530 51510 -15410
rect 51555 -15530 51675 -15410
rect 51720 -15530 51840 -15410
rect 51885 -15530 52005 -15410
rect 52060 -15530 52180 -15410
rect 52225 -15530 52345 -15410
rect 52390 -15530 52510 -15410
rect 52555 -15530 52675 -15410
rect 52730 -15530 52850 -15410
rect 52895 -15530 53015 -15410
rect 53060 -15530 53180 -15410
rect 53225 -15530 53345 -15410
<< metal5 >>
rect 30770 7200 53370 7225
rect 30770 7080 30795 7200
rect 30915 7080 30960 7200
rect 31080 7080 31125 7200
rect 31245 7080 31290 7200
rect 31410 7080 31465 7200
rect 31585 7080 31630 7200
rect 31750 7080 31795 7200
rect 31915 7080 31960 7200
rect 32080 7080 32135 7200
rect 32255 7080 32300 7200
rect 32420 7080 32465 7200
rect 32585 7080 32630 7200
rect 32750 7080 32805 7200
rect 32925 7080 32970 7200
rect 33090 7080 33135 7200
rect 33255 7080 33300 7200
rect 33420 7080 33475 7200
rect 33595 7080 33640 7200
rect 33760 7080 33805 7200
rect 33925 7080 33970 7200
rect 34090 7080 34145 7200
rect 34265 7080 34310 7200
rect 34430 7080 34475 7200
rect 34595 7080 34640 7200
rect 34760 7080 34815 7200
rect 34935 7080 34980 7200
rect 35100 7080 35145 7200
rect 35265 7080 35310 7200
rect 35430 7080 35485 7200
rect 35605 7080 35650 7200
rect 35770 7080 35815 7200
rect 35935 7080 35980 7200
rect 36100 7080 36155 7200
rect 36275 7080 36485 7200
rect 36605 7080 36650 7200
rect 36770 7080 36815 7200
rect 36935 7080 36980 7200
rect 37100 7080 37155 7200
rect 37275 7080 37320 7200
rect 37440 7080 37485 7200
rect 37605 7080 37650 7200
rect 37770 7080 37825 7200
rect 37945 7080 37990 7200
rect 38110 7080 38155 7200
rect 38275 7080 38320 7200
rect 38440 7080 38495 7200
rect 38615 7080 38660 7200
rect 38780 7080 38825 7200
rect 38945 7080 38990 7200
rect 39110 7080 39165 7200
rect 39285 7080 39330 7200
rect 39450 7080 39495 7200
rect 39615 7080 39660 7200
rect 39780 7080 39835 7200
rect 39955 7080 40000 7200
rect 40120 7080 40165 7200
rect 40285 7080 40330 7200
rect 40450 7080 40505 7200
rect 40625 7080 40670 7200
rect 40790 7080 40835 7200
rect 40955 7080 41000 7200
rect 41120 7080 41175 7200
rect 41295 7080 41340 7200
rect 41460 7080 41505 7200
rect 41625 7080 41670 7200
rect 41790 7080 41845 7200
rect 41965 7080 42175 7200
rect 42295 7080 42340 7200
rect 42460 7080 42505 7200
rect 42625 7080 42670 7200
rect 42790 7080 42845 7200
rect 42965 7080 43010 7200
rect 43130 7080 43175 7200
rect 43295 7080 43340 7200
rect 43460 7080 43515 7200
rect 43635 7080 43680 7200
rect 43800 7080 43845 7200
rect 43965 7080 44010 7200
rect 44130 7080 44185 7200
rect 44305 7080 44350 7200
rect 44470 7080 44515 7200
rect 44635 7080 44680 7200
rect 44800 7080 44855 7200
rect 44975 7080 45020 7200
rect 45140 7080 45185 7200
rect 45305 7080 45350 7200
rect 45470 7080 45525 7200
rect 45645 7080 45690 7200
rect 45810 7080 45855 7200
rect 45975 7080 46020 7200
rect 46140 7080 46195 7200
rect 46315 7080 46360 7200
rect 46480 7080 46525 7200
rect 46645 7080 46690 7200
rect 46810 7080 46865 7200
rect 46985 7080 47030 7200
rect 47150 7080 47195 7200
rect 47315 7080 47360 7200
rect 47480 7080 47535 7200
rect 47655 7080 47865 7200
rect 47985 7080 48030 7200
rect 48150 7080 48195 7200
rect 48315 7080 48360 7200
rect 48480 7080 48535 7200
rect 48655 7080 48700 7200
rect 48820 7080 48865 7200
rect 48985 7080 49030 7200
rect 49150 7080 49205 7200
rect 49325 7080 49370 7200
rect 49490 7080 49535 7200
rect 49655 7080 49700 7200
rect 49820 7080 49875 7200
rect 49995 7080 50040 7200
rect 50160 7080 50205 7200
rect 50325 7080 50370 7200
rect 50490 7080 50545 7200
rect 50665 7080 50710 7200
rect 50830 7080 50875 7200
rect 50995 7080 51040 7200
rect 51160 7080 51215 7200
rect 51335 7080 51380 7200
rect 51500 7080 51545 7200
rect 51665 7080 51710 7200
rect 51830 7080 51885 7200
rect 52005 7080 52050 7200
rect 52170 7080 52215 7200
rect 52335 7080 52380 7200
rect 52500 7080 52555 7200
rect 52675 7080 52720 7200
rect 52840 7080 52885 7200
rect 53005 7080 53050 7200
rect 53170 7080 53225 7200
rect 53345 7080 53370 7200
rect 30770 7025 53370 7080
rect 30770 6905 30795 7025
rect 30915 6905 30960 7025
rect 31080 6905 31125 7025
rect 31245 6905 31290 7025
rect 31410 6905 31465 7025
rect 31585 6905 31630 7025
rect 31750 6905 31795 7025
rect 31915 6905 31960 7025
rect 32080 6905 32135 7025
rect 32255 6905 32300 7025
rect 32420 6905 32465 7025
rect 32585 6905 32630 7025
rect 32750 6905 32805 7025
rect 32925 6905 32970 7025
rect 33090 6905 33135 7025
rect 33255 6905 33300 7025
rect 33420 6905 33475 7025
rect 33595 6905 33640 7025
rect 33760 6905 33805 7025
rect 33925 6905 33970 7025
rect 34090 6905 34145 7025
rect 34265 6905 34310 7025
rect 34430 6905 34475 7025
rect 34595 6905 34640 7025
rect 34760 6905 34815 7025
rect 34935 6905 34980 7025
rect 35100 6905 35145 7025
rect 35265 6905 35310 7025
rect 35430 6905 35485 7025
rect 35605 6905 35650 7025
rect 35770 6905 35815 7025
rect 35935 6905 35980 7025
rect 36100 6905 36155 7025
rect 36275 6905 36485 7025
rect 36605 6905 36650 7025
rect 36770 6905 36815 7025
rect 36935 6905 36980 7025
rect 37100 6905 37155 7025
rect 37275 6905 37320 7025
rect 37440 6905 37485 7025
rect 37605 6905 37650 7025
rect 37770 6905 37825 7025
rect 37945 6905 37990 7025
rect 38110 6905 38155 7025
rect 38275 6905 38320 7025
rect 38440 6905 38495 7025
rect 38615 6905 38660 7025
rect 38780 6905 38825 7025
rect 38945 6905 38990 7025
rect 39110 6905 39165 7025
rect 39285 6905 39330 7025
rect 39450 6905 39495 7025
rect 39615 6905 39660 7025
rect 39780 6905 39835 7025
rect 39955 6905 40000 7025
rect 40120 6905 40165 7025
rect 40285 6905 40330 7025
rect 40450 6905 40505 7025
rect 40625 6905 40670 7025
rect 40790 6905 40835 7025
rect 40955 6905 41000 7025
rect 41120 6905 41175 7025
rect 41295 6905 41340 7025
rect 41460 6905 41505 7025
rect 41625 6905 41670 7025
rect 41790 6905 41845 7025
rect 41965 6905 42175 7025
rect 42295 6905 42340 7025
rect 42460 6905 42505 7025
rect 42625 6905 42670 7025
rect 42790 6905 42845 7025
rect 42965 6905 43010 7025
rect 43130 6905 43175 7025
rect 43295 6905 43340 7025
rect 43460 6905 43515 7025
rect 43635 6905 43680 7025
rect 43800 6905 43845 7025
rect 43965 6905 44010 7025
rect 44130 6905 44185 7025
rect 44305 6905 44350 7025
rect 44470 6905 44515 7025
rect 44635 6905 44680 7025
rect 44800 6905 44855 7025
rect 44975 6905 45020 7025
rect 45140 6905 45185 7025
rect 45305 6905 45350 7025
rect 45470 6905 45525 7025
rect 45645 6905 45690 7025
rect 45810 6905 45855 7025
rect 45975 6905 46020 7025
rect 46140 6905 46195 7025
rect 46315 6905 46360 7025
rect 46480 6905 46525 7025
rect 46645 6905 46690 7025
rect 46810 6905 46865 7025
rect 46985 6905 47030 7025
rect 47150 6905 47195 7025
rect 47315 6905 47360 7025
rect 47480 6905 47535 7025
rect 47655 6905 47865 7025
rect 47985 6905 48030 7025
rect 48150 6905 48195 7025
rect 48315 6905 48360 7025
rect 48480 6905 48535 7025
rect 48655 6905 48700 7025
rect 48820 6905 48865 7025
rect 48985 6905 49030 7025
rect 49150 6905 49205 7025
rect 49325 6905 49370 7025
rect 49490 6905 49535 7025
rect 49655 6905 49700 7025
rect 49820 6905 49875 7025
rect 49995 6905 50040 7025
rect 50160 6905 50205 7025
rect 50325 6905 50370 7025
rect 50490 6905 50545 7025
rect 50665 6905 50710 7025
rect 50830 6905 50875 7025
rect 50995 6905 51040 7025
rect 51160 6905 51215 7025
rect 51335 6905 51380 7025
rect 51500 6905 51545 7025
rect 51665 6905 51710 7025
rect 51830 6905 51885 7025
rect 52005 6905 52050 7025
rect 52170 6905 52215 7025
rect 52335 6905 52380 7025
rect 52500 6905 52555 7025
rect 52675 6905 52720 7025
rect 52840 6905 52885 7025
rect 53005 6905 53050 7025
rect 53170 6905 53225 7025
rect 53345 6905 53370 7025
rect 30770 6860 53370 6905
rect 30770 6740 30795 6860
rect 30915 6740 30960 6860
rect 31080 6740 31125 6860
rect 31245 6740 31290 6860
rect 31410 6740 31465 6860
rect 31585 6740 31630 6860
rect 31750 6740 31795 6860
rect 31915 6740 31960 6860
rect 32080 6740 32135 6860
rect 32255 6740 32300 6860
rect 32420 6740 32465 6860
rect 32585 6740 32630 6860
rect 32750 6740 32805 6860
rect 32925 6740 32970 6860
rect 33090 6740 33135 6860
rect 33255 6740 33300 6860
rect 33420 6740 33475 6860
rect 33595 6740 33640 6860
rect 33760 6740 33805 6860
rect 33925 6740 33970 6860
rect 34090 6740 34145 6860
rect 34265 6740 34310 6860
rect 34430 6740 34475 6860
rect 34595 6740 34640 6860
rect 34760 6740 34815 6860
rect 34935 6740 34980 6860
rect 35100 6740 35145 6860
rect 35265 6740 35310 6860
rect 35430 6740 35485 6860
rect 35605 6740 35650 6860
rect 35770 6740 35815 6860
rect 35935 6740 35980 6860
rect 36100 6740 36155 6860
rect 36275 6740 36485 6860
rect 36605 6740 36650 6860
rect 36770 6740 36815 6860
rect 36935 6740 36980 6860
rect 37100 6740 37155 6860
rect 37275 6740 37320 6860
rect 37440 6740 37485 6860
rect 37605 6740 37650 6860
rect 37770 6740 37825 6860
rect 37945 6740 37990 6860
rect 38110 6740 38155 6860
rect 38275 6740 38320 6860
rect 38440 6740 38495 6860
rect 38615 6740 38660 6860
rect 38780 6740 38825 6860
rect 38945 6740 38990 6860
rect 39110 6740 39165 6860
rect 39285 6740 39330 6860
rect 39450 6740 39495 6860
rect 39615 6740 39660 6860
rect 39780 6740 39835 6860
rect 39955 6740 40000 6860
rect 40120 6740 40165 6860
rect 40285 6740 40330 6860
rect 40450 6740 40505 6860
rect 40625 6740 40670 6860
rect 40790 6740 40835 6860
rect 40955 6740 41000 6860
rect 41120 6740 41175 6860
rect 41295 6740 41340 6860
rect 41460 6740 41505 6860
rect 41625 6740 41670 6860
rect 41790 6740 41845 6860
rect 41965 6740 42175 6860
rect 42295 6740 42340 6860
rect 42460 6740 42505 6860
rect 42625 6740 42670 6860
rect 42790 6740 42845 6860
rect 42965 6740 43010 6860
rect 43130 6740 43175 6860
rect 43295 6740 43340 6860
rect 43460 6740 43515 6860
rect 43635 6740 43680 6860
rect 43800 6740 43845 6860
rect 43965 6740 44010 6860
rect 44130 6740 44185 6860
rect 44305 6740 44350 6860
rect 44470 6740 44515 6860
rect 44635 6740 44680 6860
rect 44800 6740 44855 6860
rect 44975 6740 45020 6860
rect 45140 6740 45185 6860
rect 45305 6740 45350 6860
rect 45470 6740 45525 6860
rect 45645 6740 45690 6860
rect 45810 6740 45855 6860
rect 45975 6740 46020 6860
rect 46140 6740 46195 6860
rect 46315 6740 46360 6860
rect 46480 6740 46525 6860
rect 46645 6740 46690 6860
rect 46810 6740 46865 6860
rect 46985 6740 47030 6860
rect 47150 6740 47195 6860
rect 47315 6740 47360 6860
rect 47480 6740 47535 6860
rect 47655 6740 47865 6860
rect 47985 6740 48030 6860
rect 48150 6740 48195 6860
rect 48315 6740 48360 6860
rect 48480 6740 48535 6860
rect 48655 6740 48700 6860
rect 48820 6740 48865 6860
rect 48985 6740 49030 6860
rect 49150 6740 49205 6860
rect 49325 6740 49370 6860
rect 49490 6740 49535 6860
rect 49655 6740 49700 6860
rect 49820 6740 49875 6860
rect 49995 6740 50040 6860
rect 50160 6740 50205 6860
rect 50325 6740 50370 6860
rect 50490 6740 50545 6860
rect 50665 6740 50710 6860
rect 50830 6740 50875 6860
rect 50995 6740 51040 6860
rect 51160 6740 51215 6860
rect 51335 6740 51380 6860
rect 51500 6740 51545 6860
rect 51665 6740 51710 6860
rect 51830 6740 51885 6860
rect 52005 6740 52050 6860
rect 52170 6740 52215 6860
rect 52335 6740 52380 6860
rect 52500 6740 52555 6860
rect 52675 6740 52720 6860
rect 52840 6740 52885 6860
rect 53005 6740 53050 6860
rect 53170 6740 53225 6860
rect 53345 6740 53370 6860
rect 30770 6695 53370 6740
rect 30770 6575 30795 6695
rect 30915 6575 30960 6695
rect 31080 6575 31125 6695
rect 31245 6575 31290 6695
rect 31410 6575 31465 6695
rect 31585 6575 31630 6695
rect 31750 6575 31795 6695
rect 31915 6575 31960 6695
rect 32080 6575 32135 6695
rect 32255 6575 32300 6695
rect 32420 6575 32465 6695
rect 32585 6575 32630 6695
rect 32750 6575 32805 6695
rect 32925 6575 32970 6695
rect 33090 6575 33135 6695
rect 33255 6575 33300 6695
rect 33420 6575 33475 6695
rect 33595 6575 33640 6695
rect 33760 6575 33805 6695
rect 33925 6575 33970 6695
rect 34090 6575 34145 6695
rect 34265 6575 34310 6695
rect 34430 6575 34475 6695
rect 34595 6575 34640 6695
rect 34760 6575 34815 6695
rect 34935 6575 34980 6695
rect 35100 6575 35145 6695
rect 35265 6575 35310 6695
rect 35430 6575 35485 6695
rect 35605 6575 35650 6695
rect 35770 6575 35815 6695
rect 35935 6575 35980 6695
rect 36100 6575 36155 6695
rect 36275 6575 36485 6695
rect 36605 6575 36650 6695
rect 36770 6575 36815 6695
rect 36935 6575 36980 6695
rect 37100 6575 37155 6695
rect 37275 6575 37320 6695
rect 37440 6575 37485 6695
rect 37605 6575 37650 6695
rect 37770 6575 37825 6695
rect 37945 6575 37990 6695
rect 38110 6575 38155 6695
rect 38275 6575 38320 6695
rect 38440 6575 38495 6695
rect 38615 6575 38660 6695
rect 38780 6575 38825 6695
rect 38945 6575 38990 6695
rect 39110 6575 39165 6695
rect 39285 6575 39330 6695
rect 39450 6575 39495 6695
rect 39615 6575 39660 6695
rect 39780 6575 39835 6695
rect 39955 6575 40000 6695
rect 40120 6575 40165 6695
rect 40285 6575 40330 6695
rect 40450 6575 40505 6695
rect 40625 6575 40670 6695
rect 40790 6575 40835 6695
rect 40955 6575 41000 6695
rect 41120 6575 41175 6695
rect 41295 6575 41340 6695
rect 41460 6575 41505 6695
rect 41625 6575 41670 6695
rect 41790 6575 41845 6695
rect 41965 6575 42175 6695
rect 42295 6575 42340 6695
rect 42460 6575 42505 6695
rect 42625 6575 42670 6695
rect 42790 6575 42845 6695
rect 42965 6575 43010 6695
rect 43130 6575 43175 6695
rect 43295 6575 43340 6695
rect 43460 6575 43515 6695
rect 43635 6575 43680 6695
rect 43800 6575 43845 6695
rect 43965 6575 44010 6695
rect 44130 6575 44185 6695
rect 44305 6575 44350 6695
rect 44470 6575 44515 6695
rect 44635 6575 44680 6695
rect 44800 6575 44855 6695
rect 44975 6575 45020 6695
rect 45140 6575 45185 6695
rect 45305 6575 45350 6695
rect 45470 6575 45525 6695
rect 45645 6575 45690 6695
rect 45810 6575 45855 6695
rect 45975 6575 46020 6695
rect 46140 6575 46195 6695
rect 46315 6575 46360 6695
rect 46480 6575 46525 6695
rect 46645 6575 46690 6695
rect 46810 6575 46865 6695
rect 46985 6575 47030 6695
rect 47150 6575 47195 6695
rect 47315 6575 47360 6695
rect 47480 6575 47535 6695
rect 47655 6575 47865 6695
rect 47985 6575 48030 6695
rect 48150 6575 48195 6695
rect 48315 6575 48360 6695
rect 48480 6575 48535 6695
rect 48655 6575 48700 6695
rect 48820 6575 48865 6695
rect 48985 6575 49030 6695
rect 49150 6575 49205 6695
rect 49325 6575 49370 6695
rect 49490 6575 49535 6695
rect 49655 6575 49700 6695
rect 49820 6575 49875 6695
rect 49995 6575 50040 6695
rect 50160 6575 50205 6695
rect 50325 6575 50370 6695
rect 50490 6575 50545 6695
rect 50665 6575 50710 6695
rect 50830 6575 50875 6695
rect 50995 6575 51040 6695
rect 51160 6575 51215 6695
rect 51335 6575 51380 6695
rect 51500 6575 51545 6695
rect 51665 6575 51710 6695
rect 51830 6575 51885 6695
rect 52005 6575 52050 6695
rect 52170 6575 52215 6695
rect 52335 6575 52380 6695
rect 52500 6575 52555 6695
rect 52675 6575 52720 6695
rect 52840 6575 52885 6695
rect 53005 6575 53050 6695
rect 53170 6575 53225 6695
rect 53345 6575 53370 6695
rect 30770 6530 53370 6575
rect 30770 6410 30795 6530
rect 30915 6410 30960 6530
rect 31080 6410 31125 6530
rect 31245 6410 31290 6530
rect 31410 6410 31465 6530
rect 31585 6410 31630 6530
rect 31750 6410 31795 6530
rect 31915 6410 31960 6530
rect 32080 6410 32135 6530
rect 32255 6410 32300 6530
rect 32420 6410 32465 6530
rect 32585 6410 32630 6530
rect 32750 6410 32805 6530
rect 32925 6410 32970 6530
rect 33090 6410 33135 6530
rect 33255 6410 33300 6530
rect 33420 6410 33475 6530
rect 33595 6410 33640 6530
rect 33760 6410 33805 6530
rect 33925 6410 33970 6530
rect 34090 6410 34145 6530
rect 34265 6410 34310 6530
rect 34430 6410 34475 6530
rect 34595 6410 34640 6530
rect 34760 6410 34815 6530
rect 34935 6410 34980 6530
rect 35100 6410 35145 6530
rect 35265 6410 35310 6530
rect 35430 6410 35485 6530
rect 35605 6410 35650 6530
rect 35770 6410 35815 6530
rect 35935 6410 35980 6530
rect 36100 6410 36155 6530
rect 36275 6410 36485 6530
rect 36605 6410 36650 6530
rect 36770 6410 36815 6530
rect 36935 6410 36980 6530
rect 37100 6410 37155 6530
rect 37275 6410 37320 6530
rect 37440 6410 37485 6530
rect 37605 6410 37650 6530
rect 37770 6410 37825 6530
rect 37945 6410 37990 6530
rect 38110 6410 38155 6530
rect 38275 6410 38320 6530
rect 38440 6410 38495 6530
rect 38615 6410 38660 6530
rect 38780 6410 38825 6530
rect 38945 6410 38990 6530
rect 39110 6410 39165 6530
rect 39285 6410 39330 6530
rect 39450 6410 39495 6530
rect 39615 6410 39660 6530
rect 39780 6410 39835 6530
rect 39955 6410 40000 6530
rect 40120 6410 40165 6530
rect 40285 6410 40330 6530
rect 40450 6410 40505 6530
rect 40625 6410 40670 6530
rect 40790 6410 40835 6530
rect 40955 6410 41000 6530
rect 41120 6410 41175 6530
rect 41295 6410 41340 6530
rect 41460 6410 41505 6530
rect 41625 6410 41670 6530
rect 41790 6410 41845 6530
rect 41965 6410 42175 6530
rect 42295 6410 42340 6530
rect 42460 6410 42505 6530
rect 42625 6410 42670 6530
rect 42790 6410 42845 6530
rect 42965 6410 43010 6530
rect 43130 6410 43175 6530
rect 43295 6410 43340 6530
rect 43460 6410 43515 6530
rect 43635 6410 43680 6530
rect 43800 6410 43845 6530
rect 43965 6410 44010 6530
rect 44130 6410 44185 6530
rect 44305 6410 44350 6530
rect 44470 6410 44515 6530
rect 44635 6410 44680 6530
rect 44800 6410 44855 6530
rect 44975 6410 45020 6530
rect 45140 6410 45185 6530
rect 45305 6410 45350 6530
rect 45470 6410 45525 6530
rect 45645 6410 45690 6530
rect 45810 6410 45855 6530
rect 45975 6410 46020 6530
rect 46140 6410 46195 6530
rect 46315 6410 46360 6530
rect 46480 6410 46525 6530
rect 46645 6410 46690 6530
rect 46810 6410 46865 6530
rect 46985 6410 47030 6530
rect 47150 6410 47195 6530
rect 47315 6410 47360 6530
rect 47480 6410 47535 6530
rect 47655 6410 47865 6530
rect 47985 6410 48030 6530
rect 48150 6410 48195 6530
rect 48315 6410 48360 6530
rect 48480 6410 48535 6530
rect 48655 6410 48700 6530
rect 48820 6410 48865 6530
rect 48985 6410 49030 6530
rect 49150 6410 49205 6530
rect 49325 6410 49370 6530
rect 49490 6410 49535 6530
rect 49655 6410 49700 6530
rect 49820 6410 49875 6530
rect 49995 6410 50040 6530
rect 50160 6410 50205 6530
rect 50325 6410 50370 6530
rect 50490 6410 50545 6530
rect 50665 6410 50710 6530
rect 50830 6410 50875 6530
rect 50995 6410 51040 6530
rect 51160 6410 51215 6530
rect 51335 6410 51380 6530
rect 51500 6410 51545 6530
rect 51665 6410 51710 6530
rect 51830 6410 51885 6530
rect 52005 6410 52050 6530
rect 52170 6410 52215 6530
rect 52335 6410 52380 6530
rect 52500 6410 52555 6530
rect 52675 6410 52720 6530
rect 52840 6410 52885 6530
rect 53005 6410 53050 6530
rect 53170 6410 53225 6530
rect 53345 6410 53370 6530
rect 30770 6355 53370 6410
rect 30770 6235 30795 6355
rect 30915 6235 30960 6355
rect 31080 6235 31125 6355
rect 31245 6235 31290 6355
rect 31410 6235 31465 6355
rect 31585 6235 31630 6355
rect 31750 6235 31795 6355
rect 31915 6235 31960 6355
rect 32080 6235 32135 6355
rect 32255 6235 32300 6355
rect 32420 6235 32465 6355
rect 32585 6235 32630 6355
rect 32750 6235 32805 6355
rect 32925 6235 32970 6355
rect 33090 6235 33135 6355
rect 33255 6235 33300 6355
rect 33420 6235 33475 6355
rect 33595 6235 33640 6355
rect 33760 6235 33805 6355
rect 33925 6235 33970 6355
rect 34090 6235 34145 6355
rect 34265 6235 34310 6355
rect 34430 6235 34475 6355
rect 34595 6235 34640 6355
rect 34760 6235 34815 6355
rect 34935 6235 34980 6355
rect 35100 6235 35145 6355
rect 35265 6235 35310 6355
rect 35430 6235 35485 6355
rect 35605 6235 35650 6355
rect 35770 6235 35815 6355
rect 35935 6235 35980 6355
rect 36100 6235 36155 6355
rect 36275 6235 36485 6355
rect 36605 6235 36650 6355
rect 36770 6235 36815 6355
rect 36935 6235 36980 6355
rect 37100 6235 37155 6355
rect 37275 6235 37320 6355
rect 37440 6235 37485 6355
rect 37605 6235 37650 6355
rect 37770 6235 37825 6355
rect 37945 6235 37990 6355
rect 38110 6235 38155 6355
rect 38275 6235 38320 6355
rect 38440 6235 38495 6355
rect 38615 6235 38660 6355
rect 38780 6235 38825 6355
rect 38945 6235 38990 6355
rect 39110 6235 39165 6355
rect 39285 6235 39330 6355
rect 39450 6235 39495 6355
rect 39615 6235 39660 6355
rect 39780 6235 39835 6355
rect 39955 6235 40000 6355
rect 40120 6235 40165 6355
rect 40285 6235 40330 6355
rect 40450 6235 40505 6355
rect 40625 6235 40670 6355
rect 40790 6235 40835 6355
rect 40955 6235 41000 6355
rect 41120 6235 41175 6355
rect 41295 6235 41340 6355
rect 41460 6235 41505 6355
rect 41625 6235 41670 6355
rect 41790 6235 41845 6355
rect 41965 6235 42175 6355
rect 42295 6235 42340 6355
rect 42460 6235 42505 6355
rect 42625 6235 42670 6355
rect 42790 6235 42845 6355
rect 42965 6235 43010 6355
rect 43130 6235 43175 6355
rect 43295 6235 43340 6355
rect 43460 6235 43515 6355
rect 43635 6235 43680 6355
rect 43800 6235 43845 6355
rect 43965 6235 44010 6355
rect 44130 6235 44185 6355
rect 44305 6235 44350 6355
rect 44470 6235 44515 6355
rect 44635 6235 44680 6355
rect 44800 6235 44855 6355
rect 44975 6235 45020 6355
rect 45140 6235 45185 6355
rect 45305 6235 45350 6355
rect 45470 6235 45525 6355
rect 45645 6235 45690 6355
rect 45810 6235 45855 6355
rect 45975 6235 46020 6355
rect 46140 6235 46195 6355
rect 46315 6235 46360 6355
rect 46480 6235 46525 6355
rect 46645 6235 46690 6355
rect 46810 6235 46865 6355
rect 46985 6235 47030 6355
rect 47150 6235 47195 6355
rect 47315 6235 47360 6355
rect 47480 6235 47535 6355
rect 47655 6235 47865 6355
rect 47985 6235 48030 6355
rect 48150 6235 48195 6355
rect 48315 6235 48360 6355
rect 48480 6235 48535 6355
rect 48655 6235 48700 6355
rect 48820 6235 48865 6355
rect 48985 6235 49030 6355
rect 49150 6235 49205 6355
rect 49325 6235 49370 6355
rect 49490 6235 49535 6355
rect 49655 6235 49700 6355
rect 49820 6235 49875 6355
rect 49995 6235 50040 6355
rect 50160 6235 50205 6355
rect 50325 6235 50370 6355
rect 50490 6235 50545 6355
rect 50665 6235 50710 6355
rect 50830 6235 50875 6355
rect 50995 6235 51040 6355
rect 51160 6235 51215 6355
rect 51335 6235 51380 6355
rect 51500 6235 51545 6355
rect 51665 6235 51710 6355
rect 51830 6235 51885 6355
rect 52005 6235 52050 6355
rect 52170 6235 52215 6355
rect 52335 6235 52380 6355
rect 52500 6235 52555 6355
rect 52675 6235 52720 6355
rect 52840 6235 52885 6355
rect 53005 6235 53050 6355
rect 53170 6235 53225 6355
rect 53345 6235 53370 6355
rect 30770 6190 53370 6235
rect 30770 6070 30795 6190
rect 30915 6070 30960 6190
rect 31080 6070 31125 6190
rect 31245 6070 31290 6190
rect 31410 6070 31465 6190
rect 31585 6070 31630 6190
rect 31750 6070 31795 6190
rect 31915 6070 31960 6190
rect 32080 6070 32135 6190
rect 32255 6070 32300 6190
rect 32420 6070 32465 6190
rect 32585 6070 32630 6190
rect 32750 6070 32805 6190
rect 32925 6070 32970 6190
rect 33090 6070 33135 6190
rect 33255 6070 33300 6190
rect 33420 6070 33475 6190
rect 33595 6070 33640 6190
rect 33760 6070 33805 6190
rect 33925 6070 33970 6190
rect 34090 6070 34145 6190
rect 34265 6070 34310 6190
rect 34430 6070 34475 6190
rect 34595 6070 34640 6190
rect 34760 6070 34815 6190
rect 34935 6070 34980 6190
rect 35100 6070 35145 6190
rect 35265 6070 35310 6190
rect 35430 6070 35485 6190
rect 35605 6070 35650 6190
rect 35770 6070 35815 6190
rect 35935 6070 35980 6190
rect 36100 6070 36155 6190
rect 36275 6070 36485 6190
rect 36605 6070 36650 6190
rect 36770 6070 36815 6190
rect 36935 6070 36980 6190
rect 37100 6070 37155 6190
rect 37275 6070 37320 6190
rect 37440 6070 37485 6190
rect 37605 6070 37650 6190
rect 37770 6070 37825 6190
rect 37945 6070 37990 6190
rect 38110 6070 38155 6190
rect 38275 6070 38320 6190
rect 38440 6070 38495 6190
rect 38615 6070 38660 6190
rect 38780 6070 38825 6190
rect 38945 6070 38990 6190
rect 39110 6070 39165 6190
rect 39285 6070 39330 6190
rect 39450 6070 39495 6190
rect 39615 6070 39660 6190
rect 39780 6070 39835 6190
rect 39955 6070 40000 6190
rect 40120 6070 40165 6190
rect 40285 6070 40330 6190
rect 40450 6070 40505 6190
rect 40625 6070 40670 6190
rect 40790 6070 40835 6190
rect 40955 6070 41000 6190
rect 41120 6070 41175 6190
rect 41295 6070 41340 6190
rect 41460 6070 41505 6190
rect 41625 6070 41670 6190
rect 41790 6070 41845 6190
rect 41965 6070 42175 6190
rect 42295 6070 42340 6190
rect 42460 6070 42505 6190
rect 42625 6070 42670 6190
rect 42790 6070 42845 6190
rect 42965 6070 43010 6190
rect 43130 6070 43175 6190
rect 43295 6070 43340 6190
rect 43460 6070 43515 6190
rect 43635 6070 43680 6190
rect 43800 6070 43845 6190
rect 43965 6070 44010 6190
rect 44130 6070 44185 6190
rect 44305 6070 44350 6190
rect 44470 6070 44515 6190
rect 44635 6070 44680 6190
rect 44800 6070 44855 6190
rect 44975 6070 45020 6190
rect 45140 6070 45185 6190
rect 45305 6070 45350 6190
rect 45470 6070 45525 6190
rect 45645 6070 45690 6190
rect 45810 6070 45855 6190
rect 45975 6070 46020 6190
rect 46140 6070 46195 6190
rect 46315 6070 46360 6190
rect 46480 6070 46525 6190
rect 46645 6070 46690 6190
rect 46810 6070 46865 6190
rect 46985 6070 47030 6190
rect 47150 6070 47195 6190
rect 47315 6070 47360 6190
rect 47480 6070 47535 6190
rect 47655 6070 47865 6190
rect 47985 6070 48030 6190
rect 48150 6070 48195 6190
rect 48315 6070 48360 6190
rect 48480 6070 48535 6190
rect 48655 6070 48700 6190
rect 48820 6070 48865 6190
rect 48985 6070 49030 6190
rect 49150 6070 49205 6190
rect 49325 6070 49370 6190
rect 49490 6070 49535 6190
rect 49655 6070 49700 6190
rect 49820 6070 49875 6190
rect 49995 6070 50040 6190
rect 50160 6070 50205 6190
rect 50325 6070 50370 6190
rect 50490 6070 50545 6190
rect 50665 6070 50710 6190
rect 50830 6070 50875 6190
rect 50995 6070 51040 6190
rect 51160 6070 51215 6190
rect 51335 6070 51380 6190
rect 51500 6070 51545 6190
rect 51665 6070 51710 6190
rect 51830 6070 51885 6190
rect 52005 6070 52050 6190
rect 52170 6070 52215 6190
rect 52335 6070 52380 6190
rect 52500 6070 52555 6190
rect 52675 6070 52720 6190
rect 52840 6070 52885 6190
rect 53005 6070 53050 6190
rect 53170 6070 53225 6190
rect 53345 6070 53370 6190
rect 30770 6025 53370 6070
rect 30770 5905 30795 6025
rect 30915 5905 30960 6025
rect 31080 5905 31125 6025
rect 31245 5905 31290 6025
rect 31410 5905 31465 6025
rect 31585 5905 31630 6025
rect 31750 5905 31795 6025
rect 31915 5905 31960 6025
rect 32080 5905 32135 6025
rect 32255 5905 32300 6025
rect 32420 5905 32465 6025
rect 32585 5905 32630 6025
rect 32750 5905 32805 6025
rect 32925 5905 32970 6025
rect 33090 5905 33135 6025
rect 33255 5905 33300 6025
rect 33420 5905 33475 6025
rect 33595 5905 33640 6025
rect 33760 5905 33805 6025
rect 33925 5905 33970 6025
rect 34090 5905 34145 6025
rect 34265 5905 34310 6025
rect 34430 5905 34475 6025
rect 34595 5905 34640 6025
rect 34760 5905 34815 6025
rect 34935 5905 34980 6025
rect 35100 5905 35145 6025
rect 35265 5905 35310 6025
rect 35430 5905 35485 6025
rect 35605 5905 35650 6025
rect 35770 5905 35815 6025
rect 35935 5905 35980 6025
rect 36100 5905 36155 6025
rect 36275 5905 36485 6025
rect 36605 5905 36650 6025
rect 36770 5905 36815 6025
rect 36935 5905 36980 6025
rect 37100 5905 37155 6025
rect 37275 5905 37320 6025
rect 37440 5905 37485 6025
rect 37605 5905 37650 6025
rect 37770 5905 37825 6025
rect 37945 5905 37990 6025
rect 38110 5905 38155 6025
rect 38275 5905 38320 6025
rect 38440 5905 38495 6025
rect 38615 5905 38660 6025
rect 38780 5905 38825 6025
rect 38945 5905 38990 6025
rect 39110 5905 39165 6025
rect 39285 5905 39330 6025
rect 39450 5905 39495 6025
rect 39615 5905 39660 6025
rect 39780 5905 39835 6025
rect 39955 5905 40000 6025
rect 40120 5905 40165 6025
rect 40285 5905 40330 6025
rect 40450 5905 40505 6025
rect 40625 5905 40670 6025
rect 40790 5905 40835 6025
rect 40955 5905 41000 6025
rect 41120 5905 41175 6025
rect 41295 5905 41340 6025
rect 41460 5905 41505 6025
rect 41625 5905 41670 6025
rect 41790 5905 41845 6025
rect 41965 5905 42175 6025
rect 42295 5905 42340 6025
rect 42460 5905 42505 6025
rect 42625 5905 42670 6025
rect 42790 5905 42845 6025
rect 42965 5905 43010 6025
rect 43130 5905 43175 6025
rect 43295 5905 43340 6025
rect 43460 5905 43515 6025
rect 43635 5905 43680 6025
rect 43800 5905 43845 6025
rect 43965 5905 44010 6025
rect 44130 5905 44185 6025
rect 44305 5905 44350 6025
rect 44470 5905 44515 6025
rect 44635 5905 44680 6025
rect 44800 5905 44855 6025
rect 44975 5905 45020 6025
rect 45140 5905 45185 6025
rect 45305 5905 45350 6025
rect 45470 5905 45525 6025
rect 45645 5905 45690 6025
rect 45810 5905 45855 6025
rect 45975 5905 46020 6025
rect 46140 5905 46195 6025
rect 46315 5905 46360 6025
rect 46480 5905 46525 6025
rect 46645 5905 46690 6025
rect 46810 5905 46865 6025
rect 46985 5905 47030 6025
rect 47150 5905 47195 6025
rect 47315 5905 47360 6025
rect 47480 5905 47535 6025
rect 47655 5905 47865 6025
rect 47985 5905 48030 6025
rect 48150 5905 48195 6025
rect 48315 5905 48360 6025
rect 48480 5905 48535 6025
rect 48655 5905 48700 6025
rect 48820 5905 48865 6025
rect 48985 5905 49030 6025
rect 49150 5905 49205 6025
rect 49325 5905 49370 6025
rect 49490 5905 49535 6025
rect 49655 5905 49700 6025
rect 49820 5905 49875 6025
rect 49995 5905 50040 6025
rect 50160 5905 50205 6025
rect 50325 5905 50370 6025
rect 50490 5905 50545 6025
rect 50665 5905 50710 6025
rect 50830 5905 50875 6025
rect 50995 5905 51040 6025
rect 51160 5905 51215 6025
rect 51335 5905 51380 6025
rect 51500 5905 51545 6025
rect 51665 5905 51710 6025
rect 51830 5905 51885 6025
rect 52005 5905 52050 6025
rect 52170 5905 52215 6025
rect 52335 5905 52380 6025
rect 52500 5905 52555 6025
rect 52675 5905 52720 6025
rect 52840 5905 52885 6025
rect 53005 5905 53050 6025
rect 53170 5905 53225 6025
rect 53345 5905 53370 6025
rect 30770 5860 53370 5905
rect 30770 5740 30795 5860
rect 30915 5740 30960 5860
rect 31080 5740 31125 5860
rect 31245 5740 31290 5860
rect 31410 5740 31465 5860
rect 31585 5740 31630 5860
rect 31750 5740 31795 5860
rect 31915 5740 31960 5860
rect 32080 5740 32135 5860
rect 32255 5740 32300 5860
rect 32420 5740 32465 5860
rect 32585 5740 32630 5860
rect 32750 5740 32805 5860
rect 32925 5740 32970 5860
rect 33090 5740 33135 5860
rect 33255 5740 33300 5860
rect 33420 5740 33475 5860
rect 33595 5740 33640 5860
rect 33760 5740 33805 5860
rect 33925 5740 33970 5860
rect 34090 5740 34145 5860
rect 34265 5740 34310 5860
rect 34430 5740 34475 5860
rect 34595 5740 34640 5860
rect 34760 5740 34815 5860
rect 34935 5740 34980 5860
rect 35100 5740 35145 5860
rect 35265 5740 35310 5860
rect 35430 5740 35485 5860
rect 35605 5740 35650 5860
rect 35770 5740 35815 5860
rect 35935 5740 35980 5860
rect 36100 5740 36155 5860
rect 36275 5740 36485 5860
rect 36605 5740 36650 5860
rect 36770 5740 36815 5860
rect 36935 5740 36980 5860
rect 37100 5740 37155 5860
rect 37275 5740 37320 5860
rect 37440 5740 37485 5860
rect 37605 5740 37650 5860
rect 37770 5740 37825 5860
rect 37945 5740 37990 5860
rect 38110 5740 38155 5860
rect 38275 5740 38320 5860
rect 38440 5740 38495 5860
rect 38615 5740 38660 5860
rect 38780 5740 38825 5860
rect 38945 5740 38990 5860
rect 39110 5740 39165 5860
rect 39285 5740 39330 5860
rect 39450 5740 39495 5860
rect 39615 5740 39660 5860
rect 39780 5740 39835 5860
rect 39955 5740 40000 5860
rect 40120 5740 40165 5860
rect 40285 5740 40330 5860
rect 40450 5740 40505 5860
rect 40625 5740 40670 5860
rect 40790 5740 40835 5860
rect 40955 5740 41000 5860
rect 41120 5740 41175 5860
rect 41295 5740 41340 5860
rect 41460 5740 41505 5860
rect 41625 5740 41670 5860
rect 41790 5740 41845 5860
rect 41965 5740 42175 5860
rect 42295 5740 42340 5860
rect 42460 5740 42505 5860
rect 42625 5740 42670 5860
rect 42790 5740 42845 5860
rect 42965 5740 43010 5860
rect 43130 5740 43175 5860
rect 43295 5740 43340 5860
rect 43460 5740 43515 5860
rect 43635 5740 43680 5860
rect 43800 5740 43845 5860
rect 43965 5740 44010 5860
rect 44130 5740 44185 5860
rect 44305 5740 44350 5860
rect 44470 5740 44515 5860
rect 44635 5740 44680 5860
rect 44800 5740 44855 5860
rect 44975 5740 45020 5860
rect 45140 5740 45185 5860
rect 45305 5740 45350 5860
rect 45470 5740 45525 5860
rect 45645 5740 45690 5860
rect 45810 5740 45855 5860
rect 45975 5740 46020 5860
rect 46140 5740 46195 5860
rect 46315 5740 46360 5860
rect 46480 5740 46525 5860
rect 46645 5740 46690 5860
rect 46810 5740 46865 5860
rect 46985 5740 47030 5860
rect 47150 5740 47195 5860
rect 47315 5740 47360 5860
rect 47480 5740 47535 5860
rect 47655 5740 47865 5860
rect 47985 5740 48030 5860
rect 48150 5740 48195 5860
rect 48315 5740 48360 5860
rect 48480 5740 48535 5860
rect 48655 5740 48700 5860
rect 48820 5740 48865 5860
rect 48985 5740 49030 5860
rect 49150 5740 49205 5860
rect 49325 5740 49370 5860
rect 49490 5740 49535 5860
rect 49655 5740 49700 5860
rect 49820 5740 49875 5860
rect 49995 5740 50040 5860
rect 50160 5740 50205 5860
rect 50325 5740 50370 5860
rect 50490 5740 50545 5860
rect 50665 5740 50710 5860
rect 50830 5740 50875 5860
rect 50995 5740 51040 5860
rect 51160 5740 51215 5860
rect 51335 5740 51380 5860
rect 51500 5740 51545 5860
rect 51665 5740 51710 5860
rect 51830 5740 51885 5860
rect 52005 5740 52050 5860
rect 52170 5740 52215 5860
rect 52335 5740 52380 5860
rect 52500 5740 52555 5860
rect 52675 5740 52720 5860
rect 52840 5740 52885 5860
rect 53005 5740 53050 5860
rect 53170 5740 53225 5860
rect 53345 5740 53370 5860
rect 30770 5685 53370 5740
rect 30770 5565 30795 5685
rect 30915 5565 30960 5685
rect 31080 5565 31125 5685
rect 31245 5565 31290 5685
rect 31410 5565 31465 5685
rect 31585 5565 31630 5685
rect 31750 5565 31795 5685
rect 31915 5565 31960 5685
rect 32080 5565 32135 5685
rect 32255 5565 32300 5685
rect 32420 5565 32465 5685
rect 32585 5565 32630 5685
rect 32750 5565 32805 5685
rect 32925 5565 32970 5685
rect 33090 5565 33135 5685
rect 33255 5565 33300 5685
rect 33420 5565 33475 5685
rect 33595 5565 33640 5685
rect 33760 5565 33805 5685
rect 33925 5565 33970 5685
rect 34090 5565 34145 5685
rect 34265 5565 34310 5685
rect 34430 5565 34475 5685
rect 34595 5565 34640 5685
rect 34760 5565 34815 5685
rect 34935 5565 34980 5685
rect 35100 5565 35145 5685
rect 35265 5565 35310 5685
rect 35430 5565 35485 5685
rect 35605 5565 35650 5685
rect 35770 5565 35815 5685
rect 35935 5565 35980 5685
rect 36100 5565 36155 5685
rect 36275 5565 36485 5685
rect 36605 5565 36650 5685
rect 36770 5565 36815 5685
rect 36935 5565 36980 5685
rect 37100 5565 37155 5685
rect 37275 5565 37320 5685
rect 37440 5565 37485 5685
rect 37605 5565 37650 5685
rect 37770 5565 37825 5685
rect 37945 5565 37990 5685
rect 38110 5565 38155 5685
rect 38275 5565 38320 5685
rect 38440 5565 38495 5685
rect 38615 5565 38660 5685
rect 38780 5565 38825 5685
rect 38945 5565 38990 5685
rect 39110 5565 39165 5685
rect 39285 5565 39330 5685
rect 39450 5565 39495 5685
rect 39615 5565 39660 5685
rect 39780 5565 39835 5685
rect 39955 5565 40000 5685
rect 40120 5565 40165 5685
rect 40285 5565 40330 5685
rect 40450 5565 40505 5685
rect 40625 5565 40670 5685
rect 40790 5565 40835 5685
rect 40955 5565 41000 5685
rect 41120 5565 41175 5685
rect 41295 5565 41340 5685
rect 41460 5565 41505 5685
rect 41625 5565 41670 5685
rect 41790 5565 41845 5685
rect 41965 5565 42175 5685
rect 42295 5565 42340 5685
rect 42460 5565 42505 5685
rect 42625 5565 42670 5685
rect 42790 5565 42845 5685
rect 42965 5565 43010 5685
rect 43130 5565 43175 5685
rect 43295 5565 43340 5685
rect 43460 5565 43515 5685
rect 43635 5565 43680 5685
rect 43800 5565 43845 5685
rect 43965 5565 44010 5685
rect 44130 5565 44185 5685
rect 44305 5565 44350 5685
rect 44470 5565 44515 5685
rect 44635 5565 44680 5685
rect 44800 5565 44855 5685
rect 44975 5565 45020 5685
rect 45140 5565 45185 5685
rect 45305 5565 45350 5685
rect 45470 5565 45525 5685
rect 45645 5565 45690 5685
rect 45810 5565 45855 5685
rect 45975 5565 46020 5685
rect 46140 5565 46195 5685
rect 46315 5565 46360 5685
rect 46480 5565 46525 5685
rect 46645 5565 46690 5685
rect 46810 5565 46865 5685
rect 46985 5565 47030 5685
rect 47150 5565 47195 5685
rect 47315 5565 47360 5685
rect 47480 5565 47535 5685
rect 47655 5565 47865 5685
rect 47985 5565 48030 5685
rect 48150 5565 48195 5685
rect 48315 5565 48360 5685
rect 48480 5565 48535 5685
rect 48655 5565 48700 5685
rect 48820 5565 48865 5685
rect 48985 5565 49030 5685
rect 49150 5565 49205 5685
rect 49325 5565 49370 5685
rect 49490 5565 49535 5685
rect 49655 5565 49700 5685
rect 49820 5565 49875 5685
rect 49995 5565 50040 5685
rect 50160 5565 50205 5685
rect 50325 5565 50370 5685
rect 50490 5565 50545 5685
rect 50665 5565 50710 5685
rect 50830 5565 50875 5685
rect 50995 5565 51040 5685
rect 51160 5565 51215 5685
rect 51335 5565 51380 5685
rect 51500 5565 51545 5685
rect 51665 5565 51710 5685
rect 51830 5565 51885 5685
rect 52005 5565 52050 5685
rect 52170 5565 52215 5685
rect 52335 5565 52380 5685
rect 52500 5565 52555 5685
rect 52675 5565 52720 5685
rect 52840 5565 52885 5685
rect 53005 5565 53050 5685
rect 53170 5565 53225 5685
rect 53345 5565 53370 5685
rect 30770 5520 53370 5565
rect 30770 5400 30795 5520
rect 30915 5400 30960 5520
rect 31080 5400 31125 5520
rect 31245 5400 31290 5520
rect 31410 5400 31465 5520
rect 31585 5400 31630 5520
rect 31750 5400 31795 5520
rect 31915 5400 31960 5520
rect 32080 5400 32135 5520
rect 32255 5400 32300 5520
rect 32420 5400 32465 5520
rect 32585 5400 32630 5520
rect 32750 5400 32805 5520
rect 32925 5400 32970 5520
rect 33090 5400 33135 5520
rect 33255 5400 33300 5520
rect 33420 5400 33475 5520
rect 33595 5400 33640 5520
rect 33760 5400 33805 5520
rect 33925 5400 33970 5520
rect 34090 5400 34145 5520
rect 34265 5400 34310 5520
rect 34430 5400 34475 5520
rect 34595 5400 34640 5520
rect 34760 5400 34815 5520
rect 34935 5400 34980 5520
rect 35100 5400 35145 5520
rect 35265 5400 35310 5520
rect 35430 5400 35485 5520
rect 35605 5400 35650 5520
rect 35770 5400 35815 5520
rect 35935 5400 35980 5520
rect 36100 5400 36155 5520
rect 36275 5400 36485 5520
rect 36605 5400 36650 5520
rect 36770 5400 36815 5520
rect 36935 5400 36980 5520
rect 37100 5400 37155 5520
rect 37275 5400 37320 5520
rect 37440 5400 37485 5520
rect 37605 5400 37650 5520
rect 37770 5400 37825 5520
rect 37945 5400 37990 5520
rect 38110 5400 38155 5520
rect 38275 5400 38320 5520
rect 38440 5400 38495 5520
rect 38615 5400 38660 5520
rect 38780 5400 38825 5520
rect 38945 5400 38990 5520
rect 39110 5400 39165 5520
rect 39285 5400 39330 5520
rect 39450 5400 39495 5520
rect 39615 5400 39660 5520
rect 39780 5400 39835 5520
rect 39955 5400 40000 5520
rect 40120 5400 40165 5520
rect 40285 5400 40330 5520
rect 40450 5400 40505 5520
rect 40625 5400 40670 5520
rect 40790 5400 40835 5520
rect 40955 5400 41000 5520
rect 41120 5400 41175 5520
rect 41295 5400 41340 5520
rect 41460 5400 41505 5520
rect 41625 5400 41670 5520
rect 41790 5400 41845 5520
rect 41965 5400 42175 5520
rect 42295 5400 42340 5520
rect 42460 5400 42505 5520
rect 42625 5400 42670 5520
rect 42790 5400 42845 5520
rect 42965 5400 43010 5520
rect 43130 5400 43175 5520
rect 43295 5400 43340 5520
rect 43460 5400 43515 5520
rect 43635 5400 43680 5520
rect 43800 5400 43845 5520
rect 43965 5400 44010 5520
rect 44130 5400 44185 5520
rect 44305 5400 44350 5520
rect 44470 5400 44515 5520
rect 44635 5400 44680 5520
rect 44800 5400 44855 5520
rect 44975 5400 45020 5520
rect 45140 5400 45185 5520
rect 45305 5400 45350 5520
rect 45470 5400 45525 5520
rect 45645 5400 45690 5520
rect 45810 5400 45855 5520
rect 45975 5400 46020 5520
rect 46140 5400 46195 5520
rect 46315 5400 46360 5520
rect 46480 5400 46525 5520
rect 46645 5400 46690 5520
rect 46810 5400 46865 5520
rect 46985 5400 47030 5520
rect 47150 5400 47195 5520
rect 47315 5400 47360 5520
rect 47480 5400 47535 5520
rect 47655 5400 47865 5520
rect 47985 5400 48030 5520
rect 48150 5400 48195 5520
rect 48315 5400 48360 5520
rect 48480 5400 48535 5520
rect 48655 5400 48700 5520
rect 48820 5400 48865 5520
rect 48985 5400 49030 5520
rect 49150 5400 49205 5520
rect 49325 5400 49370 5520
rect 49490 5400 49535 5520
rect 49655 5400 49700 5520
rect 49820 5400 49875 5520
rect 49995 5400 50040 5520
rect 50160 5400 50205 5520
rect 50325 5400 50370 5520
rect 50490 5400 50545 5520
rect 50665 5400 50710 5520
rect 50830 5400 50875 5520
rect 50995 5400 51040 5520
rect 51160 5400 51215 5520
rect 51335 5400 51380 5520
rect 51500 5400 51545 5520
rect 51665 5400 51710 5520
rect 51830 5400 51885 5520
rect 52005 5400 52050 5520
rect 52170 5400 52215 5520
rect 52335 5400 52380 5520
rect 52500 5400 52555 5520
rect 52675 5400 52720 5520
rect 52840 5400 52885 5520
rect 53005 5400 53050 5520
rect 53170 5400 53225 5520
rect 53345 5400 53370 5520
rect 30770 5355 53370 5400
rect 30770 5235 30795 5355
rect 30915 5235 30960 5355
rect 31080 5235 31125 5355
rect 31245 5235 31290 5355
rect 31410 5235 31465 5355
rect 31585 5235 31630 5355
rect 31750 5235 31795 5355
rect 31915 5235 31960 5355
rect 32080 5235 32135 5355
rect 32255 5235 32300 5355
rect 32420 5235 32465 5355
rect 32585 5235 32630 5355
rect 32750 5235 32805 5355
rect 32925 5235 32970 5355
rect 33090 5235 33135 5355
rect 33255 5235 33300 5355
rect 33420 5235 33475 5355
rect 33595 5235 33640 5355
rect 33760 5235 33805 5355
rect 33925 5235 33970 5355
rect 34090 5235 34145 5355
rect 34265 5235 34310 5355
rect 34430 5235 34475 5355
rect 34595 5235 34640 5355
rect 34760 5235 34815 5355
rect 34935 5235 34980 5355
rect 35100 5235 35145 5355
rect 35265 5235 35310 5355
rect 35430 5235 35485 5355
rect 35605 5235 35650 5355
rect 35770 5235 35815 5355
rect 35935 5235 35980 5355
rect 36100 5235 36155 5355
rect 36275 5235 36485 5355
rect 36605 5235 36650 5355
rect 36770 5235 36815 5355
rect 36935 5235 36980 5355
rect 37100 5235 37155 5355
rect 37275 5235 37320 5355
rect 37440 5235 37485 5355
rect 37605 5235 37650 5355
rect 37770 5235 37825 5355
rect 37945 5235 37990 5355
rect 38110 5235 38155 5355
rect 38275 5235 38320 5355
rect 38440 5235 38495 5355
rect 38615 5235 38660 5355
rect 38780 5235 38825 5355
rect 38945 5235 38990 5355
rect 39110 5235 39165 5355
rect 39285 5235 39330 5355
rect 39450 5235 39495 5355
rect 39615 5235 39660 5355
rect 39780 5235 39835 5355
rect 39955 5235 40000 5355
rect 40120 5235 40165 5355
rect 40285 5235 40330 5355
rect 40450 5235 40505 5355
rect 40625 5235 40670 5355
rect 40790 5235 40835 5355
rect 40955 5235 41000 5355
rect 41120 5235 41175 5355
rect 41295 5235 41340 5355
rect 41460 5235 41505 5355
rect 41625 5235 41670 5355
rect 41790 5235 41845 5355
rect 41965 5235 42175 5355
rect 42295 5235 42340 5355
rect 42460 5235 42505 5355
rect 42625 5235 42670 5355
rect 42790 5235 42845 5355
rect 42965 5235 43010 5355
rect 43130 5235 43175 5355
rect 43295 5235 43340 5355
rect 43460 5235 43515 5355
rect 43635 5235 43680 5355
rect 43800 5235 43845 5355
rect 43965 5235 44010 5355
rect 44130 5235 44185 5355
rect 44305 5235 44350 5355
rect 44470 5235 44515 5355
rect 44635 5235 44680 5355
rect 44800 5235 44855 5355
rect 44975 5235 45020 5355
rect 45140 5235 45185 5355
rect 45305 5235 45350 5355
rect 45470 5235 45525 5355
rect 45645 5235 45690 5355
rect 45810 5235 45855 5355
rect 45975 5235 46020 5355
rect 46140 5235 46195 5355
rect 46315 5235 46360 5355
rect 46480 5235 46525 5355
rect 46645 5235 46690 5355
rect 46810 5235 46865 5355
rect 46985 5235 47030 5355
rect 47150 5235 47195 5355
rect 47315 5235 47360 5355
rect 47480 5235 47535 5355
rect 47655 5235 47865 5355
rect 47985 5235 48030 5355
rect 48150 5235 48195 5355
rect 48315 5235 48360 5355
rect 48480 5235 48535 5355
rect 48655 5235 48700 5355
rect 48820 5235 48865 5355
rect 48985 5235 49030 5355
rect 49150 5235 49205 5355
rect 49325 5235 49370 5355
rect 49490 5235 49535 5355
rect 49655 5235 49700 5355
rect 49820 5235 49875 5355
rect 49995 5235 50040 5355
rect 50160 5235 50205 5355
rect 50325 5235 50370 5355
rect 50490 5235 50545 5355
rect 50665 5235 50710 5355
rect 50830 5235 50875 5355
rect 50995 5235 51040 5355
rect 51160 5235 51215 5355
rect 51335 5235 51380 5355
rect 51500 5235 51545 5355
rect 51665 5235 51710 5355
rect 51830 5235 51885 5355
rect 52005 5235 52050 5355
rect 52170 5235 52215 5355
rect 52335 5235 52380 5355
rect 52500 5235 52555 5355
rect 52675 5235 52720 5355
rect 52840 5235 52885 5355
rect 53005 5235 53050 5355
rect 53170 5235 53225 5355
rect 53345 5235 53370 5355
rect 30770 5190 53370 5235
rect 30770 5070 30795 5190
rect 30915 5070 30960 5190
rect 31080 5070 31125 5190
rect 31245 5070 31290 5190
rect 31410 5070 31465 5190
rect 31585 5070 31630 5190
rect 31750 5070 31795 5190
rect 31915 5070 31960 5190
rect 32080 5070 32135 5190
rect 32255 5070 32300 5190
rect 32420 5070 32465 5190
rect 32585 5070 32630 5190
rect 32750 5070 32805 5190
rect 32925 5070 32970 5190
rect 33090 5070 33135 5190
rect 33255 5070 33300 5190
rect 33420 5070 33475 5190
rect 33595 5070 33640 5190
rect 33760 5070 33805 5190
rect 33925 5070 33970 5190
rect 34090 5070 34145 5190
rect 34265 5070 34310 5190
rect 34430 5070 34475 5190
rect 34595 5070 34640 5190
rect 34760 5070 34815 5190
rect 34935 5070 34980 5190
rect 35100 5070 35145 5190
rect 35265 5070 35310 5190
rect 35430 5070 35485 5190
rect 35605 5070 35650 5190
rect 35770 5070 35815 5190
rect 35935 5070 35980 5190
rect 36100 5070 36155 5190
rect 36275 5070 36485 5190
rect 36605 5070 36650 5190
rect 36770 5070 36815 5190
rect 36935 5070 36980 5190
rect 37100 5070 37155 5190
rect 37275 5070 37320 5190
rect 37440 5070 37485 5190
rect 37605 5070 37650 5190
rect 37770 5070 37825 5190
rect 37945 5070 37990 5190
rect 38110 5070 38155 5190
rect 38275 5070 38320 5190
rect 38440 5070 38495 5190
rect 38615 5070 38660 5190
rect 38780 5070 38825 5190
rect 38945 5070 38990 5190
rect 39110 5070 39165 5190
rect 39285 5070 39330 5190
rect 39450 5070 39495 5190
rect 39615 5070 39660 5190
rect 39780 5070 39835 5190
rect 39955 5070 40000 5190
rect 40120 5070 40165 5190
rect 40285 5070 40330 5190
rect 40450 5070 40505 5190
rect 40625 5070 40670 5190
rect 40790 5070 40835 5190
rect 40955 5070 41000 5190
rect 41120 5070 41175 5190
rect 41295 5070 41340 5190
rect 41460 5070 41505 5190
rect 41625 5070 41670 5190
rect 41790 5070 41845 5190
rect 41965 5070 42175 5190
rect 42295 5070 42340 5190
rect 42460 5070 42505 5190
rect 42625 5070 42670 5190
rect 42790 5070 42845 5190
rect 42965 5070 43010 5190
rect 43130 5070 43175 5190
rect 43295 5070 43340 5190
rect 43460 5070 43515 5190
rect 43635 5070 43680 5190
rect 43800 5070 43845 5190
rect 43965 5070 44010 5190
rect 44130 5070 44185 5190
rect 44305 5070 44350 5190
rect 44470 5070 44515 5190
rect 44635 5070 44680 5190
rect 44800 5070 44855 5190
rect 44975 5070 45020 5190
rect 45140 5070 45185 5190
rect 45305 5070 45350 5190
rect 45470 5070 45525 5190
rect 45645 5070 45690 5190
rect 45810 5070 45855 5190
rect 45975 5070 46020 5190
rect 46140 5070 46195 5190
rect 46315 5070 46360 5190
rect 46480 5070 46525 5190
rect 46645 5070 46690 5190
rect 46810 5070 46865 5190
rect 46985 5070 47030 5190
rect 47150 5070 47195 5190
rect 47315 5070 47360 5190
rect 47480 5070 47535 5190
rect 47655 5070 47865 5190
rect 47985 5070 48030 5190
rect 48150 5070 48195 5190
rect 48315 5070 48360 5190
rect 48480 5070 48535 5190
rect 48655 5070 48700 5190
rect 48820 5070 48865 5190
rect 48985 5070 49030 5190
rect 49150 5070 49205 5190
rect 49325 5070 49370 5190
rect 49490 5070 49535 5190
rect 49655 5070 49700 5190
rect 49820 5070 49875 5190
rect 49995 5070 50040 5190
rect 50160 5070 50205 5190
rect 50325 5070 50370 5190
rect 50490 5070 50545 5190
rect 50665 5070 50710 5190
rect 50830 5070 50875 5190
rect 50995 5070 51040 5190
rect 51160 5070 51215 5190
rect 51335 5070 51380 5190
rect 51500 5070 51545 5190
rect 51665 5070 51710 5190
rect 51830 5070 51885 5190
rect 52005 5070 52050 5190
rect 52170 5070 52215 5190
rect 52335 5070 52380 5190
rect 52500 5070 52555 5190
rect 52675 5070 52720 5190
rect 52840 5070 52885 5190
rect 53005 5070 53050 5190
rect 53170 5070 53225 5190
rect 53345 5070 53370 5190
rect 30770 5015 53370 5070
rect 30770 4895 30795 5015
rect 30915 4895 30960 5015
rect 31080 4895 31125 5015
rect 31245 4895 31290 5015
rect 31410 4895 31465 5015
rect 31585 4895 31630 5015
rect 31750 4895 31795 5015
rect 31915 4895 31960 5015
rect 32080 4895 32135 5015
rect 32255 4895 32300 5015
rect 32420 4895 32465 5015
rect 32585 4895 32630 5015
rect 32750 4895 32805 5015
rect 32925 4895 32970 5015
rect 33090 4895 33135 5015
rect 33255 4895 33300 5015
rect 33420 4895 33475 5015
rect 33595 4895 33640 5015
rect 33760 4895 33805 5015
rect 33925 4895 33970 5015
rect 34090 4895 34145 5015
rect 34265 4895 34310 5015
rect 34430 4895 34475 5015
rect 34595 4895 34640 5015
rect 34760 4895 34815 5015
rect 34935 4895 34980 5015
rect 35100 4895 35145 5015
rect 35265 4895 35310 5015
rect 35430 4895 35485 5015
rect 35605 4895 35650 5015
rect 35770 4895 35815 5015
rect 35935 4895 35980 5015
rect 36100 4895 36155 5015
rect 36275 4895 36485 5015
rect 36605 4895 36650 5015
rect 36770 4895 36815 5015
rect 36935 4895 36980 5015
rect 37100 4895 37155 5015
rect 37275 4895 37320 5015
rect 37440 4895 37485 5015
rect 37605 4895 37650 5015
rect 37770 4895 37825 5015
rect 37945 4895 37990 5015
rect 38110 4895 38155 5015
rect 38275 4895 38320 5015
rect 38440 4895 38495 5015
rect 38615 4895 38660 5015
rect 38780 4895 38825 5015
rect 38945 4895 38990 5015
rect 39110 4895 39165 5015
rect 39285 4895 39330 5015
rect 39450 4895 39495 5015
rect 39615 4895 39660 5015
rect 39780 4895 39835 5015
rect 39955 4895 40000 5015
rect 40120 4895 40165 5015
rect 40285 4895 40330 5015
rect 40450 4895 40505 5015
rect 40625 4895 40670 5015
rect 40790 4895 40835 5015
rect 40955 4895 41000 5015
rect 41120 4895 41175 5015
rect 41295 4895 41340 5015
rect 41460 4895 41505 5015
rect 41625 4895 41670 5015
rect 41790 4895 41845 5015
rect 41965 4895 42175 5015
rect 42295 4895 42340 5015
rect 42460 4895 42505 5015
rect 42625 4895 42670 5015
rect 42790 4895 42845 5015
rect 42965 4895 43010 5015
rect 43130 4895 43175 5015
rect 43295 4895 43340 5015
rect 43460 4895 43515 5015
rect 43635 4895 43680 5015
rect 43800 4895 43845 5015
rect 43965 4895 44010 5015
rect 44130 4895 44185 5015
rect 44305 4895 44350 5015
rect 44470 4895 44515 5015
rect 44635 4895 44680 5015
rect 44800 4895 44855 5015
rect 44975 4895 45020 5015
rect 45140 4895 45185 5015
rect 45305 4895 45350 5015
rect 45470 4895 45525 5015
rect 45645 4895 45690 5015
rect 45810 4895 45855 5015
rect 45975 4895 46020 5015
rect 46140 4895 46195 5015
rect 46315 4895 46360 5015
rect 46480 4895 46525 5015
rect 46645 4895 46690 5015
rect 46810 4895 46865 5015
rect 46985 4895 47030 5015
rect 47150 4895 47195 5015
rect 47315 4895 47360 5015
rect 47480 4895 47535 5015
rect 47655 4895 47865 5015
rect 47985 4895 48030 5015
rect 48150 4895 48195 5015
rect 48315 4895 48360 5015
rect 48480 4895 48535 5015
rect 48655 4895 48700 5015
rect 48820 4895 48865 5015
rect 48985 4895 49030 5015
rect 49150 4895 49205 5015
rect 49325 4895 49370 5015
rect 49490 4895 49535 5015
rect 49655 4895 49700 5015
rect 49820 4895 49875 5015
rect 49995 4895 50040 5015
rect 50160 4895 50205 5015
rect 50325 4895 50370 5015
rect 50490 4895 50545 5015
rect 50665 4895 50710 5015
rect 50830 4895 50875 5015
rect 50995 4895 51040 5015
rect 51160 4895 51215 5015
rect 51335 4895 51380 5015
rect 51500 4895 51545 5015
rect 51665 4895 51710 5015
rect 51830 4895 51885 5015
rect 52005 4895 52050 5015
rect 52170 4895 52215 5015
rect 52335 4895 52380 5015
rect 52500 4895 52555 5015
rect 52675 4895 52720 5015
rect 52840 4895 52885 5015
rect 53005 4895 53050 5015
rect 53170 4895 53225 5015
rect 53345 4895 53370 5015
rect 30770 4850 53370 4895
rect 30770 4730 30795 4850
rect 30915 4730 30960 4850
rect 31080 4730 31125 4850
rect 31245 4730 31290 4850
rect 31410 4730 31465 4850
rect 31585 4730 31630 4850
rect 31750 4730 31795 4850
rect 31915 4730 31960 4850
rect 32080 4730 32135 4850
rect 32255 4730 32300 4850
rect 32420 4730 32465 4850
rect 32585 4730 32630 4850
rect 32750 4730 32805 4850
rect 32925 4730 32970 4850
rect 33090 4730 33135 4850
rect 33255 4730 33300 4850
rect 33420 4730 33475 4850
rect 33595 4730 33640 4850
rect 33760 4730 33805 4850
rect 33925 4730 33970 4850
rect 34090 4730 34145 4850
rect 34265 4730 34310 4850
rect 34430 4730 34475 4850
rect 34595 4730 34640 4850
rect 34760 4730 34815 4850
rect 34935 4730 34980 4850
rect 35100 4730 35145 4850
rect 35265 4730 35310 4850
rect 35430 4730 35485 4850
rect 35605 4730 35650 4850
rect 35770 4730 35815 4850
rect 35935 4730 35980 4850
rect 36100 4730 36155 4850
rect 36275 4730 36485 4850
rect 36605 4730 36650 4850
rect 36770 4730 36815 4850
rect 36935 4730 36980 4850
rect 37100 4730 37155 4850
rect 37275 4730 37320 4850
rect 37440 4730 37485 4850
rect 37605 4730 37650 4850
rect 37770 4730 37825 4850
rect 37945 4730 37990 4850
rect 38110 4730 38155 4850
rect 38275 4730 38320 4850
rect 38440 4730 38495 4850
rect 38615 4730 38660 4850
rect 38780 4730 38825 4850
rect 38945 4730 38990 4850
rect 39110 4730 39165 4850
rect 39285 4730 39330 4850
rect 39450 4730 39495 4850
rect 39615 4730 39660 4850
rect 39780 4730 39835 4850
rect 39955 4730 40000 4850
rect 40120 4730 40165 4850
rect 40285 4730 40330 4850
rect 40450 4730 40505 4850
rect 40625 4730 40670 4850
rect 40790 4730 40835 4850
rect 40955 4730 41000 4850
rect 41120 4730 41175 4850
rect 41295 4730 41340 4850
rect 41460 4730 41505 4850
rect 41625 4730 41670 4850
rect 41790 4730 41845 4850
rect 41965 4730 42175 4850
rect 42295 4730 42340 4850
rect 42460 4730 42505 4850
rect 42625 4730 42670 4850
rect 42790 4730 42845 4850
rect 42965 4730 43010 4850
rect 43130 4730 43175 4850
rect 43295 4730 43340 4850
rect 43460 4730 43515 4850
rect 43635 4730 43680 4850
rect 43800 4730 43845 4850
rect 43965 4730 44010 4850
rect 44130 4730 44185 4850
rect 44305 4730 44350 4850
rect 44470 4730 44515 4850
rect 44635 4730 44680 4850
rect 44800 4730 44855 4850
rect 44975 4730 45020 4850
rect 45140 4730 45185 4850
rect 45305 4730 45350 4850
rect 45470 4730 45525 4850
rect 45645 4730 45690 4850
rect 45810 4730 45855 4850
rect 45975 4730 46020 4850
rect 46140 4730 46195 4850
rect 46315 4730 46360 4850
rect 46480 4730 46525 4850
rect 46645 4730 46690 4850
rect 46810 4730 46865 4850
rect 46985 4730 47030 4850
rect 47150 4730 47195 4850
rect 47315 4730 47360 4850
rect 47480 4730 47535 4850
rect 47655 4730 47865 4850
rect 47985 4730 48030 4850
rect 48150 4730 48195 4850
rect 48315 4730 48360 4850
rect 48480 4730 48535 4850
rect 48655 4730 48700 4850
rect 48820 4730 48865 4850
rect 48985 4730 49030 4850
rect 49150 4730 49205 4850
rect 49325 4730 49370 4850
rect 49490 4730 49535 4850
rect 49655 4730 49700 4850
rect 49820 4730 49875 4850
rect 49995 4730 50040 4850
rect 50160 4730 50205 4850
rect 50325 4730 50370 4850
rect 50490 4730 50545 4850
rect 50665 4730 50710 4850
rect 50830 4730 50875 4850
rect 50995 4730 51040 4850
rect 51160 4730 51215 4850
rect 51335 4730 51380 4850
rect 51500 4730 51545 4850
rect 51665 4730 51710 4850
rect 51830 4730 51885 4850
rect 52005 4730 52050 4850
rect 52170 4730 52215 4850
rect 52335 4730 52380 4850
rect 52500 4730 52555 4850
rect 52675 4730 52720 4850
rect 52840 4730 52885 4850
rect 53005 4730 53050 4850
rect 53170 4730 53225 4850
rect 53345 4730 53370 4850
rect 30770 4685 53370 4730
rect 30770 4565 30795 4685
rect 30915 4565 30960 4685
rect 31080 4565 31125 4685
rect 31245 4565 31290 4685
rect 31410 4565 31465 4685
rect 31585 4565 31630 4685
rect 31750 4565 31795 4685
rect 31915 4565 31960 4685
rect 32080 4565 32135 4685
rect 32255 4565 32300 4685
rect 32420 4565 32465 4685
rect 32585 4565 32630 4685
rect 32750 4565 32805 4685
rect 32925 4565 32970 4685
rect 33090 4565 33135 4685
rect 33255 4565 33300 4685
rect 33420 4565 33475 4685
rect 33595 4565 33640 4685
rect 33760 4565 33805 4685
rect 33925 4565 33970 4685
rect 34090 4565 34145 4685
rect 34265 4565 34310 4685
rect 34430 4565 34475 4685
rect 34595 4565 34640 4685
rect 34760 4565 34815 4685
rect 34935 4565 34980 4685
rect 35100 4565 35145 4685
rect 35265 4565 35310 4685
rect 35430 4565 35485 4685
rect 35605 4565 35650 4685
rect 35770 4565 35815 4685
rect 35935 4565 35980 4685
rect 36100 4565 36155 4685
rect 36275 4565 36485 4685
rect 36605 4565 36650 4685
rect 36770 4565 36815 4685
rect 36935 4565 36980 4685
rect 37100 4565 37155 4685
rect 37275 4565 37320 4685
rect 37440 4565 37485 4685
rect 37605 4565 37650 4685
rect 37770 4565 37825 4685
rect 37945 4565 37990 4685
rect 38110 4565 38155 4685
rect 38275 4565 38320 4685
rect 38440 4565 38495 4685
rect 38615 4565 38660 4685
rect 38780 4565 38825 4685
rect 38945 4565 38990 4685
rect 39110 4565 39165 4685
rect 39285 4565 39330 4685
rect 39450 4565 39495 4685
rect 39615 4565 39660 4685
rect 39780 4565 39835 4685
rect 39955 4565 40000 4685
rect 40120 4565 40165 4685
rect 40285 4565 40330 4685
rect 40450 4565 40505 4685
rect 40625 4565 40670 4685
rect 40790 4565 40835 4685
rect 40955 4565 41000 4685
rect 41120 4565 41175 4685
rect 41295 4565 41340 4685
rect 41460 4565 41505 4685
rect 41625 4565 41670 4685
rect 41790 4565 41845 4685
rect 41965 4565 42175 4685
rect 42295 4565 42340 4685
rect 42460 4565 42505 4685
rect 42625 4565 42670 4685
rect 42790 4565 42845 4685
rect 42965 4565 43010 4685
rect 43130 4565 43175 4685
rect 43295 4565 43340 4685
rect 43460 4565 43515 4685
rect 43635 4565 43680 4685
rect 43800 4565 43845 4685
rect 43965 4565 44010 4685
rect 44130 4565 44185 4685
rect 44305 4565 44350 4685
rect 44470 4565 44515 4685
rect 44635 4565 44680 4685
rect 44800 4565 44855 4685
rect 44975 4565 45020 4685
rect 45140 4565 45185 4685
rect 45305 4565 45350 4685
rect 45470 4565 45525 4685
rect 45645 4565 45690 4685
rect 45810 4565 45855 4685
rect 45975 4565 46020 4685
rect 46140 4565 46195 4685
rect 46315 4565 46360 4685
rect 46480 4565 46525 4685
rect 46645 4565 46690 4685
rect 46810 4565 46865 4685
rect 46985 4565 47030 4685
rect 47150 4565 47195 4685
rect 47315 4565 47360 4685
rect 47480 4565 47535 4685
rect 47655 4565 47865 4685
rect 47985 4565 48030 4685
rect 48150 4565 48195 4685
rect 48315 4565 48360 4685
rect 48480 4565 48535 4685
rect 48655 4565 48700 4685
rect 48820 4565 48865 4685
rect 48985 4565 49030 4685
rect 49150 4565 49205 4685
rect 49325 4565 49370 4685
rect 49490 4565 49535 4685
rect 49655 4565 49700 4685
rect 49820 4565 49875 4685
rect 49995 4565 50040 4685
rect 50160 4565 50205 4685
rect 50325 4565 50370 4685
rect 50490 4565 50545 4685
rect 50665 4565 50710 4685
rect 50830 4565 50875 4685
rect 50995 4565 51040 4685
rect 51160 4565 51215 4685
rect 51335 4565 51380 4685
rect 51500 4565 51545 4685
rect 51665 4565 51710 4685
rect 51830 4565 51885 4685
rect 52005 4565 52050 4685
rect 52170 4565 52215 4685
rect 52335 4565 52380 4685
rect 52500 4565 52555 4685
rect 52675 4565 52720 4685
rect 52840 4565 52885 4685
rect 53005 4565 53050 4685
rect 53170 4565 53225 4685
rect 53345 4565 53370 4685
rect 30770 4520 53370 4565
rect 30770 4400 30795 4520
rect 30915 4400 30960 4520
rect 31080 4400 31125 4520
rect 31245 4400 31290 4520
rect 31410 4400 31465 4520
rect 31585 4400 31630 4520
rect 31750 4400 31795 4520
rect 31915 4400 31960 4520
rect 32080 4400 32135 4520
rect 32255 4400 32300 4520
rect 32420 4400 32465 4520
rect 32585 4400 32630 4520
rect 32750 4400 32805 4520
rect 32925 4400 32970 4520
rect 33090 4400 33135 4520
rect 33255 4400 33300 4520
rect 33420 4400 33475 4520
rect 33595 4400 33640 4520
rect 33760 4400 33805 4520
rect 33925 4400 33970 4520
rect 34090 4400 34145 4520
rect 34265 4400 34310 4520
rect 34430 4400 34475 4520
rect 34595 4400 34640 4520
rect 34760 4400 34815 4520
rect 34935 4400 34980 4520
rect 35100 4400 35145 4520
rect 35265 4400 35310 4520
rect 35430 4400 35485 4520
rect 35605 4400 35650 4520
rect 35770 4400 35815 4520
rect 35935 4400 35980 4520
rect 36100 4400 36155 4520
rect 36275 4400 36485 4520
rect 36605 4400 36650 4520
rect 36770 4400 36815 4520
rect 36935 4400 36980 4520
rect 37100 4400 37155 4520
rect 37275 4400 37320 4520
rect 37440 4400 37485 4520
rect 37605 4400 37650 4520
rect 37770 4400 37825 4520
rect 37945 4400 37990 4520
rect 38110 4400 38155 4520
rect 38275 4400 38320 4520
rect 38440 4400 38495 4520
rect 38615 4400 38660 4520
rect 38780 4400 38825 4520
rect 38945 4400 38990 4520
rect 39110 4400 39165 4520
rect 39285 4400 39330 4520
rect 39450 4400 39495 4520
rect 39615 4400 39660 4520
rect 39780 4400 39835 4520
rect 39955 4400 40000 4520
rect 40120 4400 40165 4520
rect 40285 4400 40330 4520
rect 40450 4400 40505 4520
rect 40625 4400 40670 4520
rect 40790 4400 40835 4520
rect 40955 4400 41000 4520
rect 41120 4400 41175 4520
rect 41295 4400 41340 4520
rect 41460 4400 41505 4520
rect 41625 4400 41670 4520
rect 41790 4400 41845 4520
rect 41965 4400 42175 4520
rect 42295 4400 42340 4520
rect 42460 4400 42505 4520
rect 42625 4400 42670 4520
rect 42790 4400 42845 4520
rect 42965 4400 43010 4520
rect 43130 4400 43175 4520
rect 43295 4400 43340 4520
rect 43460 4400 43515 4520
rect 43635 4400 43680 4520
rect 43800 4400 43845 4520
rect 43965 4400 44010 4520
rect 44130 4400 44185 4520
rect 44305 4400 44350 4520
rect 44470 4400 44515 4520
rect 44635 4400 44680 4520
rect 44800 4400 44855 4520
rect 44975 4400 45020 4520
rect 45140 4400 45185 4520
rect 45305 4400 45350 4520
rect 45470 4400 45525 4520
rect 45645 4400 45690 4520
rect 45810 4400 45855 4520
rect 45975 4400 46020 4520
rect 46140 4400 46195 4520
rect 46315 4400 46360 4520
rect 46480 4400 46525 4520
rect 46645 4400 46690 4520
rect 46810 4400 46865 4520
rect 46985 4400 47030 4520
rect 47150 4400 47195 4520
rect 47315 4400 47360 4520
rect 47480 4400 47535 4520
rect 47655 4400 47865 4520
rect 47985 4400 48030 4520
rect 48150 4400 48195 4520
rect 48315 4400 48360 4520
rect 48480 4400 48535 4520
rect 48655 4400 48700 4520
rect 48820 4400 48865 4520
rect 48985 4400 49030 4520
rect 49150 4400 49205 4520
rect 49325 4400 49370 4520
rect 49490 4400 49535 4520
rect 49655 4400 49700 4520
rect 49820 4400 49875 4520
rect 49995 4400 50040 4520
rect 50160 4400 50205 4520
rect 50325 4400 50370 4520
rect 50490 4400 50545 4520
rect 50665 4400 50710 4520
rect 50830 4400 50875 4520
rect 50995 4400 51040 4520
rect 51160 4400 51215 4520
rect 51335 4400 51380 4520
rect 51500 4400 51545 4520
rect 51665 4400 51710 4520
rect 51830 4400 51885 4520
rect 52005 4400 52050 4520
rect 52170 4400 52215 4520
rect 52335 4400 52380 4520
rect 52500 4400 52555 4520
rect 52675 4400 52720 4520
rect 52840 4400 52885 4520
rect 53005 4400 53050 4520
rect 53170 4400 53225 4520
rect 53345 4400 53370 4520
rect 30770 4345 53370 4400
rect 30770 4225 30795 4345
rect 30915 4225 30960 4345
rect 31080 4225 31125 4345
rect 31245 4225 31290 4345
rect 31410 4225 31465 4345
rect 31585 4225 31630 4345
rect 31750 4225 31795 4345
rect 31915 4225 31960 4345
rect 32080 4225 32135 4345
rect 32255 4225 32300 4345
rect 32420 4225 32465 4345
rect 32585 4225 32630 4345
rect 32750 4225 32805 4345
rect 32925 4225 32970 4345
rect 33090 4225 33135 4345
rect 33255 4225 33300 4345
rect 33420 4225 33475 4345
rect 33595 4225 33640 4345
rect 33760 4225 33805 4345
rect 33925 4225 33970 4345
rect 34090 4225 34145 4345
rect 34265 4225 34310 4345
rect 34430 4225 34475 4345
rect 34595 4225 34640 4345
rect 34760 4225 34815 4345
rect 34935 4225 34980 4345
rect 35100 4225 35145 4345
rect 35265 4225 35310 4345
rect 35430 4225 35485 4345
rect 35605 4225 35650 4345
rect 35770 4225 35815 4345
rect 35935 4225 35980 4345
rect 36100 4225 36155 4345
rect 36275 4225 36485 4345
rect 36605 4225 36650 4345
rect 36770 4225 36815 4345
rect 36935 4225 36980 4345
rect 37100 4225 37155 4345
rect 37275 4225 37320 4345
rect 37440 4225 37485 4345
rect 37605 4225 37650 4345
rect 37770 4225 37825 4345
rect 37945 4225 37990 4345
rect 38110 4225 38155 4345
rect 38275 4225 38320 4345
rect 38440 4225 38495 4345
rect 38615 4225 38660 4345
rect 38780 4225 38825 4345
rect 38945 4225 38990 4345
rect 39110 4225 39165 4345
rect 39285 4225 39330 4345
rect 39450 4225 39495 4345
rect 39615 4225 39660 4345
rect 39780 4225 39835 4345
rect 39955 4225 40000 4345
rect 40120 4225 40165 4345
rect 40285 4225 40330 4345
rect 40450 4225 40505 4345
rect 40625 4225 40670 4345
rect 40790 4225 40835 4345
rect 40955 4225 41000 4345
rect 41120 4225 41175 4345
rect 41295 4225 41340 4345
rect 41460 4225 41505 4345
rect 41625 4225 41670 4345
rect 41790 4225 41845 4345
rect 41965 4225 42175 4345
rect 42295 4225 42340 4345
rect 42460 4225 42505 4345
rect 42625 4225 42670 4345
rect 42790 4225 42845 4345
rect 42965 4225 43010 4345
rect 43130 4225 43175 4345
rect 43295 4225 43340 4345
rect 43460 4225 43515 4345
rect 43635 4225 43680 4345
rect 43800 4225 43845 4345
rect 43965 4225 44010 4345
rect 44130 4225 44185 4345
rect 44305 4225 44350 4345
rect 44470 4225 44515 4345
rect 44635 4225 44680 4345
rect 44800 4225 44855 4345
rect 44975 4225 45020 4345
rect 45140 4225 45185 4345
rect 45305 4225 45350 4345
rect 45470 4225 45525 4345
rect 45645 4225 45690 4345
rect 45810 4225 45855 4345
rect 45975 4225 46020 4345
rect 46140 4225 46195 4345
rect 46315 4225 46360 4345
rect 46480 4225 46525 4345
rect 46645 4225 46690 4345
rect 46810 4225 46865 4345
rect 46985 4225 47030 4345
rect 47150 4225 47195 4345
rect 47315 4225 47360 4345
rect 47480 4225 47535 4345
rect 47655 4225 47865 4345
rect 47985 4225 48030 4345
rect 48150 4225 48195 4345
rect 48315 4225 48360 4345
rect 48480 4225 48535 4345
rect 48655 4225 48700 4345
rect 48820 4225 48865 4345
rect 48985 4225 49030 4345
rect 49150 4225 49205 4345
rect 49325 4225 49370 4345
rect 49490 4225 49535 4345
rect 49655 4225 49700 4345
rect 49820 4225 49875 4345
rect 49995 4225 50040 4345
rect 50160 4225 50205 4345
rect 50325 4225 50370 4345
rect 50490 4225 50545 4345
rect 50665 4225 50710 4345
rect 50830 4225 50875 4345
rect 50995 4225 51040 4345
rect 51160 4225 51215 4345
rect 51335 4225 51380 4345
rect 51500 4225 51545 4345
rect 51665 4225 51710 4345
rect 51830 4225 51885 4345
rect 52005 4225 52050 4345
rect 52170 4225 52215 4345
rect 52335 4225 52380 4345
rect 52500 4225 52555 4345
rect 52675 4225 52720 4345
rect 52840 4225 52885 4345
rect 53005 4225 53050 4345
rect 53170 4225 53225 4345
rect 53345 4225 53370 4345
rect 30770 4180 53370 4225
rect 30770 4060 30795 4180
rect 30915 4060 30960 4180
rect 31080 4060 31125 4180
rect 31245 4060 31290 4180
rect 31410 4060 31465 4180
rect 31585 4060 31630 4180
rect 31750 4060 31795 4180
rect 31915 4060 31960 4180
rect 32080 4060 32135 4180
rect 32255 4060 32300 4180
rect 32420 4060 32465 4180
rect 32585 4060 32630 4180
rect 32750 4060 32805 4180
rect 32925 4060 32970 4180
rect 33090 4060 33135 4180
rect 33255 4060 33300 4180
rect 33420 4060 33475 4180
rect 33595 4060 33640 4180
rect 33760 4060 33805 4180
rect 33925 4060 33970 4180
rect 34090 4060 34145 4180
rect 34265 4060 34310 4180
rect 34430 4060 34475 4180
rect 34595 4060 34640 4180
rect 34760 4060 34815 4180
rect 34935 4060 34980 4180
rect 35100 4060 35145 4180
rect 35265 4060 35310 4180
rect 35430 4060 35485 4180
rect 35605 4060 35650 4180
rect 35770 4060 35815 4180
rect 35935 4060 35980 4180
rect 36100 4060 36155 4180
rect 36275 4060 36485 4180
rect 36605 4060 36650 4180
rect 36770 4060 36815 4180
rect 36935 4060 36980 4180
rect 37100 4060 37155 4180
rect 37275 4060 37320 4180
rect 37440 4060 37485 4180
rect 37605 4060 37650 4180
rect 37770 4060 37825 4180
rect 37945 4060 37990 4180
rect 38110 4060 38155 4180
rect 38275 4060 38320 4180
rect 38440 4060 38495 4180
rect 38615 4060 38660 4180
rect 38780 4060 38825 4180
rect 38945 4060 38990 4180
rect 39110 4060 39165 4180
rect 39285 4060 39330 4180
rect 39450 4060 39495 4180
rect 39615 4060 39660 4180
rect 39780 4060 39835 4180
rect 39955 4060 40000 4180
rect 40120 4060 40165 4180
rect 40285 4060 40330 4180
rect 40450 4060 40505 4180
rect 40625 4060 40670 4180
rect 40790 4060 40835 4180
rect 40955 4060 41000 4180
rect 41120 4060 41175 4180
rect 41295 4060 41340 4180
rect 41460 4060 41505 4180
rect 41625 4060 41670 4180
rect 41790 4060 41845 4180
rect 41965 4060 42175 4180
rect 42295 4060 42340 4180
rect 42460 4060 42505 4180
rect 42625 4060 42670 4180
rect 42790 4060 42845 4180
rect 42965 4060 43010 4180
rect 43130 4060 43175 4180
rect 43295 4060 43340 4180
rect 43460 4060 43515 4180
rect 43635 4060 43680 4180
rect 43800 4060 43845 4180
rect 43965 4060 44010 4180
rect 44130 4060 44185 4180
rect 44305 4060 44350 4180
rect 44470 4060 44515 4180
rect 44635 4060 44680 4180
rect 44800 4060 44855 4180
rect 44975 4060 45020 4180
rect 45140 4060 45185 4180
rect 45305 4060 45350 4180
rect 45470 4060 45525 4180
rect 45645 4060 45690 4180
rect 45810 4060 45855 4180
rect 45975 4060 46020 4180
rect 46140 4060 46195 4180
rect 46315 4060 46360 4180
rect 46480 4060 46525 4180
rect 46645 4060 46690 4180
rect 46810 4060 46865 4180
rect 46985 4060 47030 4180
rect 47150 4060 47195 4180
rect 47315 4060 47360 4180
rect 47480 4060 47535 4180
rect 47655 4060 47865 4180
rect 47985 4060 48030 4180
rect 48150 4060 48195 4180
rect 48315 4060 48360 4180
rect 48480 4060 48535 4180
rect 48655 4060 48700 4180
rect 48820 4060 48865 4180
rect 48985 4060 49030 4180
rect 49150 4060 49205 4180
rect 49325 4060 49370 4180
rect 49490 4060 49535 4180
rect 49655 4060 49700 4180
rect 49820 4060 49875 4180
rect 49995 4060 50040 4180
rect 50160 4060 50205 4180
rect 50325 4060 50370 4180
rect 50490 4060 50545 4180
rect 50665 4060 50710 4180
rect 50830 4060 50875 4180
rect 50995 4060 51040 4180
rect 51160 4060 51215 4180
rect 51335 4060 51380 4180
rect 51500 4060 51545 4180
rect 51665 4060 51710 4180
rect 51830 4060 51885 4180
rect 52005 4060 52050 4180
rect 52170 4060 52215 4180
rect 52335 4060 52380 4180
rect 52500 4060 52555 4180
rect 52675 4060 52720 4180
rect 52840 4060 52885 4180
rect 53005 4060 53050 4180
rect 53170 4060 53225 4180
rect 53345 4060 53370 4180
rect 30770 4015 53370 4060
rect 30770 3895 30795 4015
rect 30915 3895 30960 4015
rect 31080 3895 31125 4015
rect 31245 3895 31290 4015
rect 31410 3895 31465 4015
rect 31585 3895 31630 4015
rect 31750 3895 31795 4015
rect 31915 3895 31960 4015
rect 32080 3895 32135 4015
rect 32255 3895 32300 4015
rect 32420 3895 32465 4015
rect 32585 3895 32630 4015
rect 32750 3895 32805 4015
rect 32925 3895 32970 4015
rect 33090 3895 33135 4015
rect 33255 3895 33300 4015
rect 33420 3895 33475 4015
rect 33595 3895 33640 4015
rect 33760 3895 33805 4015
rect 33925 3895 33970 4015
rect 34090 3895 34145 4015
rect 34265 3895 34310 4015
rect 34430 3895 34475 4015
rect 34595 3895 34640 4015
rect 34760 3895 34815 4015
rect 34935 3895 34980 4015
rect 35100 3895 35145 4015
rect 35265 3895 35310 4015
rect 35430 3895 35485 4015
rect 35605 3895 35650 4015
rect 35770 3895 35815 4015
rect 35935 3895 35980 4015
rect 36100 3895 36155 4015
rect 36275 3895 36485 4015
rect 36605 3895 36650 4015
rect 36770 3895 36815 4015
rect 36935 3895 36980 4015
rect 37100 3895 37155 4015
rect 37275 3895 37320 4015
rect 37440 3895 37485 4015
rect 37605 3895 37650 4015
rect 37770 3895 37825 4015
rect 37945 3895 37990 4015
rect 38110 3895 38155 4015
rect 38275 3895 38320 4015
rect 38440 3895 38495 4015
rect 38615 3895 38660 4015
rect 38780 3895 38825 4015
rect 38945 3895 38990 4015
rect 39110 3895 39165 4015
rect 39285 3895 39330 4015
rect 39450 3895 39495 4015
rect 39615 3895 39660 4015
rect 39780 3895 39835 4015
rect 39955 3895 40000 4015
rect 40120 3895 40165 4015
rect 40285 3895 40330 4015
rect 40450 3895 40505 4015
rect 40625 3895 40670 4015
rect 40790 3895 40835 4015
rect 40955 3895 41000 4015
rect 41120 3895 41175 4015
rect 41295 3895 41340 4015
rect 41460 3895 41505 4015
rect 41625 3895 41670 4015
rect 41790 3895 41845 4015
rect 41965 3895 42175 4015
rect 42295 3895 42340 4015
rect 42460 3895 42505 4015
rect 42625 3895 42670 4015
rect 42790 3895 42845 4015
rect 42965 3895 43010 4015
rect 43130 3895 43175 4015
rect 43295 3895 43340 4015
rect 43460 3895 43515 4015
rect 43635 3895 43680 4015
rect 43800 3895 43845 4015
rect 43965 3895 44010 4015
rect 44130 3895 44185 4015
rect 44305 3895 44350 4015
rect 44470 3895 44515 4015
rect 44635 3895 44680 4015
rect 44800 3895 44855 4015
rect 44975 3895 45020 4015
rect 45140 3895 45185 4015
rect 45305 3895 45350 4015
rect 45470 3895 45525 4015
rect 45645 3895 45690 4015
rect 45810 3895 45855 4015
rect 45975 3895 46020 4015
rect 46140 3895 46195 4015
rect 46315 3895 46360 4015
rect 46480 3895 46525 4015
rect 46645 3895 46690 4015
rect 46810 3895 46865 4015
rect 46985 3895 47030 4015
rect 47150 3895 47195 4015
rect 47315 3895 47360 4015
rect 47480 3895 47535 4015
rect 47655 3895 47865 4015
rect 47985 3895 48030 4015
rect 48150 3895 48195 4015
rect 48315 3895 48360 4015
rect 48480 3895 48535 4015
rect 48655 3895 48700 4015
rect 48820 3895 48865 4015
rect 48985 3895 49030 4015
rect 49150 3895 49205 4015
rect 49325 3895 49370 4015
rect 49490 3895 49535 4015
rect 49655 3895 49700 4015
rect 49820 3895 49875 4015
rect 49995 3895 50040 4015
rect 50160 3895 50205 4015
rect 50325 3895 50370 4015
rect 50490 3895 50545 4015
rect 50665 3895 50710 4015
rect 50830 3895 50875 4015
rect 50995 3895 51040 4015
rect 51160 3895 51215 4015
rect 51335 3895 51380 4015
rect 51500 3895 51545 4015
rect 51665 3895 51710 4015
rect 51830 3895 51885 4015
rect 52005 3895 52050 4015
rect 52170 3895 52215 4015
rect 52335 3895 52380 4015
rect 52500 3895 52555 4015
rect 52675 3895 52720 4015
rect 52840 3895 52885 4015
rect 53005 3895 53050 4015
rect 53170 3895 53225 4015
rect 53345 3895 53370 4015
rect 30770 3850 53370 3895
rect 30770 3730 30795 3850
rect 30915 3730 30960 3850
rect 31080 3730 31125 3850
rect 31245 3730 31290 3850
rect 31410 3730 31465 3850
rect 31585 3730 31630 3850
rect 31750 3730 31795 3850
rect 31915 3730 31960 3850
rect 32080 3730 32135 3850
rect 32255 3730 32300 3850
rect 32420 3730 32465 3850
rect 32585 3730 32630 3850
rect 32750 3730 32805 3850
rect 32925 3730 32970 3850
rect 33090 3730 33135 3850
rect 33255 3730 33300 3850
rect 33420 3730 33475 3850
rect 33595 3730 33640 3850
rect 33760 3730 33805 3850
rect 33925 3730 33970 3850
rect 34090 3730 34145 3850
rect 34265 3730 34310 3850
rect 34430 3730 34475 3850
rect 34595 3730 34640 3850
rect 34760 3730 34815 3850
rect 34935 3730 34980 3850
rect 35100 3730 35145 3850
rect 35265 3730 35310 3850
rect 35430 3730 35485 3850
rect 35605 3730 35650 3850
rect 35770 3730 35815 3850
rect 35935 3730 35980 3850
rect 36100 3730 36155 3850
rect 36275 3730 36485 3850
rect 36605 3730 36650 3850
rect 36770 3730 36815 3850
rect 36935 3730 36980 3850
rect 37100 3730 37155 3850
rect 37275 3730 37320 3850
rect 37440 3730 37485 3850
rect 37605 3730 37650 3850
rect 37770 3730 37825 3850
rect 37945 3730 37990 3850
rect 38110 3730 38155 3850
rect 38275 3730 38320 3850
rect 38440 3730 38495 3850
rect 38615 3730 38660 3850
rect 38780 3730 38825 3850
rect 38945 3730 38990 3850
rect 39110 3730 39165 3850
rect 39285 3730 39330 3850
rect 39450 3730 39495 3850
rect 39615 3730 39660 3850
rect 39780 3730 39835 3850
rect 39955 3730 40000 3850
rect 40120 3730 40165 3850
rect 40285 3730 40330 3850
rect 40450 3730 40505 3850
rect 40625 3730 40670 3850
rect 40790 3730 40835 3850
rect 40955 3730 41000 3850
rect 41120 3730 41175 3850
rect 41295 3730 41340 3850
rect 41460 3730 41505 3850
rect 41625 3730 41670 3850
rect 41790 3730 41845 3850
rect 41965 3730 42175 3850
rect 42295 3730 42340 3850
rect 42460 3730 42505 3850
rect 42625 3730 42670 3850
rect 42790 3730 42845 3850
rect 42965 3730 43010 3850
rect 43130 3730 43175 3850
rect 43295 3730 43340 3850
rect 43460 3730 43515 3850
rect 43635 3730 43680 3850
rect 43800 3730 43845 3850
rect 43965 3730 44010 3850
rect 44130 3730 44185 3850
rect 44305 3730 44350 3850
rect 44470 3730 44515 3850
rect 44635 3730 44680 3850
rect 44800 3730 44855 3850
rect 44975 3730 45020 3850
rect 45140 3730 45185 3850
rect 45305 3730 45350 3850
rect 45470 3730 45525 3850
rect 45645 3730 45690 3850
rect 45810 3730 45855 3850
rect 45975 3730 46020 3850
rect 46140 3730 46195 3850
rect 46315 3730 46360 3850
rect 46480 3730 46525 3850
rect 46645 3730 46690 3850
rect 46810 3730 46865 3850
rect 46985 3730 47030 3850
rect 47150 3730 47195 3850
rect 47315 3730 47360 3850
rect 47480 3730 47535 3850
rect 47655 3730 47865 3850
rect 47985 3730 48030 3850
rect 48150 3730 48195 3850
rect 48315 3730 48360 3850
rect 48480 3730 48535 3850
rect 48655 3730 48700 3850
rect 48820 3730 48865 3850
rect 48985 3730 49030 3850
rect 49150 3730 49205 3850
rect 49325 3730 49370 3850
rect 49490 3730 49535 3850
rect 49655 3730 49700 3850
rect 49820 3730 49875 3850
rect 49995 3730 50040 3850
rect 50160 3730 50205 3850
rect 50325 3730 50370 3850
rect 50490 3730 50545 3850
rect 50665 3730 50710 3850
rect 50830 3730 50875 3850
rect 50995 3730 51040 3850
rect 51160 3730 51215 3850
rect 51335 3730 51380 3850
rect 51500 3730 51545 3850
rect 51665 3730 51710 3850
rect 51830 3730 51885 3850
rect 52005 3730 52050 3850
rect 52170 3730 52215 3850
rect 52335 3730 52380 3850
rect 52500 3730 52555 3850
rect 52675 3730 52720 3850
rect 52840 3730 52885 3850
rect 53005 3730 53050 3850
rect 53170 3730 53225 3850
rect 53345 3730 53370 3850
rect 30770 3675 53370 3730
rect 30770 3555 30795 3675
rect 30915 3555 30960 3675
rect 31080 3555 31125 3675
rect 31245 3555 31290 3675
rect 31410 3555 31465 3675
rect 31585 3555 31630 3675
rect 31750 3555 31795 3675
rect 31915 3555 31960 3675
rect 32080 3555 32135 3675
rect 32255 3555 32300 3675
rect 32420 3555 32465 3675
rect 32585 3555 32630 3675
rect 32750 3555 32805 3675
rect 32925 3555 32970 3675
rect 33090 3555 33135 3675
rect 33255 3555 33300 3675
rect 33420 3555 33475 3675
rect 33595 3555 33640 3675
rect 33760 3555 33805 3675
rect 33925 3555 33970 3675
rect 34090 3555 34145 3675
rect 34265 3555 34310 3675
rect 34430 3555 34475 3675
rect 34595 3555 34640 3675
rect 34760 3555 34815 3675
rect 34935 3555 34980 3675
rect 35100 3555 35145 3675
rect 35265 3555 35310 3675
rect 35430 3555 35485 3675
rect 35605 3555 35650 3675
rect 35770 3555 35815 3675
rect 35935 3555 35980 3675
rect 36100 3555 36155 3675
rect 36275 3555 36485 3675
rect 36605 3555 36650 3675
rect 36770 3555 36815 3675
rect 36935 3555 36980 3675
rect 37100 3555 37155 3675
rect 37275 3555 37320 3675
rect 37440 3555 37485 3675
rect 37605 3555 37650 3675
rect 37770 3555 37825 3675
rect 37945 3555 37990 3675
rect 38110 3555 38155 3675
rect 38275 3555 38320 3675
rect 38440 3555 38495 3675
rect 38615 3555 38660 3675
rect 38780 3555 38825 3675
rect 38945 3555 38990 3675
rect 39110 3555 39165 3675
rect 39285 3555 39330 3675
rect 39450 3555 39495 3675
rect 39615 3555 39660 3675
rect 39780 3555 39835 3675
rect 39955 3555 40000 3675
rect 40120 3555 40165 3675
rect 40285 3555 40330 3675
rect 40450 3555 40505 3675
rect 40625 3555 40670 3675
rect 40790 3555 40835 3675
rect 40955 3555 41000 3675
rect 41120 3555 41175 3675
rect 41295 3555 41340 3675
rect 41460 3555 41505 3675
rect 41625 3555 41670 3675
rect 41790 3555 41845 3675
rect 41965 3555 42175 3675
rect 42295 3555 42340 3675
rect 42460 3555 42505 3675
rect 42625 3555 42670 3675
rect 42790 3555 42845 3675
rect 42965 3555 43010 3675
rect 43130 3555 43175 3675
rect 43295 3555 43340 3675
rect 43460 3555 43515 3675
rect 43635 3555 43680 3675
rect 43800 3555 43845 3675
rect 43965 3555 44010 3675
rect 44130 3555 44185 3675
rect 44305 3555 44350 3675
rect 44470 3555 44515 3675
rect 44635 3555 44680 3675
rect 44800 3555 44855 3675
rect 44975 3555 45020 3675
rect 45140 3555 45185 3675
rect 45305 3555 45350 3675
rect 45470 3555 45525 3675
rect 45645 3555 45690 3675
rect 45810 3555 45855 3675
rect 45975 3555 46020 3675
rect 46140 3555 46195 3675
rect 46315 3555 46360 3675
rect 46480 3555 46525 3675
rect 46645 3555 46690 3675
rect 46810 3555 46865 3675
rect 46985 3555 47030 3675
rect 47150 3555 47195 3675
rect 47315 3555 47360 3675
rect 47480 3555 47535 3675
rect 47655 3555 47865 3675
rect 47985 3555 48030 3675
rect 48150 3555 48195 3675
rect 48315 3555 48360 3675
rect 48480 3555 48535 3675
rect 48655 3555 48700 3675
rect 48820 3555 48865 3675
rect 48985 3555 49030 3675
rect 49150 3555 49205 3675
rect 49325 3555 49370 3675
rect 49490 3555 49535 3675
rect 49655 3555 49700 3675
rect 49820 3555 49875 3675
rect 49995 3555 50040 3675
rect 50160 3555 50205 3675
rect 50325 3555 50370 3675
rect 50490 3555 50545 3675
rect 50665 3555 50710 3675
rect 50830 3555 50875 3675
rect 50995 3555 51040 3675
rect 51160 3555 51215 3675
rect 51335 3555 51380 3675
rect 51500 3555 51545 3675
rect 51665 3555 51710 3675
rect 51830 3555 51885 3675
rect 52005 3555 52050 3675
rect 52170 3555 52215 3675
rect 52335 3555 52380 3675
rect 52500 3555 52555 3675
rect 52675 3555 52720 3675
rect 52840 3555 52885 3675
rect 53005 3555 53050 3675
rect 53170 3555 53225 3675
rect 53345 3555 53370 3675
rect 30770 3510 53370 3555
rect 30770 3390 30795 3510
rect 30915 3390 30960 3510
rect 31080 3390 31125 3510
rect 31245 3390 31290 3510
rect 31410 3390 31465 3510
rect 31585 3390 31630 3510
rect 31750 3390 31795 3510
rect 31915 3390 31960 3510
rect 32080 3390 32135 3510
rect 32255 3390 32300 3510
rect 32420 3390 32465 3510
rect 32585 3390 32630 3510
rect 32750 3390 32805 3510
rect 32925 3390 32970 3510
rect 33090 3390 33135 3510
rect 33255 3390 33300 3510
rect 33420 3390 33475 3510
rect 33595 3390 33640 3510
rect 33760 3390 33805 3510
rect 33925 3390 33970 3510
rect 34090 3390 34145 3510
rect 34265 3390 34310 3510
rect 34430 3390 34475 3510
rect 34595 3390 34640 3510
rect 34760 3390 34815 3510
rect 34935 3390 34980 3510
rect 35100 3390 35145 3510
rect 35265 3390 35310 3510
rect 35430 3390 35485 3510
rect 35605 3390 35650 3510
rect 35770 3390 35815 3510
rect 35935 3390 35980 3510
rect 36100 3390 36155 3510
rect 36275 3390 36485 3510
rect 36605 3390 36650 3510
rect 36770 3390 36815 3510
rect 36935 3390 36980 3510
rect 37100 3390 37155 3510
rect 37275 3390 37320 3510
rect 37440 3390 37485 3510
rect 37605 3390 37650 3510
rect 37770 3390 37825 3510
rect 37945 3390 37990 3510
rect 38110 3390 38155 3510
rect 38275 3390 38320 3510
rect 38440 3390 38495 3510
rect 38615 3390 38660 3510
rect 38780 3390 38825 3510
rect 38945 3390 38990 3510
rect 39110 3390 39165 3510
rect 39285 3390 39330 3510
rect 39450 3390 39495 3510
rect 39615 3390 39660 3510
rect 39780 3390 39835 3510
rect 39955 3390 40000 3510
rect 40120 3390 40165 3510
rect 40285 3390 40330 3510
rect 40450 3390 40505 3510
rect 40625 3390 40670 3510
rect 40790 3390 40835 3510
rect 40955 3390 41000 3510
rect 41120 3390 41175 3510
rect 41295 3390 41340 3510
rect 41460 3390 41505 3510
rect 41625 3390 41670 3510
rect 41790 3390 41845 3510
rect 41965 3390 42175 3510
rect 42295 3390 42340 3510
rect 42460 3390 42505 3510
rect 42625 3390 42670 3510
rect 42790 3390 42845 3510
rect 42965 3390 43010 3510
rect 43130 3390 43175 3510
rect 43295 3390 43340 3510
rect 43460 3390 43515 3510
rect 43635 3390 43680 3510
rect 43800 3390 43845 3510
rect 43965 3390 44010 3510
rect 44130 3390 44185 3510
rect 44305 3390 44350 3510
rect 44470 3390 44515 3510
rect 44635 3390 44680 3510
rect 44800 3390 44855 3510
rect 44975 3390 45020 3510
rect 45140 3390 45185 3510
rect 45305 3390 45350 3510
rect 45470 3390 45525 3510
rect 45645 3390 45690 3510
rect 45810 3390 45855 3510
rect 45975 3390 46020 3510
rect 46140 3390 46195 3510
rect 46315 3390 46360 3510
rect 46480 3390 46525 3510
rect 46645 3390 46690 3510
rect 46810 3390 46865 3510
rect 46985 3390 47030 3510
rect 47150 3390 47195 3510
rect 47315 3390 47360 3510
rect 47480 3390 47535 3510
rect 47655 3390 47865 3510
rect 47985 3390 48030 3510
rect 48150 3390 48195 3510
rect 48315 3390 48360 3510
rect 48480 3390 48535 3510
rect 48655 3390 48700 3510
rect 48820 3390 48865 3510
rect 48985 3390 49030 3510
rect 49150 3390 49205 3510
rect 49325 3390 49370 3510
rect 49490 3390 49535 3510
rect 49655 3390 49700 3510
rect 49820 3390 49875 3510
rect 49995 3390 50040 3510
rect 50160 3390 50205 3510
rect 50325 3390 50370 3510
rect 50490 3390 50545 3510
rect 50665 3390 50710 3510
rect 50830 3390 50875 3510
rect 50995 3390 51040 3510
rect 51160 3390 51215 3510
rect 51335 3390 51380 3510
rect 51500 3390 51545 3510
rect 51665 3390 51710 3510
rect 51830 3390 51885 3510
rect 52005 3390 52050 3510
rect 52170 3390 52215 3510
rect 52335 3390 52380 3510
rect 52500 3390 52555 3510
rect 52675 3390 52720 3510
rect 52840 3390 52885 3510
rect 53005 3390 53050 3510
rect 53170 3390 53225 3510
rect 53345 3390 53370 3510
rect 30770 3345 53370 3390
rect 30770 3225 30795 3345
rect 30915 3225 30960 3345
rect 31080 3225 31125 3345
rect 31245 3225 31290 3345
rect 31410 3225 31465 3345
rect 31585 3225 31630 3345
rect 31750 3225 31795 3345
rect 31915 3225 31960 3345
rect 32080 3225 32135 3345
rect 32255 3225 32300 3345
rect 32420 3225 32465 3345
rect 32585 3225 32630 3345
rect 32750 3225 32805 3345
rect 32925 3225 32970 3345
rect 33090 3225 33135 3345
rect 33255 3225 33300 3345
rect 33420 3225 33475 3345
rect 33595 3225 33640 3345
rect 33760 3225 33805 3345
rect 33925 3225 33970 3345
rect 34090 3225 34145 3345
rect 34265 3225 34310 3345
rect 34430 3225 34475 3345
rect 34595 3225 34640 3345
rect 34760 3225 34815 3345
rect 34935 3225 34980 3345
rect 35100 3225 35145 3345
rect 35265 3225 35310 3345
rect 35430 3225 35485 3345
rect 35605 3225 35650 3345
rect 35770 3225 35815 3345
rect 35935 3225 35980 3345
rect 36100 3225 36155 3345
rect 36275 3225 36485 3345
rect 36605 3225 36650 3345
rect 36770 3225 36815 3345
rect 36935 3225 36980 3345
rect 37100 3225 37155 3345
rect 37275 3225 37320 3345
rect 37440 3225 37485 3345
rect 37605 3225 37650 3345
rect 37770 3225 37825 3345
rect 37945 3225 37990 3345
rect 38110 3225 38155 3345
rect 38275 3225 38320 3345
rect 38440 3225 38495 3345
rect 38615 3225 38660 3345
rect 38780 3225 38825 3345
rect 38945 3225 38990 3345
rect 39110 3225 39165 3345
rect 39285 3225 39330 3345
rect 39450 3225 39495 3345
rect 39615 3225 39660 3345
rect 39780 3225 39835 3345
rect 39955 3225 40000 3345
rect 40120 3225 40165 3345
rect 40285 3225 40330 3345
rect 40450 3225 40505 3345
rect 40625 3225 40670 3345
rect 40790 3225 40835 3345
rect 40955 3225 41000 3345
rect 41120 3225 41175 3345
rect 41295 3225 41340 3345
rect 41460 3225 41505 3345
rect 41625 3225 41670 3345
rect 41790 3225 41845 3345
rect 41965 3225 42175 3345
rect 42295 3225 42340 3345
rect 42460 3225 42505 3345
rect 42625 3225 42670 3345
rect 42790 3225 42845 3345
rect 42965 3225 43010 3345
rect 43130 3225 43175 3345
rect 43295 3225 43340 3345
rect 43460 3225 43515 3345
rect 43635 3225 43680 3345
rect 43800 3225 43845 3345
rect 43965 3225 44010 3345
rect 44130 3225 44185 3345
rect 44305 3225 44350 3345
rect 44470 3225 44515 3345
rect 44635 3225 44680 3345
rect 44800 3225 44855 3345
rect 44975 3225 45020 3345
rect 45140 3225 45185 3345
rect 45305 3225 45350 3345
rect 45470 3225 45525 3345
rect 45645 3225 45690 3345
rect 45810 3225 45855 3345
rect 45975 3225 46020 3345
rect 46140 3225 46195 3345
rect 46315 3225 46360 3345
rect 46480 3225 46525 3345
rect 46645 3225 46690 3345
rect 46810 3225 46865 3345
rect 46985 3225 47030 3345
rect 47150 3225 47195 3345
rect 47315 3225 47360 3345
rect 47480 3225 47535 3345
rect 47655 3225 47865 3345
rect 47985 3225 48030 3345
rect 48150 3225 48195 3345
rect 48315 3225 48360 3345
rect 48480 3225 48535 3345
rect 48655 3225 48700 3345
rect 48820 3225 48865 3345
rect 48985 3225 49030 3345
rect 49150 3225 49205 3345
rect 49325 3225 49370 3345
rect 49490 3225 49535 3345
rect 49655 3225 49700 3345
rect 49820 3225 49875 3345
rect 49995 3225 50040 3345
rect 50160 3225 50205 3345
rect 50325 3225 50370 3345
rect 50490 3225 50545 3345
rect 50665 3225 50710 3345
rect 50830 3225 50875 3345
rect 50995 3225 51040 3345
rect 51160 3225 51215 3345
rect 51335 3225 51380 3345
rect 51500 3225 51545 3345
rect 51665 3225 51710 3345
rect 51830 3225 51885 3345
rect 52005 3225 52050 3345
rect 52170 3225 52215 3345
rect 52335 3225 52380 3345
rect 52500 3225 52555 3345
rect 52675 3225 52720 3345
rect 52840 3225 52885 3345
rect 53005 3225 53050 3345
rect 53170 3225 53225 3345
rect 53345 3225 53370 3345
rect 30770 3180 53370 3225
rect 30770 3060 30795 3180
rect 30915 3060 30960 3180
rect 31080 3060 31125 3180
rect 31245 3060 31290 3180
rect 31410 3060 31465 3180
rect 31585 3060 31630 3180
rect 31750 3060 31795 3180
rect 31915 3060 31960 3180
rect 32080 3060 32135 3180
rect 32255 3060 32300 3180
rect 32420 3060 32465 3180
rect 32585 3060 32630 3180
rect 32750 3060 32805 3180
rect 32925 3060 32970 3180
rect 33090 3060 33135 3180
rect 33255 3060 33300 3180
rect 33420 3060 33475 3180
rect 33595 3060 33640 3180
rect 33760 3060 33805 3180
rect 33925 3060 33970 3180
rect 34090 3060 34145 3180
rect 34265 3060 34310 3180
rect 34430 3060 34475 3180
rect 34595 3060 34640 3180
rect 34760 3060 34815 3180
rect 34935 3060 34980 3180
rect 35100 3060 35145 3180
rect 35265 3060 35310 3180
rect 35430 3060 35485 3180
rect 35605 3060 35650 3180
rect 35770 3060 35815 3180
rect 35935 3060 35980 3180
rect 36100 3060 36155 3180
rect 36275 3060 36485 3180
rect 36605 3060 36650 3180
rect 36770 3060 36815 3180
rect 36935 3060 36980 3180
rect 37100 3060 37155 3180
rect 37275 3060 37320 3180
rect 37440 3060 37485 3180
rect 37605 3060 37650 3180
rect 37770 3060 37825 3180
rect 37945 3060 37990 3180
rect 38110 3060 38155 3180
rect 38275 3060 38320 3180
rect 38440 3060 38495 3180
rect 38615 3060 38660 3180
rect 38780 3060 38825 3180
rect 38945 3060 38990 3180
rect 39110 3060 39165 3180
rect 39285 3060 39330 3180
rect 39450 3060 39495 3180
rect 39615 3060 39660 3180
rect 39780 3060 39835 3180
rect 39955 3060 40000 3180
rect 40120 3060 40165 3180
rect 40285 3060 40330 3180
rect 40450 3060 40505 3180
rect 40625 3060 40670 3180
rect 40790 3060 40835 3180
rect 40955 3060 41000 3180
rect 41120 3060 41175 3180
rect 41295 3060 41340 3180
rect 41460 3060 41505 3180
rect 41625 3060 41670 3180
rect 41790 3060 41845 3180
rect 41965 3060 42175 3180
rect 42295 3060 42340 3180
rect 42460 3060 42505 3180
rect 42625 3060 42670 3180
rect 42790 3060 42845 3180
rect 42965 3060 43010 3180
rect 43130 3060 43175 3180
rect 43295 3060 43340 3180
rect 43460 3060 43515 3180
rect 43635 3060 43680 3180
rect 43800 3060 43845 3180
rect 43965 3060 44010 3180
rect 44130 3060 44185 3180
rect 44305 3060 44350 3180
rect 44470 3060 44515 3180
rect 44635 3060 44680 3180
rect 44800 3060 44855 3180
rect 44975 3060 45020 3180
rect 45140 3060 45185 3180
rect 45305 3060 45350 3180
rect 45470 3060 45525 3180
rect 45645 3060 45690 3180
rect 45810 3060 45855 3180
rect 45975 3060 46020 3180
rect 46140 3060 46195 3180
rect 46315 3060 46360 3180
rect 46480 3060 46525 3180
rect 46645 3060 46690 3180
rect 46810 3060 46865 3180
rect 46985 3060 47030 3180
rect 47150 3060 47195 3180
rect 47315 3060 47360 3180
rect 47480 3060 47535 3180
rect 47655 3060 47865 3180
rect 47985 3060 48030 3180
rect 48150 3060 48195 3180
rect 48315 3060 48360 3180
rect 48480 3060 48535 3180
rect 48655 3060 48700 3180
rect 48820 3060 48865 3180
rect 48985 3060 49030 3180
rect 49150 3060 49205 3180
rect 49325 3060 49370 3180
rect 49490 3060 49535 3180
rect 49655 3060 49700 3180
rect 49820 3060 49875 3180
rect 49995 3060 50040 3180
rect 50160 3060 50205 3180
rect 50325 3060 50370 3180
rect 50490 3060 50545 3180
rect 50665 3060 50710 3180
rect 50830 3060 50875 3180
rect 50995 3060 51040 3180
rect 51160 3060 51215 3180
rect 51335 3060 51380 3180
rect 51500 3060 51545 3180
rect 51665 3060 51710 3180
rect 51830 3060 51885 3180
rect 52005 3060 52050 3180
rect 52170 3060 52215 3180
rect 52335 3060 52380 3180
rect 52500 3060 52555 3180
rect 52675 3060 52720 3180
rect 52840 3060 52885 3180
rect 53005 3060 53050 3180
rect 53170 3060 53225 3180
rect 53345 3060 53370 3180
rect 30770 3005 53370 3060
rect 30770 2885 30795 3005
rect 30915 2885 30960 3005
rect 31080 2885 31125 3005
rect 31245 2885 31290 3005
rect 31410 2885 31465 3005
rect 31585 2885 31630 3005
rect 31750 2885 31795 3005
rect 31915 2885 31960 3005
rect 32080 2885 32135 3005
rect 32255 2885 32300 3005
rect 32420 2885 32465 3005
rect 32585 2885 32630 3005
rect 32750 2885 32805 3005
rect 32925 2885 32970 3005
rect 33090 2885 33135 3005
rect 33255 2885 33300 3005
rect 33420 2885 33475 3005
rect 33595 2885 33640 3005
rect 33760 2885 33805 3005
rect 33925 2885 33970 3005
rect 34090 2885 34145 3005
rect 34265 2885 34310 3005
rect 34430 2885 34475 3005
rect 34595 2885 34640 3005
rect 34760 2885 34815 3005
rect 34935 2885 34980 3005
rect 35100 2885 35145 3005
rect 35265 2885 35310 3005
rect 35430 2885 35485 3005
rect 35605 2885 35650 3005
rect 35770 2885 35815 3005
rect 35935 2885 35980 3005
rect 36100 2885 36155 3005
rect 36275 2885 36485 3005
rect 36605 2885 36650 3005
rect 36770 2885 36815 3005
rect 36935 2885 36980 3005
rect 37100 2885 37155 3005
rect 37275 2885 37320 3005
rect 37440 2885 37485 3005
rect 37605 2885 37650 3005
rect 37770 2885 37825 3005
rect 37945 2885 37990 3005
rect 38110 2885 38155 3005
rect 38275 2885 38320 3005
rect 38440 2885 38495 3005
rect 38615 2885 38660 3005
rect 38780 2885 38825 3005
rect 38945 2885 38990 3005
rect 39110 2885 39165 3005
rect 39285 2885 39330 3005
rect 39450 2885 39495 3005
rect 39615 2885 39660 3005
rect 39780 2885 39835 3005
rect 39955 2885 40000 3005
rect 40120 2885 40165 3005
rect 40285 2885 40330 3005
rect 40450 2885 40505 3005
rect 40625 2885 40670 3005
rect 40790 2885 40835 3005
rect 40955 2885 41000 3005
rect 41120 2885 41175 3005
rect 41295 2885 41340 3005
rect 41460 2885 41505 3005
rect 41625 2885 41670 3005
rect 41790 2885 41845 3005
rect 41965 2885 42175 3005
rect 42295 2885 42340 3005
rect 42460 2885 42505 3005
rect 42625 2885 42670 3005
rect 42790 2885 42845 3005
rect 42965 2885 43010 3005
rect 43130 2885 43175 3005
rect 43295 2885 43340 3005
rect 43460 2885 43515 3005
rect 43635 2885 43680 3005
rect 43800 2885 43845 3005
rect 43965 2885 44010 3005
rect 44130 2885 44185 3005
rect 44305 2885 44350 3005
rect 44470 2885 44515 3005
rect 44635 2885 44680 3005
rect 44800 2885 44855 3005
rect 44975 2885 45020 3005
rect 45140 2885 45185 3005
rect 45305 2885 45350 3005
rect 45470 2885 45525 3005
rect 45645 2885 45690 3005
rect 45810 2885 45855 3005
rect 45975 2885 46020 3005
rect 46140 2885 46195 3005
rect 46315 2885 46360 3005
rect 46480 2885 46525 3005
rect 46645 2885 46690 3005
rect 46810 2885 46865 3005
rect 46985 2885 47030 3005
rect 47150 2885 47195 3005
rect 47315 2885 47360 3005
rect 47480 2885 47535 3005
rect 47655 2885 47865 3005
rect 47985 2885 48030 3005
rect 48150 2885 48195 3005
rect 48315 2885 48360 3005
rect 48480 2885 48535 3005
rect 48655 2885 48700 3005
rect 48820 2885 48865 3005
rect 48985 2885 49030 3005
rect 49150 2885 49205 3005
rect 49325 2885 49370 3005
rect 49490 2885 49535 3005
rect 49655 2885 49700 3005
rect 49820 2885 49875 3005
rect 49995 2885 50040 3005
rect 50160 2885 50205 3005
rect 50325 2885 50370 3005
rect 50490 2885 50545 3005
rect 50665 2885 50710 3005
rect 50830 2885 50875 3005
rect 50995 2885 51040 3005
rect 51160 2885 51215 3005
rect 51335 2885 51380 3005
rect 51500 2885 51545 3005
rect 51665 2885 51710 3005
rect 51830 2885 51885 3005
rect 52005 2885 52050 3005
rect 52170 2885 52215 3005
rect 52335 2885 52380 3005
rect 52500 2885 52555 3005
rect 52675 2885 52720 3005
rect 52840 2885 52885 3005
rect 53005 2885 53050 3005
rect 53170 2885 53225 3005
rect 53345 2885 53370 3005
rect 30770 2840 53370 2885
rect 30770 2720 30795 2840
rect 30915 2720 30960 2840
rect 31080 2720 31125 2840
rect 31245 2720 31290 2840
rect 31410 2720 31465 2840
rect 31585 2720 31630 2840
rect 31750 2720 31795 2840
rect 31915 2720 31960 2840
rect 32080 2720 32135 2840
rect 32255 2720 32300 2840
rect 32420 2720 32465 2840
rect 32585 2720 32630 2840
rect 32750 2720 32805 2840
rect 32925 2720 32970 2840
rect 33090 2720 33135 2840
rect 33255 2720 33300 2840
rect 33420 2720 33475 2840
rect 33595 2720 33640 2840
rect 33760 2720 33805 2840
rect 33925 2720 33970 2840
rect 34090 2720 34145 2840
rect 34265 2720 34310 2840
rect 34430 2720 34475 2840
rect 34595 2720 34640 2840
rect 34760 2720 34815 2840
rect 34935 2720 34980 2840
rect 35100 2720 35145 2840
rect 35265 2720 35310 2840
rect 35430 2720 35485 2840
rect 35605 2720 35650 2840
rect 35770 2720 35815 2840
rect 35935 2720 35980 2840
rect 36100 2720 36155 2840
rect 36275 2720 36485 2840
rect 36605 2720 36650 2840
rect 36770 2720 36815 2840
rect 36935 2720 36980 2840
rect 37100 2720 37155 2840
rect 37275 2720 37320 2840
rect 37440 2720 37485 2840
rect 37605 2720 37650 2840
rect 37770 2720 37825 2840
rect 37945 2720 37990 2840
rect 38110 2720 38155 2840
rect 38275 2720 38320 2840
rect 38440 2720 38495 2840
rect 38615 2720 38660 2840
rect 38780 2720 38825 2840
rect 38945 2720 38990 2840
rect 39110 2720 39165 2840
rect 39285 2720 39330 2840
rect 39450 2720 39495 2840
rect 39615 2720 39660 2840
rect 39780 2720 39835 2840
rect 39955 2720 40000 2840
rect 40120 2720 40165 2840
rect 40285 2720 40330 2840
rect 40450 2720 40505 2840
rect 40625 2720 40670 2840
rect 40790 2720 40835 2840
rect 40955 2720 41000 2840
rect 41120 2720 41175 2840
rect 41295 2720 41340 2840
rect 41460 2720 41505 2840
rect 41625 2720 41670 2840
rect 41790 2720 41845 2840
rect 41965 2720 42175 2840
rect 42295 2720 42340 2840
rect 42460 2720 42505 2840
rect 42625 2720 42670 2840
rect 42790 2720 42845 2840
rect 42965 2720 43010 2840
rect 43130 2720 43175 2840
rect 43295 2720 43340 2840
rect 43460 2720 43515 2840
rect 43635 2720 43680 2840
rect 43800 2720 43845 2840
rect 43965 2720 44010 2840
rect 44130 2720 44185 2840
rect 44305 2720 44350 2840
rect 44470 2720 44515 2840
rect 44635 2720 44680 2840
rect 44800 2720 44855 2840
rect 44975 2720 45020 2840
rect 45140 2720 45185 2840
rect 45305 2720 45350 2840
rect 45470 2720 45525 2840
rect 45645 2720 45690 2840
rect 45810 2720 45855 2840
rect 45975 2720 46020 2840
rect 46140 2720 46195 2840
rect 46315 2720 46360 2840
rect 46480 2720 46525 2840
rect 46645 2720 46690 2840
rect 46810 2720 46865 2840
rect 46985 2720 47030 2840
rect 47150 2720 47195 2840
rect 47315 2720 47360 2840
rect 47480 2720 47535 2840
rect 47655 2720 47865 2840
rect 47985 2720 48030 2840
rect 48150 2720 48195 2840
rect 48315 2720 48360 2840
rect 48480 2720 48535 2840
rect 48655 2720 48700 2840
rect 48820 2720 48865 2840
rect 48985 2720 49030 2840
rect 49150 2720 49205 2840
rect 49325 2720 49370 2840
rect 49490 2720 49535 2840
rect 49655 2720 49700 2840
rect 49820 2720 49875 2840
rect 49995 2720 50040 2840
rect 50160 2720 50205 2840
rect 50325 2720 50370 2840
rect 50490 2720 50545 2840
rect 50665 2720 50710 2840
rect 50830 2720 50875 2840
rect 50995 2720 51040 2840
rect 51160 2720 51215 2840
rect 51335 2720 51380 2840
rect 51500 2720 51545 2840
rect 51665 2720 51710 2840
rect 51830 2720 51885 2840
rect 52005 2720 52050 2840
rect 52170 2720 52215 2840
rect 52335 2720 52380 2840
rect 52500 2720 52555 2840
rect 52675 2720 52720 2840
rect 52840 2720 52885 2840
rect 53005 2720 53050 2840
rect 53170 2720 53225 2840
rect 53345 2720 53370 2840
rect 30770 2675 53370 2720
rect 30770 2555 30795 2675
rect 30915 2555 30960 2675
rect 31080 2555 31125 2675
rect 31245 2555 31290 2675
rect 31410 2555 31465 2675
rect 31585 2555 31630 2675
rect 31750 2555 31795 2675
rect 31915 2555 31960 2675
rect 32080 2555 32135 2675
rect 32255 2555 32300 2675
rect 32420 2555 32465 2675
rect 32585 2555 32630 2675
rect 32750 2555 32805 2675
rect 32925 2555 32970 2675
rect 33090 2555 33135 2675
rect 33255 2555 33300 2675
rect 33420 2555 33475 2675
rect 33595 2555 33640 2675
rect 33760 2555 33805 2675
rect 33925 2555 33970 2675
rect 34090 2555 34145 2675
rect 34265 2555 34310 2675
rect 34430 2555 34475 2675
rect 34595 2555 34640 2675
rect 34760 2555 34815 2675
rect 34935 2555 34980 2675
rect 35100 2555 35145 2675
rect 35265 2555 35310 2675
rect 35430 2555 35485 2675
rect 35605 2555 35650 2675
rect 35770 2555 35815 2675
rect 35935 2555 35980 2675
rect 36100 2555 36155 2675
rect 36275 2555 36485 2675
rect 36605 2555 36650 2675
rect 36770 2555 36815 2675
rect 36935 2555 36980 2675
rect 37100 2555 37155 2675
rect 37275 2555 37320 2675
rect 37440 2555 37485 2675
rect 37605 2555 37650 2675
rect 37770 2555 37825 2675
rect 37945 2555 37990 2675
rect 38110 2555 38155 2675
rect 38275 2555 38320 2675
rect 38440 2555 38495 2675
rect 38615 2555 38660 2675
rect 38780 2555 38825 2675
rect 38945 2555 38990 2675
rect 39110 2555 39165 2675
rect 39285 2555 39330 2675
rect 39450 2555 39495 2675
rect 39615 2555 39660 2675
rect 39780 2555 39835 2675
rect 39955 2555 40000 2675
rect 40120 2555 40165 2675
rect 40285 2555 40330 2675
rect 40450 2555 40505 2675
rect 40625 2555 40670 2675
rect 40790 2555 40835 2675
rect 40955 2555 41000 2675
rect 41120 2555 41175 2675
rect 41295 2555 41340 2675
rect 41460 2555 41505 2675
rect 41625 2555 41670 2675
rect 41790 2555 41845 2675
rect 41965 2555 42175 2675
rect 42295 2555 42340 2675
rect 42460 2555 42505 2675
rect 42625 2555 42670 2675
rect 42790 2555 42845 2675
rect 42965 2555 43010 2675
rect 43130 2555 43175 2675
rect 43295 2555 43340 2675
rect 43460 2555 43515 2675
rect 43635 2555 43680 2675
rect 43800 2555 43845 2675
rect 43965 2555 44010 2675
rect 44130 2555 44185 2675
rect 44305 2555 44350 2675
rect 44470 2555 44515 2675
rect 44635 2555 44680 2675
rect 44800 2555 44855 2675
rect 44975 2555 45020 2675
rect 45140 2555 45185 2675
rect 45305 2555 45350 2675
rect 45470 2555 45525 2675
rect 45645 2555 45690 2675
rect 45810 2555 45855 2675
rect 45975 2555 46020 2675
rect 46140 2555 46195 2675
rect 46315 2555 46360 2675
rect 46480 2555 46525 2675
rect 46645 2555 46690 2675
rect 46810 2555 46865 2675
rect 46985 2555 47030 2675
rect 47150 2555 47195 2675
rect 47315 2555 47360 2675
rect 47480 2555 47535 2675
rect 47655 2555 47865 2675
rect 47985 2555 48030 2675
rect 48150 2555 48195 2675
rect 48315 2555 48360 2675
rect 48480 2555 48535 2675
rect 48655 2555 48700 2675
rect 48820 2555 48865 2675
rect 48985 2555 49030 2675
rect 49150 2555 49205 2675
rect 49325 2555 49370 2675
rect 49490 2555 49535 2675
rect 49655 2555 49700 2675
rect 49820 2555 49875 2675
rect 49995 2555 50040 2675
rect 50160 2555 50205 2675
rect 50325 2555 50370 2675
rect 50490 2555 50545 2675
rect 50665 2555 50710 2675
rect 50830 2555 50875 2675
rect 50995 2555 51040 2675
rect 51160 2555 51215 2675
rect 51335 2555 51380 2675
rect 51500 2555 51545 2675
rect 51665 2555 51710 2675
rect 51830 2555 51885 2675
rect 52005 2555 52050 2675
rect 52170 2555 52215 2675
rect 52335 2555 52380 2675
rect 52500 2555 52555 2675
rect 52675 2555 52720 2675
rect 52840 2555 52885 2675
rect 53005 2555 53050 2675
rect 53170 2555 53225 2675
rect 53345 2555 53370 2675
rect 30770 2510 53370 2555
rect 30770 2390 30795 2510
rect 30915 2390 30960 2510
rect 31080 2390 31125 2510
rect 31245 2390 31290 2510
rect 31410 2390 31465 2510
rect 31585 2390 31630 2510
rect 31750 2390 31795 2510
rect 31915 2390 31960 2510
rect 32080 2390 32135 2510
rect 32255 2390 32300 2510
rect 32420 2390 32465 2510
rect 32585 2390 32630 2510
rect 32750 2390 32805 2510
rect 32925 2390 32970 2510
rect 33090 2390 33135 2510
rect 33255 2390 33300 2510
rect 33420 2390 33475 2510
rect 33595 2390 33640 2510
rect 33760 2390 33805 2510
rect 33925 2390 33970 2510
rect 34090 2390 34145 2510
rect 34265 2390 34310 2510
rect 34430 2390 34475 2510
rect 34595 2390 34640 2510
rect 34760 2390 34815 2510
rect 34935 2390 34980 2510
rect 35100 2390 35145 2510
rect 35265 2390 35310 2510
rect 35430 2390 35485 2510
rect 35605 2390 35650 2510
rect 35770 2390 35815 2510
rect 35935 2390 35980 2510
rect 36100 2390 36155 2510
rect 36275 2390 36485 2510
rect 36605 2390 36650 2510
rect 36770 2390 36815 2510
rect 36935 2390 36980 2510
rect 37100 2390 37155 2510
rect 37275 2390 37320 2510
rect 37440 2390 37485 2510
rect 37605 2390 37650 2510
rect 37770 2390 37825 2510
rect 37945 2390 37990 2510
rect 38110 2390 38155 2510
rect 38275 2390 38320 2510
rect 38440 2390 38495 2510
rect 38615 2390 38660 2510
rect 38780 2390 38825 2510
rect 38945 2390 38990 2510
rect 39110 2390 39165 2510
rect 39285 2390 39330 2510
rect 39450 2390 39495 2510
rect 39615 2390 39660 2510
rect 39780 2390 39835 2510
rect 39955 2390 40000 2510
rect 40120 2390 40165 2510
rect 40285 2390 40330 2510
rect 40450 2390 40505 2510
rect 40625 2390 40670 2510
rect 40790 2390 40835 2510
rect 40955 2390 41000 2510
rect 41120 2390 41175 2510
rect 41295 2390 41340 2510
rect 41460 2390 41505 2510
rect 41625 2390 41670 2510
rect 41790 2390 41845 2510
rect 41965 2390 42175 2510
rect 42295 2390 42340 2510
rect 42460 2390 42505 2510
rect 42625 2390 42670 2510
rect 42790 2390 42845 2510
rect 42965 2390 43010 2510
rect 43130 2390 43175 2510
rect 43295 2390 43340 2510
rect 43460 2390 43515 2510
rect 43635 2390 43680 2510
rect 43800 2390 43845 2510
rect 43965 2390 44010 2510
rect 44130 2390 44185 2510
rect 44305 2390 44350 2510
rect 44470 2390 44515 2510
rect 44635 2390 44680 2510
rect 44800 2390 44855 2510
rect 44975 2390 45020 2510
rect 45140 2390 45185 2510
rect 45305 2390 45350 2510
rect 45470 2390 45525 2510
rect 45645 2390 45690 2510
rect 45810 2390 45855 2510
rect 45975 2390 46020 2510
rect 46140 2390 46195 2510
rect 46315 2390 46360 2510
rect 46480 2390 46525 2510
rect 46645 2390 46690 2510
rect 46810 2390 46865 2510
rect 46985 2390 47030 2510
rect 47150 2390 47195 2510
rect 47315 2390 47360 2510
rect 47480 2390 47535 2510
rect 47655 2390 47865 2510
rect 47985 2390 48030 2510
rect 48150 2390 48195 2510
rect 48315 2390 48360 2510
rect 48480 2390 48535 2510
rect 48655 2390 48700 2510
rect 48820 2390 48865 2510
rect 48985 2390 49030 2510
rect 49150 2390 49205 2510
rect 49325 2390 49370 2510
rect 49490 2390 49535 2510
rect 49655 2390 49700 2510
rect 49820 2390 49875 2510
rect 49995 2390 50040 2510
rect 50160 2390 50205 2510
rect 50325 2390 50370 2510
rect 50490 2390 50545 2510
rect 50665 2390 50710 2510
rect 50830 2390 50875 2510
rect 50995 2390 51040 2510
rect 51160 2390 51215 2510
rect 51335 2390 51380 2510
rect 51500 2390 51545 2510
rect 51665 2390 51710 2510
rect 51830 2390 51885 2510
rect 52005 2390 52050 2510
rect 52170 2390 52215 2510
rect 52335 2390 52380 2510
rect 52500 2390 52555 2510
rect 52675 2390 52720 2510
rect 52840 2390 52885 2510
rect 53005 2390 53050 2510
rect 53170 2390 53225 2510
rect 53345 2390 53370 2510
rect 30770 2335 53370 2390
rect 30770 2215 30795 2335
rect 30915 2215 30960 2335
rect 31080 2215 31125 2335
rect 31245 2215 31290 2335
rect 31410 2215 31465 2335
rect 31585 2215 31630 2335
rect 31750 2215 31795 2335
rect 31915 2215 31960 2335
rect 32080 2215 32135 2335
rect 32255 2215 32300 2335
rect 32420 2215 32465 2335
rect 32585 2215 32630 2335
rect 32750 2215 32805 2335
rect 32925 2215 32970 2335
rect 33090 2215 33135 2335
rect 33255 2215 33300 2335
rect 33420 2215 33475 2335
rect 33595 2215 33640 2335
rect 33760 2215 33805 2335
rect 33925 2215 33970 2335
rect 34090 2215 34145 2335
rect 34265 2215 34310 2335
rect 34430 2215 34475 2335
rect 34595 2215 34640 2335
rect 34760 2215 34815 2335
rect 34935 2215 34980 2335
rect 35100 2215 35145 2335
rect 35265 2215 35310 2335
rect 35430 2215 35485 2335
rect 35605 2215 35650 2335
rect 35770 2215 35815 2335
rect 35935 2215 35980 2335
rect 36100 2215 36155 2335
rect 36275 2215 36485 2335
rect 36605 2215 36650 2335
rect 36770 2215 36815 2335
rect 36935 2215 36980 2335
rect 37100 2215 37155 2335
rect 37275 2215 37320 2335
rect 37440 2215 37485 2335
rect 37605 2215 37650 2335
rect 37770 2215 37825 2335
rect 37945 2215 37990 2335
rect 38110 2215 38155 2335
rect 38275 2215 38320 2335
rect 38440 2215 38495 2335
rect 38615 2215 38660 2335
rect 38780 2215 38825 2335
rect 38945 2215 38990 2335
rect 39110 2215 39165 2335
rect 39285 2215 39330 2335
rect 39450 2215 39495 2335
rect 39615 2215 39660 2335
rect 39780 2215 39835 2335
rect 39955 2215 40000 2335
rect 40120 2215 40165 2335
rect 40285 2215 40330 2335
rect 40450 2215 40505 2335
rect 40625 2215 40670 2335
rect 40790 2215 40835 2335
rect 40955 2215 41000 2335
rect 41120 2215 41175 2335
rect 41295 2215 41340 2335
rect 41460 2215 41505 2335
rect 41625 2215 41670 2335
rect 41790 2215 41845 2335
rect 41965 2215 42175 2335
rect 42295 2215 42340 2335
rect 42460 2215 42505 2335
rect 42625 2215 42670 2335
rect 42790 2215 42845 2335
rect 42965 2215 43010 2335
rect 43130 2215 43175 2335
rect 43295 2215 43340 2335
rect 43460 2215 43515 2335
rect 43635 2215 43680 2335
rect 43800 2215 43845 2335
rect 43965 2215 44010 2335
rect 44130 2215 44185 2335
rect 44305 2215 44350 2335
rect 44470 2215 44515 2335
rect 44635 2215 44680 2335
rect 44800 2215 44855 2335
rect 44975 2215 45020 2335
rect 45140 2215 45185 2335
rect 45305 2215 45350 2335
rect 45470 2215 45525 2335
rect 45645 2215 45690 2335
rect 45810 2215 45855 2335
rect 45975 2215 46020 2335
rect 46140 2215 46195 2335
rect 46315 2215 46360 2335
rect 46480 2215 46525 2335
rect 46645 2215 46690 2335
rect 46810 2215 46865 2335
rect 46985 2215 47030 2335
rect 47150 2215 47195 2335
rect 47315 2215 47360 2335
rect 47480 2215 47535 2335
rect 47655 2215 47865 2335
rect 47985 2215 48030 2335
rect 48150 2215 48195 2335
rect 48315 2215 48360 2335
rect 48480 2215 48535 2335
rect 48655 2215 48700 2335
rect 48820 2215 48865 2335
rect 48985 2215 49030 2335
rect 49150 2215 49205 2335
rect 49325 2215 49370 2335
rect 49490 2215 49535 2335
rect 49655 2215 49700 2335
rect 49820 2215 49875 2335
rect 49995 2215 50040 2335
rect 50160 2215 50205 2335
rect 50325 2215 50370 2335
rect 50490 2215 50545 2335
rect 50665 2215 50710 2335
rect 50830 2215 50875 2335
rect 50995 2215 51040 2335
rect 51160 2215 51215 2335
rect 51335 2215 51380 2335
rect 51500 2215 51545 2335
rect 51665 2215 51710 2335
rect 51830 2215 51885 2335
rect 52005 2215 52050 2335
rect 52170 2215 52215 2335
rect 52335 2215 52380 2335
rect 52500 2215 52555 2335
rect 52675 2215 52720 2335
rect 52840 2215 52885 2335
rect 53005 2215 53050 2335
rect 53170 2215 53225 2335
rect 53345 2215 53370 2335
rect 30770 2170 53370 2215
rect 30770 2050 30795 2170
rect 30915 2050 30960 2170
rect 31080 2050 31125 2170
rect 31245 2050 31290 2170
rect 31410 2050 31465 2170
rect 31585 2050 31630 2170
rect 31750 2050 31795 2170
rect 31915 2050 31960 2170
rect 32080 2050 32135 2170
rect 32255 2050 32300 2170
rect 32420 2050 32465 2170
rect 32585 2050 32630 2170
rect 32750 2050 32805 2170
rect 32925 2050 32970 2170
rect 33090 2050 33135 2170
rect 33255 2050 33300 2170
rect 33420 2050 33475 2170
rect 33595 2050 33640 2170
rect 33760 2050 33805 2170
rect 33925 2050 33970 2170
rect 34090 2050 34145 2170
rect 34265 2050 34310 2170
rect 34430 2050 34475 2170
rect 34595 2050 34640 2170
rect 34760 2050 34815 2170
rect 34935 2050 34980 2170
rect 35100 2050 35145 2170
rect 35265 2050 35310 2170
rect 35430 2050 35485 2170
rect 35605 2050 35650 2170
rect 35770 2050 35815 2170
rect 35935 2050 35980 2170
rect 36100 2050 36155 2170
rect 36275 2050 36485 2170
rect 36605 2050 36650 2170
rect 36770 2050 36815 2170
rect 36935 2050 36980 2170
rect 37100 2050 37155 2170
rect 37275 2050 37320 2170
rect 37440 2050 37485 2170
rect 37605 2050 37650 2170
rect 37770 2050 37825 2170
rect 37945 2050 37990 2170
rect 38110 2050 38155 2170
rect 38275 2050 38320 2170
rect 38440 2050 38495 2170
rect 38615 2050 38660 2170
rect 38780 2050 38825 2170
rect 38945 2050 38990 2170
rect 39110 2050 39165 2170
rect 39285 2050 39330 2170
rect 39450 2050 39495 2170
rect 39615 2050 39660 2170
rect 39780 2050 39835 2170
rect 39955 2050 40000 2170
rect 40120 2050 40165 2170
rect 40285 2050 40330 2170
rect 40450 2050 40505 2170
rect 40625 2050 40670 2170
rect 40790 2050 40835 2170
rect 40955 2050 41000 2170
rect 41120 2050 41175 2170
rect 41295 2050 41340 2170
rect 41460 2050 41505 2170
rect 41625 2050 41670 2170
rect 41790 2050 41845 2170
rect 41965 2050 42175 2170
rect 42295 2050 42340 2170
rect 42460 2050 42505 2170
rect 42625 2050 42670 2170
rect 42790 2050 42845 2170
rect 42965 2050 43010 2170
rect 43130 2050 43175 2170
rect 43295 2050 43340 2170
rect 43460 2050 43515 2170
rect 43635 2050 43680 2170
rect 43800 2050 43845 2170
rect 43965 2050 44010 2170
rect 44130 2050 44185 2170
rect 44305 2050 44350 2170
rect 44470 2050 44515 2170
rect 44635 2050 44680 2170
rect 44800 2050 44855 2170
rect 44975 2050 45020 2170
rect 45140 2050 45185 2170
rect 45305 2050 45350 2170
rect 45470 2050 45525 2170
rect 45645 2050 45690 2170
rect 45810 2050 45855 2170
rect 45975 2050 46020 2170
rect 46140 2050 46195 2170
rect 46315 2050 46360 2170
rect 46480 2050 46525 2170
rect 46645 2050 46690 2170
rect 46810 2050 46865 2170
rect 46985 2050 47030 2170
rect 47150 2050 47195 2170
rect 47315 2050 47360 2170
rect 47480 2050 47535 2170
rect 47655 2050 47865 2170
rect 47985 2050 48030 2170
rect 48150 2050 48195 2170
rect 48315 2050 48360 2170
rect 48480 2050 48535 2170
rect 48655 2050 48700 2170
rect 48820 2050 48865 2170
rect 48985 2050 49030 2170
rect 49150 2050 49205 2170
rect 49325 2050 49370 2170
rect 49490 2050 49535 2170
rect 49655 2050 49700 2170
rect 49820 2050 49875 2170
rect 49995 2050 50040 2170
rect 50160 2050 50205 2170
rect 50325 2050 50370 2170
rect 50490 2050 50545 2170
rect 50665 2050 50710 2170
rect 50830 2050 50875 2170
rect 50995 2050 51040 2170
rect 51160 2050 51215 2170
rect 51335 2050 51380 2170
rect 51500 2050 51545 2170
rect 51665 2050 51710 2170
rect 51830 2050 51885 2170
rect 52005 2050 52050 2170
rect 52170 2050 52215 2170
rect 52335 2050 52380 2170
rect 52500 2050 52555 2170
rect 52675 2050 52720 2170
rect 52840 2050 52885 2170
rect 53005 2050 53050 2170
rect 53170 2050 53225 2170
rect 53345 2050 53370 2170
rect 30770 2005 53370 2050
rect 30770 1885 30795 2005
rect 30915 1885 30960 2005
rect 31080 1885 31125 2005
rect 31245 1885 31290 2005
rect 31410 1885 31465 2005
rect 31585 1885 31630 2005
rect 31750 1885 31795 2005
rect 31915 1885 31960 2005
rect 32080 1885 32135 2005
rect 32255 1885 32300 2005
rect 32420 1885 32465 2005
rect 32585 1885 32630 2005
rect 32750 1885 32805 2005
rect 32925 1885 32970 2005
rect 33090 1885 33135 2005
rect 33255 1885 33300 2005
rect 33420 1885 33475 2005
rect 33595 1885 33640 2005
rect 33760 1885 33805 2005
rect 33925 1885 33970 2005
rect 34090 1885 34145 2005
rect 34265 1885 34310 2005
rect 34430 1885 34475 2005
rect 34595 1885 34640 2005
rect 34760 1885 34815 2005
rect 34935 1885 34980 2005
rect 35100 1885 35145 2005
rect 35265 1885 35310 2005
rect 35430 1885 35485 2005
rect 35605 1885 35650 2005
rect 35770 1885 35815 2005
rect 35935 1885 35980 2005
rect 36100 1885 36155 2005
rect 36275 1885 36485 2005
rect 36605 1885 36650 2005
rect 36770 1885 36815 2005
rect 36935 1885 36980 2005
rect 37100 1885 37155 2005
rect 37275 1885 37320 2005
rect 37440 1885 37485 2005
rect 37605 1885 37650 2005
rect 37770 1885 37825 2005
rect 37945 1885 37990 2005
rect 38110 1885 38155 2005
rect 38275 1885 38320 2005
rect 38440 1885 38495 2005
rect 38615 1885 38660 2005
rect 38780 1885 38825 2005
rect 38945 1885 38990 2005
rect 39110 1885 39165 2005
rect 39285 1885 39330 2005
rect 39450 1885 39495 2005
rect 39615 1885 39660 2005
rect 39780 1885 39835 2005
rect 39955 1885 40000 2005
rect 40120 1885 40165 2005
rect 40285 1885 40330 2005
rect 40450 1885 40505 2005
rect 40625 1885 40670 2005
rect 40790 1885 40835 2005
rect 40955 1885 41000 2005
rect 41120 1885 41175 2005
rect 41295 1885 41340 2005
rect 41460 1885 41505 2005
rect 41625 1885 41670 2005
rect 41790 1885 41845 2005
rect 41965 1885 42175 2005
rect 42295 1885 42340 2005
rect 42460 1885 42505 2005
rect 42625 1885 42670 2005
rect 42790 1885 42845 2005
rect 42965 1885 43010 2005
rect 43130 1885 43175 2005
rect 43295 1885 43340 2005
rect 43460 1885 43515 2005
rect 43635 1885 43680 2005
rect 43800 1885 43845 2005
rect 43965 1885 44010 2005
rect 44130 1885 44185 2005
rect 44305 1885 44350 2005
rect 44470 1885 44515 2005
rect 44635 1885 44680 2005
rect 44800 1885 44855 2005
rect 44975 1885 45020 2005
rect 45140 1885 45185 2005
rect 45305 1885 45350 2005
rect 45470 1885 45525 2005
rect 45645 1885 45690 2005
rect 45810 1885 45855 2005
rect 45975 1885 46020 2005
rect 46140 1885 46195 2005
rect 46315 1885 46360 2005
rect 46480 1885 46525 2005
rect 46645 1885 46690 2005
rect 46810 1885 46865 2005
rect 46985 1885 47030 2005
rect 47150 1885 47195 2005
rect 47315 1885 47360 2005
rect 47480 1885 47535 2005
rect 47655 1885 47865 2005
rect 47985 1885 48030 2005
rect 48150 1885 48195 2005
rect 48315 1885 48360 2005
rect 48480 1885 48535 2005
rect 48655 1885 48700 2005
rect 48820 1885 48865 2005
rect 48985 1885 49030 2005
rect 49150 1885 49205 2005
rect 49325 1885 49370 2005
rect 49490 1885 49535 2005
rect 49655 1885 49700 2005
rect 49820 1885 49875 2005
rect 49995 1885 50040 2005
rect 50160 1885 50205 2005
rect 50325 1885 50370 2005
rect 50490 1885 50545 2005
rect 50665 1885 50710 2005
rect 50830 1885 50875 2005
rect 50995 1885 51040 2005
rect 51160 1885 51215 2005
rect 51335 1885 51380 2005
rect 51500 1885 51545 2005
rect 51665 1885 51710 2005
rect 51830 1885 51885 2005
rect 52005 1885 52050 2005
rect 52170 1885 52215 2005
rect 52335 1885 52380 2005
rect 52500 1885 52555 2005
rect 52675 1885 52720 2005
rect 52840 1885 52885 2005
rect 53005 1885 53050 2005
rect 53170 1885 53225 2005
rect 53345 1885 53370 2005
rect 30770 1840 53370 1885
rect 30770 1720 30795 1840
rect 30915 1720 30960 1840
rect 31080 1720 31125 1840
rect 31245 1720 31290 1840
rect 31410 1720 31465 1840
rect 31585 1720 31630 1840
rect 31750 1720 31795 1840
rect 31915 1720 31960 1840
rect 32080 1720 32135 1840
rect 32255 1720 32300 1840
rect 32420 1720 32465 1840
rect 32585 1720 32630 1840
rect 32750 1720 32805 1840
rect 32925 1720 32970 1840
rect 33090 1720 33135 1840
rect 33255 1720 33300 1840
rect 33420 1720 33475 1840
rect 33595 1720 33640 1840
rect 33760 1720 33805 1840
rect 33925 1720 33970 1840
rect 34090 1720 34145 1840
rect 34265 1720 34310 1840
rect 34430 1720 34475 1840
rect 34595 1720 34640 1840
rect 34760 1720 34815 1840
rect 34935 1720 34980 1840
rect 35100 1720 35145 1840
rect 35265 1720 35310 1840
rect 35430 1720 35485 1840
rect 35605 1720 35650 1840
rect 35770 1720 35815 1840
rect 35935 1720 35980 1840
rect 36100 1720 36155 1840
rect 36275 1720 36485 1840
rect 36605 1720 36650 1840
rect 36770 1720 36815 1840
rect 36935 1720 36980 1840
rect 37100 1720 37155 1840
rect 37275 1720 37320 1840
rect 37440 1720 37485 1840
rect 37605 1720 37650 1840
rect 37770 1720 37825 1840
rect 37945 1720 37990 1840
rect 38110 1720 38155 1840
rect 38275 1720 38320 1840
rect 38440 1720 38495 1840
rect 38615 1720 38660 1840
rect 38780 1720 38825 1840
rect 38945 1720 38990 1840
rect 39110 1720 39165 1840
rect 39285 1720 39330 1840
rect 39450 1720 39495 1840
rect 39615 1720 39660 1840
rect 39780 1720 39835 1840
rect 39955 1720 40000 1840
rect 40120 1720 40165 1840
rect 40285 1720 40330 1840
rect 40450 1720 40505 1840
rect 40625 1720 40670 1840
rect 40790 1720 40835 1840
rect 40955 1720 41000 1840
rect 41120 1720 41175 1840
rect 41295 1720 41340 1840
rect 41460 1720 41505 1840
rect 41625 1720 41670 1840
rect 41790 1720 41845 1840
rect 41965 1720 42175 1840
rect 42295 1720 42340 1840
rect 42460 1720 42505 1840
rect 42625 1720 42670 1840
rect 42790 1720 42845 1840
rect 42965 1720 43010 1840
rect 43130 1720 43175 1840
rect 43295 1720 43340 1840
rect 43460 1720 43515 1840
rect 43635 1720 43680 1840
rect 43800 1720 43845 1840
rect 43965 1720 44010 1840
rect 44130 1720 44185 1840
rect 44305 1720 44350 1840
rect 44470 1720 44515 1840
rect 44635 1720 44680 1840
rect 44800 1720 44855 1840
rect 44975 1720 45020 1840
rect 45140 1720 45185 1840
rect 45305 1720 45350 1840
rect 45470 1720 45525 1840
rect 45645 1720 45690 1840
rect 45810 1720 45855 1840
rect 45975 1720 46020 1840
rect 46140 1720 46195 1840
rect 46315 1720 46360 1840
rect 46480 1720 46525 1840
rect 46645 1720 46690 1840
rect 46810 1720 46865 1840
rect 46985 1720 47030 1840
rect 47150 1720 47195 1840
rect 47315 1720 47360 1840
rect 47480 1720 47535 1840
rect 47655 1720 47865 1840
rect 47985 1720 48030 1840
rect 48150 1720 48195 1840
rect 48315 1720 48360 1840
rect 48480 1720 48535 1840
rect 48655 1720 48700 1840
rect 48820 1720 48865 1840
rect 48985 1720 49030 1840
rect 49150 1720 49205 1840
rect 49325 1720 49370 1840
rect 49490 1720 49535 1840
rect 49655 1720 49700 1840
rect 49820 1720 49875 1840
rect 49995 1720 50040 1840
rect 50160 1720 50205 1840
rect 50325 1720 50370 1840
rect 50490 1720 50545 1840
rect 50665 1720 50710 1840
rect 50830 1720 50875 1840
rect 50995 1720 51040 1840
rect 51160 1720 51215 1840
rect 51335 1720 51380 1840
rect 51500 1720 51545 1840
rect 51665 1720 51710 1840
rect 51830 1720 51885 1840
rect 52005 1720 52050 1840
rect 52170 1720 52215 1840
rect 52335 1720 52380 1840
rect 52500 1720 52555 1840
rect 52675 1720 52720 1840
rect 52840 1720 52885 1840
rect 53005 1720 53050 1840
rect 53170 1720 53225 1840
rect 53345 1720 53370 1840
rect 30770 1630 53370 1720
rect 30770 1510 30835 1630
rect 30955 1510 31000 1630
rect 31120 1510 31165 1630
rect 31285 1510 31330 1630
rect 31450 1510 31495 1630
rect 31615 1510 31660 1630
rect 31780 1510 31825 1630
rect 31945 1510 31990 1630
rect 32110 1510 32155 1630
rect 32275 1510 32320 1630
rect 32440 1510 32485 1630
rect 32605 1510 32650 1630
rect 32770 1510 32815 1630
rect 32935 1510 32980 1630
rect 33100 1510 33145 1630
rect 33265 1510 33310 1630
rect 33430 1510 33475 1630
rect 33595 1510 33640 1630
rect 33760 1510 33805 1630
rect 33925 1510 33970 1630
rect 34090 1510 34135 1630
rect 34255 1510 34300 1630
rect 34420 1510 34465 1630
rect 34585 1510 34630 1630
rect 34750 1510 34795 1630
rect 34915 1510 34960 1630
rect 35080 1510 35125 1630
rect 35245 1510 35290 1630
rect 35410 1510 35455 1630
rect 35575 1510 35620 1630
rect 35740 1510 35785 1630
rect 35905 1510 35950 1630
rect 36070 1510 36115 1630
rect 36235 1510 36525 1630
rect 36645 1510 36690 1630
rect 36810 1510 36855 1630
rect 36975 1510 37020 1630
rect 37140 1510 37185 1630
rect 37305 1510 37350 1630
rect 37470 1510 37515 1630
rect 37635 1510 37680 1630
rect 37800 1510 37845 1630
rect 37965 1510 38010 1630
rect 38130 1510 38175 1630
rect 38295 1510 38340 1630
rect 38460 1510 38505 1630
rect 38625 1510 38670 1630
rect 38790 1510 38835 1630
rect 38955 1510 39000 1630
rect 39120 1510 39165 1630
rect 39285 1510 39330 1630
rect 39450 1510 39495 1630
rect 39615 1510 39660 1630
rect 39780 1510 39825 1630
rect 39945 1510 39990 1630
rect 40110 1510 40155 1630
rect 40275 1510 40320 1630
rect 40440 1510 40485 1630
rect 40605 1510 40650 1630
rect 40770 1510 40815 1630
rect 40935 1510 40980 1630
rect 41100 1510 41145 1630
rect 41265 1510 41310 1630
rect 41430 1510 41475 1630
rect 41595 1510 41640 1630
rect 41760 1510 41805 1630
rect 41925 1510 42215 1630
rect 42335 1510 42380 1630
rect 42500 1510 42545 1630
rect 42665 1510 42710 1630
rect 42830 1510 42875 1630
rect 42995 1510 43040 1630
rect 43160 1510 43205 1630
rect 43325 1510 43370 1630
rect 43490 1510 43535 1630
rect 43655 1510 43700 1630
rect 43820 1510 43865 1630
rect 43985 1510 44030 1630
rect 44150 1510 44195 1630
rect 44315 1510 44360 1630
rect 44480 1510 44525 1630
rect 44645 1510 44690 1630
rect 44810 1510 44855 1630
rect 44975 1510 45020 1630
rect 45140 1510 45185 1630
rect 45305 1510 45350 1630
rect 45470 1510 45515 1630
rect 45635 1510 45680 1630
rect 45800 1510 45845 1630
rect 45965 1510 46010 1630
rect 46130 1510 46175 1630
rect 46295 1510 46340 1630
rect 46460 1510 46505 1630
rect 46625 1510 46670 1630
rect 46790 1510 46835 1630
rect 46955 1510 47000 1630
rect 47120 1510 47165 1630
rect 47285 1510 47330 1630
rect 47450 1510 47495 1630
rect 47615 1510 47905 1630
rect 48025 1510 48070 1630
rect 48190 1510 48235 1630
rect 48355 1510 48400 1630
rect 48520 1510 48565 1630
rect 48685 1510 48730 1630
rect 48850 1510 48895 1630
rect 49015 1510 49060 1630
rect 49180 1510 49225 1630
rect 49345 1510 49390 1630
rect 49510 1510 49555 1630
rect 49675 1510 49720 1630
rect 49840 1510 49885 1630
rect 50005 1510 50050 1630
rect 50170 1510 50215 1630
rect 50335 1510 50380 1630
rect 50500 1510 50545 1630
rect 50665 1510 50710 1630
rect 50830 1510 50875 1630
rect 50995 1510 51040 1630
rect 51160 1510 51205 1630
rect 51325 1510 51370 1630
rect 51490 1510 51535 1630
rect 51655 1510 51700 1630
rect 51820 1510 51865 1630
rect 51985 1510 52030 1630
rect 52150 1510 52195 1630
rect 52315 1510 52360 1630
rect 52480 1510 52525 1630
rect 52645 1510 52690 1630
rect 52810 1510 52855 1630
rect 52975 1510 53020 1630
rect 53140 1510 53185 1630
rect 53305 1510 53370 1630
rect 30770 1420 53370 1510
rect 30770 1300 30795 1420
rect 30915 1300 30970 1420
rect 31090 1300 31135 1420
rect 31255 1300 31300 1420
rect 31420 1300 31465 1420
rect 31585 1300 31640 1420
rect 31760 1300 31805 1420
rect 31925 1300 31970 1420
rect 32090 1300 32135 1420
rect 32255 1300 32310 1420
rect 32430 1300 32475 1420
rect 32595 1300 32640 1420
rect 32760 1300 32805 1420
rect 32925 1300 32980 1420
rect 33100 1300 33145 1420
rect 33265 1300 33310 1420
rect 33430 1300 33475 1420
rect 33595 1300 33650 1420
rect 33770 1300 33815 1420
rect 33935 1300 33980 1420
rect 34100 1300 34145 1420
rect 34265 1300 34320 1420
rect 34440 1300 34485 1420
rect 34605 1300 34650 1420
rect 34770 1300 34815 1420
rect 34935 1300 34990 1420
rect 35110 1300 35155 1420
rect 35275 1300 35320 1420
rect 35440 1300 35485 1420
rect 35605 1300 35660 1420
rect 35780 1300 35825 1420
rect 35945 1300 35990 1420
rect 36110 1300 36155 1420
rect 36275 1300 36485 1420
rect 36605 1300 36660 1420
rect 36780 1300 36825 1420
rect 36945 1300 36990 1420
rect 37110 1300 37155 1420
rect 37275 1300 37330 1420
rect 37450 1300 37495 1420
rect 37615 1300 37660 1420
rect 37780 1300 37825 1420
rect 37945 1300 38000 1420
rect 38120 1300 38165 1420
rect 38285 1300 38330 1420
rect 38450 1300 38495 1420
rect 38615 1300 38670 1420
rect 38790 1300 38835 1420
rect 38955 1300 39000 1420
rect 39120 1300 39165 1420
rect 39285 1300 39340 1420
rect 39460 1300 39505 1420
rect 39625 1300 39670 1420
rect 39790 1300 39835 1420
rect 39955 1300 40010 1420
rect 40130 1300 40175 1420
rect 40295 1300 40340 1420
rect 40460 1300 40505 1420
rect 40625 1300 40680 1420
rect 40800 1300 40845 1420
rect 40965 1300 41010 1420
rect 41130 1300 41175 1420
rect 41295 1300 41350 1420
rect 41470 1300 41515 1420
rect 41635 1300 41680 1420
rect 41800 1300 41845 1420
rect 41965 1300 42175 1420
rect 42295 1300 42350 1420
rect 42470 1300 42515 1420
rect 42635 1300 42680 1420
rect 42800 1300 42845 1420
rect 42965 1300 43020 1420
rect 43140 1300 43185 1420
rect 43305 1300 43350 1420
rect 43470 1300 43515 1420
rect 43635 1300 43690 1420
rect 43810 1300 43855 1420
rect 43975 1300 44020 1420
rect 44140 1300 44185 1420
rect 44305 1300 44360 1420
rect 44480 1300 44525 1420
rect 44645 1300 44690 1420
rect 44810 1300 44855 1420
rect 44975 1300 45030 1420
rect 45150 1300 45195 1420
rect 45315 1300 45360 1420
rect 45480 1300 45525 1420
rect 45645 1300 45700 1420
rect 45820 1300 45865 1420
rect 45985 1300 46030 1420
rect 46150 1300 46195 1420
rect 46315 1300 46370 1420
rect 46490 1300 46535 1420
rect 46655 1300 46700 1420
rect 46820 1300 46865 1420
rect 46985 1300 47040 1420
rect 47160 1300 47205 1420
rect 47325 1300 47370 1420
rect 47490 1300 47535 1420
rect 47655 1300 47865 1420
rect 47985 1300 48040 1420
rect 48160 1300 48205 1420
rect 48325 1300 48370 1420
rect 48490 1300 48535 1420
rect 48655 1300 48710 1420
rect 48830 1300 48875 1420
rect 48995 1300 49040 1420
rect 49160 1300 49205 1420
rect 49325 1300 49380 1420
rect 49500 1300 49545 1420
rect 49665 1300 49710 1420
rect 49830 1300 49875 1420
rect 49995 1300 50050 1420
rect 50170 1300 50215 1420
rect 50335 1300 50380 1420
rect 50500 1300 50545 1420
rect 50665 1300 50720 1420
rect 50840 1300 50885 1420
rect 51005 1300 51050 1420
rect 51170 1300 51215 1420
rect 51335 1300 51390 1420
rect 51510 1300 51555 1420
rect 51675 1300 51720 1420
rect 51840 1300 51885 1420
rect 52005 1300 52060 1420
rect 52180 1300 52225 1420
rect 52345 1300 52390 1420
rect 52510 1300 52555 1420
rect 52675 1300 52730 1420
rect 52850 1300 52895 1420
rect 53015 1300 53060 1420
rect 53180 1300 53225 1420
rect 53345 1300 53370 1420
rect 30770 1255 53370 1300
rect 30770 1135 30795 1255
rect 30915 1135 30970 1255
rect 31090 1135 31135 1255
rect 31255 1135 31300 1255
rect 31420 1135 31465 1255
rect 31585 1135 31640 1255
rect 31760 1135 31805 1255
rect 31925 1135 31970 1255
rect 32090 1135 32135 1255
rect 32255 1135 32310 1255
rect 32430 1135 32475 1255
rect 32595 1135 32640 1255
rect 32760 1135 32805 1255
rect 32925 1135 32980 1255
rect 33100 1135 33145 1255
rect 33265 1135 33310 1255
rect 33430 1135 33475 1255
rect 33595 1135 33650 1255
rect 33770 1135 33815 1255
rect 33935 1135 33980 1255
rect 34100 1135 34145 1255
rect 34265 1135 34320 1255
rect 34440 1135 34485 1255
rect 34605 1135 34650 1255
rect 34770 1135 34815 1255
rect 34935 1135 34990 1255
rect 35110 1135 35155 1255
rect 35275 1135 35320 1255
rect 35440 1135 35485 1255
rect 35605 1135 35660 1255
rect 35780 1135 35825 1255
rect 35945 1135 35990 1255
rect 36110 1135 36155 1255
rect 36275 1135 36485 1255
rect 36605 1135 36660 1255
rect 36780 1135 36825 1255
rect 36945 1135 36990 1255
rect 37110 1135 37155 1255
rect 37275 1135 37330 1255
rect 37450 1135 37495 1255
rect 37615 1135 37660 1255
rect 37780 1135 37825 1255
rect 37945 1135 38000 1255
rect 38120 1135 38165 1255
rect 38285 1135 38330 1255
rect 38450 1135 38495 1255
rect 38615 1135 38670 1255
rect 38790 1135 38835 1255
rect 38955 1135 39000 1255
rect 39120 1135 39165 1255
rect 39285 1135 39340 1255
rect 39460 1135 39505 1255
rect 39625 1135 39670 1255
rect 39790 1135 39835 1255
rect 39955 1135 40010 1255
rect 40130 1135 40175 1255
rect 40295 1135 40340 1255
rect 40460 1135 40505 1255
rect 40625 1135 40680 1255
rect 40800 1135 40845 1255
rect 40965 1135 41010 1255
rect 41130 1135 41175 1255
rect 41295 1135 41350 1255
rect 41470 1135 41515 1255
rect 41635 1135 41680 1255
rect 41800 1135 41845 1255
rect 41965 1135 42175 1255
rect 42295 1135 42350 1255
rect 42470 1135 42515 1255
rect 42635 1135 42680 1255
rect 42800 1135 42845 1255
rect 42965 1135 43020 1255
rect 43140 1135 43185 1255
rect 43305 1135 43350 1255
rect 43470 1135 43515 1255
rect 43635 1135 43690 1255
rect 43810 1135 43855 1255
rect 43975 1135 44020 1255
rect 44140 1135 44185 1255
rect 44305 1135 44360 1255
rect 44480 1135 44525 1255
rect 44645 1135 44690 1255
rect 44810 1135 44855 1255
rect 44975 1135 45030 1255
rect 45150 1135 45195 1255
rect 45315 1135 45360 1255
rect 45480 1135 45525 1255
rect 45645 1135 45700 1255
rect 45820 1135 45865 1255
rect 45985 1135 46030 1255
rect 46150 1135 46195 1255
rect 46315 1135 46370 1255
rect 46490 1135 46535 1255
rect 46655 1135 46700 1255
rect 46820 1135 46865 1255
rect 46985 1135 47040 1255
rect 47160 1135 47205 1255
rect 47325 1135 47370 1255
rect 47490 1135 47535 1255
rect 47655 1135 47865 1255
rect 47985 1135 48040 1255
rect 48160 1135 48205 1255
rect 48325 1135 48370 1255
rect 48490 1135 48535 1255
rect 48655 1135 48710 1255
rect 48830 1135 48875 1255
rect 48995 1135 49040 1255
rect 49160 1135 49205 1255
rect 49325 1135 49380 1255
rect 49500 1135 49545 1255
rect 49665 1135 49710 1255
rect 49830 1135 49875 1255
rect 49995 1135 50050 1255
rect 50170 1135 50215 1255
rect 50335 1135 50380 1255
rect 50500 1135 50545 1255
rect 50665 1135 50720 1255
rect 50840 1135 50885 1255
rect 51005 1135 51050 1255
rect 51170 1135 51215 1255
rect 51335 1135 51390 1255
rect 51510 1135 51555 1255
rect 51675 1135 51720 1255
rect 51840 1135 51885 1255
rect 52005 1135 52060 1255
rect 52180 1135 52225 1255
rect 52345 1135 52390 1255
rect 52510 1135 52555 1255
rect 52675 1135 52730 1255
rect 52850 1135 52895 1255
rect 53015 1135 53060 1255
rect 53180 1135 53225 1255
rect 53345 1135 53370 1255
rect 30770 1090 53370 1135
rect 30770 970 30795 1090
rect 30915 970 30970 1090
rect 31090 970 31135 1090
rect 31255 970 31300 1090
rect 31420 970 31465 1090
rect 31585 970 31640 1090
rect 31760 970 31805 1090
rect 31925 970 31970 1090
rect 32090 970 32135 1090
rect 32255 970 32310 1090
rect 32430 970 32475 1090
rect 32595 970 32640 1090
rect 32760 970 32805 1090
rect 32925 970 32980 1090
rect 33100 970 33145 1090
rect 33265 970 33310 1090
rect 33430 970 33475 1090
rect 33595 970 33650 1090
rect 33770 970 33815 1090
rect 33935 970 33980 1090
rect 34100 970 34145 1090
rect 34265 970 34320 1090
rect 34440 970 34485 1090
rect 34605 970 34650 1090
rect 34770 970 34815 1090
rect 34935 970 34990 1090
rect 35110 970 35155 1090
rect 35275 970 35320 1090
rect 35440 970 35485 1090
rect 35605 970 35660 1090
rect 35780 970 35825 1090
rect 35945 970 35990 1090
rect 36110 970 36155 1090
rect 36275 970 36485 1090
rect 36605 970 36660 1090
rect 36780 970 36825 1090
rect 36945 970 36990 1090
rect 37110 970 37155 1090
rect 37275 970 37330 1090
rect 37450 970 37495 1090
rect 37615 970 37660 1090
rect 37780 970 37825 1090
rect 37945 970 38000 1090
rect 38120 970 38165 1090
rect 38285 970 38330 1090
rect 38450 970 38495 1090
rect 38615 970 38670 1090
rect 38790 970 38835 1090
rect 38955 970 39000 1090
rect 39120 970 39165 1090
rect 39285 970 39340 1090
rect 39460 970 39505 1090
rect 39625 970 39670 1090
rect 39790 970 39835 1090
rect 39955 970 40010 1090
rect 40130 970 40175 1090
rect 40295 970 40340 1090
rect 40460 970 40505 1090
rect 40625 970 40680 1090
rect 40800 970 40845 1090
rect 40965 970 41010 1090
rect 41130 970 41175 1090
rect 41295 970 41350 1090
rect 41470 970 41515 1090
rect 41635 970 41680 1090
rect 41800 970 41845 1090
rect 41965 970 42175 1090
rect 42295 970 42350 1090
rect 42470 970 42515 1090
rect 42635 970 42680 1090
rect 42800 970 42845 1090
rect 42965 970 43020 1090
rect 43140 970 43185 1090
rect 43305 970 43350 1090
rect 43470 970 43515 1090
rect 43635 970 43690 1090
rect 43810 970 43855 1090
rect 43975 970 44020 1090
rect 44140 970 44185 1090
rect 44305 970 44360 1090
rect 44480 970 44525 1090
rect 44645 970 44690 1090
rect 44810 970 44855 1090
rect 44975 970 45030 1090
rect 45150 970 45195 1090
rect 45315 970 45360 1090
rect 45480 970 45525 1090
rect 45645 970 45700 1090
rect 45820 970 45865 1090
rect 45985 970 46030 1090
rect 46150 970 46195 1090
rect 46315 970 46370 1090
rect 46490 970 46535 1090
rect 46655 970 46700 1090
rect 46820 970 46865 1090
rect 46985 970 47040 1090
rect 47160 970 47205 1090
rect 47325 970 47370 1090
rect 47490 970 47535 1090
rect 47655 970 47865 1090
rect 47985 970 48040 1090
rect 48160 970 48205 1090
rect 48325 970 48370 1090
rect 48490 970 48535 1090
rect 48655 970 48710 1090
rect 48830 970 48875 1090
rect 48995 970 49040 1090
rect 49160 970 49205 1090
rect 49325 970 49380 1090
rect 49500 970 49545 1090
rect 49665 970 49710 1090
rect 49830 970 49875 1090
rect 49995 970 50050 1090
rect 50170 970 50215 1090
rect 50335 970 50380 1090
rect 50500 970 50545 1090
rect 50665 970 50720 1090
rect 50840 970 50885 1090
rect 51005 970 51050 1090
rect 51170 970 51215 1090
rect 51335 970 51390 1090
rect 51510 970 51555 1090
rect 51675 970 51720 1090
rect 51840 970 51885 1090
rect 52005 970 52060 1090
rect 52180 970 52225 1090
rect 52345 970 52390 1090
rect 52510 970 52555 1090
rect 52675 970 52730 1090
rect 52850 970 52895 1090
rect 53015 970 53060 1090
rect 53180 970 53225 1090
rect 53345 970 53370 1090
rect 30770 925 53370 970
rect 30770 805 30795 925
rect 30915 805 30970 925
rect 31090 805 31135 925
rect 31255 805 31300 925
rect 31420 805 31465 925
rect 31585 805 31640 925
rect 31760 805 31805 925
rect 31925 805 31970 925
rect 32090 805 32135 925
rect 32255 805 32310 925
rect 32430 805 32475 925
rect 32595 805 32640 925
rect 32760 805 32805 925
rect 32925 805 32980 925
rect 33100 805 33145 925
rect 33265 805 33310 925
rect 33430 805 33475 925
rect 33595 805 33650 925
rect 33770 805 33815 925
rect 33935 805 33980 925
rect 34100 805 34145 925
rect 34265 805 34320 925
rect 34440 805 34485 925
rect 34605 805 34650 925
rect 34770 805 34815 925
rect 34935 805 34990 925
rect 35110 805 35155 925
rect 35275 805 35320 925
rect 35440 805 35485 925
rect 35605 805 35660 925
rect 35780 805 35825 925
rect 35945 805 35990 925
rect 36110 805 36155 925
rect 36275 805 36485 925
rect 36605 805 36660 925
rect 36780 805 36825 925
rect 36945 805 36990 925
rect 37110 805 37155 925
rect 37275 805 37330 925
rect 37450 805 37495 925
rect 37615 805 37660 925
rect 37780 805 37825 925
rect 37945 805 38000 925
rect 38120 805 38165 925
rect 38285 805 38330 925
rect 38450 805 38495 925
rect 38615 805 38670 925
rect 38790 805 38835 925
rect 38955 805 39000 925
rect 39120 805 39165 925
rect 39285 805 39340 925
rect 39460 805 39505 925
rect 39625 805 39670 925
rect 39790 805 39835 925
rect 39955 805 40010 925
rect 40130 805 40175 925
rect 40295 805 40340 925
rect 40460 805 40505 925
rect 40625 805 40680 925
rect 40800 805 40845 925
rect 40965 805 41010 925
rect 41130 805 41175 925
rect 41295 805 41350 925
rect 41470 805 41515 925
rect 41635 805 41680 925
rect 41800 805 41845 925
rect 41965 805 42175 925
rect 42295 805 42350 925
rect 42470 805 42515 925
rect 42635 805 42680 925
rect 42800 805 42845 925
rect 42965 805 43020 925
rect 43140 805 43185 925
rect 43305 805 43350 925
rect 43470 805 43515 925
rect 43635 805 43690 925
rect 43810 805 43855 925
rect 43975 805 44020 925
rect 44140 805 44185 925
rect 44305 805 44360 925
rect 44480 805 44525 925
rect 44645 805 44690 925
rect 44810 805 44855 925
rect 44975 805 45030 925
rect 45150 805 45195 925
rect 45315 805 45360 925
rect 45480 805 45525 925
rect 45645 805 45700 925
rect 45820 805 45865 925
rect 45985 805 46030 925
rect 46150 805 46195 925
rect 46315 805 46370 925
rect 46490 805 46535 925
rect 46655 805 46700 925
rect 46820 805 46865 925
rect 46985 805 47040 925
rect 47160 805 47205 925
rect 47325 805 47370 925
rect 47490 805 47535 925
rect 47655 805 47865 925
rect 47985 805 48040 925
rect 48160 805 48205 925
rect 48325 805 48370 925
rect 48490 805 48535 925
rect 48655 805 48710 925
rect 48830 805 48875 925
rect 48995 805 49040 925
rect 49160 805 49205 925
rect 49325 805 49380 925
rect 49500 805 49545 925
rect 49665 805 49710 925
rect 49830 805 49875 925
rect 49995 805 50050 925
rect 50170 805 50215 925
rect 50335 805 50380 925
rect 50500 805 50545 925
rect 50665 805 50720 925
rect 50840 805 50885 925
rect 51005 805 51050 925
rect 51170 805 51215 925
rect 51335 805 51390 925
rect 51510 805 51555 925
rect 51675 805 51720 925
rect 51840 805 51885 925
rect 52005 805 52060 925
rect 52180 805 52225 925
rect 52345 805 52390 925
rect 52510 805 52555 925
rect 52675 805 52730 925
rect 52850 805 52895 925
rect 53015 805 53060 925
rect 53180 805 53225 925
rect 53345 805 53370 925
rect 30770 750 53370 805
rect 30770 630 30795 750
rect 30915 630 30970 750
rect 31090 630 31135 750
rect 31255 630 31300 750
rect 31420 630 31465 750
rect 31585 630 31640 750
rect 31760 630 31805 750
rect 31925 630 31970 750
rect 32090 630 32135 750
rect 32255 630 32310 750
rect 32430 630 32475 750
rect 32595 630 32640 750
rect 32760 630 32805 750
rect 32925 630 32980 750
rect 33100 630 33145 750
rect 33265 630 33310 750
rect 33430 630 33475 750
rect 33595 630 33650 750
rect 33770 630 33815 750
rect 33935 630 33980 750
rect 34100 630 34145 750
rect 34265 630 34320 750
rect 34440 630 34485 750
rect 34605 630 34650 750
rect 34770 630 34815 750
rect 34935 630 34990 750
rect 35110 630 35155 750
rect 35275 630 35320 750
rect 35440 630 35485 750
rect 35605 630 35660 750
rect 35780 630 35825 750
rect 35945 630 35990 750
rect 36110 630 36155 750
rect 36275 630 36485 750
rect 36605 630 36660 750
rect 36780 630 36825 750
rect 36945 630 36990 750
rect 37110 630 37155 750
rect 37275 630 37330 750
rect 37450 630 37495 750
rect 37615 630 37660 750
rect 37780 630 37825 750
rect 37945 630 38000 750
rect 38120 630 38165 750
rect 38285 630 38330 750
rect 38450 630 38495 750
rect 38615 630 38670 750
rect 38790 630 38835 750
rect 38955 630 39000 750
rect 39120 630 39165 750
rect 39285 630 39340 750
rect 39460 630 39505 750
rect 39625 630 39670 750
rect 39790 630 39835 750
rect 39955 630 40010 750
rect 40130 630 40175 750
rect 40295 630 40340 750
rect 40460 630 40505 750
rect 40625 630 40680 750
rect 40800 630 40845 750
rect 40965 630 41010 750
rect 41130 630 41175 750
rect 41295 630 41350 750
rect 41470 630 41515 750
rect 41635 630 41680 750
rect 41800 630 41845 750
rect 41965 630 42175 750
rect 42295 630 42350 750
rect 42470 630 42515 750
rect 42635 630 42680 750
rect 42800 630 42845 750
rect 42965 630 43020 750
rect 43140 630 43185 750
rect 43305 630 43350 750
rect 43470 630 43515 750
rect 43635 630 43690 750
rect 43810 630 43855 750
rect 43975 630 44020 750
rect 44140 630 44185 750
rect 44305 630 44360 750
rect 44480 630 44525 750
rect 44645 630 44690 750
rect 44810 630 44855 750
rect 44975 630 45030 750
rect 45150 630 45195 750
rect 45315 630 45360 750
rect 45480 630 45525 750
rect 45645 630 45700 750
rect 45820 630 45865 750
rect 45985 630 46030 750
rect 46150 630 46195 750
rect 46315 630 46370 750
rect 46490 630 46535 750
rect 46655 630 46700 750
rect 46820 630 46865 750
rect 46985 630 47040 750
rect 47160 630 47205 750
rect 47325 630 47370 750
rect 47490 630 47535 750
rect 47655 630 47865 750
rect 47985 630 48040 750
rect 48160 630 48205 750
rect 48325 630 48370 750
rect 48490 630 48535 750
rect 48655 630 48710 750
rect 48830 630 48875 750
rect 48995 630 49040 750
rect 49160 630 49205 750
rect 49325 630 49380 750
rect 49500 630 49545 750
rect 49665 630 49710 750
rect 49830 630 49875 750
rect 49995 630 50050 750
rect 50170 630 50215 750
rect 50335 630 50380 750
rect 50500 630 50545 750
rect 50665 630 50720 750
rect 50840 630 50885 750
rect 51005 630 51050 750
rect 51170 630 51215 750
rect 51335 630 51390 750
rect 51510 630 51555 750
rect 51675 630 51720 750
rect 51840 630 51885 750
rect 52005 630 52060 750
rect 52180 630 52225 750
rect 52345 630 52390 750
rect 52510 630 52555 750
rect 52675 630 52730 750
rect 52850 630 52895 750
rect 53015 630 53060 750
rect 53180 630 53225 750
rect 53345 630 53370 750
rect 30770 585 53370 630
rect 30770 465 30795 585
rect 30915 465 30970 585
rect 31090 465 31135 585
rect 31255 465 31300 585
rect 31420 465 31465 585
rect 31585 465 31640 585
rect 31760 465 31805 585
rect 31925 465 31970 585
rect 32090 465 32135 585
rect 32255 465 32310 585
rect 32430 465 32475 585
rect 32595 465 32640 585
rect 32760 465 32805 585
rect 32925 465 32980 585
rect 33100 465 33145 585
rect 33265 465 33310 585
rect 33430 465 33475 585
rect 33595 465 33650 585
rect 33770 465 33815 585
rect 33935 465 33980 585
rect 34100 465 34145 585
rect 34265 465 34320 585
rect 34440 465 34485 585
rect 34605 465 34650 585
rect 34770 465 34815 585
rect 34935 465 34990 585
rect 35110 465 35155 585
rect 35275 465 35320 585
rect 35440 465 35485 585
rect 35605 465 35660 585
rect 35780 465 35825 585
rect 35945 465 35990 585
rect 36110 465 36155 585
rect 36275 465 36485 585
rect 36605 465 36660 585
rect 36780 465 36825 585
rect 36945 465 36990 585
rect 37110 465 37155 585
rect 37275 465 37330 585
rect 37450 465 37495 585
rect 37615 465 37660 585
rect 37780 465 37825 585
rect 37945 465 38000 585
rect 38120 465 38165 585
rect 38285 465 38330 585
rect 38450 465 38495 585
rect 38615 465 38670 585
rect 38790 465 38835 585
rect 38955 465 39000 585
rect 39120 465 39165 585
rect 39285 465 39340 585
rect 39460 465 39505 585
rect 39625 465 39670 585
rect 39790 465 39835 585
rect 39955 465 40010 585
rect 40130 465 40175 585
rect 40295 465 40340 585
rect 40460 465 40505 585
rect 40625 465 40680 585
rect 40800 465 40845 585
rect 40965 465 41010 585
rect 41130 465 41175 585
rect 41295 465 41350 585
rect 41470 465 41515 585
rect 41635 465 41680 585
rect 41800 465 41845 585
rect 41965 465 42175 585
rect 42295 465 42350 585
rect 42470 465 42515 585
rect 42635 465 42680 585
rect 42800 465 42845 585
rect 42965 465 43020 585
rect 43140 465 43185 585
rect 43305 465 43350 585
rect 43470 465 43515 585
rect 43635 465 43690 585
rect 43810 465 43855 585
rect 43975 465 44020 585
rect 44140 465 44185 585
rect 44305 465 44360 585
rect 44480 465 44525 585
rect 44645 465 44690 585
rect 44810 465 44855 585
rect 44975 465 45030 585
rect 45150 465 45195 585
rect 45315 465 45360 585
rect 45480 465 45525 585
rect 45645 465 45700 585
rect 45820 465 45865 585
rect 45985 465 46030 585
rect 46150 465 46195 585
rect 46315 465 46370 585
rect 46490 465 46535 585
rect 46655 465 46700 585
rect 46820 465 46865 585
rect 46985 465 47040 585
rect 47160 465 47205 585
rect 47325 465 47370 585
rect 47490 465 47535 585
rect 47655 465 47865 585
rect 47985 465 48040 585
rect 48160 465 48205 585
rect 48325 465 48370 585
rect 48490 465 48535 585
rect 48655 465 48710 585
rect 48830 465 48875 585
rect 48995 465 49040 585
rect 49160 465 49205 585
rect 49325 465 49380 585
rect 49500 465 49545 585
rect 49665 465 49710 585
rect 49830 465 49875 585
rect 49995 465 50050 585
rect 50170 465 50215 585
rect 50335 465 50380 585
rect 50500 465 50545 585
rect 50665 465 50720 585
rect 50840 465 50885 585
rect 51005 465 51050 585
rect 51170 465 51215 585
rect 51335 465 51390 585
rect 51510 465 51555 585
rect 51675 465 51720 585
rect 51840 465 51885 585
rect 52005 465 52060 585
rect 52180 465 52225 585
rect 52345 465 52390 585
rect 52510 465 52555 585
rect 52675 465 52730 585
rect 52850 465 52895 585
rect 53015 465 53060 585
rect 53180 465 53225 585
rect 53345 465 53370 585
rect 30770 420 53370 465
rect 30770 300 30795 420
rect 30915 300 30970 420
rect 31090 300 31135 420
rect 31255 300 31300 420
rect 31420 300 31465 420
rect 31585 300 31640 420
rect 31760 300 31805 420
rect 31925 300 31970 420
rect 32090 300 32135 420
rect 32255 300 32310 420
rect 32430 300 32475 420
rect 32595 300 32640 420
rect 32760 300 32805 420
rect 32925 300 32980 420
rect 33100 300 33145 420
rect 33265 300 33310 420
rect 33430 300 33475 420
rect 33595 300 33650 420
rect 33770 300 33815 420
rect 33935 300 33980 420
rect 34100 300 34145 420
rect 34265 300 34320 420
rect 34440 300 34485 420
rect 34605 300 34650 420
rect 34770 300 34815 420
rect 34935 300 34990 420
rect 35110 300 35155 420
rect 35275 300 35320 420
rect 35440 300 35485 420
rect 35605 300 35660 420
rect 35780 300 35825 420
rect 35945 300 35990 420
rect 36110 300 36155 420
rect 36275 300 36485 420
rect 36605 300 36660 420
rect 36780 300 36825 420
rect 36945 300 36990 420
rect 37110 300 37155 420
rect 37275 300 37330 420
rect 37450 300 37495 420
rect 37615 300 37660 420
rect 37780 300 37825 420
rect 37945 300 38000 420
rect 38120 300 38165 420
rect 38285 300 38330 420
rect 38450 300 38495 420
rect 38615 300 38670 420
rect 38790 300 38835 420
rect 38955 300 39000 420
rect 39120 300 39165 420
rect 39285 300 39340 420
rect 39460 300 39505 420
rect 39625 300 39670 420
rect 39790 300 39835 420
rect 39955 300 40010 420
rect 40130 300 40175 420
rect 40295 300 40340 420
rect 40460 300 40505 420
rect 40625 300 40680 420
rect 40800 300 40845 420
rect 40965 300 41010 420
rect 41130 300 41175 420
rect 41295 300 41350 420
rect 41470 300 41515 420
rect 41635 300 41680 420
rect 41800 300 41845 420
rect 41965 300 42175 420
rect 42295 300 42350 420
rect 42470 300 42515 420
rect 42635 300 42680 420
rect 42800 300 42845 420
rect 42965 300 43020 420
rect 43140 300 43185 420
rect 43305 300 43350 420
rect 43470 300 43515 420
rect 43635 300 43690 420
rect 43810 300 43855 420
rect 43975 300 44020 420
rect 44140 300 44185 420
rect 44305 300 44360 420
rect 44480 300 44525 420
rect 44645 300 44690 420
rect 44810 300 44855 420
rect 44975 300 45030 420
rect 45150 300 45195 420
rect 45315 300 45360 420
rect 45480 300 45525 420
rect 45645 300 45700 420
rect 45820 300 45865 420
rect 45985 300 46030 420
rect 46150 300 46195 420
rect 46315 300 46370 420
rect 46490 300 46535 420
rect 46655 300 46700 420
rect 46820 300 46865 420
rect 46985 300 47040 420
rect 47160 300 47205 420
rect 47325 300 47370 420
rect 47490 300 47535 420
rect 47655 300 47865 420
rect 47985 300 48040 420
rect 48160 300 48205 420
rect 48325 300 48370 420
rect 48490 300 48535 420
rect 48655 300 48710 420
rect 48830 300 48875 420
rect 48995 300 49040 420
rect 49160 300 49205 420
rect 49325 300 49380 420
rect 49500 300 49545 420
rect 49665 300 49710 420
rect 49830 300 49875 420
rect 49995 300 50050 420
rect 50170 300 50215 420
rect 50335 300 50380 420
rect 50500 300 50545 420
rect 50665 300 50720 420
rect 50840 300 50885 420
rect 51005 300 51050 420
rect 51170 300 51215 420
rect 51335 300 51390 420
rect 51510 300 51555 420
rect 51675 300 51720 420
rect 51840 300 51885 420
rect 52005 300 52060 420
rect 52180 300 52225 420
rect 52345 300 52390 420
rect 52510 300 52555 420
rect 52675 300 52730 420
rect 52850 300 52895 420
rect 53015 300 53060 420
rect 53180 300 53225 420
rect 53345 300 53370 420
rect 30770 255 53370 300
rect 30770 135 30795 255
rect 30915 135 30970 255
rect 31090 135 31135 255
rect 31255 135 31300 255
rect 31420 135 31465 255
rect 31585 135 31640 255
rect 31760 135 31805 255
rect 31925 135 31970 255
rect 32090 135 32135 255
rect 32255 135 32310 255
rect 32430 135 32475 255
rect 32595 135 32640 255
rect 32760 135 32805 255
rect 32925 135 32980 255
rect 33100 135 33145 255
rect 33265 135 33310 255
rect 33430 135 33475 255
rect 33595 135 33650 255
rect 33770 135 33815 255
rect 33935 135 33980 255
rect 34100 135 34145 255
rect 34265 135 34320 255
rect 34440 135 34485 255
rect 34605 135 34650 255
rect 34770 135 34815 255
rect 34935 135 34990 255
rect 35110 135 35155 255
rect 35275 135 35320 255
rect 35440 135 35485 255
rect 35605 135 35660 255
rect 35780 135 35825 255
rect 35945 135 35990 255
rect 36110 135 36155 255
rect 36275 135 36485 255
rect 36605 135 36660 255
rect 36780 135 36825 255
rect 36945 135 36990 255
rect 37110 135 37155 255
rect 37275 135 37330 255
rect 37450 135 37495 255
rect 37615 135 37660 255
rect 37780 135 37825 255
rect 37945 135 38000 255
rect 38120 135 38165 255
rect 38285 135 38330 255
rect 38450 135 38495 255
rect 38615 135 38670 255
rect 38790 135 38835 255
rect 38955 135 39000 255
rect 39120 135 39165 255
rect 39285 135 39340 255
rect 39460 135 39505 255
rect 39625 135 39670 255
rect 39790 135 39835 255
rect 39955 135 40010 255
rect 40130 135 40175 255
rect 40295 135 40340 255
rect 40460 135 40505 255
rect 40625 135 40680 255
rect 40800 135 40845 255
rect 40965 135 41010 255
rect 41130 135 41175 255
rect 41295 135 41350 255
rect 41470 135 41515 255
rect 41635 135 41680 255
rect 41800 135 41845 255
rect 41965 135 42175 255
rect 42295 135 42350 255
rect 42470 135 42515 255
rect 42635 135 42680 255
rect 42800 135 42845 255
rect 42965 135 43020 255
rect 43140 135 43185 255
rect 43305 135 43350 255
rect 43470 135 43515 255
rect 43635 135 43690 255
rect 43810 135 43855 255
rect 43975 135 44020 255
rect 44140 135 44185 255
rect 44305 135 44360 255
rect 44480 135 44525 255
rect 44645 135 44690 255
rect 44810 135 44855 255
rect 44975 135 45030 255
rect 45150 135 45195 255
rect 45315 135 45360 255
rect 45480 135 45525 255
rect 45645 135 45700 255
rect 45820 135 45865 255
rect 45985 135 46030 255
rect 46150 135 46195 255
rect 46315 135 46370 255
rect 46490 135 46535 255
rect 46655 135 46700 255
rect 46820 135 46865 255
rect 46985 135 47040 255
rect 47160 135 47205 255
rect 47325 135 47370 255
rect 47490 135 47535 255
rect 47655 135 47865 255
rect 47985 135 48040 255
rect 48160 135 48205 255
rect 48325 135 48370 255
rect 48490 135 48535 255
rect 48655 135 48710 255
rect 48830 135 48875 255
rect 48995 135 49040 255
rect 49160 135 49205 255
rect 49325 135 49380 255
rect 49500 135 49545 255
rect 49665 135 49710 255
rect 49830 135 49875 255
rect 49995 135 50050 255
rect 50170 135 50215 255
rect 50335 135 50380 255
rect 50500 135 50545 255
rect 50665 135 50720 255
rect 50840 135 50885 255
rect 51005 135 51050 255
rect 51170 135 51215 255
rect 51335 135 51390 255
rect 51510 135 51555 255
rect 51675 135 51720 255
rect 51840 135 51885 255
rect 52005 135 52060 255
rect 52180 135 52225 255
rect 52345 135 52390 255
rect 52510 135 52555 255
rect 52675 135 52730 255
rect 52850 135 52895 255
rect 53015 135 53060 255
rect 53180 135 53225 255
rect 53345 135 53370 255
rect 30770 80 53370 135
rect 30770 -40 30795 80
rect 30915 -40 30970 80
rect 31090 -40 31135 80
rect 31255 -40 31300 80
rect 31420 -40 31465 80
rect 31585 -40 31640 80
rect 31760 -40 31805 80
rect 31925 -40 31970 80
rect 32090 -40 32135 80
rect 32255 -40 32310 80
rect 32430 -40 32475 80
rect 32595 -40 32640 80
rect 32760 -40 32805 80
rect 32925 -40 32980 80
rect 33100 -40 33145 80
rect 33265 -40 33310 80
rect 33430 -40 33475 80
rect 33595 -40 33650 80
rect 33770 -40 33815 80
rect 33935 -40 33980 80
rect 34100 -40 34145 80
rect 34265 -40 34320 80
rect 34440 -40 34485 80
rect 34605 -40 34650 80
rect 34770 -40 34815 80
rect 34935 -40 34990 80
rect 35110 -40 35155 80
rect 35275 -40 35320 80
rect 35440 -40 35485 80
rect 35605 -40 35660 80
rect 35780 -40 35825 80
rect 35945 -40 35990 80
rect 36110 -40 36155 80
rect 36275 -40 36485 80
rect 36605 -40 36660 80
rect 36780 -40 36825 80
rect 36945 -40 36990 80
rect 37110 -40 37155 80
rect 37275 -40 37330 80
rect 37450 -40 37495 80
rect 37615 -40 37660 80
rect 37780 -40 37825 80
rect 37945 -40 38000 80
rect 38120 -40 38165 80
rect 38285 -40 38330 80
rect 38450 -40 38495 80
rect 38615 -40 38670 80
rect 38790 -40 38835 80
rect 38955 -40 39000 80
rect 39120 -40 39165 80
rect 39285 -40 39340 80
rect 39460 -40 39505 80
rect 39625 -40 39670 80
rect 39790 -40 39835 80
rect 39955 -40 40010 80
rect 40130 -40 40175 80
rect 40295 -40 40340 80
rect 40460 -40 40505 80
rect 40625 -40 40680 80
rect 40800 -40 40845 80
rect 40965 -40 41010 80
rect 41130 -40 41175 80
rect 41295 -40 41350 80
rect 41470 -40 41515 80
rect 41635 -40 41680 80
rect 41800 -40 41845 80
rect 41965 -40 42175 80
rect 42295 -40 42350 80
rect 42470 -40 42515 80
rect 42635 -40 42680 80
rect 42800 -40 42845 80
rect 42965 -40 43020 80
rect 43140 -40 43185 80
rect 43305 -40 43350 80
rect 43470 -40 43515 80
rect 43635 -40 43690 80
rect 43810 -40 43855 80
rect 43975 -40 44020 80
rect 44140 -40 44185 80
rect 44305 -40 44360 80
rect 44480 -40 44525 80
rect 44645 -40 44690 80
rect 44810 -40 44855 80
rect 44975 -40 45030 80
rect 45150 -40 45195 80
rect 45315 -40 45360 80
rect 45480 -40 45525 80
rect 45645 -40 45700 80
rect 45820 -40 45865 80
rect 45985 -40 46030 80
rect 46150 -40 46195 80
rect 46315 -40 46370 80
rect 46490 -40 46535 80
rect 46655 -40 46700 80
rect 46820 -40 46865 80
rect 46985 -40 47040 80
rect 47160 -40 47205 80
rect 47325 -40 47370 80
rect 47490 -40 47535 80
rect 47655 -40 47865 80
rect 47985 -40 48040 80
rect 48160 -40 48205 80
rect 48325 -40 48370 80
rect 48490 -40 48535 80
rect 48655 -40 48710 80
rect 48830 -40 48875 80
rect 48995 -40 49040 80
rect 49160 -40 49205 80
rect 49325 -40 49380 80
rect 49500 -40 49545 80
rect 49665 -40 49710 80
rect 49830 -40 49875 80
rect 49995 -40 50050 80
rect 50170 -40 50215 80
rect 50335 -40 50380 80
rect 50500 -40 50545 80
rect 50665 -40 50720 80
rect 50840 -40 50885 80
rect 51005 -40 51050 80
rect 51170 -40 51215 80
rect 51335 -40 51390 80
rect 51510 -40 51555 80
rect 51675 -40 51720 80
rect 51840 -40 51885 80
rect 52005 -40 52060 80
rect 52180 -40 52225 80
rect 52345 -40 52390 80
rect 52510 -40 52555 80
rect 52675 -40 52730 80
rect 52850 -40 52895 80
rect 53015 -40 53060 80
rect 53180 -40 53225 80
rect 53345 -40 53370 80
rect 30770 -85 53370 -40
rect 30770 -205 30795 -85
rect 30915 -205 30970 -85
rect 31090 -205 31135 -85
rect 31255 -205 31300 -85
rect 31420 -205 31465 -85
rect 31585 -205 31640 -85
rect 31760 -205 31805 -85
rect 31925 -205 31970 -85
rect 32090 -205 32135 -85
rect 32255 -205 32310 -85
rect 32430 -205 32475 -85
rect 32595 -205 32640 -85
rect 32760 -205 32805 -85
rect 32925 -205 32980 -85
rect 33100 -205 33145 -85
rect 33265 -205 33310 -85
rect 33430 -205 33475 -85
rect 33595 -205 33650 -85
rect 33770 -205 33815 -85
rect 33935 -205 33980 -85
rect 34100 -205 34145 -85
rect 34265 -205 34320 -85
rect 34440 -205 34485 -85
rect 34605 -205 34650 -85
rect 34770 -205 34815 -85
rect 34935 -205 34990 -85
rect 35110 -205 35155 -85
rect 35275 -205 35320 -85
rect 35440 -205 35485 -85
rect 35605 -205 35660 -85
rect 35780 -205 35825 -85
rect 35945 -205 35990 -85
rect 36110 -205 36155 -85
rect 36275 -205 36485 -85
rect 36605 -205 36660 -85
rect 36780 -205 36825 -85
rect 36945 -205 36990 -85
rect 37110 -205 37155 -85
rect 37275 -205 37330 -85
rect 37450 -205 37495 -85
rect 37615 -205 37660 -85
rect 37780 -205 37825 -85
rect 37945 -205 38000 -85
rect 38120 -205 38165 -85
rect 38285 -205 38330 -85
rect 38450 -205 38495 -85
rect 38615 -205 38670 -85
rect 38790 -205 38835 -85
rect 38955 -205 39000 -85
rect 39120 -205 39165 -85
rect 39285 -205 39340 -85
rect 39460 -205 39505 -85
rect 39625 -205 39670 -85
rect 39790 -205 39835 -85
rect 39955 -205 40010 -85
rect 40130 -205 40175 -85
rect 40295 -205 40340 -85
rect 40460 -205 40505 -85
rect 40625 -205 40680 -85
rect 40800 -205 40845 -85
rect 40965 -205 41010 -85
rect 41130 -205 41175 -85
rect 41295 -205 41350 -85
rect 41470 -205 41515 -85
rect 41635 -205 41680 -85
rect 41800 -205 41845 -85
rect 41965 -205 42175 -85
rect 42295 -205 42350 -85
rect 42470 -205 42515 -85
rect 42635 -205 42680 -85
rect 42800 -205 42845 -85
rect 42965 -205 43020 -85
rect 43140 -205 43185 -85
rect 43305 -205 43350 -85
rect 43470 -205 43515 -85
rect 43635 -205 43690 -85
rect 43810 -205 43855 -85
rect 43975 -205 44020 -85
rect 44140 -205 44185 -85
rect 44305 -205 44360 -85
rect 44480 -205 44525 -85
rect 44645 -205 44690 -85
rect 44810 -205 44855 -85
rect 44975 -205 45030 -85
rect 45150 -205 45195 -85
rect 45315 -205 45360 -85
rect 45480 -205 45525 -85
rect 45645 -205 45700 -85
rect 45820 -205 45865 -85
rect 45985 -205 46030 -85
rect 46150 -205 46195 -85
rect 46315 -205 46370 -85
rect 46490 -205 46535 -85
rect 46655 -205 46700 -85
rect 46820 -205 46865 -85
rect 46985 -205 47040 -85
rect 47160 -205 47205 -85
rect 47325 -205 47370 -85
rect 47490 -205 47535 -85
rect 47655 -205 47865 -85
rect 47985 -205 48040 -85
rect 48160 -205 48205 -85
rect 48325 -205 48370 -85
rect 48490 -205 48535 -85
rect 48655 -205 48710 -85
rect 48830 -205 48875 -85
rect 48995 -205 49040 -85
rect 49160 -205 49205 -85
rect 49325 -205 49380 -85
rect 49500 -205 49545 -85
rect 49665 -205 49710 -85
rect 49830 -205 49875 -85
rect 49995 -205 50050 -85
rect 50170 -205 50215 -85
rect 50335 -205 50380 -85
rect 50500 -205 50545 -85
rect 50665 -205 50720 -85
rect 50840 -205 50885 -85
rect 51005 -205 51050 -85
rect 51170 -205 51215 -85
rect 51335 -205 51390 -85
rect 51510 -205 51555 -85
rect 51675 -205 51720 -85
rect 51840 -205 51885 -85
rect 52005 -205 52060 -85
rect 52180 -205 52225 -85
rect 52345 -205 52390 -85
rect 52510 -205 52555 -85
rect 52675 -205 52730 -85
rect 52850 -205 52895 -85
rect 53015 -205 53060 -85
rect 53180 -205 53225 -85
rect 53345 -205 53370 -85
rect 30770 -250 53370 -205
rect 30770 -370 30795 -250
rect 30915 -370 30970 -250
rect 31090 -370 31135 -250
rect 31255 -370 31300 -250
rect 31420 -370 31465 -250
rect 31585 -370 31640 -250
rect 31760 -370 31805 -250
rect 31925 -370 31970 -250
rect 32090 -370 32135 -250
rect 32255 -370 32310 -250
rect 32430 -370 32475 -250
rect 32595 -370 32640 -250
rect 32760 -370 32805 -250
rect 32925 -370 32980 -250
rect 33100 -370 33145 -250
rect 33265 -370 33310 -250
rect 33430 -370 33475 -250
rect 33595 -370 33650 -250
rect 33770 -370 33815 -250
rect 33935 -370 33980 -250
rect 34100 -370 34145 -250
rect 34265 -370 34320 -250
rect 34440 -370 34485 -250
rect 34605 -370 34650 -250
rect 34770 -370 34815 -250
rect 34935 -370 34990 -250
rect 35110 -370 35155 -250
rect 35275 -370 35320 -250
rect 35440 -370 35485 -250
rect 35605 -370 35660 -250
rect 35780 -370 35825 -250
rect 35945 -370 35990 -250
rect 36110 -370 36155 -250
rect 36275 -370 36485 -250
rect 36605 -370 36660 -250
rect 36780 -370 36825 -250
rect 36945 -370 36990 -250
rect 37110 -370 37155 -250
rect 37275 -370 37330 -250
rect 37450 -370 37495 -250
rect 37615 -370 37660 -250
rect 37780 -370 37825 -250
rect 37945 -370 38000 -250
rect 38120 -370 38165 -250
rect 38285 -370 38330 -250
rect 38450 -370 38495 -250
rect 38615 -370 38670 -250
rect 38790 -370 38835 -250
rect 38955 -370 39000 -250
rect 39120 -370 39165 -250
rect 39285 -370 39340 -250
rect 39460 -370 39505 -250
rect 39625 -370 39670 -250
rect 39790 -370 39835 -250
rect 39955 -370 40010 -250
rect 40130 -370 40175 -250
rect 40295 -370 40340 -250
rect 40460 -370 40505 -250
rect 40625 -370 40680 -250
rect 40800 -370 40845 -250
rect 40965 -370 41010 -250
rect 41130 -370 41175 -250
rect 41295 -370 41350 -250
rect 41470 -370 41515 -250
rect 41635 -370 41680 -250
rect 41800 -370 41845 -250
rect 41965 -370 42175 -250
rect 42295 -370 42350 -250
rect 42470 -370 42515 -250
rect 42635 -370 42680 -250
rect 42800 -370 42845 -250
rect 42965 -370 43020 -250
rect 43140 -370 43185 -250
rect 43305 -370 43350 -250
rect 43470 -370 43515 -250
rect 43635 -370 43690 -250
rect 43810 -370 43855 -250
rect 43975 -370 44020 -250
rect 44140 -370 44185 -250
rect 44305 -370 44360 -250
rect 44480 -370 44525 -250
rect 44645 -370 44690 -250
rect 44810 -370 44855 -250
rect 44975 -370 45030 -250
rect 45150 -370 45195 -250
rect 45315 -370 45360 -250
rect 45480 -370 45525 -250
rect 45645 -370 45700 -250
rect 45820 -370 45865 -250
rect 45985 -370 46030 -250
rect 46150 -370 46195 -250
rect 46315 -370 46370 -250
rect 46490 -370 46535 -250
rect 46655 -370 46700 -250
rect 46820 -370 46865 -250
rect 46985 -370 47040 -250
rect 47160 -370 47205 -250
rect 47325 -370 47370 -250
rect 47490 -370 47535 -250
rect 47655 -370 47865 -250
rect 47985 -370 48040 -250
rect 48160 -370 48205 -250
rect 48325 -370 48370 -250
rect 48490 -370 48535 -250
rect 48655 -370 48710 -250
rect 48830 -370 48875 -250
rect 48995 -370 49040 -250
rect 49160 -370 49205 -250
rect 49325 -370 49380 -250
rect 49500 -370 49545 -250
rect 49665 -370 49710 -250
rect 49830 -370 49875 -250
rect 49995 -370 50050 -250
rect 50170 -370 50215 -250
rect 50335 -370 50380 -250
rect 50500 -370 50545 -250
rect 50665 -370 50720 -250
rect 50840 -370 50885 -250
rect 51005 -370 51050 -250
rect 51170 -370 51215 -250
rect 51335 -370 51390 -250
rect 51510 -370 51555 -250
rect 51675 -370 51720 -250
rect 51840 -370 51885 -250
rect 52005 -370 52060 -250
rect 52180 -370 52225 -250
rect 52345 -370 52390 -250
rect 52510 -370 52555 -250
rect 52675 -370 52730 -250
rect 52850 -370 52895 -250
rect 53015 -370 53060 -250
rect 53180 -370 53225 -250
rect 53345 -370 53370 -250
rect 30770 -415 53370 -370
rect 30770 -535 30795 -415
rect 30915 -535 30970 -415
rect 31090 -535 31135 -415
rect 31255 -535 31300 -415
rect 31420 -535 31465 -415
rect 31585 -535 31640 -415
rect 31760 -535 31805 -415
rect 31925 -535 31970 -415
rect 32090 -535 32135 -415
rect 32255 -535 32310 -415
rect 32430 -535 32475 -415
rect 32595 -535 32640 -415
rect 32760 -535 32805 -415
rect 32925 -535 32980 -415
rect 33100 -535 33145 -415
rect 33265 -535 33310 -415
rect 33430 -535 33475 -415
rect 33595 -535 33650 -415
rect 33770 -535 33815 -415
rect 33935 -535 33980 -415
rect 34100 -535 34145 -415
rect 34265 -535 34320 -415
rect 34440 -535 34485 -415
rect 34605 -535 34650 -415
rect 34770 -535 34815 -415
rect 34935 -535 34990 -415
rect 35110 -535 35155 -415
rect 35275 -535 35320 -415
rect 35440 -535 35485 -415
rect 35605 -535 35660 -415
rect 35780 -535 35825 -415
rect 35945 -535 35990 -415
rect 36110 -535 36155 -415
rect 36275 -535 36485 -415
rect 36605 -535 36660 -415
rect 36780 -535 36825 -415
rect 36945 -535 36990 -415
rect 37110 -535 37155 -415
rect 37275 -535 37330 -415
rect 37450 -535 37495 -415
rect 37615 -535 37660 -415
rect 37780 -535 37825 -415
rect 37945 -535 38000 -415
rect 38120 -535 38165 -415
rect 38285 -535 38330 -415
rect 38450 -535 38495 -415
rect 38615 -535 38670 -415
rect 38790 -535 38835 -415
rect 38955 -535 39000 -415
rect 39120 -535 39165 -415
rect 39285 -535 39340 -415
rect 39460 -535 39505 -415
rect 39625 -535 39670 -415
rect 39790 -535 39835 -415
rect 39955 -535 40010 -415
rect 40130 -535 40175 -415
rect 40295 -535 40340 -415
rect 40460 -535 40505 -415
rect 40625 -535 40680 -415
rect 40800 -535 40845 -415
rect 40965 -535 41010 -415
rect 41130 -535 41175 -415
rect 41295 -535 41350 -415
rect 41470 -535 41515 -415
rect 41635 -535 41680 -415
rect 41800 -535 41845 -415
rect 41965 -535 42175 -415
rect 42295 -535 42350 -415
rect 42470 -535 42515 -415
rect 42635 -535 42680 -415
rect 42800 -535 42845 -415
rect 42965 -535 43020 -415
rect 43140 -535 43185 -415
rect 43305 -535 43350 -415
rect 43470 -535 43515 -415
rect 43635 -535 43690 -415
rect 43810 -535 43855 -415
rect 43975 -535 44020 -415
rect 44140 -535 44185 -415
rect 44305 -535 44360 -415
rect 44480 -535 44525 -415
rect 44645 -535 44690 -415
rect 44810 -535 44855 -415
rect 44975 -535 45030 -415
rect 45150 -535 45195 -415
rect 45315 -535 45360 -415
rect 45480 -535 45525 -415
rect 45645 -535 45700 -415
rect 45820 -535 45865 -415
rect 45985 -535 46030 -415
rect 46150 -535 46195 -415
rect 46315 -535 46370 -415
rect 46490 -535 46535 -415
rect 46655 -535 46700 -415
rect 46820 -535 46865 -415
rect 46985 -535 47040 -415
rect 47160 -535 47205 -415
rect 47325 -535 47370 -415
rect 47490 -535 47535 -415
rect 47655 -535 47865 -415
rect 47985 -535 48040 -415
rect 48160 -535 48205 -415
rect 48325 -535 48370 -415
rect 48490 -535 48535 -415
rect 48655 -535 48710 -415
rect 48830 -535 48875 -415
rect 48995 -535 49040 -415
rect 49160 -535 49205 -415
rect 49325 -535 49380 -415
rect 49500 -535 49545 -415
rect 49665 -535 49710 -415
rect 49830 -535 49875 -415
rect 49995 -535 50050 -415
rect 50170 -535 50215 -415
rect 50335 -535 50380 -415
rect 50500 -535 50545 -415
rect 50665 -535 50720 -415
rect 50840 -535 50885 -415
rect 51005 -535 51050 -415
rect 51170 -535 51215 -415
rect 51335 -535 51390 -415
rect 51510 -535 51555 -415
rect 51675 -535 51720 -415
rect 51840 -535 51885 -415
rect 52005 -535 52060 -415
rect 52180 -535 52225 -415
rect 52345 -535 52390 -415
rect 52510 -535 52555 -415
rect 52675 -535 52730 -415
rect 52850 -535 52895 -415
rect 53015 -535 53060 -415
rect 53180 -535 53225 -415
rect 53345 -535 53370 -415
rect 30770 -590 53370 -535
rect 30770 -710 30795 -590
rect 30915 -710 30970 -590
rect 31090 -710 31135 -590
rect 31255 -710 31300 -590
rect 31420 -710 31465 -590
rect 31585 -710 31640 -590
rect 31760 -710 31805 -590
rect 31925 -710 31970 -590
rect 32090 -710 32135 -590
rect 32255 -710 32310 -590
rect 32430 -710 32475 -590
rect 32595 -710 32640 -590
rect 32760 -710 32805 -590
rect 32925 -710 32980 -590
rect 33100 -710 33145 -590
rect 33265 -710 33310 -590
rect 33430 -710 33475 -590
rect 33595 -710 33650 -590
rect 33770 -710 33815 -590
rect 33935 -710 33980 -590
rect 34100 -710 34145 -590
rect 34265 -710 34320 -590
rect 34440 -710 34485 -590
rect 34605 -710 34650 -590
rect 34770 -710 34815 -590
rect 34935 -710 34990 -590
rect 35110 -710 35155 -590
rect 35275 -710 35320 -590
rect 35440 -710 35485 -590
rect 35605 -710 35660 -590
rect 35780 -710 35825 -590
rect 35945 -710 35990 -590
rect 36110 -710 36155 -590
rect 36275 -710 36485 -590
rect 36605 -710 36660 -590
rect 36780 -710 36825 -590
rect 36945 -710 36990 -590
rect 37110 -710 37155 -590
rect 37275 -710 37330 -590
rect 37450 -710 37495 -590
rect 37615 -710 37660 -590
rect 37780 -710 37825 -590
rect 37945 -710 38000 -590
rect 38120 -710 38165 -590
rect 38285 -710 38330 -590
rect 38450 -710 38495 -590
rect 38615 -710 38670 -590
rect 38790 -710 38835 -590
rect 38955 -710 39000 -590
rect 39120 -710 39165 -590
rect 39285 -710 39340 -590
rect 39460 -710 39505 -590
rect 39625 -710 39670 -590
rect 39790 -710 39835 -590
rect 39955 -710 40010 -590
rect 40130 -710 40175 -590
rect 40295 -710 40340 -590
rect 40460 -710 40505 -590
rect 40625 -710 40680 -590
rect 40800 -710 40845 -590
rect 40965 -710 41010 -590
rect 41130 -710 41175 -590
rect 41295 -710 41350 -590
rect 41470 -710 41515 -590
rect 41635 -710 41680 -590
rect 41800 -710 41845 -590
rect 41965 -710 42175 -590
rect 42295 -710 42350 -590
rect 42470 -710 42515 -590
rect 42635 -710 42680 -590
rect 42800 -710 42845 -590
rect 42965 -710 43020 -590
rect 43140 -710 43185 -590
rect 43305 -710 43350 -590
rect 43470 -710 43515 -590
rect 43635 -710 43690 -590
rect 43810 -710 43855 -590
rect 43975 -710 44020 -590
rect 44140 -710 44185 -590
rect 44305 -710 44360 -590
rect 44480 -710 44525 -590
rect 44645 -710 44690 -590
rect 44810 -710 44855 -590
rect 44975 -710 45030 -590
rect 45150 -710 45195 -590
rect 45315 -710 45360 -590
rect 45480 -710 45525 -590
rect 45645 -710 45700 -590
rect 45820 -710 45865 -590
rect 45985 -710 46030 -590
rect 46150 -710 46195 -590
rect 46315 -710 46370 -590
rect 46490 -710 46535 -590
rect 46655 -710 46700 -590
rect 46820 -710 46865 -590
rect 46985 -710 47040 -590
rect 47160 -710 47205 -590
rect 47325 -710 47370 -590
rect 47490 -710 47535 -590
rect 47655 -710 47865 -590
rect 47985 -710 48040 -590
rect 48160 -710 48205 -590
rect 48325 -710 48370 -590
rect 48490 -710 48535 -590
rect 48655 -710 48710 -590
rect 48830 -710 48875 -590
rect 48995 -710 49040 -590
rect 49160 -710 49205 -590
rect 49325 -710 49380 -590
rect 49500 -710 49545 -590
rect 49665 -710 49710 -590
rect 49830 -710 49875 -590
rect 49995 -710 50050 -590
rect 50170 -710 50215 -590
rect 50335 -710 50380 -590
rect 50500 -710 50545 -590
rect 50665 -710 50720 -590
rect 50840 -710 50885 -590
rect 51005 -710 51050 -590
rect 51170 -710 51215 -590
rect 51335 -710 51390 -590
rect 51510 -710 51555 -590
rect 51675 -710 51720 -590
rect 51840 -710 51885 -590
rect 52005 -710 52060 -590
rect 52180 -710 52225 -590
rect 52345 -710 52390 -590
rect 52510 -710 52555 -590
rect 52675 -710 52730 -590
rect 52850 -710 52895 -590
rect 53015 -710 53060 -590
rect 53180 -710 53225 -590
rect 53345 -710 53370 -590
rect 30770 -755 53370 -710
rect 30770 -875 30795 -755
rect 30915 -875 30970 -755
rect 31090 -875 31135 -755
rect 31255 -875 31300 -755
rect 31420 -875 31465 -755
rect 31585 -875 31640 -755
rect 31760 -875 31805 -755
rect 31925 -875 31970 -755
rect 32090 -875 32135 -755
rect 32255 -875 32310 -755
rect 32430 -875 32475 -755
rect 32595 -875 32640 -755
rect 32760 -875 32805 -755
rect 32925 -875 32980 -755
rect 33100 -875 33145 -755
rect 33265 -875 33310 -755
rect 33430 -875 33475 -755
rect 33595 -875 33650 -755
rect 33770 -875 33815 -755
rect 33935 -875 33980 -755
rect 34100 -875 34145 -755
rect 34265 -875 34320 -755
rect 34440 -875 34485 -755
rect 34605 -875 34650 -755
rect 34770 -875 34815 -755
rect 34935 -875 34990 -755
rect 35110 -875 35155 -755
rect 35275 -875 35320 -755
rect 35440 -875 35485 -755
rect 35605 -875 35660 -755
rect 35780 -875 35825 -755
rect 35945 -875 35990 -755
rect 36110 -875 36155 -755
rect 36275 -875 36485 -755
rect 36605 -875 36660 -755
rect 36780 -875 36825 -755
rect 36945 -875 36990 -755
rect 37110 -875 37155 -755
rect 37275 -875 37330 -755
rect 37450 -875 37495 -755
rect 37615 -875 37660 -755
rect 37780 -875 37825 -755
rect 37945 -875 38000 -755
rect 38120 -875 38165 -755
rect 38285 -875 38330 -755
rect 38450 -875 38495 -755
rect 38615 -875 38670 -755
rect 38790 -875 38835 -755
rect 38955 -875 39000 -755
rect 39120 -875 39165 -755
rect 39285 -875 39340 -755
rect 39460 -875 39505 -755
rect 39625 -875 39670 -755
rect 39790 -875 39835 -755
rect 39955 -875 40010 -755
rect 40130 -875 40175 -755
rect 40295 -875 40340 -755
rect 40460 -875 40505 -755
rect 40625 -875 40680 -755
rect 40800 -875 40845 -755
rect 40965 -875 41010 -755
rect 41130 -875 41175 -755
rect 41295 -875 41350 -755
rect 41470 -875 41515 -755
rect 41635 -875 41680 -755
rect 41800 -875 41845 -755
rect 41965 -875 42175 -755
rect 42295 -875 42350 -755
rect 42470 -875 42515 -755
rect 42635 -875 42680 -755
rect 42800 -875 42845 -755
rect 42965 -875 43020 -755
rect 43140 -875 43185 -755
rect 43305 -875 43350 -755
rect 43470 -875 43515 -755
rect 43635 -875 43690 -755
rect 43810 -875 43855 -755
rect 43975 -875 44020 -755
rect 44140 -875 44185 -755
rect 44305 -875 44360 -755
rect 44480 -875 44525 -755
rect 44645 -875 44690 -755
rect 44810 -875 44855 -755
rect 44975 -875 45030 -755
rect 45150 -875 45195 -755
rect 45315 -875 45360 -755
rect 45480 -875 45525 -755
rect 45645 -875 45700 -755
rect 45820 -875 45865 -755
rect 45985 -875 46030 -755
rect 46150 -875 46195 -755
rect 46315 -875 46370 -755
rect 46490 -875 46535 -755
rect 46655 -875 46700 -755
rect 46820 -875 46865 -755
rect 46985 -875 47040 -755
rect 47160 -875 47205 -755
rect 47325 -875 47370 -755
rect 47490 -875 47535 -755
rect 47655 -875 47865 -755
rect 47985 -875 48040 -755
rect 48160 -875 48205 -755
rect 48325 -875 48370 -755
rect 48490 -875 48535 -755
rect 48655 -875 48710 -755
rect 48830 -875 48875 -755
rect 48995 -875 49040 -755
rect 49160 -875 49205 -755
rect 49325 -875 49380 -755
rect 49500 -875 49545 -755
rect 49665 -875 49710 -755
rect 49830 -875 49875 -755
rect 49995 -875 50050 -755
rect 50170 -875 50215 -755
rect 50335 -875 50380 -755
rect 50500 -875 50545 -755
rect 50665 -875 50720 -755
rect 50840 -875 50885 -755
rect 51005 -875 51050 -755
rect 51170 -875 51215 -755
rect 51335 -875 51390 -755
rect 51510 -875 51555 -755
rect 51675 -875 51720 -755
rect 51840 -875 51885 -755
rect 52005 -875 52060 -755
rect 52180 -875 52225 -755
rect 52345 -875 52390 -755
rect 52510 -875 52555 -755
rect 52675 -875 52730 -755
rect 52850 -875 52895 -755
rect 53015 -875 53060 -755
rect 53180 -875 53225 -755
rect 53345 -875 53370 -755
rect 30770 -920 53370 -875
rect 30770 -1040 30795 -920
rect 30915 -1040 30970 -920
rect 31090 -1040 31135 -920
rect 31255 -1040 31300 -920
rect 31420 -1040 31465 -920
rect 31585 -1040 31640 -920
rect 31760 -1040 31805 -920
rect 31925 -1040 31970 -920
rect 32090 -1040 32135 -920
rect 32255 -1040 32310 -920
rect 32430 -1040 32475 -920
rect 32595 -1040 32640 -920
rect 32760 -1040 32805 -920
rect 32925 -1040 32980 -920
rect 33100 -1040 33145 -920
rect 33265 -1040 33310 -920
rect 33430 -1040 33475 -920
rect 33595 -1040 33650 -920
rect 33770 -1040 33815 -920
rect 33935 -1040 33980 -920
rect 34100 -1040 34145 -920
rect 34265 -1040 34320 -920
rect 34440 -1040 34485 -920
rect 34605 -1040 34650 -920
rect 34770 -1040 34815 -920
rect 34935 -1040 34990 -920
rect 35110 -1040 35155 -920
rect 35275 -1040 35320 -920
rect 35440 -1040 35485 -920
rect 35605 -1040 35660 -920
rect 35780 -1040 35825 -920
rect 35945 -1040 35990 -920
rect 36110 -1040 36155 -920
rect 36275 -1040 36485 -920
rect 36605 -1040 36660 -920
rect 36780 -1040 36825 -920
rect 36945 -1040 36990 -920
rect 37110 -1040 37155 -920
rect 37275 -1040 37330 -920
rect 37450 -1040 37495 -920
rect 37615 -1040 37660 -920
rect 37780 -1040 37825 -920
rect 37945 -1040 38000 -920
rect 38120 -1040 38165 -920
rect 38285 -1040 38330 -920
rect 38450 -1040 38495 -920
rect 38615 -1040 38670 -920
rect 38790 -1040 38835 -920
rect 38955 -1040 39000 -920
rect 39120 -1040 39165 -920
rect 39285 -1040 39340 -920
rect 39460 -1040 39505 -920
rect 39625 -1040 39670 -920
rect 39790 -1040 39835 -920
rect 39955 -1040 40010 -920
rect 40130 -1040 40175 -920
rect 40295 -1040 40340 -920
rect 40460 -1040 40505 -920
rect 40625 -1040 40680 -920
rect 40800 -1040 40845 -920
rect 40965 -1040 41010 -920
rect 41130 -1040 41175 -920
rect 41295 -1040 41350 -920
rect 41470 -1040 41515 -920
rect 41635 -1040 41680 -920
rect 41800 -1040 41845 -920
rect 41965 -1040 42175 -920
rect 42295 -1040 42350 -920
rect 42470 -1040 42515 -920
rect 42635 -1040 42680 -920
rect 42800 -1040 42845 -920
rect 42965 -1040 43020 -920
rect 43140 -1040 43185 -920
rect 43305 -1040 43350 -920
rect 43470 -1040 43515 -920
rect 43635 -1040 43690 -920
rect 43810 -1040 43855 -920
rect 43975 -1040 44020 -920
rect 44140 -1040 44185 -920
rect 44305 -1040 44360 -920
rect 44480 -1040 44525 -920
rect 44645 -1040 44690 -920
rect 44810 -1040 44855 -920
rect 44975 -1040 45030 -920
rect 45150 -1040 45195 -920
rect 45315 -1040 45360 -920
rect 45480 -1040 45525 -920
rect 45645 -1040 45700 -920
rect 45820 -1040 45865 -920
rect 45985 -1040 46030 -920
rect 46150 -1040 46195 -920
rect 46315 -1040 46370 -920
rect 46490 -1040 46535 -920
rect 46655 -1040 46700 -920
rect 46820 -1040 46865 -920
rect 46985 -1040 47040 -920
rect 47160 -1040 47205 -920
rect 47325 -1040 47370 -920
rect 47490 -1040 47535 -920
rect 47655 -1040 47865 -920
rect 47985 -1040 48040 -920
rect 48160 -1040 48205 -920
rect 48325 -1040 48370 -920
rect 48490 -1040 48535 -920
rect 48655 -1040 48710 -920
rect 48830 -1040 48875 -920
rect 48995 -1040 49040 -920
rect 49160 -1040 49205 -920
rect 49325 -1040 49380 -920
rect 49500 -1040 49545 -920
rect 49665 -1040 49710 -920
rect 49830 -1040 49875 -920
rect 49995 -1040 50050 -920
rect 50170 -1040 50215 -920
rect 50335 -1040 50380 -920
rect 50500 -1040 50545 -920
rect 50665 -1040 50720 -920
rect 50840 -1040 50885 -920
rect 51005 -1040 51050 -920
rect 51170 -1040 51215 -920
rect 51335 -1040 51390 -920
rect 51510 -1040 51555 -920
rect 51675 -1040 51720 -920
rect 51840 -1040 51885 -920
rect 52005 -1040 52060 -920
rect 52180 -1040 52225 -920
rect 52345 -1040 52390 -920
rect 52510 -1040 52555 -920
rect 52675 -1040 52730 -920
rect 52850 -1040 52895 -920
rect 53015 -1040 53060 -920
rect 53180 -1040 53225 -920
rect 53345 -1040 53370 -920
rect 30770 -1085 53370 -1040
rect 30770 -1205 30795 -1085
rect 30915 -1205 30970 -1085
rect 31090 -1205 31135 -1085
rect 31255 -1205 31300 -1085
rect 31420 -1205 31465 -1085
rect 31585 -1205 31640 -1085
rect 31760 -1205 31805 -1085
rect 31925 -1205 31970 -1085
rect 32090 -1205 32135 -1085
rect 32255 -1205 32310 -1085
rect 32430 -1205 32475 -1085
rect 32595 -1205 32640 -1085
rect 32760 -1205 32805 -1085
rect 32925 -1205 32980 -1085
rect 33100 -1205 33145 -1085
rect 33265 -1205 33310 -1085
rect 33430 -1205 33475 -1085
rect 33595 -1205 33650 -1085
rect 33770 -1205 33815 -1085
rect 33935 -1205 33980 -1085
rect 34100 -1205 34145 -1085
rect 34265 -1205 34320 -1085
rect 34440 -1205 34485 -1085
rect 34605 -1205 34650 -1085
rect 34770 -1205 34815 -1085
rect 34935 -1205 34990 -1085
rect 35110 -1205 35155 -1085
rect 35275 -1205 35320 -1085
rect 35440 -1205 35485 -1085
rect 35605 -1205 35660 -1085
rect 35780 -1205 35825 -1085
rect 35945 -1205 35990 -1085
rect 36110 -1205 36155 -1085
rect 36275 -1205 36485 -1085
rect 36605 -1205 36660 -1085
rect 36780 -1205 36825 -1085
rect 36945 -1205 36990 -1085
rect 37110 -1205 37155 -1085
rect 37275 -1205 37330 -1085
rect 37450 -1205 37495 -1085
rect 37615 -1205 37660 -1085
rect 37780 -1205 37825 -1085
rect 37945 -1205 38000 -1085
rect 38120 -1205 38165 -1085
rect 38285 -1205 38330 -1085
rect 38450 -1205 38495 -1085
rect 38615 -1205 38670 -1085
rect 38790 -1205 38835 -1085
rect 38955 -1205 39000 -1085
rect 39120 -1205 39165 -1085
rect 39285 -1205 39340 -1085
rect 39460 -1205 39505 -1085
rect 39625 -1205 39670 -1085
rect 39790 -1205 39835 -1085
rect 39955 -1205 40010 -1085
rect 40130 -1205 40175 -1085
rect 40295 -1205 40340 -1085
rect 40460 -1205 40505 -1085
rect 40625 -1205 40680 -1085
rect 40800 -1205 40845 -1085
rect 40965 -1205 41010 -1085
rect 41130 -1205 41175 -1085
rect 41295 -1205 41350 -1085
rect 41470 -1205 41515 -1085
rect 41635 -1205 41680 -1085
rect 41800 -1205 41845 -1085
rect 41965 -1205 42175 -1085
rect 42295 -1205 42350 -1085
rect 42470 -1205 42515 -1085
rect 42635 -1205 42680 -1085
rect 42800 -1205 42845 -1085
rect 42965 -1205 43020 -1085
rect 43140 -1205 43185 -1085
rect 43305 -1205 43350 -1085
rect 43470 -1205 43515 -1085
rect 43635 -1205 43690 -1085
rect 43810 -1205 43855 -1085
rect 43975 -1205 44020 -1085
rect 44140 -1205 44185 -1085
rect 44305 -1205 44360 -1085
rect 44480 -1205 44525 -1085
rect 44645 -1205 44690 -1085
rect 44810 -1205 44855 -1085
rect 44975 -1205 45030 -1085
rect 45150 -1205 45195 -1085
rect 45315 -1205 45360 -1085
rect 45480 -1205 45525 -1085
rect 45645 -1205 45700 -1085
rect 45820 -1205 45865 -1085
rect 45985 -1205 46030 -1085
rect 46150 -1205 46195 -1085
rect 46315 -1205 46370 -1085
rect 46490 -1205 46535 -1085
rect 46655 -1205 46700 -1085
rect 46820 -1205 46865 -1085
rect 46985 -1205 47040 -1085
rect 47160 -1205 47205 -1085
rect 47325 -1205 47370 -1085
rect 47490 -1205 47535 -1085
rect 47655 -1205 47865 -1085
rect 47985 -1205 48040 -1085
rect 48160 -1205 48205 -1085
rect 48325 -1205 48370 -1085
rect 48490 -1205 48535 -1085
rect 48655 -1205 48710 -1085
rect 48830 -1205 48875 -1085
rect 48995 -1205 49040 -1085
rect 49160 -1205 49205 -1085
rect 49325 -1205 49380 -1085
rect 49500 -1205 49545 -1085
rect 49665 -1205 49710 -1085
rect 49830 -1205 49875 -1085
rect 49995 -1205 50050 -1085
rect 50170 -1205 50215 -1085
rect 50335 -1205 50380 -1085
rect 50500 -1205 50545 -1085
rect 50665 -1205 50720 -1085
rect 50840 -1205 50885 -1085
rect 51005 -1205 51050 -1085
rect 51170 -1205 51215 -1085
rect 51335 -1205 51390 -1085
rect 51510 -1205 51555 -1085
rect 51675 -1205 51720 -1085
rect 51840 -1205 51885 -1085
rect 52005 -1205 52060 -1085
rect 52180 -1205 52225 -1085
rect 52345 -1205 52390 -1085
rect 52510 -1205 52555 -1085
rect 52675 -1205 52730 -1085
rect 52850 -1205 52895 -1085
rect 53015 -1205 53060 -1085
rect 53180 -1205 53225 -1085
rect 53345 -1205 53370 -1085
rect 30770 -1260 53370 -1205
rect 30770 -1380 30795 -1260
rect 30915 -1380 30970 -1260
rect 31090 -1380 31135 -1260
rect 31255 -1380 31300 -1260
rect 31420 -1380 31465 -1260
rect 31585 -1380 31640 -1260
rect 31760 -1380 31805 -1260
rect 31925 -1380 31970 -1260
rect 32090 -1380 32135 -1260
rect 32255 -1380 32310 -1260
rect 32430 -1380 32475 -1260
rect 32595 -1380 32640 -1260
rect 32760 -1380 32805 -1260
rect 32925 -1380 32980 -1260
rect 33100 -1380 33145 -1260
rect 33265 -1380 33310 -1260
rect 33430 -1380 33475 -1260
rect 33595 -1380 33650 -1260
rect 33770 -1380 33815 -1260
rect 33935 -1380 33980 -1260
rect 34100 -1380 34145 -1260
rect 34265 -1380 34320 -1260
rect 34440 -1380 34485 -1260
rect 34605 -1380 34650 -1260
rect 34770 -1380 34815 -1260
rect 34935 -1380 34990 -1260
rect 35110 -1380 35155 -1260
rect 35275 -1380 35320 -1260
rect 35440 -1380 35485 -1260
rect 35605 -1380 35660 -1260
rect 35780 -1380 35825 -1260
rect 35945 -1380 35990 -1260
rect 36110 -1380 36155 -1260
rect 36275 -1380 36485 -1260
rect 36605 -1380 36660 -1260
rect 36780 -1380 36825 -1260
rect 36945 -1380 36990 -1260
rect 37110 -1380 37155 -1260
rect 37275 -1380 37330 -1260
rect 37450 -1380 37495 -1260
rect 37615 -1380 37660 -1260
rect 37780 -1380 37825 -1260
rect 37945 -1380 38000 -1260
rect 38120 -1380 38165 -1260
rect 38285 -1380 38330 -1260
rect 38450 -1380 38495 -1260
rect 38615 -1380 38670 -1260
rect 38790 -1380 38835 -1260
rect 38955 -1380 39000 -1260
rect 39120 -1380 39165 -1260
rect 39285 -1380 39340 -1260
rect 39460 -1380 39505 -1260
rect 39625 -1380 39670 -1260
rect 39790 -1380 39835 -1260
rect 39955 -1380 40010 -1260
rect 40130 -1380 40175 -1260
rect 40295 -1380 40340 -1260
rect 40460 -1380 40505 -1260
rect 40625 -1380 40680 -1260
rect 40800 -1380 40845 -1260
rect 40965 -1380 41010 -1260
rect 41130 -1380 41175 -1260
rect 41295 -1380 41350 -1260
rect 41470 -1380 41515 -1260
rect 41635 -1380 41680 -1260
rect 41800 -1380 41845 -1260
rect 41965 -1380 42175 -1260
rect 42295 -1380 42350 -1260
rect 42470 -1380 42515 -1260
rect 42635 -1380 42680 -1260
rect 42800 -1380 42845 -1260
rect 42965 -1380 43020 -1260
rect 43140 -1380 43185 -1260
rect 43305 -1380 43350 -1260
rect 43470 -1380 43515 -1260
rect 43635 -1380 43690 -1260
rect 43810 -1380 43855 -1260
rect 43975 -1380 44020 -1260
rect 44140 -1380 44185 -1260
rect 44305 -1380 44360 -1260
rect 44480 -1380 44525 -1260
rect 44645 -1380 44690 -1260
rect 44810 -1380 44855 -1260
rect 44975 -1380 45030 -1260
rect 45150 -1380 45195 -1260
rect 45315 -1380 45360 -1260
rect 45480 -1380 45525 -1260
rect 45645 -1380 45700 -1260
rect 45820 -1380 45865 -1260
rect 45985 -1380 46030 -1260
rect 46150 -1380 46195 -1260
rect 46315 -1380 46370 -1260
rect 46490 -1380 46535 -1260
rect 46655 -1380 46700 -1260
rect 46820 -1380 46865 -1260
rect 46985 -1380 47040 -1260
rect 47160 -1380 47205 -1260
rect 47325 -1380 47370 -1260
rect 47490 -1380 47535 -1260
rect 47655 -1380 47865 -1260
rect 47985 -1380 48040 -1260
rect 48160 -1380 48205 -1260
rect 48325 -1380 48370 -1260
rect 48490 -1380 48535 -1260
rect 48655 -1380 48710 -1260
rect 48830 -1380 48875 -1260
rect 48995 -1380 49040 -1260
rect 49160 -1380 49205 -1260
rect 49325 -1380 49380 -1260
rect 49500 -1380 49545 -1260
rect 49665 -1380 49710 -1260
rect 49830 -1380 49875 -1260
rect 49995 -1380 50050 -1260
rect 50170 -1380 50215 -1260
rect 50335 -1380 50380 -1260
rect 50500 -1380 50545 -1260
rect 50665 -1380 50720 -1260
rect 50840 -1380 50885 -1260
rect 51005 -1380 51050 -1260
rect 51170 -1380 51215 -1260
rect 51335 -1380 51390 -1260
rect 51510 -1380 51555 -1260
rect 51675 -1380 51720 -1260
rect 51840 -1380 51885 -1260
rect 52005 -1380 52060 -1260
rect 52180 -1380 52225 -1260
rect 52345 -1380 52390 -1260
rect 52510 -1380 52555 -1260
rect 52675 -1380 52730 -1260
rect 52850 -1380 52895 -1260
rect 53015 -1380 53060 -1260
rect 53180 -1380 53225 -1260
rect 53345 -1380 53370 -1260
rect 30770 -1425 53370 -1380
rect 30770 -1545 30795 -1425
rect 30915 -1545 30970 -1425
rect 31090 -1545 31135 -1425
rect 31255 -1545 31300 -1425
rect 31420 -1545 31465 -1425
rect 31585 -1545 31640 -1425
rect 31760 -1545 31805 -1425
rect 31925 -1545 31970 -1425
rect 32090 -1545 32135 -1425
rect 32255 -1545 32310 -1425
rect 32430 -1545 32475 -1425
rect 32595 -1545 32640 -1425
rect 32760 -1545 32805 -1425
rect 32925 -1545 32980 -1425
rect 33100 -1545 33145 -1425
rect 33265 -1545 33310 -1425
rect 33430 -1545 33475 -1425
rect 33595 -1545 33650 -1425
rect 33770 -1545 33815 -1425
rect 33935 -1545 33980 -1425
rect 34100 -1545 34145 -1425
rect 34265 -1545 34320 -1425
rect 34440 -1545 34485 -1425
rect 34605 -1545 34650 -1425
rect 34770 -1545 34815 -1425
rect 34935 -1545 34990 -1425
rect 35110 -1545 35155 -1425
rect 35275 -1545 35320 -1425
rect 35440 -1545 35485 -1425
rect 35605 -1545 35660 -1425
rect 35780 -1545 35825 -1425
rect 35945 -1545 35990 -1425
rect 36110 -1545 36155 -1425
rect 36275 -1545 36485 -1425
rect 36605 -1545 36660 -1425
rect 36780 -1545 36825 -1425
rect 36945 -1545 36990 -1425
rect 37110 -1545 37155 -1425
rect 37275 -1545 37330 -1425
rect 37450 -1545 37495 -1425
rect 37615 -1545 37660 -1425
rect 37780 -1545 37825 -1425
rect 37945 -1545 38000 -1425
rect 38120 -1545 38165 -1425
rect 38285 -1545 38330 -1425
rect 38450 -1545 38495 -1425
rect 38615 -1545 38670 -1425
rect 38790 -1545 38835 -1425
rect 38955 -1545 39000 -1425
rect 39120 -1545 39165 -1425
rect 39285 -1545 39340 -1425
rect 39460 -1545 39505 -1425
rect 39625 -1545 39670 -1425
rect 39790 -1545 39835 -1425
rect 39955 -1545 40010 -1425
rect 40130 -1545 40175 -1425
rect 40295 -1545 40340 -1425
rect 40460 -1545 40505 -1425
rect 40625 -1545 40680 -1425
rect 40800 -1545 40845 -1425
rect 40965 -1545 41010 -1425
rect 41130 -1545 41175 -1425
rect 41295 -1545 41350 -1425
rect 41470 -1545 41515 -1425
rect 41635 -1545 41680 -1425
rect 41800 -1545 41845 -1425
rect 41965 -1545 42175 -1425
rect 42295 -1545 42350 -1425
rect 42470 -1545 42515 -1425
rect 42635 -1545 42680 -1425
rect 42800 -1545 42845 -1425
rect 42965 -1545 43020 -1425
rect 43140 -1545 43185 -1425
rect 43305 -1545 43350 -1425
rect 43470 -1545 43515 -1425
rect 43635 -1545 43690 -1425
rect 43810 -1545 43855 -1425
rect 43975 -1545 44020 -1425
rect 44140 -1545 44185 -1425
rect 44305 -1545 44360 -1425
rect 44480 -1545 44525 -1425
rect 44645 -1545 44690 -1425
rect 44810 -1545 44855 -1425
rect 44975 -1545 45030 -1425
rect 45150 -1545 45195 -1425
rect 45315 -1545 45360 -1425
rect 45480 -1545 45525 -1425
rect 45645 -1545 45700 -1425
rect 45820 -1545 45865 -1425
rect 45985 -1545 46030 -1425
rect 46150 -1545 46195 -1425
rect 46315 -1545 46370 -1425
rect 46490 -1545 46535 -1425
rect 46655 -1545 46700 -1425
rect 46820 -1545 46865 -1425
rect 46985 -1545 47040 -1425
rect 47160 -1545 47205 -1425
rect 47325 -1545 47370 -1425
rect 47490 -1545 47535 -1425
rect 47655 -1545 47865 -1425
rect 47985 -1545 48040 -1425
rect 48160 -1545 48205 -1425
rect 48325 -1545 48370 -1425
rect 48490 -1545 48535 -1425
rect 48655 -1545 48710 -1425
rect 48830 -1545 48875 -1425
rect 48995 -1545 49040 -1425
rect 49160 -1545 49205 -1425
rect 49325 -1545 49380 -1425
rect 49500 -1545 49545 -1425
rect 49665 -1545 49710 -1425
rect 49830 -1545 49875 -1425
rect 49995 -1545 50050 -1425
rect 50170 -1545 50215 -1425
rect 50335 -1545 50380 -1425
rect 50500 -1545 50545 -1425
rect 50665 -1545 50720 -1425
rect 50840 -1545 50885 -1425
rect 51005 -1545 51050 -1425
rect 51170 -1545 51215 -1425
rect 51335 -1545 51390 -1425
rect 51510 -1545 51555 -1425
rect 51675 -1545 51720 -1425
rect 51840 -1545 51885 -1425
rect 52005 -1545 52060 -1425
rect 52180 -1545 52225 -1425
rect 52345 -1545 52390 -1425
rect 52510 -1545 52555 -1425
rect 52675 -1545 52730 -1425
rect 52850 -1545 52895 -1425
rect 53015 -1545 53060 -1425
rect 53180 -1545 53225 -1425
rect 53345 -1545 53370 -1425
rect 30770 -1590 53370 -1545
rect 30770 -1710 30795 -1590
rect 30915 -1710 30970 -1590
rect 31090 -1710 31135 -1590
rect 31255 -1710 31300 -1590
rect 31420 -1710 31465 -1590
rect 31585 -1710 31640 -1590
rect 31760 -1710 31805 -1590
rect 31925 -1710 31970 -1590
rect 32090 -1710 32135 -1590
rect 32255 -1710 32310 -1590
rect 32430 -1710 32475 -1590
rect 32595 -1710 32640 -1590
rect 32760 -1710 32805 -1590
rect 32925 -1710 32980 -1590
rect 33100 -1710 33145 -1590
rect 33265 -1710 33310 -1590
rect 33430 -1710 33475 -1590
rect 33595 -1710 33650 -1590
rect 33770 -1710 33815 -1590
rect 33935 -1710 33980 -1590
rect 34100 -1710 34145 -1590
rect 34265 -1710 34320 -1590
rect 34440 -1710 34485 -1590
rect 34605 -1710 34650 -1590
rect 34770 -1710 34815 -1590
rect 34935 -1710 34990 -1590
rect 35110 -1710 35155 -1590
rect 35275 -1710 35320 -1590
rect 35440 -1710 35485 -1590
rect 35605 -1710 35660 -1590
rect 35780 -1710 35825 -1590
rect 35945 -1710 35990 -1590
rect 36110 -1710 36155 -1590
rect 36275 -1710 36485 -1590
rect 36605 -1710 36660 -1590
rect 36780 -1710 36825 -1590
rect 36945 -1710 36990 -1590
rect 37110 -1710 37155 -1590
rect 37275 -1710 37330 -1590
rect 37450 -1710 37495 -1590
rect 37615 -1710 37660 -1590
rect 37780 -1710 37825 -1590
rect 37945 -1710 38000 -1590
rect 38120 -1710 38165 -1590
rect 38285 -1710 38330 -1590
rect 38450 -1710 38495 -1590
rect 38615 -1710 38670 -1590
rect 38790 -1710 38835 -1590
rect 38955 -1710 39000 -1590
rect 39120 -1710 39165 -1590
rect 39285 -1710 39340 -1590
rect 39460 -1710 39505 -1590
rect 39625 -1710 39670 -1590
rect 39790 -1710 39835 -1590
rect 39955 -1710 40010 -1590
rect 40130 -1710 40175 -1590
rect 40295 -1710 40340 -1590
rect 40460 -1710 40505 -1590
rect 40625 -1710 40680 -1590
rect 40800 -1710 40845 -1590
rect 40965 -1710 41010 -1590
rect 41130 -1710 41175 -1590
rect 41295 -1710 41350 -1590
rect 41470 -1710 41515 -1590
rect 41635 -1710 41680 -1590
rect 41800 -1710 41845 -1590
rect 41965 -1710 42175 -1590
rect 42295 -1710 42350 -1590
rect 42470 -1710 42515 -1590
rect 42635 -1710 42680 -1590
rect 42800 -1710 42845 -1590
rect 42965 -1710 43020 -1590
rect 43140 -1710 43185 -1590
rect 43305 -1710 43350 -1590
rect 43470 -1710 43515 -1590
rect 43635 -1710 43690 -1590
rect 43810 -1710 43855 -1590
rect 43975 -1710 44020 -1590
rect 44140 -1710 44185 -1590
rect 44305 -1710 44360 -1590
rect 44480 -1710 44525 -1590
rect 44645 -1710 44690 -1590
rect 44810 -1710 44855 -1590
rect 44975 -1710 45030 -1590
rect 45150 -1710 45195 -1590
rect 45315 -1710 45360 -1590
rect 45480 -1710 45525 -1590
rect 45645 -1710 45700 -1590
rect 45820 -1710 45865 -1590
rect 45985 -1710 46030 -1590
rect 46150 -1710 46195 -1590
rect 46315 -1710 46370 -1590
rect 46490 -1710 46535 -1590
rect 46655 -1710 46700 -1590
rect 46820 -1710 46865 -1590
rect 46985 -1710 47040 -1590
rect 47160 -1710 47205 -1590
rect 47325 -1710 47370 -1590
rect 47490 -1710 47535 -1590
rect 47655 -1710 47865 -1590
rect 47985 -1710 48040 -1590
rect 48160 -1710 48205 -1590
rect 48325 -1710 48370 -1590
rect 48490 -1710 48535 -1590
rect 48655 -1710 48710 -1590
rect 48830 -1710 48875 -1590
rect 48995 -1710 49040 -1590
rect 49160 -1710 49205 -1590
rect 49325 -1710 49380 -1590
rect 49500 -1710 49545 -1590
rect 49665 -1710 49710 -1590
rect 49830 -1710 49875 -1590
rect 49995 -1710 50050 -1590
rect 50170 -1710 50215 -1590
rect 50335 -1710 50380 -1590
rect 50500 -1710 50545 -1590
rect 50665 -1710 50720 -1590
rect 50840 -1710 50885 -1590
rect 51005 -1710 51050 -1590
rect 51170 -1710 51215 -1590
rect 51335 -1710 51390 -1590
rect 51510 -1710 51555 -1590
rect 51675 -1710 51720 -1590
rect 51840 -1710 51885 -1590
rect 52005 -1710 52060 -1590
rect 52180 -1710 52225 -1590
rect 52345 -1710 52390 -1590
rect 52510 -1710 52555 -1590
rect 52675 -1710 52730 -1590
rect 52850 -1710 52895 -1590
rect 53015 -1710 53060 -1590
rect 53180 -1710 53225 -1590
rect 53345 -1710 53370 -1590
rect 30770 -1755 53370 -1710
rect 30770 -1875 30795 -1755
rect 30915 -1875 30970 -1755
rect 31090 -1875 31135 -1755
rect 31255 -1875 31300 -1755
rect 31420 -1875 31465 -1755
rect 31585 -1875 31640 -1755
rect 31760 -1875 31805 -1755
rect 31925 -1875 31970 -1755
rect 32090 -1875 32135 -1755
rect 32255 -1875 32310 -1755
rect 32430 -1875 32475 -1755
rect 32595 -1875 32640 -1755
rect 32760 -1875 32805 -1755
rect 32925 -1875 32980 -1755
rect 33100 -1875 33145 -1755
rect 33265 -1875 33310 -1755
rect 33430 -1875 33475 -1755
rect 33595 -1875 33650 -1755
rect 33770 -1875 33815 -1755
rect 33935 -1875 33980 -1755
rect 34100 -1875 34145 -1755
rect 34265 -1875 34320 -1755
rect 34440 -1875 34485 -1755
rect 34605 -1875 34650 -1755
rect 34770 -1875 34815 -1755
rect 34935 -1875 34990 -1755
rect 35110 -1875 35155 -1755
rect 35275 -1875 35320 -1755
rect 35440 -1875 35485 -1755
rect 35605 -1875 35660 -1755
rect 35780 -1875 35825 -1755
rect 35945 -1875 35990 -1755
rect 36110 -1875 36155 -1755
rect 36275 -1875 36485 -1755
rect 36605 -1875 36660 -1755
rect 36780 -1875 36825 -1755
rect 36945 -1875 36990 -1755
rect 37110 -1875 37155 -1755
rect 37275 -1875 37330 -1755
rect 37450 -1875 37495 -1755
rect 37615 -1875 37660 -1755
rect 37780 -1875 37825 -1755
rect 37945 -1875 38000 -1755
rect 38120 -1875 38165 -1755
rect 38285 -1875 38330 -1755
rect 38450 -1875 38495 -1755
rect 38615 -1875 38670 -1755
rect 38790 -1875 38835 -1755
rect 38955 -1875 39000 -1755
rect 39120 -1875 39165 -1755
rect 39285 -1875 39340 -1755
rect 39460 -1875 39505 -1755
rect 39625 -1875 39670 -1755
rect 39790 -1875 39835 -1755
rect 39955 -1875 40010 -1755
rect 40130 -1875 40175 -1755
rect 40295 -1875 40340 -1755
rect 40460 -1875 40505 -1755
rect 40625 -1875 40680 -1755
rect 40800 -1875 40845 -1755
rect 40965 -1875 41010 -1755
rect 41130 -1875 41175 -1755
rect 41295 -1875 41350 -1755
rect 41470 -1875 41515 -1755
rect 41635 -1875 41680 -1755
rect 41800 -1875 41845 -1755
rect 41965 -1875 42175 -1755
rect 42295 -1875 42350 -1755
rect 42470 -1875 42515 -1755
rect 42635 -1875 42680 -1755
rect 42800 -1875 42845 -1755
rect 42965 -1875 43020 -1755
rect 43140 -1875 43185 -1755
rect 43305 -1875 43350 -1755
rect 43470 -1875 43515 -1755
rect 43635 -1875 43690 -1755
rect 43810 -1875 43855 -1755
rect 43975 -1875 44020 -1755
rect 44140 -1875 44185 -1755
rect 44305 -1875 44360 -1755
rect 44480 -1875 44525 -1755
rect 44645 -1875 44690 -1755
rect 44810 -1875 44855 -1755
rect 44975 -1875 45030 -1755
rect 45150 -1875 45195 -1755
rect 45315 -1875 45360 -1755
rect 45480 -1875 45525 -1755
rect 45645 -1875 45700 -1755
rect 45820 -1875 45865 -1755
rect 45985 -1875 46030 -1755
rect 46150 -1875 46195 -1755
rect 46315 -1875 46370 -1755
rect 46490 -1875 46535 -1755
rect 46655 -1875 46700 -1755
rect 46820 -1875 46865 -1755
rect 46985 -1875 47040 -1755
rect 47160 -1875 47205 -1755
rect 47325 -1875 47370 -1755
rect 47490 -1875 47535 -1755
rect 47655 -1875 47865 -1755
rect 47985 -1875 48040 -1755
rect 48160 -1875 48205 -1755
rect 48325 -1875 48370 -1755
rect 48490 -1875 48535 -1755
rect 48655 -1875 48710 -1755
rect 48830 -1875 48875 -1755
rect 48995 -1875 49040 -1755
rect 49160 -1875 49205 -1755
rect 49325 -1875 49380 -1755
rect 49500 -1875 49545 -1755
rect 49665 -1875 49710 -1755
rect 49830 -1875 49875 -1755
rect 49995 -1875 50050 -1755
rect 50170 -1875 50215 -1755
rect 50335 -1875 50380 -1755
rect 50500 -1875 50545 -1755
rect 50665 -1875 50720 -1755
rect 50840 -1875 50885 -1755
rect 51005 -1875 51050 -1755
rect 51170 -1875 51215 -1755
rect 51335 -1875 51390 -1755
rect 51510 -1875 51555 -1755
rect 51675 -1875 51720 -1755
rect 51840 -1875 51885 -1755
rect 52005 -1875 52060 -1755
rect 52180 -1875 52225 -1755
rect 52345 -1875 52390 -1755
rect 52510 -1875 52555 -1755
rect 52675 -1875 52730 -1755
rect 52850 -1875 52895 -1755
rect 53015 -1875 53060 -1755
rect 53180 -1875 53225 -1755
rect 53345 -1875 53370 -1755
rect 30770 -1930 53370 -1875
rect 30770 -2050 30795 -1930
rect 30915 -2050 30970 -1930
rect 31090 -2050 31135 -1930
rect 31255 -2050 31300 -1930
rect 31420 -2050 31465 -1930
rect 31585 -2050 31640 -1930
rect 31760 -2050 31805 -1930
rect 31925 -2050 31970 -1930
rect 32090 -2050 32135 -1930
rect 32255 -2050 32310 -1930
rect 32430 -2050 32475 -1930
rect 32595 -2050 32640 -1930
rect 32760 -2050 32805 -1930
rect 32925 -2050 32980 -1930
rect 33100 -2050 33145 -1930
rect 33265 -2050 33310 -1930
rect 33430 -2050 33475 -1930
rect 33595 -2050 33650 -1930
rect 33770 -2050 33815 -1930
rect 33935 -2050 33980 -1930
rect 34100 -2050 34145 -1930
rect 34265 -2050 34320 -1930
rect 34440 -2050 34485 -1930
rect 34605 -2050 34650 -1930
rect 34770 -2050 34815 -1930
rect 34935 -2050 34990 -1930
rect 35110 -2050 35155 -1930
rect 35275 -2050 35320 -1930
rect 35440 -2050 35485 -1930
rect 35605 -2050 35660 -1930
rect 35780 -2050 35825 -1930
rect 35945 -2050 35990 -1930
rect 36110 -2050 36155 -1930
rect 36275 -2050 36485 -1930
rect 36605 -2050 36660 -1930
rect 36780 -2050 36825 -1930
rect 36945 -2050 36990 -1930
rect 37110 -2050 37155 -1930
rect 37275 -2050 37330 -1930
rect 37450 -2050 37495 -1930
rect 37615 -2050 37660 -1930
rect 37780 -2050 37825 -1930
rect 37945 -2050 38000 -1930
rect 38120 -2050 38165 -1930
rect 38285 -2050 38330 -1930
rect 38450 -2050 38495 -1930
rect 38615 -2050 38670 -1930
rect 38790 -2050 38835 -1930
rect 38955 -2050 39000 -1930
rect 39120 -2050 39165 -1930
rect 39285 -2050 39340 -1930
rect 39460 -2050 39505 -1930
rect 39625 -2050 39670 -1930
rect 39790 -2050 39835 -1930
rect 39955 -2050 40010 -1930
rect 40130 -2050 40175 -1930
rect 40295 -2050 40340 -1930
rect 40460 -2050 40505 -1930
rect 40625 -2050 40680 -1930
rect 40800 -2050 40845 -1930
rect 40965 -2050 41010 -1930
rect 41130 -2050 41175 -1930
rect 41295 -2050 41350 -1930
rect 41470 -2050 41515 -1930
rect 41635 -2050 41680 -1930
rect 41800 -2050 41845 -1930
rect 41965 -2050 42175 -1930
rect 42295 -2050 42350 -1930
rect 42470 -2050 42515 -1930
rect 42635 -2050 42680 -1930
rect 42800 -2050 42845 -1930
rect 42965 -2050 43020 -1930
rect 43140 -2050 43185 -1930
rect 43305 -2050 43350 -1930
rect 43470 -2050 43515 -1930
rect 43635 -2050 43690 -1930
rect 43810 -2050 43855 -1930
rect 43975 -2050 44020 -1930
rect 44140 -2050 44185 -1930
rect 44305 -2050 44360 -1930
rect 44480 -2050 44525 -1930
rect 44645 -2050 44690 -1930
rect 44810 -2050 44855 -1930
rect 44975 -2050 45030 -1930
rect 45150 -2050 45195 -1930
rect 45315 -2050 45360 -1930
rect 45480 -2050 45525 -1930
rect 45645 -2050 45700 -1930
rect 45820 -2050 45865 -1930
rect 45985 -2050 46030 -1930
rect 46150 -2050 46195 -1930
rect 46315 -2050 46370 -1930
rect 46490 -2050 46535 -1930
rect 46655 -2050 46700 -1930
rect 46820 -2050 46865 -1930
rect 46985 -2050 47040 -1930
rect 47160 -2050 47205 -1930
rect 47325 -2050 47370 -1930
rect 47490 -2050 47535 -1930
rect 47655 -2050 47865 -1930
rect 47985 -2050 48040 -1930
rect 48160 -2050 48205 -1930
rect 48325 -2050 48370 -1930
rect 48490 -2050 48535 -1930
rect 48655 -2050 48710 -1930
rect 48830 -2050 48875 -1930
rect 48995 -2050 49040 -1930
rect 49160 -2050 49205 -1930
rect 49325 -2050 49380 -1930
rect 49500 -2050 49545 -1930
rect 49665 -2050 49710 -1930
rect 49830 -2050 49875 -1930
rect 49995 -2050 50050 -1930
rect 50170 -2050 50215 -1930
rect 50335 -2050 50380 -1930
rect 50500 -2050 50545 -1930
rect 50665 -2050 50720 -1930
rect 50840 -2050 50885 -1930
rect 51005 -2050 51050 -1930
rect 51170 -2050 51215 -1930
rect 51335 -2050 51390 -1930
rect 51510 -2050 51555 -1930
rect 51675 -2050 51720 -1930
rect 51840 -2050 51885 -1930
rect 52005 -2050 52060 -1930
rect 52180 -2050 52225 -1930
rect 52345 -2050 52390 -1930
rect 52510 -2050 52555 -1930
rect 52675 -2050 52730 -1930
rect 52850 -2050 52895 -1930
rect 53015 -2050 53060 -1930
rect 53180 -2050 53225 -1930
rect 53345 -2050 53370 -1930
rect 30770 -2095 53370 -2050
rect 30770 -2215 30795 -2095
rect 30915 -2215 30970 -2095
rect 31090 -2215 31135 -2095
rect 31255 -2215 31300 -2095
rect 31420 -2215 31465 -2095
rect 31585 -2215 31640 -2095
rect 31760 -2215 31805 -2095
rect 31925 -2215 31970 -2095
rect 32090 -2215 32135 -2095
rect 32255 -2215 32310 -2095
rect 32430 -2215 32475 -2095
rect 32595 -2215 32640 -2095
rect 32760 -2215 32805 -2095
rect 32925 -2215 32980 -2095
rect 33100 -2215 33145 -2095
rect 33265 -2215 33310 -2095
rect 33430 -2215 33475 -2095
rect 33595 -2215 33650 -2095
rect 33770 -2215 33815 -2095
rect 33935 -2215 33980 -2095
rect 34100 -2215 34145 -2095
rect 34265 -2215 34320 -2095
rect 34440 -2215 34485 -2095
rect 34605 -2215 34650 -2095
rect 34770 -2215 34815 -2095
rect 34935 -2215 34990 -2095
rect 35110 -2215 35155 -2095
rect 35275 -2215 35320 -2095
rect 35440 -2215 35485 -2095
rect 35605 -2215 35660 -2095
rect 35780 -2215 35825 -2095
rect 35945 -2215 35990 -2095
rect 36110 -2215 36155 -2095
rect 36275 -2215 36485 -2095
rect 36605 -2215 36660 -2095
rect 36780 -2215 36825 -2095
rect 36945 -2215 36990 -2095
rect 37110 -2215 37155 -2095
rect 37275 -2215 37330 -2095
rect 37450 -2215 37495 -2095
rect 37615 -2215 37660 -2095
rect 37780 -2215 37825 -2095
rect 37945 -2215 38000 -2095
rect 38120 -2215 38165 -2095
rect 38285 -2215 38330 -2095
rect 38450 -2215 38495 -2095
rect 38615 -2215 38670 -2095
rect 38790 -2215 38835 -2095
rect 38955 -2215 39000 -2095
rect 39120 -2215 39165 -2095
rect 39285 -2215 39340 -2095
rect 39460 -2215 39505 -2095
rect 39625 -2215 39670 -2095
rect 39790 -2215 39835 -2095
rect 39955 -2215 40010 -2095
rect 40130 -2215 40175 -2095
rect 40295 -2215 40340 -2095
rect 40460 -2215 40505 -2095
rect 40625 -2215 40680 -2095
rect 40800 -2215 40845 -2095
rect 40965 -2215 41010 -2095
rect 41130 -2215 41175 -2095
rect 41295 -2215 41350 -2095
rect 41470 -2215 41515 -2095
rect 41635 -2215 41680 -2095
rect 41800 -2215 41845 -2095
rect 41965 -2215 42175 -2095
rect 42295 -2215 42350 -2095
rect 42470 -2215 42515 -2095
rect 42635 -2215 42680 -2095
rect 42800 -2215 42845 -2095
rect 42965 -2215 43020 -2095
rect 43140 -2215 43185 -2095
rect 43305 -2215 43350 -2095
rect 43470 -2215 43515 -2095
rect 43635 -2215 43690 -2095
rect 43810 -2215 43855 -2095
rect 43975 -2215 44020 -2095
rect 44140 -2215 44185 -2095
rect 44305 -2215 44360 -2095
rect 44480 -2215 44525 -2095
rect 44645 -2215 44690 -2095
rect 44810 -2215 44855 -2095
rect 44975 -2215 45030 -2095
rect 45150 -2215 45195 -2095
rect 45315 -2215 45360 -2095
rect 45480 -2215 45525 -2095
rect 45645 -2215 45700 -2095
rect 45820 -2215 45865 -2095
rect 45985 -2215 46030 -2095
rect 46150 -2215 46195 -2095
rect 46315 -2215 46370 -2095
rect 46490 -2215 46535 -2095
rect 46655 -2215 46700 -2095
rect 46820 -2215 46865 -2095
rect 46985 -2215 47040 -2095
rect 47160 -2215 47205 -2095
rect 47325 -2215 47370 -2095
rect 47490 -2215 47535 -2095
rect 47655 -2215 47865 -2095
rect 47985 -2215 48040 -2095
rect 48160 -2215 48205 -2095
rect 48325 -2215 48370 -2095
rect 48490 -2215 48535 -2095
rect 48655 -2215 48710 -2095
rect 48830 -2215 48875 -2095
rect 48995 -2215 49040 -2095
rect 49160 -2215 49205 -2095
rect 49325 -2215 49380 -2095
rect 49500 -2215 49545 -2095
rect 49665 -2215 49710 -2095
rect 49830 -2215 49875 -2095
rect 49995 -2215 50050 -2095
rect 50170 -2215 50215 -2095
rect 50335 -2215 50380 -2095
rect 50500 -2215 50545 -2095
rect 50665 -2215 50720 -2095
rect 50840 -2215 50885 -2095
rect 51005 -2215 51050 -2095
rect 51170 -2215 51215 -2095
rect 51335 -2215 51390 -2095
rect 51510 -2215 51555 -2095
rect 51675 -2215 51720 -2095
rect 51840 -2215 51885 -2095
rect 52005 -2215 52060 -2095
rect 52180 -2215 52225 -2095
rect 52345 -2215 52390 -2095
rect 52510 -2215 52555 -2095
rect 52675 -2215 52730 -2095
rect 52850 -2215 52895 -2095
rect 53015 -2215 53060 -2095
rect 53180 -2215 53225 -2095
rect 53345 -2215 53370 -2095
rect 30770 -2260 53370 -2215
rect 30770 -2380 30795 -2260
rect 30915 -2380 30970 -2260
rect 31090 -2380 31135 -2260
rect 31255 -2380 31300 -2260
rect 31420 -2380 31465 -2260
rect 31585 -2380 31640 -2260
rect 31760 -2380 31805 -2260
rect 31925 -2380 31970 -2260
rect 32090 -2380 32135 -2260
rect 32255 -2380 32310 -2260
rect 32430 -2380 32475 -2260
rect 32595 -2380 32640 -2260
rect 32760 -2380 32805 -2260
rect 32925 -2380 32980 -2260
rect 33100 -2380 33145 -2260
rect 33265 -2380 33310 -2260
rect 33430 -2380 33475 -2260
rect 33595 -2380 33650 -2260
rect 33770 -2380 33815 -2260
rect 33935 -2380 33980 -2260
rect 34100 -2380 34145 -2260
rect 34265 -2380 34320 -2260
rect 34440 -2380 34485 -2260
rect 34605 -2380 34650 -2260
rect 34770 -2380 34815 -2260
rect 34935 -2380 34990 -2260
rect 35110 -2380 35155 -2260
rect 35275 -2380 35320 -2260
rect 35440 -2380 35485 -2260
rect 35605 -2380 35660 -2260
rect 35780 -2380 35825 -2260
rect 35945 -2380 35990 -2260
rect 36110 -2380 36155 -2260
rect 36275 -2380 36485 -2260
rect 36605 -2380 36660 -2260
rect 36780 -2380 36825 -2260
rect 36945 -2380 36990 -2260
rect 37110 -2380 37155 -2260
rect 37275 -2380 37330 -2260
rect 37450 -2380 37495 -2260
rect 37615 -2380 37660 -2260
rect 37780 -2380 37825 -2260
rect 37945 -2380 38000 -2260
rect 38120 -2380 38165 -2260
rect 38285 -2380 38330 -2260
rect 38450 -2380 38495 -2260
rect 38615 -2380 38670 -2260
rect 38790 -2380 38835 -2260
rect 38955 -2380 39000 -2260
rect 39120 -2380 39165 -2260
rect 39285 -2380 39340 -2260
rect 39460 -2380 39505 -2260
rect 39625 -2380 39670 -2260
rect 39790 -2380 39835 -2260
rect 39955 -2380 40010 -2260
rect 40130 -2380 40175 -2260
rect 40295 -2380 40340 -2260
rect 40460 -2380 40505 -2260
rect 40625 -2380 40680 -2260
rect 40800 -2380 40845 -2260
rect 40965 -2380 41010 -2260
rect 41130 -2380 41175 -2260
rect 41295 -2380 41350 -2260
rect 41470 -2380 41515 -2260
rect 41635 -2380 41680 -2260
rect 41800 -2380 41845 -2260
rect 41965 -2380 42175 -2260
rect 42295 -2380 42350 -2260
rect 42470 -2380 42515 -2260
rect 42635 -2380 42680 -2260
rect 42800 -2380 42845 -2260
rect 42965 -2380 43020 -2260
rect 43140 -2380 43185 -2260
rect 43305 -2380 43350 -2260
rect 43470 -2380 43515 -2260
rect 43635 -2380 43690 -2260
rect 43810 -2380 43855 -2260
rect 43975 -2380 44020 -2260
rect 44140 -2380 44185 -2260
rect 44305 -2380 44360 -2260
rect 44480 -2380 44525 -2260
rect 44645 -2380 44690 -2260
rect 44810 -2380 44855 -2260
rect 44975 -2380 45030 -2260
rect 45150 -2380 45195 -2260
rect 45315 -2380 45360 -2260
rect 45480 -2380 45525 -2260
rect 45645 -2380 45700 -2260
rect 45820 -2380 45865 -2260
rect 45985 -2380 46030 -2260
rect 46150 -2380 46195 -2260
rect 46315 -2380 46370 -2260
rect 46490 -2380 46535 -2260
rect 46655 -2380 46700 -2260
rect 46820 -2380 46865 -2260
rect 46985 -2380 47040 -2260
rect 47160 -2380 47205 -2260
rect 47325 -2380 47370 -2260
rect 47490 -2380 47535 -2260
rect 47655 -2380 47865 -2260
rect 47985 -2380 48040 -2260
rect 48160 -2380 48205 -2260
rect 48325 -2380 48370 -2260
rect 48490 -2380 48535 -2260
rect 48655 -2380 48710 -2260
rect 48830 -2380 48875 -2260
rect 48995 -2380 49040 -2260
rect 49160 -2380 49205 -2260
rect 49325 -2380 49380 -2260
rect 49500 -2380 49545 -2260
rect 49665 -2380 49710 -2260
rect 49830 -2380 49875 -2260
rect 49995 -2380 50050 -2260
rect 50170 -2380 50215 -2260
rect 50335 -2380 50380 -2260
rect 50500 -2380 50545 -2260
rect 50665 -2380 50720 -2260
rect 50840 -2380 50885 -2260
rect 51005 -2380 51050 -2260
rect 51170 -2380 51215 -2260
rect 51335 -2380 51390 -2260
rect 51510 -2380 51555 -2260
rect 51675 -2380 51720 -2260
rect 51840 -2380 51885 -2260
rect 52005 -2380 52060 -2260
rect 52180 -2380 52225 -2260
rect 52345 -2380 52390 -2260
rect 52510 -2380 52555 -2260
rect 52675 -2380 52730 -2260
rect 52850 -2380 52895 -2260
rect 53015 -2380 53060 -2260
rect 53180 -2380 53225 -2260
rect 53345 -2380 53370 -2260
rect 30770 -2425 53370 -2380
rect 30770 -2545 30795 -2425
rect 30915 -2545 30970 -2425
rect 31090 -2545 31135 -2425
rect 31255 -2545 31300 -2425
rect 31420 -2545 31465 -2425
rect 31585 -2545 31640 -2425
rect 31760 -2545 31805 -2425
rect 31925 -2545 31970 -2425
rect 32090 -2545 32135 -2425
rect 32255 -2545 32310 -2425
rect 32430 -2545 32475 -2425
rect 32595 -2545 32640 -2425
rect 32760 -2545 32805 -2425
rect 32925 -2545 32980 -2425
rect 33100 -2545 33145 -2425
rect 33265 -2545 33310 -2425
rect 33430 -2545 33475 -2425
rect 33595 -2545 33650 -2425
rect 33770 -2545 33815 -2425
rect 33935 -2545 33980 -2425
rect 34100 -2545 34145 -2425
rect 34265 -2545 34320 -2425
rect 34440 -2545 34485 -2425
rect 34605 -2545 34650 -2425
rect 34770 -2545 34815 -2425
rect 34935 -2545 34990 -2425
rect 35110 -2545 35155 -2425
rect 35275 -2545 35320 -2425
rect 35440 -2545 35485 -2425
rect 35605 -2545 35660 -2425
rect 35780 -2545 35825 -2425
rect 35945 -2545 35990 -2425
rect 36110 -2545 36155 -2425
rect 36275 -2545 36485 -2425
rect 36605 -2545 36660 -2425
rect 36780 -2545 36825 -2425
rect 36945 -2545 36990 -2425
rect 37110 -2545 37155 -2425
rect 37275 -2545 37330 -2425
rect 37450 -2545 37495 -2425
rect 37615 -2545 37660 -2425
rect 37780 -2545 37825 -2425
rect 37945 -2545 38000 -2425
rect 38120 -2545 38165 -2425
rect 38285 -2545 38330 -2425
rect 38450 -2545 38495 -2425
rect 38615 -2545 38670 -2425
rect 38790 -2545 38835 -2425
rect 38955 -2545 39000 -2425
rect 39120 -2545 39165 -2425
rect 39285 -2545 39340 -2425
rect 39460 -2545 39505 -2425
rect 39625 -2545 39670 -2425
rect 39790 -2545 39835 -2425
rect 39955 -2545 40010 -2425
rect 40130 -2545 40175 -2425
rect 40295 -2545 40340 -2425
rect 40460 -2545 40505 -2425
rect 40625 -2545 40680 -2425
rect 40800 -2545 40845 -2425
rect 40965 -2545 41010 -2425
rect 41130 -2545 41175 -2425
rect 41295 -2545 41350 -2425
rect 41470 -2545 41515 -2425
rect 41635 -2545 41680 -2425
rect 41800 -2545 41845 -2425
rect 41965 -2545 42175 -2425
rect 42295 -2545 42350 -2425
rect 42470 -2545 42515 -2425
rect 42635 -2545 42680 -2425
rect 42800 -2545 42845 -2425
rect 42965 -2545 43020 -2425
rect 43140 -2545 43185 -2425
rect 43305 -2545 43350 -2425
rect 43470 -2545 43515 -2425
rect 43635 -2545 43690 -2425
rect 43810 -2545 43855 -2425
rect 43975 -2545 44020 -2425
rect 44140 -2545 44185 -2425
rect 44305 -2545 44360 -2425
rect 44480 -2545 44525 -2425
rect 44645 -2545 44690 -2425
rect 44810 -2545 44855 -2425
rect 44975 -2545 45030 -2425
rect 45150 -2545 45195 -2425
rect 45315 -2545 45360 -2425
rect 45480 -2545 45525 -2425
rect 45645 -2545 45700 -2425
rect 45820 -2545 45865 -2425
rect 45985 -2545 46030 -2425
rect 46150 -2545 46195 -2425
rect 46315 -2545 46370 -2425
rect 46490 -2545 46535 -2425
rect 46655 -2545 46700 -2425
rect 46820 -2545 46865 -2425
rect 46985 -2545 47040 -2425
rect 47160 -2545 47205 -2425
rect 47325 -2545 47370 -2425
rect 47490 -2545 47535 -2425
rect 47655 -2545 47865 -2425
rect 47985 -2545 48040 -2425
rect 48160 -2545 48205 -2425
rect 48325 -2545 48370 -2425
rect 48490 -2545 48535 -2425
rect 48655 -2545 48710 -2425
rect 48830 -2545 48875 -2425
rect 48995 -2545 49040 -2425
rect 49160 -2545 49205 -2425
rect 49325 -2545 49380 -2425
rect 49500 -2545 49545 -2425
rect 49665 -2545 49710 -2425
rect 49830 -2545 49875 -2425
rect 49995 -2545 50050 -2425
rect 50170 -2545 50215 -2425
rect 50335 -2545 50380 -2425
rect 50500 -2545 50545 -2425
rect 50665 -2545 50720 -2425
rect 50840 -2545 50885 -2425
rect 51005 -2545 51050 -2425
rect 51170 -2545 51215 -2425
rect 51335 -2545 51390 -2425
rect 51510 -2545 51555 -2425
rect 51675 -2545 51720 -2425
rect 51840 -2545 51885 -2425
rect 52005 -2545 52060 -2425
rect 52180 -2545 52225 -2425
rect 52345 -2545 52390 -2425
rect 52510 -2545 52555 -2425
rect 52675 -2545 52730 -2425
rect 52850 -2545 52895 -2425
rect 53015 -2545 53060 -2425
rect 53180 -2545 53225 -2425
rect 53345 -2545 53370 -2425
rect 30770 -2600 53370 -2545
rect 30770 -2720 30795 -2600
rect 30915 -2720 30970 -2600
rect 31090 -2720 31135 -2600
rect 31255 -2720 31300 -2600
rect 31420 -2720 31465 -2600
rect 31585 -2720 31640 -2600
rect 31760 -2720 31805 -2600
rect 31925 -2720 31970 -2600
rect 32090 -2720 32135 -2600
rect 32255 -2720 32310 -2600
rect 32430 -2720 32475 -2600
rect 32595 -2720 32640 -2600
rect 32760 -2720 32805 -2600
rect 32925 -2720 32980 -2600
rect 33100 -2720 33145 -2600
rect 33265 -2720 33310 -2600
rect 33430 -2720 33475 -2600
rect 33595 -2720 33650 -2600
rect 33770 -2720 33815 -2600
rect 33935 -2720 33980 -2600
rect 34100 -2720 34145 -2600
rect 34265 -2720 34320 -2600
rect 34440 -2720 34485 -2600
rect 34605 -2720 34650 -2600
rect 34770 -2720 34815 -2600
rect 34935 -2720 34990 -2600
rect 35110 -2720 35155 -2600
rect 35275 -2720 35320 -2600
rect 35440 -2720 35485 -2600
rect 35605 -2720 35660 -2600
rect 35780 -2720 35825 -2600
rect 35945 -2720 35990 -2600
rect 36110 -2720 36155 -2600
rect 36275 -2720 36485 -2600
rect 36605 -2720 36660 -2600
rect 36780 -2720 36825 -2600
rect 36945 -2720 36990 -2600
rect 37110 -2720 37155 -2600
rect 37275 -2720 37330 -2600
rect 37450 -2720 37495 -2600
rect 37615 -2720 37660 -2600
rect 37780 -2720 37825 -2600
rect 37945 -2720 38000 -2600
rect 38120 -2720 38165 -2600
rect 38285 -2720 38330 -2600
rect 38450 -2720 38495 -2600
rect 38615 -2720 38670 -2600
rect 38790 -2720 38835 -2600
rect 38955 -2720 39000 -2600
rect 39120 -2720 39165 -2600
rect 39285 -2720 39340 -2600
rect 39460 -2720 39505 -2600
rect 39625 -2720 39670 -2600
rect 39790 -2720 39835 -2600
rect 39955 -2720 40010 -2600
rect 40130 -2720 40175 -2600
rect 40295 -2720 40340 -2600
rect 40460 -2720 40505 -2600
rect 40625 -2720 40680 -2600
rect 40800 -2720 40845 -2600
rect 40965 -2720 41010 -2600
rect 41130 -2720 41175 -2600
rect 41295 -2720 41350 -2600
rect 41470 -2720 41515 -2600
rect 41635 -2720 41680 -2600
rect 41800 -2720 41845 -2600
rect 41965 -2720 42175 -2600
rect 42295 -2720 42350 -2600
rect 42470 -2720 42515 -2600
rect 42635 -2720 42680 -2600
rect 42800 -2720 42845 -2600
rect 42965 -2720 43020 -2600
rect 43140 -2720 43185 -2600
rect 43305 -2720 43350 -2600
rect 43470 -2720 43515 -2600
rect 43635 -2720 43690 -2600
rect 43810 -2720 43855 -2600
rect 43975 -2720 44020 -2600
rect 44140 -2720 44185 -2600
rect 44305 -2720 44360 -2600
rect 44480 -2720 44525 -2600
rect 44645 -2720 44690 -2600
rect 44810 -2720 44855 -2600
rect 44975 -2720 45030 -2600
rect 45150 -2720 45195 -2600
rect 45315 -2720 45360 -2600
rect 45480 -2720 45525 -2600
rect 45645 -2720 45700 -2600
rect 45820 -2720 45865 -2600
rect 45985 -2720 46030 -2600
rect 46150 -2720 46195 -2600
rect 46315 -2720 46370 -2600
rect 46490 -2720 46535 -2600
rect 46655 -2720 46700 -2600
rect 46820 -2720 46865 -2600
rect 46985 -2720 47040 -2600
rect 47160 -2720 47205 -2600
rect 47325 -2720 47370 -2600
rect 47490 -2720 47535 -2600
rect 47655 -2720 47865 -2600
rect 47985 -2720 48040 -2600
rect 48160 -2720 48205 -2600
rect 48325 -2720 48370 -2600
rect 48490 -2720 48535 -2600
rect 48655 -2720 48710 -2600
rect 48830 -2720 48875 -2600
rect 48995 -2720 49040 -2600
rect 49160 -2720 49205 -2600
rect 49325 -2720 49380 -2600
rect 49500 -2720 49545 -2600
rect 49665 -2720 49710 -2600
rect 49830 -2720 49875 -2600
rect 49995 -2720 50050 -2600
rect 50170 -2720 50215 -2600
rect 50335 -2720 50380 -2600
rect 50500 -2720 50545 -2600
rect 50665 -2720 50720 -2600
rect 50840 -2720 50885 -2600
rect 51005 -2720 51050 -2600
rect 51170 -2720 51215 -2600
rect 51335 -2720 51390 -2600
rect 51510 -2720 51555 -2600
rect 51675 -2720 51720 -2600
rect 51840 -2720 51885 -2600
rect 52005 -2720 52060 -2600
rect 52180 -2720 52225 -2600
rect 52345 -2720 52390 -2600
rect 52510 -2720 52555 -2600
rect 52675 -2720 52730 -2600
rect 52850 -2720 52895 -2600
rect 53015 -2720 53060 -2600
rect 53180 -2720 53225 -2600
rect 53345 -2720 53370 -2600
rect 30770 -2765 53370 -2720
rect 30770 -2885 30795 -2765
rect 30915 -2885 30970 -2765
rect 31090 -2885 31135 -2765
rect 31255 -2885 31300 -2765
rect 31420 -2885 31465 -2765
rect 31585 -2885 31640 -2765
rect 31760 -2885 31805 -2765
rect 31925 -2885 31970 -2765
rect 32090 -2885 32135 -2765
rect 32255 -2885 32310 -2765
rect 32430 -2885 32475 -2765
rect 32595 -2885 32640 -2765
rect 32760 -2885 32805 -2765
rect 32925 -2885 32980 -2765
rect 33100 -2885 33145 -2765
rect 33265 -2885 33310 -2765
rect 33430 -2885 33475 -2765
rect 33595 -2885 33650 -2765
rect 33770 -2885 33815 -2765
rect 33935 -2885 33980 -2765
rect 34100 -2885 34145 -2765
rect 34265 -2885 34320 -2765
rect 34440 -2885 34485 -2765
rect 34605 -2885 34650 -2765
rect 34770 -2885 34815 -2765
rect 34935 -2885 34990 -2765
rect 35110 -2885 35155 -2765
rect 35275 -2885 35320 -2765
rect 35440 -2885 35485 -2765
rect 35605 -2885 35660 -2765
rect 35780 -2885 35825 -2765
rect 35945 -2885 35990 -2765
rect 36110 -2885 36155 -2765
rect 36275 -2885 36485 -2765
rect 36605 -2885 36660 -2765
rect 36780 -2885 36825 -2765
rect 36945 -2885 36990 -2765
rect 37110 -2885 37155 -2765
rect 37275 -2885 37330 -2765
rect 37450 -2885 37495 -2765
rect 37615 -2885 37660 -2765
rect 37780 -2885 37825 -2765
rect 37945 -2885 38000 -2765
rect 38120 -2885 38165 -2765
rect 38285 -2885 38330 -2765
rect 38450 -2885 38495 -2765
rect 38615 -2885 38670 -2765
rect 38790 -2885 38835 -2765
rect 38955 -2885 39000 -2765
rect 39120 -2885 39165 -2765
rect 39285 -2885 39340 -2765
rect 39460 -2885 39505 -2765
rect 39625 -2885 39670 -2765
rect 39790 -2885 39835 -2765
rect 39955 -2885 40010 -2765
rect 40130 -2885 40175 -2765
rect 40295 -2885 40340 -2765
rect 40460 -2885 40505 -2765
rect 40625 -2885 40680 -2765
rect 40800 -2885 40845 -2765
rect 40965 -2885 41010 -2765
rect 41130 -2885 41175 -2765
rect 41295 -2885 41350 -2765
rect 41470 -2885 41515 -2765
rect 41635 -2885 41680 -2765
rect 41800 -2885 41845 -2765
rect 41965 -2885 42175 -2765
rect 42295 -2885 42350 -2765
rect 42470 -2885 42515 -2765
rect 42635 -2885 42680 -2765
rect 42800 -2885 42845 -2765
rect 42965 -2885 43020 -2765
rect 43140 -2885 43185 -2765
rect 43305 -2885 43350 -2765
rect 43470 -2885 43515 -2765
rect 43635 -2885 43690 -2765
rect 43810 -2885 43855 -2765
rect 43975 -2885 44020 -2765
rect 44140 -2885 44185 -2765
rect 44305 -2885 44360 -2765
rect 44480 -2885 44525 -2765
rect 44645 -2885 44690 -2765
rect 44810 -2885 44855 -2765
rect 44975 -2885 45030 -2765
rect 45150 -2885 45195 -2765
rect 45315 -2885 45360 -2765
rect 45480 -2885 45525 -2765
rect 45645 -2885 45700 -2765
rect 45820 -2885 45865 -2765
rect 45985 -2885 46030 -2765
rect 46150 -2885 46195 -2765
rect 46315 -2885 46370 -2765
rect 46490 -2885 46535 -2765
rect 46655 -2885 46700 -2765
rect 46820 -2885 46865 -2765
rect 46985 -2885 47040 -2765
rect 47160 -2885 47205 -2765
rect 47325 -2885 47370 -2765
rect 47490 -2885 47535 -2765
rect 47655 -2885 47865 -2765
rect 47985 -2885 48040 -2765
rect 48160 -2885 48205 -2765
rect 48325 -2885 48370 -2765
rect 48490 -2885 48535 -2765
rect 48655 -2885 48710 -2765
rect 48830 -2885 48875 -2765
rect 48995 -2885 49040 -2765
rect 49160 -2885 49205 -2765
rect 49325 -2885 49380 -2765
rect 49500 -2885 49545 -2765
rect 49665 -2885 49710 -2765
rect 49830 -2885 49875 -2765
rect 49995 -2885 50050 -2765
rect 50170 -2885 50215 -2765
rect 50335 -2885 50380 -2765
rect 50500 -2885 50545 -2765
rect 50665 -2885 50720 -2765
rect 50840 -2885 50885 -2765
rect 51005 -2885 51050 -2765
rect 51170 -2885 51215 -2765
rect 51335 -2885 51390 -2765
rect 51510 -2885 51555 -2765
rect 51675 -2885 51720 -2765
rect 51840 -2885 51885 -2765
rect 52005 -2885 52060 -2765
rect 52180 -2885 52225 -2765
rect 52345 -2885 52390 -2765
rect 52510 -2885 52555 -2765
rect 52675 -2885 52730 -2765
rect 52850 -2885 52895 -2765
rect 53015 -2885 53060 -2765
rect 53180 -2885 53225 -2765
rect 53345 -2885 53370 -2765
rect 30770 -2930 53370 -2885
rect 30770 -3050 30795 -2930
rect 30915 -3050 30970 -2930
rect 31090 -3050 31135 -2930
rect 31255 -3050 31300 -2930
rect 31420 -3050 31465 -2930
rect 31585 -3050 31640 -2930
rect 31760 -3050 31805 -2930
rect 31925 -3050 31970 -2930
rect 32090 -3050 32135 -2930
rect 32255 -3050 32310 -2930
rect 32430 -3050 32475 -2930
rect 32595 -3050 32640 -2930
rect 32760 -3050 32805 -2930
rect 32925 -3050 32980 -2930
rect 33100 -3050 33145 -2930
rect 33265 -3050 33310 -2930
rect 33430 -3050 33475 -2930
rect 33595 -3050 33650 -2930
rect 33770 -3050 33815 -2930
rect 33935 -3050 33980 -2930
rect 34100 -3050 34145 -2930
rect 34265 -3050 34320 -2930
rect 34440 -3050 34485 -2930
rect 34605 -3050 34650 -2930
rect 34770 -3050 34815 -2930
rect 34935 -3050 34990 -2930
rect 35110 -3050 35155 -2930
rect 35275 -3050 35320 -2930
rect 35440 -3050 35485 -2930
rect 35605 -3050 35660 -2930
rect 35780 -3050 35825 -2930
rect 35945 -3050 35990 -2930
rect 36110 -3050 36155 -2930
rect 36275 -3050 36485 -2930
rect 36605 -3050 36660 -2930
rect 36780 -3050 36825 -2930
rect 36945 -3050 36990 -2930
rect 37110 -3050 37155 -2930
rect 37275 -3050 37330 -2930
rect 37450 -3050 37495 -2930
rect 37615 -3050 37660 -2930
rect 37780 -3050 37825 -2930
rect 37945 -3050 38000 -2930
rect 38120 -3050 38165 -2930
rect 38285 -3050 38330 -2930
rect 38450 -3050 38495 -2930
rect 38615 -3050 38670 -2930
rect 38790 -3050 38835 -2930
rect 38955 -3050 39000 -2930
rect 39120 -3050 39165 -2930
rect 39285 -3050 39340 -2930
rect 39460 -3050 39505 -2930
rect 39625 -3050 39670 -2930
rect 39790 -3050 39835 -2930
rect 39955 -3050 40010 -2930
rect 40130 -3050 40175 -2930
rect 40295 -3050 40340 -2930
rect 40460 -3050 40505 -2930
rect 40625 -3050 40680 -2930
rect 40800 -3050 40845 -2930
rect 40965 -3050 41010 -2930
rect 41130 -3050 41175 -2930
rect 41295 -3050 41350 -2930
rect 41470 -3050 41515 -2930
rect 41635 -3050 41680 -2930
rect 41800 -3050 41845 -2930
rect 41965 -3050 42175 -2930
rect 42295 -3050 42350 -2930
rect 42470 -3050 42515 -2930
rect 42635 -3050 42680 -2930
rect 42800 -3050 42845 -2930
rect 42965 -3050 43020 -2930
rect 43140 -3050 43185 -2930
rect 43305 -3050 43350 -2930
rect 43470 -3050 43515 -2930
rect 43635 -3050 43690 -2930
rect 43810 -3050 43855 -2930
rect 43975 -3050 44020 -2930
rect 44140 -3050 44185 -2930
rect 44305 -3050 44360 -2930
rect 44480 -3050 44525 -2930
rect 44645 -3050 44690 -2930
rect 44810 -3050 44855 -2930
rect 44975 -3050 45030 -2930
rect 45150 -3050 45195 -2930
rect 45315 -3050 45360 -2930
rect 45480 -3050 45525 -2930
rect 45645 -3050 45700 -2930
rect 45820 -3050 45865 -2930
rect 45985 -3050 46030 -2930
rect 46150 -3050 46195 -2930
rect 46315 -3050 46370 -2930
rect 46490 -3050 46535 -2930
rect 46655 -3050 46700 -2930
rect 46820 -3050 46865 -2930
rect 46985 -3050 47040 -2930
rect 47160 -3050 47205 -2930
rect 47325 -3050 47370 -2930
rect 47490 -3050 47535 -2930
rect 47655 -3050 47865 -2930
rect 47985 -3050 48040 -2930
rect 48160 -3050 48205 -2930
rect 48325 -3050 48370 -2930
rect 48490 -3050 48535 -2930
rect 48655 -3050 48710 -2930
rect 48830 -3050 48875 -2930
rect 48995 -3050 49040 -2930
rect 49160 -3050 49205 -2930
rect 49325 -3050 49380 -2930
rect 49500 -3050 49545 -2930
rect 49665 -3050 49710 -2930
rect 49830 -3050 49875 -2930
rect 49995 -3050 50050 -2930
rect 50170 -3050 50215 -2930
rect 50335 -3050 50380 -2930
rect 50500 -3050 50545 -2930
rect 50665 -3050 50720 -2930
rect 50840 -3050 50885 -2930
rect 51005 -3050 51050 -2930
rect 51170 -3050 51215 -2930
rect 51335 -3050 51390 -2930
rect 51510 -3050 51555 -2930
rect 51675 -3050 51720 -2930
rect 51840 -3050 51885 -2930
rect 52005 -3050 52060 -2930
rect 52180 -3050 52225 -2930
rect 52345 -3050 52390 -2930
rect 52510 -3050 52555 -2930
rect 52675 -3050 52730 -2930
rect 52850 -3050 52895 -2930
rect 53015 -3050 53060 -2930
rect 53180 -3050 53225 -2930
rect 53345 -3050 53370 -2930
rect 30770 -3095 53370 -3050
rect 30770 -3215 30795 -3095
rect 30915 -3215 30970 -3095
rect 31090 -3215 31135 -3095
rect 31255 -3215 31300 -3095
rect 31420 -3215 31465 -3095
rect 31585 -3215 31640 -3095
rect 31760 -3215 31805 -3095
rect 31925 -3215 31970 -3095
rect 32090 -3215 32135 -3095
rect 32255 -3215 32310 -3095
rect 32430 -3215 32475 -3095
rect 32595 -3215 32640 -3095
rect 32760 -3215 32805 -3095
rect 32925 -3215 32980 -3095
rect 33100 -3215 33145 -3095
rect 33265 -3215 33310 -3095
rect 33430 -3215 33475 -3095
rect 33595 -3215 33650 -3095
rect 33770 -3215 33815 -3095
rect 33935 -3215 33980 -3095
rect 34100 -3215 34145 -3095
rect 34265 -3215 34320 -3095
rect 34440 -3215 34485 -3095
rect 34605 -3215 34650 -3095
rect 34770 -3215 34815 -3095
rect 34935 -3215 34990 -3095
rect 35110 -3215 35155 -3095
rect 35275 -3215 35320 -3095
rect 35440 -3215 35485 -3095
rect 35605 -3215 35660 -3095
rect 35780 -3215 35825 -3095
rect 35945 -3215 35990 -3095
rect 36110 -3215 36155 -3095
rect 36275 -3215 36485 -3095
rect 36605 -3215 36660 -3095
rect 36780 -3215 36825 -3095
rect 36945 -3215 36990 -3095
rect 37110 -3215 37155 -3095
rect 37275 -3215 37330 -3095
rect 37450 -3215 37495 -3095
rect 37615 -3215 37660 -3095
rect 37780 -3215 37825 -3095
rect 37945 -3215 38000 -3095
rect 38120 -3215 38165 -3095
rect 38285 -3215 38330 -3095
rect 38450 -3215 38495 -3095
rect 38615 -3215 38670 -3095
rect 38790 -3215 38835 -3095
rect 38955 -3215 39000 -3095
rect 39120 -3215 39165 -3095
rect 39285 -3215 39340 -3095
rect 39460 -3215 39505 -3095
rect 39625 -3215 39670 -3095
rect 39790 -3215 39835 -3095
rect 39955 -3215 40010 -3095
rect 40130 -3215 40175 -3095
rect 40295 -3215 40340 -3095
rect 40460 -3215 40505 -3095
rect 40625 -3215 40680 -3095
rect 40800 -3215 40845 -3095
rect 40965 -3215 41010 -3095
rect 41130 -3215 41175 -3095
rect 41295 -3215 41350 -3095
rect 41470 -3215 41515 -3095
rect 41635 -3215 41680 -3095
rect 41800 -3215 41845 -3095
rect 41965 -3215 42175 -3095
rect 42295 -3215 42350 -3095
rect 42470 -3215 42515 -3095
rect 42635 -3215 42680 -3095
rect 42800 -3215 42845 -3095
rect 42965 -3215 43020 -3095
rect 43140 -3215 43185 -3095
rect 43305 -3215 43350 -3095
rect 43470 -3215 43515 -3095
rect 43635 -3215 43690 -3095
rect 43810 -3215 43855 -3095
rect 43975 -3215 44020 -3095
rect 44140 -3215 44185 -3095
rect 44305 -3215 44360 -3095
rect 44480 -3215 44525 -3095
rect 44645 -3215 44690 -3095
rect 44810 -3215 44855 -3095
rect 44975 -3215 45030 -3095
rect 45150 -3215 45195 -3095
rect 45315 -3215 45360 -3095
rect 45480 -3215 45525 -3095
rect 45645 -3215 45700 -3095
rect 45820 -3215 45865 -3095
rect 45985 -3215 46030 -3095
rect 46150 -3215 46195 -3095
rect 46315 -3215 46370 -3095
rect 46490 -3215 46535 -3095
rect 46655 -3215 46700 -3095
rect 46820 -3215 46865 -3095
rect 46985 -3215 47040 -3095
rect 47160 -3215 47205 -3095
rect 47325 -3215 47370 -3095
rect 47490 -3215 47535 -3095
rect 47655 -3215 47865 -3095
rect 47985 -3215 48040 -3095
rect 48160 -3215 48205 -3095
rect 48325 -3215 48370 -3095
rect 48490 -3215 48535 -3095
rect 48655 -3215 48710 -3095
rect 48830 -3215 48875 -3095
rect 48995 -3215 49040 -3095
rect 49160 -3215 49205 -3095
rect 49325 -3215 49380 -3095
rect 49500 -3215 49545 -3095
rect 49665 -3215 49710 -3095
rect 49830 -3215 49875 -3095
rect 49995 -3215 50050 -3095
rect 50170 -3215 50215 -3095
rect 50335 -3215 50380 -3095
rect 50500 -3215 50545 -3095
rect 50665 -3215 50720 -3095
rect 50840 -3215 50885 -3095
rect 51005 -3215 51050 -3095
rect 51170 -3215 51215 -3095
rect 51335 -3215 51390 -3095
rect 51510 -3215 51555 -3095
rect 51675 -3215 51720 -3095
rect 51840 -3215 51885 -3095
rect 52005 -3215 52060 -3095
rect 52180 -3215 52225 -3095
rect 52345 -3215 52390 -3095
rect 52510 -3215 52555 -3095
rect 52675 -3215 52730 -3095
rect 52850 -3215 52895 -3095
rect 53015 -3215 53060 -3095
rect 53180 -3215 53225 -3095
rect 53345 -3215 53370 -3095
rect 30770 -3270 53370 -3215
rect 30770 -3390 30795 -3270
rect 30915 -3390 30970 -3270
rect 31090 -3390 31135 -3270
rect 31255 -3390 31300 -3270
rect 31420 -3390 31465 -3270
rect 31585 -3390 31640 -3270
rect 31760 -3390 31805 -3270
rect 31925 -3390 31970 -3270
rect 32090 -3390 32135 -3270
rect 32255 -3390 32310 -3270
rect 32430 -3390 32475 -3270
rect 32595 -3390 32640 -3270
rect 32760 -3390 32805 -3270
rect 32925 -3390 32980 -3270
rect 33100 -3390 33145 -3270
rect 33265 -3390 33310 -3270
rect 33430 -3390 33475 -3270
rect 33595 -3390 33650 -3270
rect 33770 -3390 33815 -3270
rect 33935 -3390 33980 -3270
rect 34100 -3390 34145 -3270
rect 34265 -3390 34320 -3270
rect 34440 -3390 34485 -3270
rect 34605 -3390 34650 -3270
rect 34770 -3390 34815 -3270
rect 34935 -3390 34990 -3270
rect 35110 -3390 35155 -3270
rect 35275 -3390 35320 -3270
rect 35440 -3390 35485 -3270
rect 35605 -3390 35660 -3270
rect 35780 -3390 35825 -3270
rect 35945 -3390 35990 -3270
rect 36110 -3390 36155 -3270
rect 36275 -3390 36485 -3270
rect 36605 -3390 36660 -3270
rect 36780 -3390 36825 -3270
rect 36945 -3390 36990 -3270
rect 37110 -3390 37155 -3270
rect 37275 -3390 37330 -3270
rect 37450 -3390 37495 -3270
rect 37615 -3390 37660 -3270
rect 37780 -3390 37825 -3270
rect 37945 -3390 38000 -3270
rect 38120 -3390 38165 -3270
rect 38285 -3390 38330 -3270
rect 38450 -3390 38495 -3270
rect 38615 -3390 38670 -3270
rect 38790 -3390 38835 -3270
rect 38955 -3390 39000 -3270
rect 39120 -3390 39165 -3270
rect 39285 -3390 39340 -3270
rect 39460 -3390 39505 -3270
rect 39625 -3390 39670 -3270
rect 39790 -3390 39835 -3270
rect 39955 -3390 40010 -3270
rect 40130 -3390 40175 -3270
rect 40295 -3390 40340 -3270
rect 40460 -3390 40505 -3270
rect 40625 -3390 40680 -3270
rect 40800 -3390 40845 -3270
rect 40965 -3390 41010 -3270
rect 41130 -3390 41175 -3270
rect 41295 -3390 41350 -3270
rect 41470 -3390 41515 -3270
rect 41635 -3390 41680 -3270
rect 41800 -3390 41845 -3270
rect 41965 -3390 42175 -3270
rect 42295 -3390 42350 -3270
rect 42470 -3390 42515 -3270
rect 42635 -3390 42680 -3270
rect 42800 -3390 42845 -3270
rect 42965 -3390 43020 -3270
rect 43140 -3390 43185 -3270
rect 43305 -3390 43350 -3270
rect 43470 -3390 43515 -3270
rect 43635 -3390 43690 -3270
rect 43810 -3390 43855 -3270
rect 43975 -3390 44020 -3270
rect 44140 -3390 44185 -3270
rect 44305 -3390 44360 -3270
rect 44480 -3390 44525 -3270
rect 44645 -3390 44690 -3270
rect 44810 -3390 44855 -3270
rect 44975 -3390 45030 -3270
rect 45150 -3390 45195 -3270
rect 45315 -3390 45360 -3270
rect 45480 -3390 45525 -3270
rect 45645 -3390 45700 -3270
rect 45820 -3390 45865 -3270
rect 45985 -3390 46030 -3270
rect 46150 -3390 46195 -3270
rect 46315 -3390 46370 -3270
rect 46490 -3390 46535 -3270
rect 46655 -3390 46700 -3270
rect 46820 -3390 46865 -3270
rect 46985 -3390 47040 -3270
rect 47160 -3390 47205 -3270
rect 47325 -3390 47370 -3270
rect 47490 -3390 47535 -3270
rect 47655 -3390 47865 -3270
rect 47985 -3390 48040 -3270
rect 48160 -3390 48205 -3270
rect 48325 -3390 48370 -3270
rect 48490 -3390 48535 -3270
rect 48655 -3390 48710 -3270
rect 48830 -3390 48875 -3270
rect 48995 -3390 49040 -3270
rect 49160 -3390 49205 -3270
rect 49325 -3390 49380 -3270
rect 49500 -3390 49545 -3270
rect 49665 -3390 49710 -3270
rect 49830 -3390 49875 -3270
rect 49995 -3390 50050 -3270
rect 50170 -3390 50215 -3270
rect 50335 -3390 50380 -3270
rect 50500 -3390 50545 -3270
rect 50665 -3390 50720 -3270
rect 50840 -3390 50885 -3270
rect 51005 -3390 51050 -3270
rect 51170 -3390 51215 -3270
rect 51335 -3390 51390 -3270
rect 51510 -3390 51555 -3270
rect 51675 -3390 51720 -3270
rect 51840 -3390 51885 -3270
rect 52005 -3390 52060 -3270
rect 52180 -3390 52225 -3270
rect 52345 -3390 52390 -3270
rect 52510 -3390 52555 -3270
rect 52675 -3390 52730 -3270
rect 52850 -3390 52895 -3270
rect 53015 -3390 53060 -3270
rect 53180 -3390 53225 -3270
rect 53345 -3390 53370 -3270
rect 30770 -3435 53370 -3390
rect 30770 -3555 30795 -3435
rect 30915 -3555 30970 -3435
rect 31090 -3555 31135 -3435
rect 31255 -3555 31300 -3435
rect 31420 -3555 31465 -3435
rect 31585 -3555 31640 -3435
rect 31760 -3555 31805 -3435
rect 31925 -3555 31970 -3435
rect 32090 -3555 32135 -3435
rect 32255 -3555 32310 -3435
rect 32430 -3555 32475 -3435
rect 32595 -3555 32640 -3435
rect 32760 -3555 32805 -3435
rect 32925 -3555 32980 -3435
rect 33100 -3555 33145 -3435
rect 33265 -3555 33310 -3435
rect 33430 -3555 33475 -3435
rect 33595 -3555 33650 -3435
rect 33770 -3555 33815 -3435
rect 33935 -3555 33980 -3435
rect 34100 -3555 34145 -3435
rect 34265 -3555 34320 -3435
rect 34440 -3555 34485 -3435
rect 34605 -3555 34650 -3435
rect 34770 -3555 34815 -3435
rect 34935 -3555 34990 -3435
rect 35110 -3555 35155 -3435
rect 35275 -3555 35320 -3435
rect 35440 -3555 35485 -3435
rect 35605 -3555 35660 -3435
rect 35780 -3555 35825 -3435
rect 35945 -3555 35990 -3435
rect 36110 -3555 36155 -3435
rect 36275 -3555 36485 -3435
rect 36605 -3555 36660 -3435
rect 36780 -3555 36825 -3435
rect 36945 -3555 36990 -3435
rect 37110 -3555 37155 -3435
rect 37275 -3555 37330 -3435
rect 37450 -3555 37495 -3435
rect 37615 -3555 37660 -3435
rect 37780 -3555 37825 -3435
rect 37945 -3555 38000 -3435
rect 38120 -3555 38165 -3435
rect 38285 -3555 38330 -3435
rect 38450 -3555 38495 -3435
rect 38615 -3555 38670 -3435
rect 38790 -3555 38835 -3435
rect 38955 -3555 39000 -3435
rect 39120 -3555 39165 -3435
rect 39285 -3555 39340 -3435
rect 39460 -3555 39505 -3435
rect 39625 -3555 39670 -3435
rect 39790 -3555 39835 -3435
rect 39955 -3555 40010 -3435
rect 40130 -3555 40175 -3435
rect 40295 -3555 40340 -3435
rect 40460 -3555 40505 -3435
rect 40625 -3555 40680 -3435
rect 40800 -3555 40845 -3435
rect 40965 -3555 41010 -3435
rect 41130 -3555 41175 -3435
rect 41295 -3555 41350 -3435
rect 41470 -3555 41515 -3435
rect 41635 -3555 41680 -3435
rect 41800 -3555 41845 -3435
rect 41965 -3555 42175 -3435
rect 42295 -3555 42350 -3435
rect 42470 -3555 42515 -3435
rect 42635 -3555 42680 -3435
rect 42800 -3555 42845 -3435
rect 42965 -3555 43020 -3435
rect 43140 -3555 43185 -3435
rect 43305 -3555 43350 -3435
rect 43470 -3555 43515 -3435
rect 43635 -3555 43690 -3435
rect 43810 -3555 43855 -3435
rect 43975 -3555 44020 -3435
rect 44140 -3555 44185 -3435
rect 44305 -3555 44360 -3435
rect 44480 -3555 44525 -3435
rect 44645 -3555 44690 -3435
rect 44810 -3555 44855 -3435
rect 44975 -3555 45030 -3435
rect 45150 -3555 45195 -3435
rect 45315 -3555 45360 -3435
rect 45480 -3555 45525 -3435
rect 45645 -3555 45700 -3435
rect 45820 -3555 45865 -3435
rect 45985 -3555 46030 -3435
rect 46150 -3555 46195 -3435
rect 46315 -3555 46370 -3435
rect 46490 -3555 46535 -3435
rect 46655 -3555 46700 -3435
rect 46820 -3555 46865 -3435
rect 46985 -3555 47040 -3435
rect 47160 -3555 47205 -3435
rect 47325 -3555 47370 -3435
rect 47490 -3555 47535 -3435
rect 47655 -3555 47865 -3435
rect 47985 -3555 48040 -3435
rect 48160 -3555 48205 -3435
rect 48325 -3555 48370 -3435
rect 48490 -3555 48535 -3435
rect 48655 -3555 48710 -3435
rect 48830 -3555 48875 -3435
rect 48995 -3555 49040 -3435
rect 49160 -3555 49205 -3435
rect 49325 -3555 49380 -3435
rect 49500 -3555 49545 -3435
rect 49665 -3555 49710 -3435
rect 49830 -3555 49875 -3435
rect 49995 -3555 50050 -3435
rect 50170 -3555 50215 -3435
rect 50335 -3555 50380 -3435
rect 50500 -3555 50545 -3435
rect 50665 -3555 50720 -3435
rect 50840 -3555 50885 -3435
rect 51005 -3555 51050 -3435
rect 51170 -3555 51215 -3435
rect 51335 -3555 51390 -3435
rect 51510 -3555 51555 -3435
rect 51675 -3555 51720 -3435
rect 51840 -3555 51885 -3435
rect 52005 -3555 52060 -3435
rect 52180 -3555 52225 -3435
rect 52345 -3555 52390 -3435
rect 52510 -3555 52555 -3435
rect 52675 -3555 52730 -3435
rect 52850 -3555 52895 -3435
rect 53015 -3555 53060 -3435
rect 53180 -3555 53225 -3435
rect 53345 -3555 53370 -3435
rect 30770 -3600 53370 -3555
rect 30770 -3720 30795 -3600
rect 30915 -3720 30970 -3600
rect 31090 -3720 31135 -3600
rect 31255 -3720 31300 -3600
rect 31420 -3720 31465 -3600
rect 31585 -3720 31640 -3600
rect 31760 -3720 31805 -3600
rect 31925 -3720 31970 -3600
rect 32090 -3720 32135 -3600
rect 32255 -3720 32310 -3600
rect 32430 -3720 32475 -3600
rect 32595 -3720 32640 -3600
rect 32760 -3720 32805 -3600
rect 32925 -3720 32980 -3600
rect 33100 -3720 33145 -3600
rect 33265 -3720 33310 -3600
rect 33430 -3720 33475 -3600
rect 33595 -3720 33650 -3600
rect 33770 -3720 33815 -3600
rect 33935 -3720 33980 -3600
rect 34100 -3720 34145 -3600
rect 34265 -3720 34320 -3600
rect 34440 -3720 34485 -3600
rect 34605 -3720 34650 -3600
rect 34770 -3720 34815 -3600
rect 34935 -3720 34990 -3600
rect 35110 -3720 35155 -3600
rect 35275 -3720 35320 -3600
rect 35440 -3720 35485 -3600
rect 35605 -3720 35660 -3600
rect 35780 -3720 35825 -3600
rect 35945 -3720 35990 -3600
rect 36110 -3720 36155 -3600
rect 36275 -3720 36485 -3600
rect 36605 -3720 36660 -3600
rect 36780 -3720 36825 -3600
rect 36945 -3720 36990 -3600
rect 37110 -3720 37155 -3600
rect 37275 -3720 37330 -3600
rect 37450 -3720 37495 -3600
rect 37615 -3720 37660 -3600
rect 37780 -3720 37825 -3600
rect 37945 -3720 38000 -3600
rect 38120 -3720 38165 -3600
rect 38285 -3720 38330 -3600
rect 38450 -3720 38495 -3600
rect 38615 -3720 38670 -3600
rect 38790 -3720 38835 -3600
rect 38955 -3720 39000 -3600
rect 39120 -3720 39165 -3600
rect 39285 -3720 39340 -3600
rect 39460 -3720 39505 -3600
rect 39625 -3720 39670 -3600
rect 39790 -3720 39835 -3600
rect 39955 -3720 40010 -3600
rect 40130 -3720 40175 -3600
rect 40295 -3720 40340 -3600
rect 40460 -3720 40505 -3600
rect 40625 -3720 40680 -3600
rect 40800 -3720 40845 -3600
rect 40965 -3720 41010 -3600
rect 41130 -3720 41175 -3600
rect 41295 -3720 41350 -3600
rect 41470 -3720 41515 -3600
rect 41635 -3720 41680 -3600
rect 41800 -3720 41845 -3600
rect 41965 -3720 42175 -3600
rect 42295 -3720 42350 -3600
rect 42470 -3720 42515 -3600
rect 42635 -3720 42680 -3600
rect 42800 -3720 42845 -3600
rect 42965 -3720 43020 -3600
rect 43140 -3720 43185 -3600
rect 43305 -3720 43350 -3600
rect 43470 -3720 43515 -3600
rect 43635 -3720 43690 -3600
rect 43810 -3720 43855 -3600
rect 43975 -3720 44020 -3600
rect 44140 -3720 44185 -3600
rect 44305 -3720 44360 -3600
rect 44480 -3720 44525 -3600
rect 44645 -3720 44690 -3600
rect 44810 -3720 44855 -3600
rect 44975 -3720 45030 -3600
rect 45150 -3720 45195 -3600
rect 45315 -3720 45360 -3600
rect 45480 -3720 45525 -3600
rect 45645 -3720 45700 -3600
rect 45820 -3720 45865 -3600
rect 45985 -3720 46030 -3600
rect 46150 -3720 46195 -3600
rect 46315 -3720 46370 -3600
rect 46490 -3720 46535 -3600
rect 46655 -3720 46700 -3600
rect 46820 -3720 46865 -3600
rect 46985 -3720 47040 -3600
rect 47160 -3720 47205 -3600
rect 47325 -3720 47370 -3600
rect 47490 -3720 47535 -3600
rect 47655 -3720 47865 -3600
rect 47985 -3720 48040 -3600
rect 48160 -3720 48205 -3600
rect 48325 -3720 48370 -3600
rect 48490 -3720 48535 -3600
rect 48655 -3720 48710 -3600
rect 48830 -3720 48875 -3600
rect 48995 -3720 49040 -3600
rect 49160 -3720 49205 -3600
rect 49325 -3720 49380 -3600
rect 49500 -3720 49545 -3600
rect 49665 -3720 49710 -3600
rect 49830 -3720 49875 -3600
rect 49995 -3720 50050 -3600
rect 50170 -3720 50215 -3600
rect 50335 -3720 50380 -3600
rect 50500 -3720 50545 -3600
rect 50665 -3720 50720 -3600
rect 50840 -3720 50885 -3600
rect 51005 -3720 51050 -3600
rect 51170 -3720 51215 -3600
rect 51335 -3720 51390 -3600
rect 51510 -3720 51555 -3600
rect 51675 -3720 51720 -3600
rect 51840 -3720 51885 -3600
rect 52005 -3720 52060 -3600
rect 52180 -3720 52225 -3600
rect 52345 -3720 52390 -3600
rect 52510 -3720 52555 -3600
rect 52675 -3720 52730 -3600
rect 52850 -3720 52895 -3600
rect 53015 -3720 53060 -3600
rect 53180 -3720 53225 -3600
rect 53345 -3720 53370 -3600
rect 30770 -3765 53370 -3720
rect 30770 -3885 30795 -3765
rect 30915 -3885 30970 -3765
rect 31090 -3885 31135 -3765
rect 31255 -3885 31300 -3765
rect 31420 -3885 31465 -3765
rect 31585 -3885 31640 -3765
rect 31760 -3885 31805 -3765
rect 31925 -3885 31970 -3765
rect 32090 -3885 32135 -3765
rect 32255 -3885 32310 -3765
rect 32430 -3885 32475 -3765
rect 32595 -3885 32640 -3765
rect 32760 -3885 32805 -3765
rect 32925 -3885 32980 -3765
rect 33100 -3885 33145 -3765
rect 33265 -3885 33310 -3765
rect 33430 -3885 33475 -3765
rect 33595 -3885 33650 -3765
rect 33770 -3885 33815 -3765
rect 33935 -3885 33980 -3765
rect 34100 -3885 34145 -3765
rect 34265 -3885 34320 -3765
rect 34440 -3885 34485 -3765
rect 34605 -3885 34650 -3765
rect 34770 -3885 34815 -3765
rect 34935 -3885 34990 -3765
rect 35110 -3885 35155 -3765
rect 35275 -3885 35320 -3765
rect 35440 -3885 35485 -3765
rect 35605 -3885 35660 -3765
rect 35780 -3885 35825 -3765
rect 35945 -3885 35990 -3765
rect 36110 -3885 36155 -3765
rect 36275 -3885 36485 -3765
rect 36605 -3885 36660 -3765
rect 36780 -3885 36825 -3765
rect 36945 -3885 36990 -3765
rect 37110 -3885 37155 -3765
rect 37275 -3885 37330 -3765
rect 37450 -3885 37495 -3765
rect 37615 -3885 37660 -3765
rect 37780 -3885 37825 -3765
rect 37945 -3885 38000 -3765
rect 38120 -3885 38165 -3765
rect 38285 -3885 38330 -3765
rect 38450 -3885 38495 -3765
rect 38615 -3885 38670 -3765
rect 38790 -3885 38835 -3765
rect 38955 -3885 39000 -3765
rect 39120 -3885 39165 -3765
rect 39285 -3885 39340 -3765
rect 39460 -3885 39505 -3765
rect 39625 -3885 39670 -3765
rect 39790 -3885 39835 -3765
rect 39955 -3885 40010 -3765
rect 40130 -3885 40175 -3765
rect 40295 -3885 40340 -3765
rect 40460 -3885 40505 -3765
rect 40625 -3885 40680 -3765
rect 40800 -3885 40845 -3765
rect 40965 -3885 41010 -3765
rect 41130 -3885 41175 -3765
rect 41295 -3885 41350 -3765
rect 41470 -3885 41515 -3765
rect 41635 -3885 41680 -3765
rect 41800 -3885 41845 -3765
rect 41965 -3885 42175 -3765
rect 42295 -3885 42350 -3765
rect 42470 -3885 42515 -3765
rect 42635 -3885 42680 -3765
rect 42800 -3885 42845 -3765
rect 42965 -3885 43020 -3765
rect 43140 -3885 43185 -3765
rect 43305 -3885 43350 -3765
rect 43470 -3885 43515 -3765
rect 43635 -3885 43690 -3765
rect 43810 -3885 43855 -3765
rect 43975 -3885 44020 -3765
rect 44140 -3885 44185 -3765
rect 44305 -3885 44360 -3765
rect 44480 -3885 44525 -3765
rect 44645 -3885 44690 -3765
rect 44810 -3885 44855 -3765
rect 44975 -3885 45030 -3765
rect 45150 -3885 45195 -3765
rect 45315 -3885 45360 -3765
rect 45480 -3885 45525 -3765
rect 45645 -3885 45700 -3765
rect 45820 -3885 45865 -3765
rect 45985 -3885 46030 -3765
rect 46150 -3885 46195 -3765
rect 46315 -3885 46370 -3765
rect 46490 -3885 46535 -3765
rect 46655 -3885 46700 -3765
rect 46820 -3885 46865 -3765
rect 46985 -3885 47040 -3765
rect 47160 -3885 47205 -3765
rect 47325 -3885 47370 -3765
rect 47490 -3885 47535 -3765
rect 47655 -3885 47865 -3765
rect 47985 -3885 48040 -3765
rect 48160 -3885 48205 -3765
rect 48325 -3885 48370 -3765
rect 48490 -3885 48535 -3765
rect 48655 -3885 48710 -3765
rect 48830 -3885 48875 -3765
rect 48995 -3885 49040 -3765
rect 49160 -3885 49205 -3765
rect 49325 -3885 49380 -3765
rect 49500 -3885 49545 -3765
rect 49665 -3885 49710 -3765
rect 49830 -3885 49875 -3765
rect 49995 -3885 50050 -3765
rect 50170 -3885 50215 -3765
rect 50335 -3885 50380 -3765
rect 50500 -3885 50545 -3765
rect 50665 -3885 50720 -3765
rect 50840 -3885 50885 -3765
rect 51005 -3885 51050 -3765
rect 51170 -3885 51215 -3765
rect 51335 -3885 51390 -3765
rect 51510 -3885 51555 -3765
rect 51675 -3885 51720 -3765
rect 51840 -3885 51885 -3765
rect 52005 -3885 52060 -3765
rect 52180 -3885 52225 -3765
rect 52345 -3885 52390 -3765
rect 52510 -3885 52555 -3765
rect 52675 -3885 52730 -3765
rect 52850 -3885 52895 -3765
rect 53015 -3885 53060 -3765
rect 53180 -3885 53225 -3765
rect 53345 -3885 53370 -3765
rect 30770 -3940 53370 -3885
rect 30770 -4060 30795 -3940
rect 30915 -4060 30970 -3940
rect 31090 -4060 31135 -3940
rect 31255 -4060 31300 -3940
rect 31420 -4060 31465 -3940
rect 31585 -4060 31640 -3940
rect 31760 -4060 31805 -3940
rect 31925 -4060 31970 -3940
rect 32090 -4060 32135 -3940
rect 32255 -4060 32310 -3940
rect 32430 -4060 32475 -3940
rect 32595 -4060 32640 -3940
rect 32760 -4060 32805 -3940
rect 32925 -4060 32980 -3940
rect 33100 -4060 33145 -3940
rect 33265 -4060 33310 -3940
rect 33430 -4060 33475 -3940
rect 33595 -4060 33650 -3940
rect 33770 -4060 33815 -3940
rect 33935 -4060 33980 -3940
rect 34100 -4060 34145 -3940
rect 34265 -4060 34320 -3940
rect 34440 -4060 34485 -3940
rect 34605 -4060 34650 -3940
rect 34770 -4060 34815 -3940
rect 34935 -4060 34990 -3940
rect 35110 -4060 35155 -3940
rect 35275 -4060 35320 -3940
rect 35440 -4060 35485 -3940
rect 35605 -4060 35660 -3940
rect 35780 -4060 35825 -3940
rect 35945 -4060 35990 -3940
rect 36110 -4060 36155 -3940
rect 36275 -4060 36485 -3940
rect 36605 -4060 36660 -3940
rect 36780 -4060 36825 -3940
rect 36945 -4060 36990 -3940
rect 37110 -4060 37155 -3940
rect 37275 -4060 37330 -3940
rect 37450 -4060 37495 -3940
rect 37615 -4060 37660 -3940
rect 37780 -4060 37825 -3940
rect 37945 -4060 38000 -3940
rect 38120 -4060 38165 -3940
rect 38285 -4060 38330 -3940
rect 38450 -4060 38495 -3940
rect 38615 -4060 38670 -3940
rect 38790 -4060 38835 -3940
rect 38955 -4060 39000 -3940
rect 39120 -4060 39165 -3940
rect 39285 -4060 39340 -3940
rect 39460 -4060 39505 -3940
rect 39625 -4060 39670 -3940
rect 39790 -4060 39835 -3940
rect 39955 -4060 40010 -3940
rect 40130 -4060 40175 -3940
rect 40295 -4060 40340 -3940
rect 40460 -4060 40505 -3940
rect 40625 -4060 40680 -3940
rect 40800 -4060 40845 -3940
rect 40965 -4060 41010 -3940
rect 41130 -4060 41175 -3940
rect 41295 -4060 41350 -3940
rect 41470 -4060 41515 -3940
rect 41635 -4060 41680 -3940
rect 41800 -4060 41845 -3940
rect 41965 -4060 42175 -3940
rect 42295 -4060 42350 -3940
rect 42470 -4060 42515 -3940
rect 42635 -4060 42680 -3940
rect 42800 -4060 42845 -3940
rect 42965 -4060 43020 -3940
rect 43140 -4060 43185 -3940
rect 43305 -4060 43350 -3940
rect 43470 -4060 43515 -3940
rect 43635 -4060 43690 -3940
rect 43810 -4060 43855 -3940
rect 43975 -4060 44020 -3940
rect 44140 -4060 44185 -3940
rect 44305 -4060 44360 -3940
rect 44480 -4060 44525 -3940
rect 44645 -4060 44690 -3940
rect 44810 -4060 44855 -3940
rect 44975 -4060 45030 -3940
rect 45150 -4060 45195 -3940
rect 45315 -4060 45360 -3940
rect 45480 -4060 45525 -3940
rect 45645 -4060 45700 -3940
rect 45820 -4060 45865 -3940
rect 45985 -4060 46030 -3940
rect 46150 -4060 46195 -3940
rect 46315 -4060 46370 -3940
rect 46490 -4060 46535 -3940
rect 46655 -4060 46700 -3940
rect 46820 -4060 46865 -3940
rect 46985 -4060 47040 -3940
rect 47160 -4060 47205 -3940
rect 47325 -4060 47370 -3940
rect 47490 -4060 47535 -3940
rect 47655 -4060 47865 -3940
rect 47985 -4060 48040 -3940
rect 48160 -4060 48205 -3940
rect 48325 -4060 48370 -3940
rect 48490 -4060 48535 -3940
rect 48655 -4060 48710 -3940
rect 48830 -4060 48875 -3940
rect 48995 -4060 49040 -3940
rect 49160 -4060 49205 -3940
rect 49325 -4060 49380 -3940
rect 49500 -4060 49545 -3940
rect 49665 -4060 49710 -3940
rect 49830 -4060 49875 -3940
rect 49995 -4060 50050 -3940
rect 50170 -4060 50215 -3940
rect 50335 -4060 50380 -3940
rect 50500 -4060 50545 -3940
rect 50665 -4060 50720 -3940
rect 50840 -4060 50885 -3940
rect 51005 -4060 51050 -3940
rect 51170 -4060 51215 -3940
rect 51335 -4060 51390 -3940
rect 51510 -4060 51555 -3940
rect 51675 -4060 51720 -3940
rect 51840 -4060 51885 -3940
rect 52005 -4060 52060 -3940
rect 52180 -4060 52225 -3940
rect 52345 -4060 52390 -3940
rect 52510 -4060 52555 -3940
rect 52675 -4060 52730 -3940
rect 52850 -4060 52895 -3940
rect 53015 -4060 53060 -3940
rect 53180 -4060 53225 -3940
rect 53345 -4060 53370 -3940
rect 30770 -4270 53370 -4060
rect 30770 -4390 30795 -4270
rect 30915 -4390 30960 -4270
rect 31080 -4390 31125 -4270
rect 31245 -4390 31290 -4270
rect 31410 -4390 31465 -4270
rect 31585 -4390 31630 -4270
rect 31750 -4390 31795 -4270
rect 31915 -4390 31960 -4270
rect 32080 -4390 32135 -4270
rect 32255 -4390 32300 -4270
rect 32420 -4390 32465 -4270
rect 32585 -4390 32630 -4270
rect 32750 -4390 32805 -4270
rect 32925 -4390 32970 -4270
rect 33090 -4390 33135 -4270
rect 33255 -4390 33300 -4270
rect 33420 -4390 33475 -4270
rect 33595 -4390 33640 -4270
rect 33760 -4390 33805 -4270
rect 33925 -4390 33970 -4270
rect 34090 -4390 34145 -4270
rect 34265 -4390 34310 -4270
rect 34430 -4390 34475 -4270
rect 34595 -4390 34640 -4270
rect 34760 -4390 34815 -4270
rect 34935 -4390 34980 -4270
rect 35100 -4390 35145 -4270
rect 35265 -4390 35310 -4270
rect 35430 -4390 35485 -4270
rect 35605 -4390 35650 -4270
rect 35770 -4390 35815 -4270
rect 35935 -4390 35980 -4270
rect 36100 -4390 36155 -4270
rect 36275 -4390 36485 -4270
rect 36605 -4390 36650 -4270
rect 36770 -4390 36815 -4270
rect 36935 -4390 36980 -4270
rect 37100 -4390 37155 -4270
rect 37275 -4390 37320 -4270
rect 37440 -4390 37485 -4270
rect 37605 -4390 37650 -4270
rect 37770 -4390 37825 -4270
rect 37945 -4390 37990 -4270
rect 38110 -4390 38155 -4270
rect 38275 -4390 38320 -4270
rect 38440 -4390 38495 -4270
rect 38615 -4390 38660 -4270
rect 38780 -4390 38825 -4270
rect 38945 -4390 38990 -4270
rect 39110 -4390 39165 -4270
rect 39285 -4390 39330 -4270
rect 39450 -4390 39495 -4270
rect 39615 -4390 39660 -4270
rect 39780 -4390 39835 -4270
rect 39955 -4390 40000 -4270
rect 40120 -4390 40165 -4270
rect 40285 -4390 40330 -4270
rect 40450 -4390 40505 -4270
rect 40625 -4390 40670 -4270
rect 40790 -4390 40835 -4270
rect 40955 -4390 41000 -4270
rect 41120 -4390 41175 -4270
rect 41295 -4390 41340 -4270
rect 41460 -4390 41505 -4270
rect 41625 -4390 41670 -4270
rect 41790 -4390 41845 -4270
rect 41965 -4390 42175 -4270
rect 42295 -4390 42340 -4270
rect 42460 -4390 42505 -4270
rect 42625 -4390 42670 -4270
rect 42790 -4390 42845 -4270
rect 42965 -4390 43010 -4270
rect 43130 -4390 43175 -4270
rect 43295 -4390 43340 -4270
rect 43460 -4390 43515 -4270
rect 43635 -4390 43680 -4270
rect 43800 -4390 43845 -4270
rect 43965 -4390 44010 -4270
rect 44130 -4390 44185 -4270
rect 44305 -4390 44350 -4270
rect 44470 -4390 44515 -4270
rect 44635 -4390 44680 -4270
rect 44800 -4390 44855 -4270
rect 44975 -4390 45020 -4270
rect 45140 -4390 45185 -4270
rect 45305 -4390 45350 -4270
rect 45470 -4390 45525 -4270
rect 45645 -4390 45690 -4270
rect 45810 -4390 45855 -4270
rect 45975 -4390 46020 -4270
rect 46140 -4390 46195 -4270
rect 46315 -4390 46360 -4270
rect 46480 -4390 46525 -4270
rect 46645 -4390 46690 -4270
rect 46810 -4390 46865 -4270
rect 46985 -4390 47030 -4270
rect 47150 -4390 47195 -4270
rect 47315 -4390 47360 -4270
rect 47480 -4390 47535 -4270
rect 47655 -4390 47865 -4270
rect 47985 -4390 48030 -4270
rect 48150 -4390 48195 -4270
rect 48315 -4390 48360 -4270
rect 48480 -4390 48535 -4270
rect 48655 -4390 48700 -4270
rect 48820 -4390 48865 -4270
rect 48985 -4390 49030 -4270
rect 49150 -4390 49205 -4270
rect 49325 -4390 49370 -4270
rect 49490 -4390 49535 -4270
rect 49655 -4390 49700 -4270
rect 49820 -4390 49875 -4270
rect 49995 -4390 50040 -4270
rect 50160 -4390 50205 -4270
rect 50325 -4390 50370 -4270
rect 50490 -4390 50545 -4270
rect 50665 -4390 50710 -4270
rect 50830 -4390 50875 -4270
rect 50995 -4390 51040 -4270
rect 51160 -4390 51215 -4270
rect 51335 -4390 51380 -4270
rect 51500 -4390 51545 -4270
rect 51665 -4390 51710 -4270
rect 51830 -4390 51885 -4270
rect 52005 -4390 52050 -4270
rect 52170 -4390 52215 -4270
rect 52335 -4390 52380 -4270
rect 52500 -4390 52555 -4270
rect 52675 -4390 52720 -4270
rect 52840 -4390 52885 -4270
rect 53005 -4390 53050 -4270
rect 53170 -4390 53225 -4270
rect 53345 -4390 53370 -4270
rect 30770 -4445 53370 -4390
rect 30770 -4565 30795 -4445
rect 30915 -4565 30960 -4445
rect 31080 -4565 31125 -4445
rect 31245 -4565 31290 -4445
rect 31410 -4565 31465 -4445
rect 31585 -4565 31630 -4445
rect 31750 -4565 31795 -4445
rect 31915 -4565 31960 -4445
rect 32080 -4565 32135 -4445
rect 32255 -4565 32300 -4445
rect 32420 -4565 32465 -4445
rect 32585 -4565 32630 -4445
rect 32750 -4565 32805 -4445
rect 32925 -4565 32970 -4445
rect 33090 -4565 33135 -4445
rect 33255 -4565 33300 -4445
rect 33420 -4565 33475 -4445
rect 33595 -4565 33640 -4445
rect 33760 -4565 33805 -4445
rect 33925 -4565 33970 -4445
rect 34090 -4565 34145 -4445
rect 34265 -4565 34310 -4445
rect 34430 -4565 34475 -4445
rect 34595 -4565 34640 -4445
rect 34760 -4565 34815 -4445
rect 34935 -4565 34980 -4445
rect 35100 -4565 35145 -4445
rect 35265 -4565 35310 -4445
rect 35430 -4565 35485 -4445
rect 35605 -4565 35650 -4445
rect 35770 -4565 35815 -4445
rect 35935 -4565 35980 -4445
rect 36100 -4565 36155 -4445
rect 36275 -4565 36485 -4445
rect 36605 -4565 36650 -4445
rect 36770 -4565 36815 -4445
rect 36935 -4565 36980 -4445
rect 37100 -4565 37155 -4445
rect 37275 -4565 37320 -4445
rect 37440 -4565 37485 -4445
rect 37605 -4565 37650 -4445
rect 37770 -4565 37825 -4445
rect 37945 -4565 37990 -4445
rect 38110 -4565 38155 -4445
rect 38275 -4565 38320 -4445
rect 38440 -4565 38495 -4445
rect 38615 -4565 38660 -4445
rect 38780 -4565 38825 -4445
rect 38945 -4565 38990 -4445
rect 39110 -4565 39165 -4445
rect 39285 -4565 39330 -4445
rect 39450 -4565 39495 -4445
rect 39615 -4565 39660 -4445
rect 39780 -4565 39835 -4445
rect 39955 -4565 40000 -4445
rect 40120 -4565 40165 -4445
rect 40285 -4565 40330 -4445
rect 40450 -4565 40505 -4445
rect 40625 -4565 40670 -4445
rect 40790 -4565 40835 -4445
rect 40955 -4565 41000 -4445
rect 41120 -4565 41175 -4445
rect 41295 -4565 41340 -4445
rect 41460 -4565 41505 -4445
rect 41625 -4565 41670 -4445
rect 41790 -4565 41845 -4445
rect 41965 -4565 42175 -4445
rect 42295 -4565 42340 -4445
rect 42460 -4565 42505 -4445
rect 42625 -4565 42670 -4445
rect 42790 -4565 42845 -4445
rect 42965 -4565 43010 -4445
rect 43130 -4565 43175 -4445
rect 43295 -4565 43340 -4445
rect 43460 -4565 43515 -4445
rect 43635 -4565 43680 -4445
rect 43800 -4565 43845 -4445
rect 43965 -4565 44010 -4445
rect 44130 -4565 44185 -4445
rect 44305 -4565 44350 -4445
rect 44470 -4565 44515 -4445
rect 44635 -4565 44680 -4445
rect 44800 -4565 44855 -4445
rect 44975 -4565 45020 -4445
rect 45140 -4565 45185 -4445
rect 45305 -4565 45350 -4445
rect 45470 -4565 45525 -4445
rect 45645 -4565 45690 -4445
rect 45810 -4565 45855 -4445
rect 45975 -4565 46020 -4445
rect 46140 -4565 46195 -4445
rect 46315 -4565 46360 -4445
rect 46480 -4565 46525 -4445
rect 46645 -4565 46690 -4445
rect 46810 -4565 46865 -4445
rect 46985 -4565 47030 -4445
rect 47150 -4565 47195 -4445
rect 47315 -4565 47360 -4445
rect 47480 -4565 47535 -4445
rect 47655 -4565 47865 -4445
rect 47985 -4565 48030 -4445
rect 48150 -4565 48195 -4445
rect 48315 -4565 48360 -4445
rect 48480 -4565 48535 -4445
rect 48655 -4565 48700 -4445
rect 48820 -4565 48865 -4445
rect 48985 -4565 49030 -4445
rect 49150 -4565 49205 -4445
rect 49325 -4565 49370 -4445
rect 49490 -4565 49535 -4445
rect 49655 -4565 49700 -4445
rect 49820 -4565 49875 -4445
rect 49995 -4565 50040 -4445
rect 50160 -4565 50205 -4445
rect 50325 -4565 50370 -4445
rect 50490 -4565 50545 -4445
rect 50665 -4565 50710 -4445
rect 50830 -4565 50875 -4445
rect 50995 -4565 51040 -4445
rect 51160 -4565 51215 -4445
rect 51335 -4565 51380 -4445
rect 51500 -4565 51545 -4445
rect 51665 -4565 51710 -4445
rect 51830 -4565 51885 -4445
rect 52005 -4565 52050 -4445
rect 52170 -4565 52215 -4445
rect 52335 -4565 52380 -4445
rect 52500 -4565 52555 -4445
rect 52675 -4565 52720 -4445
rect 52840 -4565 52885 -4445
rect 53005 -4565 53050 -4445
rect 53170 -4565 53225 -4445
rect 53345 -4565 53370 -4445
rect 30770 -4610 53370 -4565
rect 30770 -4730 30795 -4610
rect 30915 -4730 30960 -4610
rect 31080 -4730 31125 -4610
rect 31245 -4730 31290 -4610
rect 31410 -4730 31465 -4610
rect 31585 -4730 31630 -4610
rect 31750 -4730 31795 -4610
rect 31915 -4730 31960 -4610
rect 32080 -4730 32135 -4610
rect 32255 -4730 32300 -4610
rect 32420 -4730 32465 -4610
rect 32585 -4730 32630 -4610
rect 32750 -4730 32805 -4610
rect 32925 -4730 32970 -4610
rect 33090 -4730 33135 -4610
rect 33255 -4730 33300 -4610
rect 33420 -4730 33475 -4610
rect 33595 -4730 33640 -4610
rect 33760 -4730 33805 -4610
rect 33925 -4730 33970 -4610
rect 34090 -4730 34145 -4610
rect 34265 -4730 34310 -4610
rect 34430 -4730 34475 -4610
rect 34595 -4730 34640 -4610
rect 34760 -4730 34815 -4610
rect 34935 -4730 34980 -4610
rect 35100 -4730 35145 -4610
rect 35265 -4730 35310 -4610
rect 35430 -4730 35485 -4610
rect 35605 -4730 35650 -4610
rect 35770 -4730 35815 -4610
rect 35935 -4730 35980 -4610
rect 36100 -4730 36155 -4610
rect 36275 -4730 36485 -4610
rect 36605 -4730 36650 -4610
rect 36770 -4730 36815 -4610
rect 36935 -4730 36980 -4610
rect 37100 -4730 37155 -4610
rect 37275 -4730 37320 -4610
rect 37440 -4730 37485 -4610
rect 37605 -4730 37650 -4610
rect 37770 -4730 37825 -4610
rect 37945 -4730 37990 -4610
rect 38110 -4730 38155 -4610
rect 38275 -4730 38320 -4610
rect 38440 -4730 38495 -4610
rect 38615 -4730 38660 -4610
rect 38780 -4730 38825 -4610
rect 38945 -4730 38990 -4610
rect 39110 -4730 39165 -4610
rect 39285 -4730 39330 -4610
rect 39450 -4730 39495 -4610
rect 39615 -4730 39660 -4610
rect 39780 -4730 39835 -4610
rect 39955 -4730 40000 -4610
rect 40120 -4730 40165 -4610
rect 40285 -4730 40330 -4610
rect 40450 -4730 40505 -4610
rect 40625 -4730 40670 -4610
rect 40790 -4730 40835 -4610
rect 40955 -4730 41000 -4610
rect 41120 -4730 41175 -4610
rect 41295 -4730 41340 -4610
rect 41460 -4730 41505 -4610
rect 41625 -4730 41670 -4610
rect 41790 -4730 41845 -4610
rect 41965 -4730 42175 -4610
rect 42295 -4730 42340 -4610
rect 42460 -4730 42505 -4610
rect 42625 -4730 42670 -4610
rect 42790 -4730 42845 -4610
rect 42965 -4730 43010 -4610
rect 43130 -4730 43175 -4610
rect 43295 -4730 43340 -4610
rect 43460 -4730 43515 -4610
rect 43635 -4730 43680 -4610
rect 43800 -4730 43845 -4610
rect 43965 -4730 44010 -4610
rect 44130 -4730 44185 -4610
rect 44305 -4730 44350 -4610
rect 44470 -4730 44515 -4610
rect 44635 -4730 44680 -4610
rect 44800 -4730 44855 -4610
rect 44975 -4730 45020 -4610
rect 45140 -4730 45185 -4610
rect 45305 -4730 45350 -4610
rect 45470 -4730 45525 -4610
rect 45645 -4730 45690 -4610
rect 45810 -4730 45855 -4610
rect 45975 -4730 46020 -4610
rect 46140 -4730 46195 -4610
rect 46315 -4730 46360 -4610
rect 46480 -4730 46525 -4610
rect 46645 -4730 46690 -4610
rect 46810 -4730 46865 -4610
rect 46985 -4730 47030 -4610
rect 47150 -4730 47195 -4610
rect 47315 -4730 47360 -4610
rect 47480 -4730 47535 -4610
rect 47655 -4730 47865 -4610
rect 47985 -4730 48030 -4610
rect 48150 -4730 48195 -4610
rect 48315 -4730 48360 -4610
rect 48480 -4730 48535 -4610
rect 48655 -4730 48700 -4610
rect 48820 -4730 48865 -4610
rect 48985 -4730 49030 -4610
rect 49150 -4730 49205 -4610
rect 49325 -4730 49370 -4610
rect 49490 -4730 49535 -4610
rect 49655 -4730 49700 -4610
rect 49820 -4730 49875 -4610
rect 49995 -4730 50040 -4610
rect 50160 -4730 50205 -4610
rect 50325 -4730 50370 -4610
rect 50490 -4730 50545 -4610
rect 50665 -4730 50710 -4610
rect 50830 -4730 50875 -4610
rect 50995 -4730 51040 -4610
rect 51160 -4730 51215 -4610
rect 51335 -4730 51380 -4610
rect 51500 -4730 51545 -4610
rect 51665 -4730 51710 -4610
rect 51830 -4730 51885 -4610
rect 52005 -4730 52050 -4610
rect 52170 -4730 52215 -4610
rect 52335 -4730 52380 -4610
rect 52500 -4730 52555 -4610
rect 52675 -4730 52720 -4610
rect 52840 -4730 52885 -4610
rect 53005 -4730 53050 -4610
rect 53170 -4730 53225 -4610
rect 53345 -4730 53370 -4610
rect 30770 -4775 53370 -4730
rect 30770 -4895 30795 -4775
rect 30915 -4895 30960 -4775
rect 31080 -4895 31125 -4775
rect 31245 -4895 31290 -4775
rect 31410 -4895 31465 -4775
rect 31585 -4895 31630 -4775
rect 31750 -4895 31795 -4775
rect 31915 -4895 31960 -4775
rect 32080 -4895 32135 -4775
rect 32255 -4895 32300 -4775
rect 32420 -4895 32465 -4775
rect 32585 -4895 32630 -4775
rect 32750 -4895 32805 -4775
rect 32925 -4895 32970 -4775
rect 33090 -4895 33135 -4775
rect 33255 -4895 33300 -4775
rect 33420 -4895 33475 -4775
rect 33595 -4895 33640 -4775
rect 33760 -4895 33805 -4775
rect 33925 -4895 33970 -4775
rect 34090 -4895 34145 -4775
rect 34265 -4895 34310 -4775
rect 34430 -4895 34475 -4775
rect 34595 -4895 34640 -4775
rect 34760 -4895 34815 -4775
rect 34935 -4895 34980 -4775
rect 35100 -4895 35145 -4775
rect 35265 -4895 35310 -4775
rect 35430 -4895 35485 -4775
rect 35605 -4895 35650 -4775
rect 35770 -4895 35815 -4775
rect 35935 -4895 35980 -4775
rect 36100 -4895 36155 -4775
rect 36275 -4895 36485 -4775
rect 36605 -4895 36650 -4775
rect 36770 -4895 36815 -4775
rect 36935 -4895 36980 -4775
rect 37100 -4895 37155 -4775
rect 37275 -4895 37320 -4775
rect 37440 -4895 37485 -4775
rect 37605 -4895 37650 -4775
rect 37770 -4895 37825 -4775
rect 37945 -4895 37990 -4775
rect 38110 -4895 38155 -4775
rect 38275 -4895 38320 -4775
rect 38440 -4895 38495 -4775
rect 38615 -4895 38660 -4775
rect 38780 -4895 38825 -4775
rect 38945 -4895 38990 -4775
rect 39110 -4895 39165 -4775
rect 39285 -4895 39330 -4775
rect 39450 -4895 39495 -4775
rect 39615 -4895 39660 -4775
rect 39780 -4895 39835 -4775
rect 39955 -4895 40000 -4775
rect 40120 -4895 40165 -4775
rect 40285 -4895 40330 -4775
rect 40450 -4895 40505 -4775
rect 40625 -4895 40670 -4775
rect 40790 -4895 40835 -4775
rect 40955 -4895 41000 -4775
rect 41120 -4895 41175 -4775
rect 41295 -4895 41340 -4775
rect 41460 -4895 41505 -4775
rect 41625 -4895 41670 -4775
rect 41790 -4895 41845 -4775
rect 41965 -4895 42175 -4775
rect 42295 -4895 42340 -4775
rect 42460 -4895 42505 -4775
rect 42625 -4895 42670 -4775
rect 42790 -4895 42845 -4775
rect 42965 -4895 43010 -4775
rect 43130 -4895 43175 -4775
rect 43295 -4895 43340 -4775
rect 43460 -4895 43515 -4775
rect 43635 -4895 43680 -4775
rect 43800 -4895 43845 -4775
rect 43965 -4895 44010 -4775
rect 44130 -4895 44185 -4775
rect 44305 -4895 44350 -4775
rect 44470 -4895 44515 -4775
rect 44635 -4895 44680 -4775
rect 44800 -4895 44855 -4775
rect 44975 -4895 45020 -4775
rect 45140 -4895 45185 -4775
rect 45305 -4895 45350 -4775
rect 45470 -4895 45525 -4775
rect 45645 -4895 45690 -4775
rect 45810 -4895 45855 -4775
rect 45975 -4895 46020 -4775
rect 46140 -4895 46195 -4775
rect 46315 -4895 46360 -4775
rect 46480 -4895 46525 -4775
rect 46645 -4895 46690 -4775
rect 46810 -4895 46865 -4775
rect 46985 -4895 47030 -4775
rect 47150 -4895 47195 -4775
rect 47315 -4895 47360 -4775
rect 47480 -4895 47535 -4775
rect 47655 -4895 47865 -4775
rect 47985 -4895 48030 -4775
rect 48150 -4895 48195 -4775
rect 48315 -4895 48360 -4775
rect 48480 -4895 48535 -4775
rect 48655 -4895 48700 -4775
rect 48820 -4895 48865 -4775
rect 48985 -4895 49030 -4775
rect 49150 -4895 49205 -4775
rect 49325 -4895 49370 -4775
rect 49490 -4895 49535 -4775
rect 49655 -4895 49700 -4775
rect 49820 -4895 49875 -4775
rect 49995 -4895 50040 -4775
rect 50160 -4895 50205 -4775
rect 50325 -4895 50370 -4775
rect 50490 -4895 50545 -4775
rect 50665 -4895 50710 -4775
rect 50830 -4895 50875 -4775
rect 50995 -4895 51040 -4775
rect 51160 -4895 51215 -4775
rect 51335 -4895 51380 -4775
rect 51500 -4895 51545 -4775
rect 51665 -4895 51710 -4775
rect 51830 -4895 51885 -4775
rect 52005 -4895 52050 -4775
rect 52170 -4895 52215 -4775
rect 52335 -4895 52380 -4775
rect 52500 -4895 52555 -4775
rect 52675 -4895 52720 -4775
rect 52840 -4895 52885 -4775
rect 53005 -4895 53050 -4775
rect 53170 -4895 53225 -4775
rect 53345 -4895 53370 -4775
rect 30770 -4940 53370 -4895
rect 30770 -5060 30795 -4940
rect 30915 -5060 30960 -4940
rect 31080 -5060 31125 -4940
rect 31245 -5060 31290 -4940
rect 31410 -5060 31465 -4940
rect 31585 -5060 31630 -4940
rect 31750 -5060 31795 -4940
rect 31915 -5060 31960 -4940
rect 32080 -5060 32135 -4940
rect 32255 -5060 32300 -4940
rect 32420 -5060 32465 -4940
rect 32585 -5060 32630 -4940
rect 32750 -5060 32805 -4940
rect 32925 -5060 32970 -4940
rect 33090 -5060 33135 -4940
rect 33255 -5060 33300 -4940
rect 33420 -5060 33475 -4940
rect 33595 -5060 33640 -4940
rect 33760 -5060 33805 -4940
rect 33925 -5060 33970 -4940
rect 34090 -5060 34145 -4940
rect 34265 -5060 34310 -4940
rect 34430 -5060 34475 -4940
rect 34595 -5060 34640 -4940
rect 34760 -5060 34815 -4940
rect 34935 -5060 34980 -4940
rect 35100 -5060 35145 -4940
rect 35265 -5060 35310 -4940
rect 35430 -5060 35485 -4940
rect 35605 -5060 35650 -4940
rect 35770 -5060 35815 -4940
rect 35935 -5060 35980 -4940
rect 36100 -5060 36155 -4940
rect 36275 -5060 36485 -4940
rect 36605 -5060 36650 -4940
rect 36770 -5060 36815 -4940
rect 36935 -5060 36980 -4940
rect 37100 -5060 37155 -4940
rect 37275 -5060 37320 -4940
rect 37440 -5060 37485 -4940
rect 37605 -5060 37650 -4940
rect 37770 -5060 37825 -4940
rect 37945 -5060 37990 -4940
rect 38110 -5060 38155 -4940
rect 38275 -5060 38320 -4940
rect 38440 -5060 38495 -4940
rect 38615 -5060 38660 -4940
rect 38780 -5060 38825 -4940
rect 38945 -5060 38990 -4940
rect 39110 -5060 39165 -4940
rect 39285 -5060 39330 -4940
rect 39450 -5060 39495 -4940
rect 39615 -5060 39660 -4940
rect 39780 -5060 39835 -4940
rect 39955 -5060 40000 -4940
rect 40120 -5060 40165 -4940
rect 40285 -5060 40330 -4940
rect 40450 -5060 40505 -4940
rect 40625 -5060 40670 -4940
rect 40790 -5060 40835 -4940
rect 40955 -5060 41000 -4940
rect 41120 -5060 41175 -4940
rect 41295 -5060 41340 -4940
rect 41460 -5060 41505 -4940
rect 41625 -5060 41670 -4940
rect 41790 -5060 41845 -4940
rect 41965 -5060 42175 -4940
rect 42295 -5060 42340 -4940
rect 42460 -5060 42505 -4940
rect 42625 -5060 42670 -4940
rect 42790 -5060 42845 -4940
rect 42965 -5060 43010 -4940
rect 43130 -5060 43175 -4940
rect 43295 -5060 43340 -4940
rect 43460 -5060 43515 -4940
rect 43635 -5060 43680 -4940
rect 43800 -5060 43845 -4940
rect 43965 -5060 44010 -4940
rect 44130 -5060 44185 -4940
rect 44305 -5060 44350 -4940
rect 44470 -5060 44515 -4940
rect 44635 -5060 44680 -4940
rect 44800 -5060 44855 -4940
rect 44975 -5060 45020 -4940
rect 45140 -5060 45185 -4940
rect 45305 -5060 45350 -4940
rect 45470 -5060 45525 -4940
rect 45645 -5060 45690 -4940
rect 45810 -5060 45855 -4940
rect 45975 -5060 46020 -4940
rect 46140 -5060 46195 -4940
rect 46315 -5060 46360 -4940
rect 46480 -5060 46525 -4940
rect 46645 -5060 46690 -4940
rect 46810 -5060 46865 -4940
rect 46985 -5060 47030 -4940
rect 47150 -5060 47195 -4940
rect 47315 -5060 47360 -4940
rect 47480 -5060 47535 -4940
rect 47655 -5060 47865 -4940
rect 47985 -5060 48030 -4940
rect 48150 -5060 48195 -4940
rect 48315 -5060 48360 -4940
rect 48480 -5060 48535 -4940
rect 48655 -5060 48700 -4940
rect 48820 -5060 48865 -4940
rect 48985 -5060 49030 -4940
rect 49150 -5060 49205 -4940
rect 49325 -5060 49370 -4940
rect 49490 -5060 49535 -4940
rect 49655 -5060 49700 -4940
rect 49820 -5060 49875 -4940
rect 49995 -5060 50040 -4940
rect 50160 -5060 50205 -4940
rect 50325 -5060 50370 -4940
rect 50490 -5060 50545 -4940
rect 50665 -5060 50710 -4940
rect 50830 -5060 50875 -4940
rect 50995 -5060 51040 -4940
rect 51160 -5060 51215 -4940
rect 51335 -5060 51380 -4940
rect 51500 -5060 51545 -4940
rect 51665 -5060 51710 -4940
rect 51830 -5060 51885 -4940
rect 52005 -5060 52050 -4940
rect 52170 -5060 52215 -4940
rect 52335 -5060 52380 -4940
rect 52500 -5060 52555 -4940
rect 52675 -5060 52720 -4940
rect 52840 -5060 52885 -4940
rect 53005 -5060 53050 -4940
rect 53170 -5060 53225 -4940
rect 53345 -5060 53370 -4940
rect 30770 -5115 53370 -5060
rect 30770 -5235 30795 -5115
rect 30915 -5235 30960 -5115
rect 31080 -5235 31125 -5115
rect 31245 -5235 31290 -5115
rect 31410 -5235 31465 -5115
rect 31585 -5235 31630 -5115
rect 31750 -5235 31795 -5115
rect 31915 -5235 31960 -5115
rect 32080 -5235 32135 -5115
rect 32255 -5235 32300 -5115
rect 32420 -5235 32465 -5115
rect 32585 -5235 32630 -5115
rect 32750 -5235 32805 -5115
rect 32925 -5235 32970 -5115
rect 33090 -5235 33135 -5115
rect 33255 -5235 33300 -5115
rect 33420 -5235 33475 -5115
rect 33595 -5235 33640 -5115
rect 33760 -5235 33805 -5115
rect 33925 -5235 33970 -5115
rect 34090 -5235 34145 -5115
rect 34265 -5235 34310 -5115
rect 34430 -5235 34475 -5115
rect 34595 -5235 34640 -5115
rect 34760 -5235 34815 -5115
rect 34935 -5235 34980 -5115
rect 35100 -5235 35145 -5115
rect 35265 -5235 35310 -5115
rect 35430 -5235 35485 -5115
rect 35605 -5235 35650 -5115
rect 35770 -5235 35815 -5115
rect 35935 -5235 35980 -5115
rect 36100 -5235 36155 -5115
rect 36275 -5235 36485 -5115
rect 36605 -5235 36650 -5115
rect 36770 -5235 36815 -5115
rect 36935 -5235 36980 -5115
rect 37100 -5235 37155 -5115
rect 37275 -5235 37320 -5115
rect 37440 -5235 37485 -5115
rect 37605 -5235 37650 -5115
rect 37770 -5235 37825 -5115
rect 37945 -5235 37990 -5115
rect 38110 -5235 38155 -5115
rect 38275 -5235 38320 -5115
rect 38440 -5235 38495 -5115
rect 38615 -5235 38660 -5115
rect 38780 -5235 38825 -5115
rect 38945 -5235 38990 -5115
rect 39110 -5235 39165 -5115
rect 39285 -5235 39330 -5115
rect 39450 -5235 39495 -5115
rect 39615 -5235 39660 -5115
rect 39780 -5235 39835 -5115
rect 39955 -5235 40000 -5115
rect 40120 -5235 40165 -5115
rect 40285 -5235 40330 -5115
rect 40450 -5235 40505 -5115
rect 40625 -5235 40670 -5115
rect 40790 -5235 40835 -5115
rect 40955 -5235 41000 -5115
rect 41120 -5235 41175 -5115
rect 41295 -5235 41340 -5115
rect 41460 -5235 41505 -5115
rect 41625 -5235 41670 -5115
rect 41790 -5235 41845 -5115
rect 41965 -5235 42175 -5115
rect 42295 -5235 42340 -5115
rect 42460 -5235 42505 -5115
rect 42625 -5235 42670 -5115
rect 42790 -5235 42845 -5115
rect 42965 -5235 43010 -5115
rect 43130 -5235 43175 -5115
rect 43295 -5235 43340 -5115
rect 43460 -5235 43515 -5115
rect 43635 -5235 43680 -5115
rect 43800 -5235 43845 -5115
rect 43965 -5235 44010 -5115
rect 44130 -5235 44185 -5115
rect 44305 -5235 44350 -5115
rect 44470 -5235 44515 -5115
rect 44635 -5235 44680 -5115
rect 44800 -5235 44855 -5115
rect 44975 -5235 45020 -5115
rect 45140 -5235 45185 -5115
rect 45305 -5235 45350 -5115
rect 45470 -5235 45525 -5115
rect 45645 -5235 45690 -5115
rect 45810 -5235 45855 -5115
rect 45975 -5235 46020 -5115
rect 46140 -5235 46195 -5115
rect 46315 -5235 46360 -5115
rect 46480 -5235 46525 -5115
rect 46645 -5235 46690 -5115
rect 46810 -5235 46865 -5115
rect 46985 -5235 47030 -5115
rect 47150 -5235 47195 -5115
rect 47315 -5235 47360 -5115
rect 47480 -5235 47535 -5115
rect 47655 -5235 47865 -5115
rect 47985 -5235 48030 -5115
rect 48150 -5235 48195 -5115
rect 48315 -5235 48360 -5115
rect 48480 -5235 48535 -5115
rect 48655 -5235 48700 -5115
rect 48820 -5235 48865 -5115
rect 48985 -5235 49030 -5115
rect 49150 -5235 49205 -5115
rect 49325 -5235 49370 -5115
rect 49490 -5235 49535 -5115
rect 49655 -5235 49700 -5115
rect 49820 -5235 49875 -5115
rect 49995 -5235 50040 -5115
rect 50160 -5235 50205 -5115
rect 50325 -5235 50370 -5115
rect 50490 -5235 50545 -5115
rect 50665 -5235 50710 -5115
rect 50830 -5235 50875 -5115
rect 50995 -5235 51040 -5115
rect 51160 -5235 51215 -5115
rect 51335 -5235 51380 -5115
rect 51500 -5235 51545 -5115
rect 51665 -5235 51710 -5115
rect 51830 -5235 51885 -5115
rect 52005 -5235 52050 -5115
rect 52170 -5235 52215 -5115
rect 52335 -5235 52380 -5115
rect 52500 -5235 52555 -5115
rect 52675 -5235 52720 -5115
rect 52840 -5235 52885 -5115
rect 53005 -5235 53050 -5115
rect 53170 -5235 53225 -5115
rect 53345 -5235 53370 -5115
rect 30770 -5280 53370 -5235
rect 30770 -5400 30795 -5280
rect 30915 -5400 30960 -5280
rect 31080 -5400 31125 -5280
rect 31245 -5400 31290 -5280
rect 31410 -5400 31465 -5280
rect 31585 -5400 31630 -5280
rect 31750 -5400 31795 -5280
rect 31915 -5400 31960 -5280
rect 32080 -5400 32135 -5280
rect 32255 -5400 32300 -5280
rect 32420 -5400 32465 -5280
rect 32585 -5400 32630 -5280
rect 32750 -5400 32805 -5280
rect 32925 -5400 32970 -5280
rect 33090 -5400 33135 -5280
rect 33255 -5400 33300 -5280
rect 33420 -5400 33475 -5280
rect 33595 -5400 33640 -5280
rect 33760 -5400 33805 -5280
rect 33925 -5400 33970 -5280
rect 34090 -5400 34145 -5280
rect 34265 -5400 34310 -5280
rect 34430 -5400 34475 -5280
rect 34595 -5400 34640 -5280
rect 34760 -5400 34815 -5280
rect 34935 -5400 34980 -5280
rect 35100 -5400 35145 -5280
rect 35265 -5400 35310 -5280
rect 35430 -5400 35485 -5280
rect 35605 -5400 35650 -5280
rect 35770 -5400 35815 -5280
rect 35935 -5400 35980 -5280
rect 36100 -5400 36155 -5280
rect 36275 -5400 36485 -5280
rect 36605 -5400 36650 -5280
rect 36770 -5400 36815 -5280
rect 36935 -5400 36980 -5280
rect 37100 -5400 37155 -5280
rect 37275 -5400 37320 -5280
rect 37440 -5400 37485 -5280
rect 37605 -5400 37650 -5280
rect 37770 -5400 37825 -5280
rect 37945 -5400 37990 -5280
rect 38110 -5400 38155 -5280
rect 38275 -5400 38320 -5280
rect 38440 -5400 38495 -5280
rect 38615 -5400 38660 -5280
rect 38780 -5400 38825 -5280
rect 38945 -5400 38990 -5280
rect 39110 -5400 39165 -5280
rect 39285 -5400 39330 -5280
rect 39450 -5400 39495 -5280
rect 39615 -5400 39660 -5280
rect 39780 -5400 39835 -5280
rect 39955 -5400 40000 -5280
rect 40120 -5400 40165 -5280
rect 40285 -5400 40330 -5280
rect 40450 -5400 40505 -5280
rect 40625 -5400 40670 -5280
rect 40790 -5400 40835 -5280
rect 40955 -5400 41000 -5280
rect 41120 -5400 41175 -5280
rect 41295 -5400 41340 -5280
rect 41460 -5400 41505 -5280
rect 41625 -5400 41670 -5280
rect 41790 -5400 41845 -5280
rect 41965 -5400 42175 -5280
rect 42295 -5400 42340 -5280
rect 42460 -5400 42505 -5280
rect 42625 -5400 42670 -5280
rect 42790 -5400 42845 -5280
rect 42965 -5400 43010 -5280
rect 43130 -5400 43175 -5280
rect 43295 -5400 43340 -5280
rect 43460 -5400 43515 -5280
rect 43635 -5400 43680 -5280
rect 43800 -5400 43845 -5280
rect 43965 -5400 44010 -5280
rect 44130 -5400 44185 -5280
rect 44305 -5400 44350 -5280
rect 44470 -5400 44515 -5280
rect 44635 -5400 44680 -5280
rect 44800 -5400 44855 -5280
rect 44975 -5400 45020 -5280
rect 45140 -5400 45185 -5280
rect 45305 -5400 45350 -5280
rect 45470 -5400 45525 -5280
rect 45645 -5400 45690 -5280
rect 45810 -5400 45855 -5280
rect 45975 -5400 46020 -5280
rect 46140 -5400 46195 -5280
rect 46315 -5400 46360 -5280
rect 46480 -5400 46525 -5280
rect 46645 -5400 46690 -5280
rect 46810 -5400 46865 -5280
rect 46985 -5400 47030 -5280
rect 47150 -5400 47195 -5280
rect 47315 -5400 47360 -5280
rect 47480 -5400 47535 -5280
rect 47655 -5400 47865 -5280
rect 47985 -5400 48030 -5280
rect 48150 -5400 48195 -5280
rect 48315 -5400 48360 -5280
rect 48480 -5400 48535 -5280
rect 48655 -5400 48700 -5280
rect 48820 -5400 48865 -5280
rect 48985 -5400 49030 -5280
rect 49150 -5400 49205 -5280
rect 49325 -5400 49370 -5280
rect 49490 -5400 49535 -5280
rect 49655 -5400 49700 -5280
rect 49820 -5400 49875 -5280
rect 49995 -5400 50040 -5280
rect 50160 -5400 50205 -5280
rect 50325 -5400 50370 -5280
rect 50490 -5400 50545 -5280
rect 50665 -5400 50710 -5280
rect 50830 -5400 50875 -5280
rect 50995 -5400 51040 -5280
rect 51160 -5400 51215 -5280
rect 51335 -5400 51380 -5280
rect 51500 -5400 51545 -5280
rect 51665 -5400 51710 -5280
rect 51830 -5400 51885 -5280
rect 52005 -5400 52050 -5280
rect 52170 -5400 52215 -5280
rect 52335 -5400 52380 -5280
rect 52500 -5400 52555 -5280
rect 52675 -5400 52720 -5280
rect 52840 -5400 52885 -5280
rect 53005 -5400 53050 -5280
rect 53170 -5400 53225 -5280
rect 53345 -5400 53370 -5280
rect 30770 -5445 53370 -5400
rect 30770 -5565 30795 -5445
rect 30915 -5565 30960 -5445
rect 31080 -5565 31125 -5445
rect 31245 -5565 31290 -5445
rect 31410 -5565 31465 -5445
rect 31585 -5565 31630 -5445
rect 31750 -5565 31795 -5445
rect 31915 -5565 31960 -5445
rect 32080 -5565 32135 -5445
rect 32255 -5565 32300 -5445
rect 32420 -5565 32465 -5445
rect 32585 -5565 32630 -5445
rect 32750 -5565 32805 -5445
rect 32925 -5565 32970 -5445
rect 33090 -5565 33135 -5445
rect 33255 -5565 33300 -5445
rect 33420 -5565 33475 -5445
rect 33595 -5565 33640 -5445
rect 33760 -5565 33805 -5445
rect 33925 -5565 33970 -5445
rect 34090 -5565 34145 -5445
rect 34265 -5565 34310 -5445
rect 34430 -5565 34475 -5445
rect 34595 -5565 34640 -5445
rect 34760 -5565 34815 -5445
rect 34935 -5565 34980 -5445
rect 35100 -5565 35145 -5445
rect 35265 -5565 35310 -5445
rect 35430 -5565 35485 -5445
rect 35605 -5565 35650 -5445
rect 35770 -5565 35815 -5445
rect 35935 -5565 35980 -5445
rect 36100 -5565 36155 -5445
rect 36275 -5565 36485 -5445
rect 36605 -5565 36650 -5445
rect 36770 -5565 36815 -5445
rect 36935 -5565 36980 -5445
rect 37100 -5565 37155 -5445
rect 37275 -5565 37320 -5445
rect 37440 -5565 37485 -5445
rect 37605 -5565 37650 -5445
rect 37770 -5565 37825 -5445
rect 37945 -5565 37990 -5445
rect 38110 -5565 38155 -5445
rect 38275 -5565 38320 -5445
rect 38440 -5565 38495 -5445
rect 38615 -5565 38660 -5445
rect 38780 -5565 38825 -5445
rect 38945 -5565 38990 -5445
rect 39110 -5565 39165 -5445
rect 39285 -5565 39330 -5445
rect 39450 -5565 39495 -5445
rect 39615 -5565 39660 -5445
rect 39780 -5565 39835 -5445
rect 39955 -5565 40000 -5445
rect 40120 -5565 40165 -5445
rect 40285 -5565 40330 -5445
rect 40450 -5565 40505 -5445
rect 40625 -5565 40670 -5445
rect 40790 -5565 40835 -5445
rect 40955 -5565 41000 -5445
rect 41120 -5565 41175 -5445
rect 41295 -5565 41340 -5445
rect 41460 -5565 41505 -5445
rect 41625 -5565 41670 -5445
rect 41790 -5565 41845 -5445
rect 41965 -5565 42175 -5445
rect 42295 -5565 42340 -5445
rect 42460 -5565 42505 -5445
rect 42625 -5565 42670 -5445
rect 42790 -5565 42845 -5445
rect 42965 -5565 43010 -5445
rect 43130 -5565 43175 -5445
rect 43295 -5565 43340 -5445
rect 43460 -5565 43515 -5445
rect 43635 -5565 43680 -5445
rect 43800 -5565 43845 -5445
rect 43965 -5565 44010 -5445
rect 44130 -5565 44185 -5445
rect 44305 -5565 44350 -5445
rect 44470 -5565 44515 -5445
rect 44635 -5565 44680 -5445
rect 44800 -5565 44855 -5445
rect 44975 -5565 45020 -5445
rect 45140 -5565 45185 -5445
rect 45305 -5565 45350 -5445
rect 45470 -5565 45525 -5445
rect 45645 -5565 45690 -5445
rect 45810 -5565 45855 -5445
rect 45975 -5565 46020 -5445
rect 46140 -5565 46195 -5445
rect 46315 -5565 46360 -5445
rect 46480 -5565 46525 -5445
rect 46645 -5565 46690 -5445
rect 46810 -5565 46865 -5445
rect 46985 -5565 47030 -5445
rect 47150 -5565 47195 -5445
rect 47315 -5565 47360 -5445
rect 47480 -5565 47535 -5445
rect 47655 -5565 47865 -5445
rect 47985 -5565 48030 -5445
rect 48150 -5565 48195 -5445
rect 48315 -5565 48360 -5445
rect 48480 -5565 48535 -5445
rect 48655 -5565 48700 -5445
rect 48820 -5565 48865 -5445
rect 48985 -5565 49030 -5445
rect 49150 -5565 49205 -5445
rect 49325 -5565 49370 -5445
rect 49490 -5565 49535 -5445
rect 49655 -5565 49700 -5445
rect 49820 -5565 49875 -5445
rect 49995 -5565 50040 -5445
rect 50160 -5565 50205 -5445
rect 50325 -5565 50370 -5445
rect 50490 -5565 50545 -5445
rect 50665 -5565 50710 -5445
rect 50830 -5565 50875 -5445
rect 50995 -5565 51040 -5445
rect 51160 -5565 51215 -5445
rect 51335 -5565 51380 -5445
rect 51500 -5565 51545 -5445
rect 51665 -5565 51710 -5445
rect 51830 -5565 51885 -5445
rect 52005 -5565 52050 -5445
rect 52170 -5565 52215 -5445
rect 52335 -5565 52380 -5445
rect 52500 -5565 52555 -5445
rect 52675 -5565 52720 -5445
rect 52840 -5565 52885 -5445
rect 53005 -5565 53050 -5445
rect 53170 -5565 53225 -5445
rect 53345 -5565 53370 -5445
rect 30770 -5610 53370 -5565
rect 30770 -5730 30795 -5610
rect 30915 -5730 30960 -5610
rect 31080 -5730 31125 -5610
rect 31245 -5730 31290 -5610
rect 31410 -5730 31465 -5610
rect 31585 -5730 31630 -5610
rect 31750 -5730 31795 -5610
rect 31915 -5730 31960 -5610
rect 32080 -5730 32135 -5610
rect 32255 -5730 32300 -5610
rect 32420 -5730 32465 -5610
rect 32585 -5730 32630 -5610
rect 32750 -5730 32805 -5610
rect 32925 -5730 32970 -5610
rect 33090 -5730 33135 -5610
rect 33255 -5730 33300 -5610
rect 33420 -5730 33475 -5610
rect 33595 -5730 33640 -5610
rect 33760 -5730 33805 -5610
rect 33925 -5730 33970 -5610
rect 34090 -5730 34145 -5610
rect 34265 -5730 34310 -5610
rect 34430 -5730 34475 -5610
rect 34595 -5730 34640 -5610
rect 34760 -5730 34815 -5610
rect 34935 -5730 34980 -5610
rect 35100 -5730 35145 -5610
rect 35265 -5730 35310 -5610
rect 35430 -5730 35485 -5610
rect 35605 -5730 35650 -5610
rect 35770 -5730 35815 -5610
rect 35935 -5730 35980 -5610
rect 36100 -5730 36155 -5610
rect 36275 -5730 36485 -5610
rect 36605 -5730 36650 -5610
rect 36770 -5730 36815 -5610
rect 36935 -5730 36980 -5610
rect 37100 -5730 37155 -5610
rect 37275 -5730 37320 -5610
rect 37440 -5730 37485 -5610
rect 37605 -5730 37650 -5610
rect 37770 -5730 37825 -5610
rect 37945 -5730 37990 -5610
rect 38110 -5730 38155 -5610
rect 38275 -5730 38320 -5610
rect 38440 -5730 38495 -5610
rect 38615 -5730 38660 -5610
rect 38780 -5730 38825 -5610
rect 38945 -5730 38990 -5610
rect 39110 -5730 39165 -5610
rect 39285 -5730 39330 -5610
rect 39450 -5730 39495 -5610
rect 39615 -5730 39660 -5610
rect 39780 -5730 39835 -5610
rect 39955 -5730 40000 -5610
rect 40120 -5730 40165 -5610
rect 40285 -5730 40330 -5610
rect 40450 -5730 40505 -5610
rect 40625 -5730 40670 -5610
rect 40790 -5730 40835 -5610
rect 40955 -5730 41000 -5610
rect 41120 -5730 41175 -5610
rect 41295 -5730 41340 -5610
rect 41460 -5730 41505 -5610
rect 41625 -5730 41670 -5610
rect 41790 -5730 41845 -5610
rect 41965 -5730 42175 -5610
rect 42295 -5730 42340 -5610
rect 42460 -5730 42505 -5610
rect 42625 -5730 42670 -5610
rect 42790 -5730 42845 -5610
rect 42965 -5730 43010 -5610
rect 43130 -5730 43175 -5610
rect 43295 -5730 43340 -5610
rect 43460 -5730 43515 -5610
rect 43635 -5730 43680 -5610
rect 43800 -5730 43845 -5610
rect 43965 -5730 44010 -5610
rect 44130 -5730 44185 -5610
rect 44305 -5730 44350 -5610
rect 44470 -5730 44515 -5610
rect 44635 -5730 44680 -5610
rect 44800 -5730 44855 -5610
rect 44975 -5730 45020 -5610
rect 45140 -5730 45185 -5610
rect 45305 -5730 45350 -5610
rect 45470 -5730 45525 -5610
rect 45645 -5730 45690 -5610
rect 45810 -5730 45855 -5610
rect 45975 -5730 46020 -5610
rect 46140 -5730 46195 -5610
rect 46315 -5730 46360 -5610
rect 46480 -5730 46525 -5610
rect 46645 -5730 46690 -5610
rect 46810 -5730 46865 -5610
rect 46985 -5730 47030 -5610
rect 47150 -5730 47195 -5610
rect 47315 -5730 47360 -5610
rect 47480 -5730 47535 -5610
rect 47655 -5730 47865 -5610
rect 47985 -5730 48030 -5610
rect 48150 -5730 48195 -5610
rect 48315 -5730 48360 -5610
rect 48480 -5730 48535 -5610
rect 48655 -5730 48700 -5610
rect 48820 -5730 48865 -5610
rect 48985 -5730 49030 -5610
rect 49150 -5730 49205 -5610
rect 49325 -5730 49370 -5610
rect 49490 -5730 49535 -5610
rect 49655 -5730 49700 -5610
rect 49820 -5730 49875 -5610
rect 49995 -5730 50040 -5610
rect 50160 -5730 50205 -5610
rect 50325 -5730 50370 -5610
rect 50490 -5730 50545 -5610
rect 50665 -5730 50710 -5610
rect 50830 -5730 50875 -5610
rect 50995 -5730 51040 -5610
rect 51160 -5730 51215 -5610
rect 51335 -5730 51380 -5610
rect 51500 -5730 51545 -5610
rect 51665 -5730 51710 -5610
rect 51830 -5730 51885 -5610
rect 52005 -5730 52050 -5610
rect 52170 -5730 52215 -5610
rect 52335 -5730 52380 -5610
rect 52500 -5730 52555 -5610
rect 52675 -5730 52720 -5610
rect 52840 -5730 52885 -5610
rect 53005 -5730 53050 -5610
rect 53170 -5730 53225 -5610
rect 53345 -5730 53370 -5610
rect 30770 -5785 53370 -5730
rect 30770 -5905 30795 -5785
rect 30915 -5905 30960 -5785
rect 31080 -5905 31125 -5785
rect 31245 -5905 31290 -5785
rect 31410 -5905 31465 -5785
rect 31585 -5905 31630 -5785
rect 31750 -5905 31795 -5785
rect 31915 -5905 31960 -5785
rect 32080 -5905 32135 -5785
rect 32255 -5905 32300 -5785
rect 32420 -5905 32465 -5785
rect 32585 -5905 32630 -5785
rect 32750 -5905 32805 -5785
rect 32925 -5905 32970 -5785
rect 33090 -5905 33135 -5785
rect 33255 -5905 33300 -5785
rect 33420 -5905 33475 -5785
rect 33595 -5905 33640 -5785
rect 33760 -5905 33805 -5785
rect 33925 -5905 33970 -5785
rect 34090 -5905 34145 -5785
rect 34265 -5905 34310 -5785
rect 34430 -5905 34475 -5785
rect 34595 -5905 34640 -5785
rect 34760 -5905 34815 -5785
rect 34935 -5905 34980 -5785
rect 35100 -5905 35145 -5785
rect 35265 -5905 35310 -5785
rect 35430 -5905 35485 -5785
rect 35605 -5905 35650 -5785
rect 35770 -5905 35815 -5785
rect 35935 -5905 35980 -5785
rect 36100 -5905 36155 -5785
rect 36275 -5905 36485 -5785
rect 36605 -5905 36650 -5785
rect 36770 -5905 36815 -5785
rect 36935 -5905 36980 -5785
rect 37100 -5905 37155 -5785
rect 37275 -5905 37320 -5785
rect 37440 -5905 37485 -5785
rect 37605 -5905 37650 -5785
rect 37770 -5905 37825 -5785
rect 37945 -5905 37990 -5785
rect 38110 -5905 38155 -5785
rect 38275 -5905 38320 -5785
rect 38440 -5905 38495 -5785
rect 38615 -5905 38660 -5785
rect 38780 -5905 38825 -5785
rect 38945 -5905 38990 -5785
rect 39110 -5905 39165 -5785
rect 39285 -5905 39330 -5785
rect 39450 -5905 39495 -5785
rect 39615 -5905 39660 -5785
rect 39780 -5905 39835 -5785
rect 39955 -5905 40000 -5785
rect 40120 -5905 40165 -5785
rect 40285 -5905 40330 -5785
rect 40450 -5905 40505 -5785
rect 40625 -5905 40670 -5785
rect 40790 -5905 40835 -5785
rect 40955 -5905 41000 -5785
rect 41120 -5905 41175 -5785
rect 41295 -5905 41340 -5785
rect 41460 -5905 41505 -5785
rect 41625 -5905 41670 -5785
rect 41790 -5905 41845 -5785
rect 41965 -5905 42175 -5785
rect 42295 -5905 42340 -5785
rect 42460 -5905 42505 -5785
rect 42625 -5905 42670 -5785
rect 42790 -5905 42845 -5785
rect 42965 -5905 43010 -5785
rect 43130 -5905 43175 -5785
rect 43295 -5905 43340 -5785
rect 43460 -5905 43515 -5785
rect 43635 -5905 43680 -5785
rect 43800 -5905 43845 -5785
rect 43965 -5905 44010 -5785
rect 44130 -5905 44185 -5785
rect 44305 -5905 44350 -5785
rect 44470 -5905 44515 -5785
rect 44635 -5905 44680 -5785
rect 44800 -5905 44855 -5785
rect 44975 -5905 45020 -5785
rect 45140 -5905 45185 -5785
rect 45305 -5905 45350 -5785
rect 45470 -5905 45525 -5785
rect 45645 -5905 45690 -5785
rect 45810 -5905 45855 -5785
rect 45975 -5905 46020 -5785
rect 46140 -5905 46195 -5785
rect 46315 -5905 46360 -5785
rect 46480 -5905 46525 -5785
rect 46645 -5905 46690 -5785
rect 46810 -5905 46865 -5785
rect 46985 -5905 47030 -5785
rect 47150 -5905 47195 -5785
rect 47315 -5905 47360 -5785
rect 47480 -5905 47535 -5785
rect 47655 -5905 47865 -5785
rect 47985 -5905 48030 -5785
rect 48150 -5905 48195 -5785
rect 48315 -5905 48360 -5785
rect 48480 -5905 48535 -5785
rect 48655 -5905 48700 -5785
rect 48820 -5905 48865 -5785
rect 48985 -5905 49030 -5785
rect 49150 -5905 49205 -5785
rect 49325 -5905 49370 -5785
rect 49490 -5905 49535 -5785
rect 49655 -5905 49700 -5785
rect 49820 -5905 49875 -5785
rect 49995 -5905 50040 -5785
rect 50160 -5905 50205 -5785
rect 50325 -5905 50370 -5785
rect 50490 -5905 50545 -5785
rect 50665 -5905 50710 -5785
rect 50830 -5905 50875 -5785
rect 50995 -5905 51040 -5785
rect 51160 -5905 51215 -5785
rect 51335 -5905 51380 -5785
rect 51500 -5905 51545 -5785
rect 51665 -5905 51710 -5785
rect 51830 -5905 51885 -5785
rect 52005 -5905 52050 -5785
rect 52170 -5905 52215 -5785
rect 52335 -5905 52380 -5785
rect 52500 -5905 52555 -5785
rect 52675 -5905 52720 -5785
rect 52840 -5905 52885 -5785
rect 53005 -5905 53050 -5785
rect 53170 -5905 53225 -5785
rect 53345 -5905 53370 -5785
rect 30770 -5950 53370 -5905
rect 30770 -6070 30795 -5950
rect 30915 -6070 30960 -5950
rect 31080 -6070 31125 -5950
rect 31245 -6070 31290 -5950
rect 31410 -6070 31465 -5950
rect 31585 -6070 31630 -5950
rect 31750 -6070 31795 -5950
rect 31915 -6070 31960 -5950
rect 32080 -6070 32135 -5950
rect 32255 -6070 32300 -5950
rect 32420 -6070 32465 -5950
rect 32585 -6070 32630 -5950
rect 32750 -6070 32805 -5950
rect 32925 -6070 32970 -5950
rect 33090 -6070 33135 -5950
rect 33255 -6070 33300 -5950
rect 33420 -6070 33475 -5950
rect 33595 -6070 33640 -5950
rect 33760 -6070 33805 -5950
rect 33925 -6070 33970 -5950
rect 34090 -6070 34145 -5950
rect 34265 -6070 34310 -5950
rect 34430 -6070 34475 -5950
rect 34595 -6070 34640 -5950
rect 34760 -6070 34815 -5950
rect 34935 -6070 34980 -5950
rect 35100 -6070 35145 -5950
rect 35265 -6070 35310 -5950
rect 35430 -6070 35485 -5950
rect 35605 -6070 35650 -5950
rect 35770 -6070 35815 -5950
rect 35935 -6070 35980 -5950
rect 36100 -6070 36155 -5950
rect 36275 -6070 36485 -5950
rect 36605 -6070 36650 -5950
rect 36770 -6070 36815 -5950
rect 36935 -6070 36980 -5950
rect 37100 -6070 37155 -5950
rect 37275 -6070 37320 -5950
rect 37440 -6070 37485 -5950
rect 37605 -6070 37650 -5950
rect 37770 -6070 37825 -5950
rect 37945 -6070 37990 -5950
rect 38110 -6070 38155 -5950
rect 38275 -6070 38320 -5950
rect 38440 -6070 38495 -5950
rect 38615 -6070 38660 -5950
rect 38780 -6070 38825 -5950
rect 38945 -6070 38990 -5950
rect 39110 -6070 39165 -5950
rect 39285 -6070 39330 -5950
rect 39450 -6070 39495 -5950
rect 39615 -6070 39660 -5950
rect 39780 -6070 39835 -5950
rect 39955 -6070 40000 -5950
rect 40120 -6070 40165 -5950
rect 40285 -6070 40330 -5950
rect 40450 -6070 40505 -5950
rect 40625 -6070 40670 -5950
rect 40790 -6070 40835 -5950
rect 40955 -6070 41000 -5950
rect 41120 -6070 41175 -5950
rect 41295 -6070 41340 -5950
rect 41460 -6070 41505 -5950
rect 41625 -6070 41670 -5950
rect 41790 -6070 41845 -5950
rect 41965 -6070 42175 -5950
rect 42295 -6070 42340 -5950
rect 42460 -6070 42505 -5950
rect 42625 -6070 42670 -5950
rect 42790 -6070 42845 -5950
rect 42965 -6070 43010 -5950
rect 43130 -6070 43175 -5950
rect 43295 -6070 43340 -5950
rect 43460 -6070 43515 -5950
rect 43635 -6070 43680 -5950
rect 43800 -6070 43845 -5950
rect 43965 -6070 44010 -5950
rect 44130 -6070 44185 -5950
rect 44305 -6070 44350 -5950
rect 44470 -6070 44515 -5950
rect 44635 -6070 44680 -5950
rect 44800 -6070 44855 -5950
rect 44975 -6070 45020 -5950
rect 45140 -6070 45185 -5950
rect 45305 -6070 45350 -5950
rect 45470 -6070 45525 -5950
rect 45645 -6070 45690 -5950
rect 45810 -6070 45855 -5950
rect 45975 -6070 46020 -5950
rect 46140 -6070 46195 -5950
rect 46315 -6070 46360 -5950
rect 46480 -6070 46525 -5950
rect 46645 -6070 46690 -5950
rect 46810 -6070 46865 -5950
rect 46985 -6070 47030 -5950
rect 47150 -6070 47195 -5950
rect 47315 -6070 47360 -5950
rect 47480 -6070 47535 -5950
rect 47655 -6070 47865 -5950
rect 47985 -6070 48030 -5950
rect 48150 -6070 48195 -5950
rect 48315 -6070 48360 -5950
rect 48480 -6070 48535 -5950
rect 48655 -6070 48700 -5950
rect 48820 -6070 48865 -5950
rect 48985 -6070 49030 -5950
rect 49150 -6070 49205 -5950
rect 49325 -6070 49370 -5950
rect 49490 -6070 49535 -5950
rect 49655 -6070 49700 -5950
rect 49820 -6070 49875 -5950
rect 49995 -6070 50040 -5950
rect 50160 -6070 50205 -5950
rect 50325 -6070 50370 -5950
rect 50490 -6070 50545 -5950
rect 50665 -6070 50710 -5950
rect 50830 -6070 50875 -5950
rect 50995 -6070 51040 -5950
rect 51160 -6070 51215 -5950
rect 51335 -6070 51380 -5950
rect 51500 -6070 51545 -5950
rect 51665 -6070 51710 -5950
rect 51830 -6070 51885 -5950
rect 52005 -6070 52050 -5950
rect 52170 -6070 52215 -5950
rect 52335 -6070 52380 -5950
rect 52500 -6070 52555 -5950
rect 52675 -6070 52720 -5950
rect 52840 -6070 52885 -5950
rect 53005 -6070 53050 -5950
rect 53170 -6070 53225 -5950
rect 53345 -6070 53370 -5950
rect 30770 -6115 53370 -6070
rect 30770 -6235 30795 -6115
rect 30915 -6235 30960 -6115
rect 31080 -6235 31125 -6115
rect 31245 -6235 31290 -6115
rect 31410 -6235 31465 -6115
rect 31585 -6235 31630 -6115
rect 31750 -6235 31795 -6115
rect 31915 -6235 31960 -6115
rect 32080 -6235 32135 -6115
rect 32255 -6235 32300 -6115
rect 32420 -6235 32465 -6115
rect 32585 -6235 32630 -6115
rect 32750 -6235 32805 -6115
rect 32925 -6235 32970 -6115
rect 33090 -6235 33135 -6115
rect 33255 -6235 33300 -6115
rect 33420 -6235 33475 -6115
rect 33595 -6235 33640 -6115
rect 33760 -6235 33805 -6115
rect 33925 -6235 33970 -6115
rect 34090 -6235 34145 -6115
rect 34265 -6235 34310 -6115
rect 34430 -6235 34475 -6115
rect 34595 -6235 34640 -6115
rect 34760 -6235 34815 -6115
rect 34935 -6235 34980 -6115
rect 35100 -6235 35145 -6115
rect 35265 -6235 35310 -6115
rect 35430 -6235 35485 -6115
rect 35605 -6235 35650 -6115
rect 35770 -6235 35815 -6115
rect 35935 -6235 35980 -6115
rect 36100 -6235 36155 -6115
rect 36275 -6235 36485 -6115
rect 36605 -6235 36650 -6115
rect 36770 -6235 36815 -6115
rect 36935 -6235 36980 -6115
rect 37100 -6235 37155 -6115
rect 37275 -6235 37320 -6115
rect 37440 -6235 37485 -6115
rect 37605 -6235 37650 -6115
rect 37770 -6235 37825 -6115
rect 37945 -6235 37990 -6115
rect 38110 -6235 38155 -6115
rect 38275 -6235 38320 -6115
rect 38440 -6235 38495 -6115
rect 38615 -6235 38660 -6115
rect 38780 -6235 38825 -6115
rect 38945 -6235 38990 -6115
rect 39110 -6235 39165 -6115
rect 39285 -6235 39330 -6115
rect 39450 -6235 39495 -6115
rect 39615 -6235 39660 -6115
rect 39780 -6235 39835 -6115
rect 39955 -6235 40000 -6115
rect 40120 -6235 40165 -6115
rect 40285 -6235 40330 -6115
rect 40450 -6235 40505 -6115
rect 40625 -6235 40670 -6115
rect 40790 -6235 40835 -6115
rect 40955 -6235 41000 -6115
rect 41120 -6235 41175 -6115
rect 41295 -6235 41340 -6115
rect 41460 -6235 41505 -6115
rect 41625 -6235 41670 -6115
rect 41790 -6235 41845 -6115
rect 41965 -6235 42175 -6115
rect 42295 -6235 42340 -6115
rect 42460 -6235 42505 -6115
rect 42625 -6235 42670 -6115
rect 42790 -6235 42845 -6115
rect 42965 -6235 43010 -6115
rect 43130 -6235 43175 -6115
rect 43295 -6235 43340 -6115
rect 43460 -6235 43515 -6115
rect 43635 -6235 43680 -6115
rect 43800 -6235 43845 -6115
rect 43965 -6235 44010 -6115
rect 44130 -6235 44185 -6115
rect 44305 -6235 44350 -6115
rect 44470 -6235 44515 -6115
rect 44635 -6235 44680 -6115
rect 44800 -6235 44855 -6115
rect 44975 -6235 45020 -6115
rect 45140 -6235 45185 -6115
rect 45305 -6235 45350 -6115
rect 45470 -6235 45525 -6115
rect 45645 -6235 45690 -6115
rect 45810 -6235 45855 -6115
rect 45975 -6235 46020 -6115
rect 46140 -6235 46195 -6115
rect 46315 -6235 46360 -6115
rect 46480 -6235 46525 -6115
rect 46645 -6235 46690 -6115
rect 46810 -6235 46865 -6115
rect 46985 -6235 47030 -6115
rect 47150 -6235 47195 -6115
rect 47315 -6235 47360 -6115
rect 47480 -6235 47535 -6115
rect 47655 -6235 47865 -6115
rect 47985 -6235 48030 -6115
rect 48150 -6235 48195 -6115
rect 48315 -6235 48360 -6115
rect 48480 -6235 48535 -6115
rect 48655 -6235 48700 -6115
rect 48820 -6235 48865 -6115
rect 48985 -6235 49030 -6115
rect 49150 -6235 49205 -6115
rect 49325 -6235 49370 -6115
rect 49490 -6235 49535 -6115
rect 49655 -6235 49700 -6115
rect 49820 -6235 49875 -6115
rect 49995 -6235 50040 -6115
rect 50160 -6235 50205 -6115
rect 50325 -6235 50370 -6115
rect 50490 -6235 50545 -6115
rect 50665 -6235 50710 -6115
rect 50830 -6235 50875 -6115
rect 50995 -6235 51040 -6115
rect 51160 -6235 51215 -6115
rect 51335 -6235 51380 -6115
rect 51500 -6235 51545 -6115
rect 51665 -6235 51710 -6115
rect 51830 -6235 51885 -6115
rect 52005 -6235 52050 -6115
rect 52170 -6235 52215 -6115
rect 52335 -6235 52380 -6115
rect 52500 -6235 52555 -6115
rect 52675 -6235 52720 -6115
rect 52840 -6235 52885 -6115
rect 53005 -6235 53050 -6115
rect 53170 -6235 53225 -6115
rect 53345 -6235 53370 -6115
rect 30770 -6280 53370 -6235
rect 30770 -6400 30795 -6280
rect 30915 -6400 30960 -6280
rect 31080 -6400 31125 -6280
rect 31245 -6400 31290 -6280
rect 31410 -6400 31465 -6280
rect 31585 -6400 31630 -6280
rect 31750 -6400 31795 -6280
rect 31915 -6400 31960 -6280
rect 32080 -6400 32135 -6280
rect 32255 -6400 32300 -6280
rect 32420 -6400 32465 -6280
rect 32585 -6400 32630 -6280
rect 32750 -6400 32805 -6280
rect 32925 -6400 32970 -6280
rect 33090 -6400 33135 -6280
rect 33255 -6400 33300 -6280
rect 33420 -6400 33475 -6280
rect 33595 -6400 33640 -6280
rect 33760 -6400 33805 -6280
rect 33925 -6400 33970 -6280
rect 34090 -6400 34145 -6280
rect 34265 -6400 34310 -6280
rect 34430 -6400 34475 -6280
rect 34595 -6400 34640 -6280
rect 34760 -6400 34815 -6280
rect 34935 -6400 34980 -6280
rect 35100 -6400 35145 -6280
rect 35265 -6400 35310 -6280
rect 35430 -6400 35485 -6280
rect 35605 -6400 35650 -6280
rect 35770 -6400 35815 -6280
rect 35935 -6400 35980 -6280
rect 36100 -6400 36155 -6280
rect 36275 -6400 36485 -6280
rect 36605 -6400 36650 -6280
rect 36770 -6400 36815 -6280
rect 36935 -6400 36980 -6280
rect 37100 -6400 37155 -6280
rect 37275 -6400 37320 -6280
rect 37440 -6400 37485 -6280
rect 37605 -6400 37650 -6280
rect 37770 -6400 37825 -6280
rect 37945 -6400 37990 -6280
rect 38110 -6400 38155 -6280
rect 38275 -6400 38320 -6280
rect 38440 -6400 38495 -6280
rect 38615 -6400 38660 -6280
rect 38780 -6400 38825 -6280
rect 38945 -6400 38990 -6280
rect 39110 -6400 39165 -6280
rect 39285 -6400 39330 -6280
rect 39450 -6400 39495 -6280
rect 39615 -6400 39660 -6280
rect 39780 -6400 39835 -6280
rect 39955 -6400 40000 -6280
rect 40120 -6400 40165 -6280
rect 40285 -6400 40330 -6280
rect 40450 -6400 40505 -6280
rect 40625 -6400 40670 -6280
rect 40790 -6400 40835 -6280
rect 40955 -6400 41000 -6280
rect 41120 -6400 41175 -6280
rect 41295 -6400 41340 -6280
rect 41460 -6400 41505 -6280
rect 41625 -6400 41670 -6280
rect 41790 -6400 41845 -6280
rect 41965 -6400 42175 -6280
rect 42295 -6400 42340 -6280
rect 42460 -6400 42505 -6280
rect 42625 -6400 42670 -6280
rect 42790 -6400 42845 -6280
rect 42965 -6400 43010 -6280
rect 43130 -6400 43175 -6280
rect 43295 -6400 43340 -6280
rect 43460 -6400 43515 -6280
rect 43635 -6400 43680 -6280
rect 43800 -6400 43845 -6280
rect 43965 -6400 44010 -6280
rect 44130 -6400 44185 -6280
rect 44305 -6400 44350 -6280
rect 44470 -6400 44515 -6280
rect 44635 -6400 44680 -6280
rect 44800 -6400 44855 -6280
rect 44975 -6400 45020 -6280
rect 45140 -6400 45185 -6280
rect 45305 -6400 45350 -6280
rect 45470 -6400 45525 -6280
rect 45645 -6400 45690 -6280
rect 45810 -6400 45855 -6280
rect 45975 -6400 46020 -6280
rect 46140 -6400 46195 -6280
rect 46315 -6400 46360 -6280
rect 46480 -6400 46525 -6280
rect 46645 -6400 46690 -6280
rect 46810 -6400 46865 -6280
rect 46985 -6400 47030 -6280
rect 47150 -6400 47195 -6280
rect 47315 -6400 47360 -6280
rect 47480 -6400 47535 -6280
rect 47655 -6400 47865 -6280
rect 47985 -6400 48030 -6280
rect 48150 -6400 48195 -6280
rect 48315 -6400 48360 -6280
rect 48480 -6400 48535 -6280
rect 48655 -6400 48700 -6280
rect 48820 -6400 48865 -6280
rect 48985 -6400 49030 -6280
rect 49150 -6400 49205 -6280
rect 49325 -6400 49370 -6280
rect 49490 -6400 49535 -6280
rect 49655 -6400 49700 -6280
rect 49820 -6400 49875 -6280
rect 49995 -6400 50040 -6280
rect 50160 -6400 50205 -6280
rect 50325 -6400 50370 -6280
rect 50490 -6400 50545 -6280
rect 50665 -6400 50710 -6280
rect 50830 -6400 50875 -6280
rect 50995 -6400 51040 -6280
rect 51160 -6400 51215 -6280
rect 51335 -6400 51380 -6280
rect 51500 -6400 51545 -6280
rect 51665 -6400 51710 -6280
rect 51830 -6400 51885 -6280
rect 52005 -6400 52050 -6280
rect 52170 -6400 52215 -6280
rect 52335 -6400 52380 -6280
rect 52500 -6400 52555 -6280
rect 52675 -6400 52720 -6280
rect 52840 -6400 52885 -6280
rect 53005 -6400 53050 -6280
rect 53170 -6400 53225 -6280
rect 53345 -6400 53370 -6280
rect 30770 -6455 53370 -6400
rect 30770 -6575 30795 -6455
rect 30915 -6575 30960 -6455
rect 31080 -6575 31125 -6455
rect 31245 -6575 31290 -6455
rect 31410 -6575 31465 -6455
rect 31585 -6575 31630 -6455
rect 31750 -6575 31795 -6455
rect 31915 -6575 31960 -6455
rect 32080 -6575 32135 -6455
rect 32255 -6575 32300 -6455
rect 32420 -6575 32465 -6455
rect 32585 -6575 32630 -6455
rect 32750 -6575 32805 -6455
rect 32925 -6575 32970 -6455
rect 33090 -6575 33135 -6455
rect 33255 -6575 33300 -6455
rect 33420 -6575 33475 -6455
rect 33595 -6575 33640 -6455
rect 33760 -6575 33805 -6455
rect 33925 -6575 33970 -6455
rect 34090 -6575 34145 -6455
rect 34265 -6575 34310 -6455
rect 34430 -6575 34475 -6455
rect 34595 -6575 34640 -6455
rect 34760 -6575 34815 -6455
rect 34935 -6575 34980 -6455
rect 35100 -6575 35145 -6455
rect 35265 -6575 35310 -6455
rect 35430 -6575 35485 -6455
rect 35605 -6575 35650 -6455
rect 35770 -6575 35815 -6455
rect 35935 -6575 35980 -6455
rect 36100 -6575 36155 -6455
rect 36275 -6575 36485 -6455
rect 36605 -6575 36650 -6455
rect 36770 -6575 36815 -6455
rect 36935 -6575 36980 -6455
rect 37100 -6575 37155 -6455
rect 37275 -6575 37320 -6455
rect 37440 -6575 37485 -6455
rect 37605 -6575 37650 -6455
rect 37770 -6575 37825 -6455
rect 37945 -6575 37990 -6455
rect 38110 -6575 38155 -6455
rect 38275 -6575 38320 -6455
rect 38440 -6575 38495 -6455
rect 38615 -6575 38660 -6455
rect 38780 -6575 38825 -6455
rect 38945 -6575 38990 -6455
rect 39110 -6575 39165 -6455
rect 39285 -6575 39330 -6455
rect 39450 -6575 39495 -6455
rect 39615 -6575 39660 -6455
rect 39780 -6575 39835 -6455
rect 39955 -6575 40000 -6455
rect 40120 -6575 40165 -6455
rect 40285 -6575 40330 -6455
rect 40450 -6575 40505 -6455
rect 40625 -6575 40670 -6455
rect 40790 -6575 40835 -6455
rect 40955 -6575 41000 -6455
rect 41120 -6575 41175 -6455
rect 41295 -6575 41340 -6455
rect 41460 -6575 41505 -6455
rect 41625 -6575 41670 -6455
rect 41790 -6575 41845 -6455
rect 41965 -6575 42175 -6455
rect 42295 -6575 42340 -6455
rect 42460 -6575 42505 -6455
rect 42625 -6575 42670 -6455
rect 42790 -6575 42845 -6455
rect 42965 -6575 43010 -6455
rect 43130 -6575 43175 -6455
rect 43295 -6575 43340 -6455
rect 43460 -6575 43515 -6455
rect 43635 -6575 43680 -6455
rect 43800 -6575 43845 -6455
rect 43965 -6575 44010 -6455
rect 44130 -6575 44185 -6455
rect 44305 -6575 44350 -6455
rect 44470 -6575 44515 -6455
rect 44635 -6575 44680 -6455
rect 44800 -6575 44855 -6455
rect 44975 -6575 45020 -6455
rect 45140 -6575 45185 -6455
rect 45305 -6575 45350 -6455
rect 45470 -6575 45525 -6455
rect 45645 -6575 45690 -6455
rect 45810 -6575 45855 -6455
rect 45975 -6575 46020 -6455
rect 46140 -6575 46195 -6455
rect 46315 -6575 46360 -6455
rect 46480 -6575 46525 -6455
rect 46645 -6575 46690 -6455
rect 46810 -6575 46865 -6455
rect 46985 -6575 47030 -6455
rect 47150 -6575 47195 -6455
rect 47315 -6575 47360 -6455
rect 47480 -6575 47535 -6455
rect 47655 -6575 47865 -6455
rect 47985 -6575 48030 -6455
rect 48150 -6575 48195 -6455
rect 48315 -6575 48360 -6455
rect 48480 -6575 48535 -6455
rect 48655 -6575 48700 -6455
rect 48820 -6575 48865 -6455
rect 48985 -6575 49030 -6455
rect 49150 -6575 49205 -6455
rect 49325 -6575 49370 -6455
rect 49490 -6575 49535 -6455
rect 49655 -6575 49700 -6455
rect 49820 -6575 49875 -6455
rect 49995 -6575 50040 -6455
rect 50160 -6575 50205 -6455
rect 50325 -6575 50370 -6455
rect 50490 -6575 50545 -6455
rect 50665 -6575 50710 -6455
rect 50830 -6575 50875 -6455
rect 50995 -6575 51040 -6455
rect 51160 -6575 51215 -6455
rect 51335 -6575 51380 -6455
rect 51500 -6575 51545 -6455
rect 51665 -6575 51710 -6455
rect 51830 -6575 51885 -6455
rect 52005 -6575 52050 -6455
rect 52170 -6575 52215 -6455
rect 52335 -6575 52380 -6455
rect 52500 -6575 52555 -6455
rect 52675 -6575 52720 -6455
rect 52840 -6575 52885 -6455
rect 53005 -6575 53050 -6455
rect 53170 -6575 53225 -6455
rect 53345 -6575 53370 -6455
rect 30770 -6620 53370 -6575
rect 30770 -6740 30795 -6620
rect 30915 -6740 30960 -6620
rect 31080 -6740 31125 -6620
rect 31245 -6740 31290 -6620
rect 31410 -6740 31465 -6620
rect 31585 -6740 31630 -6620
rect 31750 -6740 31795 -6620
rect 31915 -6740 31960 -6620
rect 32080 -6740 32135 -6620
rect 32255 -6740 32300 -6620
rect 32420 -6740 32465 -6620
rect 32585 -6740 32630 -6620
rect 32750 -6740 32805 -6620
rect 32925 -6740 32970 -6620
rect 33090 -6740 33135 -6620
rect 33255 -6740 33300 -6620
rect 33420 -6740 33475 -6620
rect 33595 -6740 33640 -6620
rect 33760 -6740 33805 -6620
rect 33925 -6740 33970 -6620
rect 34090 -6740 34145 -6620
rect 34265 -6740 34310 -6620
rect 34430 -6740 34475 -6620
rect 34595 -6740 34640 -6620
rect 34760 -6740 34815 -6620
rect 34935 -6740 34980 -6620
rect 35100 -6740 35145 -6620
rect 35265 -6740 35310 -6620
rect 35430 -6740 35485 -6620
rect 35605 -6740 35650 -6620
rect 35770 -6740 35815 -6620
rect 35935 -6740 35980 -6620
rect 36100 -6740 36155 -6620
rect 36275 -6740 36485 -6620
rect 36605 -6740 36650 -6620
rect 36770 -6740 36815 -6620
rect 36935 -6740 36980 -6620
rect 37100 -6740 37155 -6620
rect 37275 -6740 37320 -6620
rect 37440 -6740 37485 -6620
rect 37605 -6740 37650 -6620
rect 37770 -6740 37825 -6620
rect 37945 -6740 37990 -6620
rect 38110 -6740 38155 -6620
rect 38275 -6740 38320 -6620
rect 38440 -6740 38495 -6620
rect 38615 -6740 38660 -6620
rect 38780 -6740 38825 -6620
rect 38945 -6740 38990 -6620
rect 39110 -6740 39165 -6620
rect 39285 -6740 39330 -6620
rect 39450 -6740 39495 -6620
rect 39615 -6740 39660 -6620
rect 39780 -6740 39835 -6620
rect 39955 -6740 40000 -6620
rect 40120 -6740 40165 -6620
rect 40285 -6740 40330 -6620
rect 40450 -6740 40505 -6620
rect 40625 -6740 40670 -6620
rect 40790 -6740 40835 -6620
rect 40955 -6740 41000 -6620
rect 41120 -6740 41175 -6620
rect 41295 -6740 41340 -6620
rect 41460 -6740 41505 -6620
rect 41625 -6740 41670 -6620
rect 41790 -6740 41845 -6620
rect 41965 -6740 42175 -6620
rect 42295 -6740 42340 -6620
rect 42460 -6740 42505 -6620
rect 42625 -6740 42670 -6620
rect 42790 -6740 42845 -6620
rect 42965 -6740 43010 -6620
rect 43130 -6740 43175 -6620
rect 43295 -6740 43340 -6620
rect 43460 -6740 43515 -6620
rect 43635 -6740 43680 -6620
rect 43800 -6740 43845 -6620
rect 43965 -6740 44010 -6620
rect 44130 -6740 44185 -6620
rect 44305 -6740 44350 -6620
rect 44470 -6740 44515 -6620
rect 44635 -6740 44680 -6620
rect 44800 -6740 44855 -6620
rect 44975 -6740 45020 -6620
rect 45140 -6740 45185 -6620
rect 45305 -6740 45350 -6620
rect 45470 -6740 45525 -6620
rect 45645 -6740 45690 -6620
rect 45810 -6740 45855 -6620
rect 45975 -6740 46020 -6620
rect 46140 -6740 46195 -6620
rect 46315 -6740 46360 -6620
rect 46480 -6740 46525 -6620
rect 46645 -6740 46690 -6620
rect 46810 -6740 46865 -6620
rect 46985 -6740 47030 -6620
rect 47150 -6740 47195 -6620
rect 47315 -6740 47360 -6620
rect 47480 -6740 47535 -6620
rect 47655 -6740 47865 -6620
rect 47985 -6740 48030 -6620
rect 48150 -6740 48195 -6620
rect 48315 -6740 48360 -6620
rect 48480 -6740 48535 -6620
rect 48655 -6740 48700 -6620
rect 48820 -6740 48865 -6620
rect 48985 -6740 49030 -6620
rect 49150 -6740 49205 -6620
rect 49325 -6740 49370 -6620
rect 49490 -6740 49535 -6620
rect 49655 -6740 49700 -6620
rect 49820 -6740 49875 -6620
rect 49995 -6740 50040 -6620
rect 50160 -6740 50205 -6620
rect 50325 -6740 50370 -6620
rect 50490 -6740 50545 -6620
rect 50665 -6740 50710 -6620
rect 50830 -6740 50875 -6620
rect 50995 -6740 51040 -6620
rect 51160 -6740 51215 -6620
rect 51335 -6740 51380 -6620
rect 51500 -6740 51545 -6620
rect 51665 -6740 51710 -6620
rect 51830 -6740 51885 -6620
rect 52005 -6740 52050 -6620
rect 52170 -6740 52215 -6620
rect 52335 -6740 52380 -6620
rect 52500 -6740 52555 -6620
rect 52675 -6740 52720 -6620
rect 52840 -6740 52885 -6620
rect 53005 -6740 53050 -6620
rect 53170 -6740 53225 -6620
rect 53345 -6740 53370 -6620
rect 30770 -6785 53370 -6740
rect 30770 -6905 30795 -6785
rect 30915 -6905 30960 -6785
rect 31080 -6905 31125 -6785
rect 31245 -6905 31290 -6785
rect 31410 -6905 31465 -6785
rect 31585 -6905 31630 -6785
rect 31750 -6905 31795 -6785
rect 31915 -6905 31960 -6785
rect 32080 -6905 32135 -6785
rect 32255 -6905 32300 -6785
rect 32420 -6905 32465 -6785
rect 32585 -6905 32630 -6785
rect 32750 -6905 32805 -6785
rect 32925 -6905 32970 -6785
rect 33090 -6905 33135 -6785
rect 33255 -6905 33300 -6785
rect 33420 -6905 33475 -6785
rect 33595 -6905 33640 -6785
rect 33760 -6905 33805 -6785
rect 33925 -6905 33970 -6785
rect 34090 -6905 34145 -6785
rect 34265 -6905 34310 -6785
rect 34430 -6905 34475 -6785
rect 34595 -6905 34640 -6785
rect 34760 -6905 34815 -6785
rect 34935 -6905 34980 -6785
rect 35100 -6905 35145 -6785
rect 35265 -6905 35310 -6785
rect 35430 -6905 35485 -6785
rect 35605 -6905 35650 -6785
rect 35770 -6905 35815 -6785
rect 35935 -6905 35980 -6785
rect 36100 -6905 36155 -6785
rect 36275 -6905 36485 -6785
rect 36605 -6905 36650 -6785
rect 36770 -6905 36815 -6785
rect 36935 -6905 36980 -6785
rect 37100 -6905 37155 -6785
rect 37275 -6905 37320 -6785
rect 37440 -6905 37485 -6785
rect 37605 -6905 37650 -6785
rect 37770 -6905 37825 -6785
rect 37945 -6905 37990 -6785
rect 38110 -6905 38155 -6785
rect 38275 -6905 38320 -6785
rect 38440 -6905 38495 -6785
rect 38615 -6905 38660 -6785
rect 38780 -6905 38825 -6785
rect 38945 -6905 38990 -6785
rect 39110 -6905 39165 -6785
rect 39285 -6905 39330 -6785
rect 39450 -6905 39495 -6785
rect 39615 -6905 39660 -6785
rect 39780 -6905 39835 -6785
rect 39955 -6905 40000 -6785
rect 40120 -6905 40165 -6785
rect 40285 -6905 40330 -6785
rect 40450 -6905 40505 -6785
rect 40625 -6905 40670 -6785
rect 40790 -6905 40835 -6785
rect 40955 -6905 41000 -6785
rect 41120 -6905 41175 -6785
rect 41295 -6905 41340 -6785
rect 41460 -6905 41505 -6785
rect 41625 -6905 41670 -6785
rect 41790 -6905 41845 -6785
rect 41965 -6905 42175 -6785
rect 42295 -6905 42340 -6785
rect 42460 -6905 42505 -6785
rect 42625 -6905 42670 -6785
rect 42790 -6905 42845 -6785
rect 42965 -6905 43010 -6785
rect 43130 -6905 43175 -6785
rect 43295 -6905 43340 -6785
rect 43460 -6905 43515 -6785
rect 43635 -6905 43680 -6785
rect 43800 -6905 43845 -6785
rect 43965 -6905 44010 -6785
rect 44130 -6905 44185 -6785
rect 44305 -6905 44350 -6785
rect 44470 -6905 44515 -6785
rect 44635 -6905 44680 -6785
rect 44800 -6905 44855 -6785
rect 44975 -6905 45020 -6785
rect 45140 -6905 45185 -6785
rect 45305 -6905 45350 -6785
rect 45470 -6905 45525 -6785
rect 45645 -6905 45690 -6785
rect 45810 -6905 45855 -6785
rect 45975 -6905 46020 -6785
rect 46140 -6905 46195 -6785
rect 46315 -6905 46360 -6785
rect 46480 -6905 46525 -6785
rect 46645 -6905 46690 -6785
rect 46810 -6905 46865 -6785
rect 46985 -6905 47030 -6785
rect 47150 -6905 47195 -6785
rect 47315 -6905 47360 -6785
rect 47480 -6905 47535 -6785
rect 47655 -6905 47865 -6785
rect 47985 -6905 48030 -6785
rect 48150 -6905 48195 -6785
rect 48315 -6905 48360 -6785
rect 48480 -6905 48535 -6785
rect 48655 -6905 48700 -6785
rect 48820 -6905 48865 -6785
rect 48985 -6905 49030 -6785
rect 49150 -6905 49205 -6785
rect 49325 -6905 49370 -6785
rect 49490 -6905 49535 -6785
rect 49655 -6905 49700 -6785
rect 49820 -6905 49875 -6785
rect 49995 -6905 50040 -6785
rect 50160 -6905 50205 -6785
rect 50325 -6905 50370 -6785
rect 50490 -6905 50545 -6785
rect 50665 -6905 50710 -6785
rect 50830 -6905 50875 -6785
rect 50995 -6905 51040 -6785
rect 51160 -6905 51215 -6785
rect 51335 -6905 51380 -6785
rect 51500 -6905 51545 -6785
rect 51665 -6905 51710 -6785
rect 51830 -6905 51885 -6785
rect 52005 -6905 52050 -6785
rect 52170 -6905 52215 -6785
rect 52335 -6905 52380 -6785
rect 52500 -6905 52555 -6785
rect 52675 -6905 52720 -6785
rect 52840 -6905 52885 -6785
rect 53005 -6905 53050 -6785
rect 53170 -6905 53225 -6785
rect 53345 -6905 53370 -6785
rect 30770 -6950 53370 -6905
rect 30770 -7070 30795 -6950
rect 30915 -7070 30960 -6950
rect 31080 -7070 31125 -6950
rect 31245 -7070 31290 -6950
rect 31410 -7070 31465 -6950
rect 31585 -7070 31630 -6950
rect 31750 -7070 31795 -6950
rect 31915 -7070 31960 -6950
rect 32080 -7070 32135 -6950
rect 32255 -7070 32300 -6950
rect 32420 -7070 32465 -6950
rect 32585 -7070 32630 -6950
rect 32750 -7070 32805 -6950
rect 32925 -7070 32970 -6950
rect 33090 -7070 33135 -6950
rect 33255 -7070 33300 -6950
rect 33420 -7070 33475 -6950
rect 33595 -7070 33640 -6950
rect 33760 -7070 33805 -6950
rect 33925 -7070 33970 -6950
rect 34090 -7070 34145 -6950
rect 34265 -7070 34310 -6950
rect 34430 -7070 34475 -6950
rect 34595 -7070 34640 -6950
rect 34760 -7070 34815 -6950
rect 34935 -7070 34980 -6950
rect 35100 -7070 35145 -6950
rect 35265 -7070 35310 -6950
rect 35430 -7070 35485 -6950
rect 35605 -7070 35650 -6950
rect 35770 -7070 35815 -6950
rect 35935 -7070 35980 -6950
rect 36100 -7070 36155 -6950
rect 36275 -7070 36485 -6950
rect 36605 -7070 36650 -6950
rect 36770 -7070 36815 -6950
rect 36935 -7070 36980 -6950
rect 37100 -7070 37155 -6950
rect 37275 -7070 37320 -6950
rect 37440 -7070 37485 -6950
rect 37605 -7070 37650 -6950
rect 37770 -7070 37825 -6950
rect 37945 -7070 37990 -6950
rect 38110 -7070 38155 -6950
rect 38275 -7070 38320 -6950
rect 38440 -7070 38495 -6950
rect 38615 -7070 38660 -6950
rect 38780 -7070 38825 -6950
rect 38945 -7070 38990 -6950
rect 39110 -7070 39165 -6950
rect 39285 -7070 39330 -6950
rect 39450 -7070 39495 -6950
rect 39615 -7070 39660 -6950
rect 39780 -7070 39835 -6950
rect 39955 -7070 40000 -6950
rect 40120 -7070 40165 -6950
rect 40285 -7070 40330 -6950
rect 40450 -7070 40505 -6950
rect 40625 -7070 40670 -6950
rect 40790 -7070 40835 -6950
rect 40955 -7070 41000 -6950
rect 41120 -7070 41175 -6950
rect 41295 -7070 41340 -6950
rect 41460 -7070 41505 -6950
rect 41625 -7070 41670 -6950
rect 41790 -7070 41845 -6950
rect 41965 -7070 42175 -6950
rect 42295 -7070 42340 -6950
rect 42460 -7070 42505 -6950
rect 42625 -7070 42670 -6950
rect 42790 -7070 42845 -6950
rect 42965 -7070 43010 -6950
rect 43130 -7070 43175 -6950
rect 43295 -7070 43340 -6950
rect 43460 -7070 43515 -6950
rect 43635 -7070 43680 -6950
rect 43800 -7070 43845 -6950
rect 43965 -7070 44010 -6950
rect 44130 -7070 44185 -6950
rect 44305 -7070 44350 -6950
rect 44470 -7070 44515 -6950
rect 44635 -7070 44680 -6950
rect 44800 -7070 44855 -6950
rect 44975 -7070 45020 -6950
rect 45140 -7070 45185 -6950
rect 45305 -7070 45350 -6950
rect 45470 -7070 45525 -6950
rect 45645 -7070 45690 -6950
rect 45810 -7070 45855 -6950
rect 45975 -7070 46020 -6950
rect 46140 -7070 46195 -6950
rect 46315 -7070 46360 -6950
rect 46480 -7070 46525 -6950
rect 46645 -7070 46690 -6950
rect 46810 -7070 46865 -6950
rect 46985 -7070 47030 -6950
rect 47150 -7070 47195 -6950
rect 47315 -7070 47360 -6950
rect 47480 -7070 47535 -6950
rect 47655 -7070 47865 -6950
rect 47985 -7070 48030 -6950
rect 48150 -7070 48195 -6950
rect 48315 -7070 48360 -6950
rect 48480 -7070 48535 -6950
rect 48655 -7070 48700 -6950
rect 48820 -7070 48865 -6950
rect 48985 -7070 49030 -6950
rect 49150 -7070 49205 -6950
rect 49325 -7070 49370 -6950
rect 49490 -7070 49535 -6950
rect 49655 -7070 49700 -6950
rect 49820 -7070 49875 -6950
rect 49995 -7070 50040 -6950
rect 50160 -7070 50205 -6950
rect 50325 -7070 50370 -6950
rect 50490 -7070 50545 -6950
rect 50665 -7070 50710 -6950
rect 50830 -7070 50875 -6950
rect 50995 -7070 51040 -6950
rect 51160 -7070 51215 -6950
rect 51335 -7070 51380 -6950
rect 51500 -7070 51545 -6950
rect 51665 -7070 51710 -6950
rect 51830 -7070 51885 -6950
rect 52005 -7070 52050 -6950
rect 52170 -7070 52215 -6950
rect 52335 -7070 52380 -6950
rect 52500 -7070 52555 -6950
rect 52675 -7070 52720 -6950
rect 52840 -7070 52885 -6950
rect 53005 -7070 53050 -6950
rect 53170 -7070 53225 -6950
rect 53345 -7070 53370 -6950
rect 30770 -7125 53370 -7070
rect 30770 -7245 30795 -7125
rect 30915 -7245 30960 -7125
rect 31080 -7245 31125 -7125
rect 31245 -7245 31290 -7125
rect 31410 -7245 31465 -7125
rect 31585 -7245 31630 -7125
rect 31750 -7245 31795 -7125
rect 31915 -7245 31960 -7125
rect 32080 -7245 32135 -7125
rect 32255 -7245 32300 -7125
rect 32420 -7245 32465 -7125
rect 32585 -7245 32630 -7125
rect 32750 -7245 32805 -7125
rect 32925 -7245 32970 -7125
rect 33090 -7245 33135 -7125
rect 33255 -7245 33300 -7125
rect 33420 -7245 33475 -7125
rect 33595 -7245 33640 -7125
rect 33760 -7245 33805 -7125
rect 33925 -7245 33970 -7125
rect 34090 -7245 34145 -7125
rect 34265 -7245 34310 -7125
rect 34430 -7245 34475 -7125
rect 34595 -7245 34640 -7125
rect 34760 -7245 34815 -7125
rect 34935 -7245 34980 -7125
rect 35100 -7245 35145 -7125
rect 35265 -7245 35310 -7125
rect 35430 -7245 35485 -7125
rect 35605 -7245 35650 -7125
rect 35770 -7245 35815 -7125
rect 35935 -7245 35980 -7125
rect 36100 -7245 36155 -7125
rect 36275 -7245 36485 -7125
rect 36605 -7245 36650 -7125
rect 36770 -7245 36815 -7125
rect 36935 -7245 36980 -7125
rect 37100 -7245 37155 -7125
rect 37275 -7245 37320 -7125
rect 37440 -7245 37485 -7125
rect 37605 -7245 37650 -7125
rect 37770 -7245 37825 -7125
rect 37945 -7245 37990 -7125
rect 38110 -7245 38155 -7125
rect 38275 -7245 38320 -7125
rect 38440 -7245 38495 -7125
rect 38615 -7245 38660 -7125
rect 38780 -7245 38825 -7125
rect 38945 -7245 38990 -7125
rect 39110 -7245 39165 -7125
rect 39285 -7245 39330 -7125
rect 39450 -7245 39495 -7125
rect 39615 -7245 39660 -7125
rect 39780 -7245 39835 -7125
rect 39955 -7245 40000 -7125
rect 40120 -7245 40165 -7125
rect 40285 -7245 40330 -7125
rect 40450 -7245 40505 -7125
rect 40625 -7245 40670 -7125
rect 40790 -7245 40835 -7125
rect 40955 -7245 41000 -7125
rect 41120 -7245 41175 -7125
rect 41295 -7245 41340 -7125
rect 41460 -7245 41505 -7125
rect 41625 -7245 41670 -7125
rect 41790 -7245 41845 -7125
rect 41965 -7245 42175 -7125
rect 42295 -7245 42340 -7125
rect 42460 -7245 42505 -7125
rect 42625 -7245 42670 -7125
rect 42790 -7245 42845 -7125
rect 42965 -7245 43010 -7125
rect 43130 -7245 43175 -7125
rect 43295 -7245 43340 -7125
rect 43460 -7245 43515 -7125
rect 43635 -7245 43680 -7125
rect 43800 -7245 43845 -7125
rect 43965 -7245 44010 -7125
rect 44130 -7245 44185 -7125
rect 44305 -7245 44350 -7125
rect 44470 -7245 44515 -7125
rect 44635 -7245 44680 -7125
rect 44800 -7245 44855 -7125
rect 44975 -7245 45020 -7125
rect 45140 -7245 45185 -7125
rect 45305 -7245 45350 -7125
rect 45470 -7245 45525 -7125
rect 45645 -7245 45690 -7125
rect 45810 -7245 45855 -7125
rect 45975 -7245 46020 -7125
rect 46140 -7245 46195 -7125
rect 46315 -7245 46360 -7125
rect 46480 -7245 46525 -7125
rect 46645 -7245 46690 -7125
rect 46810 -7245 46865 -7125
rect 46985 -7245 47030 -7125
rect 47150 -7245 47195 -7125
rect 47315 -7245 47360 -7125
rect 47480 -7245 47535 -7125
rect 47655 -7245 47865 -7125
rect 47985 -7245 48030 -7125
rect 48150 -7245 48195 -7125
rect 48315 -7245 48360 -7125
rect 48480 -7245 48535 -7125
rect 48655 -7245 48700 -7125
rect 48820 -7245 48865 -7125
rect 48985 -7245 49030 -7125
rect 49150 -7245 49205 -7125
rect 49325 -7245 49370 -7125
rect 49490 -7245 49535 -7125
rect 49655 -7245 49700 -7125
rect 49820 -7245 49875 -7125
rect 49995 -7245 50040 -7125
rect 50160 -7245 50205 -7125
rect 50325 -7245 50370 -7125
rect 50490 -7245 50545 -7125
rect 50665 -7245 50710 -7125
rect 50830 -7245 50875 -7125
rect 50995 -7245 51040 -7125
rect 51160 -7245 51215 -7125
rect 51335 -7245 51380 -7125
rect 51500 -7245 51545 -7125
rect 51665 -7245 51710 -7125
rect 51830 -7245 51885 -7125
rect 52005 -7245 52050 -7125
rect 52170 -7245 52215 -7125
rect 52335 -7245 52380 -7125
rect 52500 -7245 52555 -7125
rect 52675 -7245 52720 -7125
rect 52840 -7245 52885 -7125
rect 53005 -7245 53050 -7125
rect 53170 -7245 53225 -7125
rect 53345 -7245 53370 -7125
rect 30770 -7290 53370 -7245
rect 30770 -7410 30795 -7290
rect 30915 -7410 30960 -7290
rect 31080 -7410 31125 -7290
rect 31245 -7410 31290 -7290
rect 31410 -7410 31465 -7290
rect 31585 -7410 31630 -7290
rect 31750 -7410 31795 -7290
rect 31915 -7410 31960 -7290
rect 32080 -7410 32135 -7290
rect 32255 -7410 32300 -7290
rect 32420 -7410 32465 -7290
rect 32585 -7410 32630 -7290
rect 32750 -7410 32805 -7290
rect 32925 -7410 32970 -7290
rect 33090 -7410 33135 -7290
rect 33255 -7410 33300 -7290
rect 33420 -7410 33475 -7290
rect 33595 -7410 33640 -7290
rect 33760 -7410 33805 -7290
rect 33925 -7410 33970 -7290
rect 34090 -7410 34145 -7290
rect 34265 -7410 34310 -7290
rect 34430 -7410 34475 -7290
rect 34595 -7410 34640 -7290
rect 34760 -7410 34815 -7290
rect 34935 -7410 34980 -7290
rect 35100 -7410 35145 -7290
rect 35265 -7410 35310 -7290
rect 35430 -7410 35485 -7290
rect 35605 -7410 35650 -7290
rect 35770 -7410 35815 -7290
rect 35935 -7410 35980 -7290
rect 36100 -7410 36155 -7290
rect 36275 -7410 36485 -7290
rect 36605 -7410 36650 -7290
rect 36770 -7410 36815 -7290
rect 36935 -7410 36980 -7290
rect 37100 -7410 37155 -7290
rect 37275 -7410 37320 -7290
rect 37440 -7410 37485 -7290
rect 37605 -7410 37650 -7290
rect 37770 -7410 37825 -7290
rect 37945 -7410 37990 -7290
rect 38110 -7410 38155 -7290
rect 38275 -7410 38320 -7290
rect 38440 -7410 38495 -7290
rect 38615 -7410 38660 -7290
rect 38780 -7410 38825 -7290
rect 38945 -7410 38990 -7290
rect 39110 -7410 39165 -7290
rect 39285 -7410 39330 -7290
rect 39450 -7410 39495 -7290
rect 39615 -7410 39660 -7290
rect 39780 -7410 39835 -7290
rect 39955 -7410 40000 -7290
rect 40120 -7410 40165 -7290
rect 40285 -7410 40330 -7290
rect 40450 -7410 40505 -7290
rect 40625 -7410 40670 -7290
rect 40790 -7410 40835 -7290
rect 40955 -7410 41000 -7290
rect 41120 -7410 41175 -7290
rect 41295 -7410 41340 -7290
rect 41460 -7410 41505 -7290
rect 41625 -7410 41670 -7290
rect 41790 -7410 41845 -7290
rect 41965 -7410 42175 -7290
rect 42295 -7410 42340 -7290
rect 42460 -7410 42505 -7290
rect 42625 -7410 42670 -7290
rect 42790 -7410 42845 -7290
rect 42965 -7410 43010 -7290
rect 43130 -7410 43175 -7290
rect 43295 -7410 43340 -7290
rect 43460 -7410 43515 -7290
rect 43635 -7410 43680 -7290
rect 43800 -7410 43845 -7290
rect 43965 -7410 44010 -7290
rect 44130 -7410 44185 -7290
rect 44305 -7410 44350 -7290
rect 44470 -7410 44515 -7290
rect 44635 -7410 44680 -7290
rect 44800 -7410 44855 -7290
rect 44975 -7410 45020 -7290
rect 45140 -7410 45185 -7290
rect 45305 -7410 45350 -7290
rect 45470 -7410 45525 -7290
rect 45645 -7410 45690 -7290
rect 45810 -7410 45855 -7290
rect 45975 -7410 46020 -7290
rect 46140 -7410 46195 -7290
rect 46315 -7410 46360 -7290
rect 46480 -7410 46525 -7290
rect 46645 -7410 46690 -7290
rect 46810 -7410 46865 -7290
rect 46985 -7410 47030 -7290
rect 47150 -7410 47195 -7290
rect 47315 -7410 47360 -7290
rect 47480 -7410 47535 -7290
rect 47655 -7410 47865 -7290
rect 47985 -7410 48030 -7290
rect 48150 -7410 48195 -7290
rect 48315 -7410 48360 -7290
rect 48480 -7410 48535 -7290
rect 48655 -7410 48700 -7290
rect 48820 -7410 48865 -7290
rect 48985 -7410 49030 -7290
rect 49150 -7410 49205 -7290
rect 49325 -7410 49370 -7290
rect 49490 -7410 49535 -7290
rect 49655 -7410 49700 -7290
rect 49820 -7410 49875 -7290
rect 49995 -7410 50040 -7290
rect 50160 -7410 50205 -7290
rect 50325 -7410 50370 -7290
rect 50490 -7410 50545 -7290
rect 50665 -7410 50710 -7290
rect 50830 -7410 50875 -7290
rect 50995 -7410 51040 -7290
rect 51160 -7410 51215 -7290
rect 51335 -7410 51380 -7290
rect 51500 -7410 51545 -7290
rect 51665 -7410 51710 -7290
rect 51830 -7410 51885 -7290
rect 52005 -7410 52050 -7290
rect 52170 -7410 52215 -7290
rect 52335 -7410 52380 -7290
rect 52500 -7410 52555 -7290
rect 52675 -7410 52720 -7290
rect 52840 -7410 52885 -7290
rect 53005 -7410 53050 -7290
rect 53170 -7410 53225 -7290
rect 53345 -7410 53370 -7290
rect 30770 -7455 53370 -7410
rect 30770 -7575 30795 -7455
rect 30915 -7575 30960 -7455
rect 31080 -7575 31125 -7455
rect 31245 -7575 31290 -7455
rect 31410 -7575 31465 -7455
rect 31585 -7575 31630 -7455
rect 31750 -7575 31795 -7455
rect 31915 -7575 31960 -7455
rect 32080 -7575 32135 -7455
rect 32255 -7575 32300 -7455
rect 32420 -7575 32465 -7455
rect 32585 -7575 32630 -7455
rect 32750 -7575 32805 -7455
rect 32925 -7575 32970 -7455
rect 33090 -7575 33135 -7455
rect 33255 -7575 33300 -7455
rect 33420 -7575 33475 -7455
rect 33595 -7575 33640 -7455
rect 33760 -7575 33805 -7455
rect 33925 -7575 33970 -7455
rect 34090 -7575 34145 -7455
rect 34265 -7575 34310 -7455
rect 34430 -7575 34475 -7455
rect 34595 -7575 34640 -7455
rect 34760 -7575 34815 -7455
rect 34935 -7575 34980 -7455
rect 35100 -7575 35145 -7455
rect 35265 -7575 35310 -7455
rect 35430 -7575 35485 -7455
rect 35605 -7575 35650 -7455
rect 35770 -7575 35815 -7455
rect 35935 -7575 35980 -7455
rect 36100 -7575 36155 -7455
rect 36275 -7575 36485 -7455
rect 36605 -7575 36650 -7455
rect 36770 -7575 36815 -7455
rect 36935 -7575 36980 -7455
rect 37100 -7575 37155 -7455
rect 37275 -7575 37320 -7455
rect 37440 -7575 37485 -7455
rect 37605 -7575 37650 -7455
rect 37770 -7575 37825 -7455
rect 37945 -7575 37990 -7455
rect 38110 -7575 38155 -7455
rect 38275 -7575 38320 -7455
rect 38440 -7575 38495 -7455
rect 38615 -7575 38660 -7455
rect 38780 -7575 38825 -7455
rect 38945 -7575 38990 -7455
rect 39110 -7575 39165 -7455
rect 39285 -7575 39330 -7455
rect 39450 -7575 39495 -7455
rect 39615 -7575 39660 -7455
rect 39780 -7575 39835 -7455
rect 39955 -7575 40000 -7455
rect 40120 -7575 40165 -7455
rect 40285 -7575 40330 -7455
rect 40450 -7575 40505 -7455
rect 40625 -7575 40670 -7455
rect 40790 -7575 40835 -7455
rect 40955 -7575 41000 -7455
rect 41120 -7575 41175 -7455
rect 41295 -7575 41340 -7455
rect 41460 -7575 41505 -7455
rect 41625 -7575 41670 -7455
rect 41790 -7575 41845 -7455
rect 41965 -7575 42175 -7455
rect 42295 -7575 42340 -7455
rect 42460 -7575 42505 -7455
rect 42625 -7575 42670 -7455
rect 42790 -7575 42845 -7455
rect 42965 -7575 43010 -7455
rect 43130 -7575 43175 -7455
rect 43295 -7575 43340 -7455
rect 43460 -7575 43515 -7455
rect 43635 -7575 43680 -7455
rect 43800 -7575 43845 -7455
rect 43965 -7575 44010 -7455
rect 44130 -7575 44185 -7455
rect 44305 -7575 44350 -7455
rect 44470 -7575 44515 -7455
rect 44635 -7575 44680 -7455
rect 44800 -7575 44855 -7455
rect 44975 -7575 45020 -7455
rect 45140 -7575 45185 -7455
rect 45305 -7575 45350 -7455
rect 45470 -7575 45525 -7455
rect 45645 -7575 45690 -7455
rect 45810 -7575 45855 -7455
rect 45975 -7575 46020 -7455
rect 46140 -7575 46195 -7455
rect 46315 -7575 46360 -7455
rect 46480 -7575 46525 -7455
rect 46645 -7575 46690 -7455
rect 46810 -7575 46865 -7455
rect 46985 -7575 47030 -7455
rect 47150 -7575 47195 -7455
rect 47315 -7575 47360 -7455
rect 47480 -7575 47535 -7455
rect 47655 -7575 47865 -7455
rect 47985 -7575 48030 -7455
rect 48150 -7575 48195 -7455
rect 48315 -7575 48360 -7455
rect 48480 -7575 48535 -7455
rect 48655 -7575 48700 -7455
rect 48820 -7575 48865 -7455
rect 48985 -7575 49030 -7455
rect 49150 -7575 49205 -7455
rect 49325 -7575 49370 -7455
rect 49490 -7575 49535 -7455
rect 49655 -7575 49700 -7455
rect 49820 -7575 49875 -7455
rect 49995 -7575 50040 -7455
rect 50160 -7575 50205 -7455
rect 50325 -7575 50370 -7455
rect 50490 -7575 50545 -7455
rect 50665 -7575 50710 -7455
rect 50830 -7575 50875 -7455
rect 50995 -7575 51040 -7455
rect 51160 -7575 51215 -7455
rect 51335 -7575 51380 -7455
rect 51500 -7575 51545 -7455
rect 51665 -7575 51710 -7455
rect 51830 -7575 51885 -7455
rect 52005 -7575 52050 -7455
rect 52170 -7575 52215 -7455
rect 52335 -7575 52380 -7455
rect 52500 -7575 52555 -7455
rect 52675 -7575 52720 -7455
rect 52840 -7575 52885 -7455
rect 53005 -7575 53050 -7455
rect 53170 -7575 53225 -7455
rect 53345 -7575 53370 -7455
rect 30770 -7620 53370 -7575
rect 30770 -7740 30795 -7620
rect 30915 -7740 30960 -7620
rect 31080 -7740 31125 -7620
rect 31245 -7740 31290 -7620
rect 31410 -7740 31465 -7620
rect 31585 -7740 31630 -7620
rect 31750 -7740 31795 -7620
rect 31915 -7740 31960 -7620
rect 32080 -7740 32135 -7620
rect 32255 -7740 32300 -7620
rect 32420 -7740 32465 -7620
rect 32585 -7740 32630 -7620
rect 32750 -7740 32805 -7620
rect 32925 -7740 32970 -7620
rect 33090 -7740 33135 -7620
rect 33255 -7740 33300 -7620
rect 33420 -7740 33475 -7620
rect 33595 -7740 33640 -7620
rect 33760 -7740 33805 -7620
rect 33925 -7740 33970 -7620
rect 34090 -7740 34145 -7620
rect 34265 -7740 34310 -7620
rect 34430 -7740 34475 -7620
rect 34595 -7740 34640 -7620
rect 34760 -7740 34815 -7620
rect 34935 -7740 34980 -7620
rect 35100 -7740 35145 -7620
rect 35265 -7740 35310 -7620
rect 35430 -7740 35485 -7620
rect 35605 -7740 35650 -7620
rect 35770 -7740 35815 -7620
rect 35935 -7740 35980 -7620
rect 36100 -7740 36155 -7620
rect 36275 -7740 36485 -7620
rect 36605 -7740 36650 -7620
rect 36770 -7740 36815 -7620
rect 36935 -7740 36980 -7620
rect 37100 -7740 37155 -7620
rect 37275 -7740 37320 -7620
rect 37440 -7740 37485 -7620
rect 37605 -7740 37650 -7620
rect 37770 -7740 37825 -7620
rect 37945 -7740 37990 -7620
rect 38110 -7740 38155 -7620
rect 38275 -7740 38320 -7620
rect 38440 -7740 38495 -7620
rect 38615 -7740 38660 -7620
rect 38780 -7740 38825 -7620
rect 38945 -7740 38990 -7620
rect 39110 -7740 39165 -7620
rect 39285 -7740 39330 -7620
rect 39450 -7740 39495 -7620
rect 39615 -7740 39660 -7620
rect 39780 -7740 39835 -7620
rect 39955 -7740 40000 -7620
rect 40120 -7740 40165 -7620
rect 40285 -7740 40330 -7620
rect 40450 -7740 40505 -7620
rect 40625 -7740 40670 -7620
rect 40790 -7740 40835 -7620
rect 40955 -7740 41000 -7620
rect 41120 -7740 41175 -7620
rect 41295 -7740 41340 -7620
rect 41460 -7740 41505 -7620
rect 41625 -7740 41670 -7620
rect 41790 -7740 41845 -7620
rect 41965 -7740 42175 -7620
rect 42295 -7740 42340 -7620
rect 42460 -7740 42505 -7620
rect 42625 -7740 42670 -7620
rect 42790 -7740 42845 -7620
rect 42965 -7740 43010 -7620
rect 43130 -7740 43175 -7620
rect 43295 -7740 43340 -7620
rect 43460 -7740 43515 -7620
rect 43635 -7740 43680 -7620
rect 43800 -7740 43845 -7620
rect 43965 -7740 44010 -7620
rect 44130 -7740 44185 -7620
rect 44305 -7740 44350 -7620
rect 44470 -7740 44515 -7620
rect 44635 -7740 44680 -7620
rect 44800 -7740 44855 -7620
rect 44975 -7740 45020 -7620
rect 45140 -7740 45185 -7620
rect 45305 -7740 45350 -7620
rect 45470 -7740 45525 -7620
rect 45645 -7740 45690 -7620
rect 45810 -7740 45855 -7620
rect 45975 -7740 46020 -7620
rect 46140 -7740 46195 -7620
rect 46315 -7740 46360 -7620
rect 46480 -7740 46525 -7620
rect 46645 -7740 46690 -7620
rect 46810 -7740 46865 -7620
rect 46985 -7740 47030 -7620
rect 47150 -7740 47195 -7620
rect 47315 -7740 47360 -7620
rect 47480 -7740 47535 -7620
rect 47655 -7740 47865 -7620
rect 47985 -7740 48030 -7620
rect 48150 -7740 48195 -7620
rect 48315 -7740 48360 -7620
rect 48480 -7740 48535 -7620
rect 48655 -7740 48700 -7620
rect 48820 -7740 48865 -7620
rect 48985 -7740 49030 -7620
rect 49150 -7740 49205 -7620
rect 49325 -7740 49370 -7620
rect 49490 -7740 49535 -7620
rect 49655 -7740 49700 -7620
rect 49820 -7740 49875 -7620
rect 49995 -7740 50040 -7620
rect 50160 -7740 50205 -7620
rect 50325 -7740 50370 -7620
rect 50490 -7740 50545 -7620
rect 50665 -7740 50710 -7620
rect 50830 -7740 50875 -7620
rect 50995 -7740 51040 -7620
rect 51160 -7740 51215 -7620
rect 51335 -7740 51380 -7620
rect 51500 -7740 51545 -7620
rect 51665 -7740 51710 -7620
rect 51830 -7740 51885 -7620
rect 52005 -7740 52050 -7620
rect 52170 -7740 52215 -7620
rect 52335 -7740 52380 -7620
rect 52500 -7740 52555 -7620
rect 52675 -7740 52720 -7620
rect 52840 -7740 52885 -7620
rect 53005 -7740 53050 -7620
rect 53170 -7740 53225 -7620
rect 53345 -7740 53370 -7620
rect 30770 -7795 53370 -7740
rect 30770 -7915 30795 -7795
rect 30915 -7915 30960 -7795
rect 31080 -7915 31125 -7795
rect 31245 -7915 31290 -7795
rect 31410 -7915 31465 -7795
rect 31585 -7915 31630 -7795
rect 31750 -7915 31795 -7795
rect 31915 -7915 31960 -7795
rect 32080 -7915 32135 -7795
rect 32255 -7915 32300 -7795
rect 32420 -7915 32465 -7795
rect 32585 -7915 32630 -7795
rect 32750 -7915 32805 -7795
rect 32925 -7915 32970 -7795
rect 33090 -7915 33135 -7795
rect 33255 -7915 33300 -7795
rect 33420 -7915 33475 -7795
rect 33595 -7915 33640 -7795
rect 33760 -7915 33805 -7795
rect 33925 -7915 33970 -7795
rect 34090 -7915 34145 -7795
rect 34265 -7915 34310 -7795
rect 34430 -7915 34475 -7795
rect 34595 -7915 34640 -7795
rect 34760 -7915 34815 -7795
rect 34935 -7915 34980 -7795
rect 35100 -7915 35145 -7795
rect 35265 -7915 35310 -7795
rect 35430 -7915 35485 -7795
rect 35605 -7915 35650 -7795
rect 35770 -7915 35815 -7795
rect 35935 -7915 35980 -7795
rect 36100 -7915 36155 -7795
rect 36275 -7915 36485 -7795
rect 36605 -7915 36650 -7795
rect 36770 -7915 36815 -7795
rect 36935 -7915 36980 -7795
rect 37100 -7915 37155 -7795
rect 37275 -7915 37320 -7795
rect 37440 -7915 37485 -7795
rect 37605 -7915 37650 -7795
rect 37770 -7915 37825 -7795
rect 37945 -7915 37990 -7795
rect 38110 -7915 38155 -7795
rect 38275 -7915 38320 -7795
rect 38440 -7915 38495 -7795
rect 38615 -7915 38660 -7795
rect 38780 -7915 38825 -7795
rect 38945 -7915 38990 -7795
rect 39110 -7915 39165 -7795
rect 39285 -7915 39330 -7795
rect 39450 -7915 39495 -7795
rect 39615 -7915 39660 -7795
rect 39780 -7915 39835 -7795
rect 39955 -7915 40000 -7795
rect 40120 -7915 40165 -7795
rect 40285 -7915 40330 -7795
rect 40450 -7915 40505 -7795
rect 40625 -7915 40670 -7795
rect 40790 -7915 40835 -7795
rect 40955 -7915 41000 -7795
rect 41120 -7915 41175 -7795
rect 41295 -7915 41340 -7795
rect 41460 -7915 41505 -7795
rect 41625 -7915 41670 -7795
rect 41790 -7915 41845 -7795
rect 41965 -7915 42175 -7795
rect 42295 -7915 42340 -7795
rect 42460 -7915 42505 -7795
rect 42625 -7915 42670 -7795
rect 42790 -7915 42845 -7795
rect 42965 -7915 43010 -7795
rect 43130 -7915 43175 -7795
rect 43295 -7915 43340 -7795
rect 43460 -7915 43515 -7795
rect 43635 -7915 43680 -7795
rect 43800 -7915 43845 -7795
rect 43965 -7915 44010 -7795
rect 44130 -7915 44185 -7795
rect 44305 -7915 44350 -7795
rect 44470 -7915 44515 -7795
rect 44635 -7915 44680 -7795
rect 44800 -7915 44855 -7795
rect 44975 -7915 45020 -7795
rect 45140 -7915 45185 -7795
rect 45305 -7915 45350 -7795
rect 45470 -7915 45525 -7795
rect 45645 -7915 45690 -7795
rect 45810 -7915 45855 -7795
rect 45975 -7915 46020 -7795
rect 46140 -7915 46195 -7795
rect 46315 -7915 46360 -7795
rect 46480 -7915 46525 -7795
rect 46645 -7915 46690 -7795
rect 46810 -7915 46865 -7795
rect 46985 -7915 47030 -7795
rect 47150 -7915 47195 -7795
rect 47315 -7915 47360 -7795
rect 47480 -7915 47535 -7795
rect 47655 -7915 47865 -7795
rect 47985 -7915 48030 -7795
rect 48150 -7915 48195 -7795
rect 48315 -7915 48360 -7795
rect 48480 -7915 48535 -7795
rect 48655 -7915 48700 -7795
rect 48820 -7915 48865 -7795
rect 48985 -7915 49030 -7795
rect 49150 -7915 49205 -7795
rect 49325 -7915 49370 -7795
rect 49490 -7915 49535 -7795
rect 49655 -7915 49700 -7795
rect 49820 -7915 49875 -7795
rect 49995 -7915 50040 -7795
rect 50160 -7915 50205 -7795
rect 50325 -7915 50370 -7795
rect 50490 -7915 50545 -7795
rect 50665 -7915 50710 -7795
rect 50830 -7915 50875 -7795
rect 50995 -7915 51040 -7795
rect 51160 -7915 51215 -7795
rect 51335 -7915 51380 -7795
rect 51500 -7915 51545 -7795
rect 51665 -7915 51710 -7795
rect 51830 -7915 51885 -7795
rect 52005 -7915 52050 -7795
rect 52170 -7915 52215 -7795
rect 52335 -7915 52380 -7795
rect 52500 -7915 52555 -7795
rect 52675 -7915 52720 -7795
rect 52840 -7915 52885 -7795
rect 53005 -7915 53050 -7795
rect 53170 -7915 53225 -7795
rect 53345 -7915 53370 -7795
rect 30770 -7960 53370 -7915
rect 30770 -8080 30795 -7960
rect 30915 -8080 30960 -7960
rect 31080 -8080 31125 -7960
rect 31245 -8080 31290 -7960
rect 31410 -8080 31465 -7960
rect 31585 -8080 31630 -7960
rect 31750 -8080 31795 -7960
rect 31915 -8080 31960 -7960
rect 32080 -8080 32135 -7960
rect 32255 -8080 32300 -7960
rect 32420 -8080 32465 -7960
rect 32585 -8080 32630 -7960
rect 32750 -8080 32805 -7960
rect 32925 -8080 32970 -7960
rect 33090 -8080 33135 -7960
rect 33255 -8080 33300 -7960
rect 33420 -8080 33475 -7960
rect 33595 -8080 33640 -7960
rect 33760 -8080 33805 -7960
rect 33925 -8080 33970 -7960
rect 34090 -8080 34145 -7960
rect 34265 -8080 34310 -7960
rect 34430 -8080 34475 -7960
rect 34595 -8080 34640 -7960
rect 34760 -8080 34815 -7960
rect 34935 -8080 34980 -7960
rect 35100 -8080 35145 -7960
rect 35265 -8080 35310 -7960
rect 35430 -8080 35485 -7960
rect 35605 -8080 35650 -7960
rect 35770 -8080 35815 -7960
rect 35935 -8080 35980 -7960
rect 36100 -8080 36155 -7960
rect 36275 -8080 36485 -7960
rect 36605 -8080 36650 -7960
rect 36770 -8080 36815 -7960
rect 36935 -8080 36980 -7960
rect 37100 -8080 37155 -7960
rect 37275 -8080 37320 -7960
rect 37440 -8080 37485 -7960
rect 37605 -8080 37650 -7960
rect 37770 -8080 37825 -7960
rect 37945 -8080 37990 -7960
rect 38110 -8080 38155 -7960
rect 38275 -8080 38320 -7960
rect 38440 -8080 38495 -7960
rect 38615 -8080 38660 -7960
rect 38780 -8080 38825 -7960
rect 38945 -8080 38990 -7960
rect 39110 -8080 39165 -7960
rect 39285 -8080 39330 -7960
rect 39450 -8080 39495 -7960
rect 39615 -8080 39660 -7960
rect 39780 -8080 39835 -7960
rect 39955 -8080 40000 -7960
rect 40120 -8080 40165 -7960
rect 40285 -8080 40330 -7960
rect 40450 -8080 40505 -7960
rect 40625 -8080 40670 -7960
rect 40790 -8080 40835 -7960
rect 40955 -8080 41000 -7960
rect 41120 -8080 41175 -7960
rect 41295 -8080 41340 -7960
rect 41460 -8080 41505 -7960
rect 41625 -8080 41670 -7960
rect 41790 -8080 41845 -7960
rect 41965 -8080 42175 -7960
rect 42295 -8080 42340 -7960
rect 42460 -8080 42505 -7960
rect 42625 -8080 42670 -7960
rect 42790 -8080 42845 -7960
rect 42965 -8080 43010 -7960
rect 43130 -8080 43175 -7960
rect 43295 -8080 43340 -7960
rect 43460 -8080 43515 -7960
rect 43635 -8080 43680 -7960
rect 43800 -8080 43845 -7960
rect 43965 -8080 44010 -7960
rect 44130 -8080 44185 -7960
rect 44305 -8080 44350 -7960
rect 44470 -8080 44515 -7960
rect 44635 -8080 44680 -7960
rect 44800 -8080 44855 -7960
rect 44975 -8080 45020 -7960
rect 45140 -8080 45185 -7960
rect 45305 -8080 45350 -7960
rect 45470 -8080 45525 -7960
rect 45645 -8080 45690 -7960
rect 45810 -8080 45855 -7960
rect 45975 -8080 46020 -7960
rect 46140 -8080 46195 -7960
rect 46315 -8080 46360 -7960
rect 46480 -8080 46525 -7960
rect 46645 -8080 46690 -7960
rect 46810 -8080 46865 -7960
rect 46985 -8080 47030 -7960
rect 47150 -8080 47195 -7960
rect 47315 -8080 47360 -7960
rect 47480 -8080 47535 -7960
rect 47655 -8080 47865 -7960
rect 47985 -8080 48030 -7960
rect 48150 -8080 48195 -7960
rect 48315 -8080 48360 -7960
rect 48480 -8080 48535 -7960
rect 48655 -8080 48700 -7960
rect 48820 -8080 48865 -7960
rect 48985 -8080 49030 -7960
rect 49150 -8080 49205 -7960
rect 49325 -8080 49370 -7960
rect 49490 -8080 49535 -7960
rect 49655 -8080 49700 -7960
rect 49820 -8080 49875 -7960
rect 49995 -8080 50040 -7960
rect 50160 -8080 50205 -7960
rect 50325 -8080 50370 -7960
rect 50490 -8080 50545 -7960
rect 50665 -8080 50710 -7960
rect 50830 -8080 50875 -7960
rect 50995 -8080 51040 -7960
rect 51160 -8080 51215 -7960
rect 51335 -8080 51380 -7960
rect 51500 -8080 51545 -7960
rect 51665 -8080 51710 -7960
rect 51830 -8080 51885 -7960
rect 52005 -8080 52050 -7960
rect 52170 -8080 52215 -7960
rect 52335 -8080 52380 -7960
rect 52500 -8080 52555 -7960
rect 52675 -8080 52720 -7960
rect 52840 -8080 52885 -7960
rect 53005 -8080 53050 -7960
rect 53170 -8080 53225 -7960
rect 53345 -8080 53370 -7960
rect 30770 -8125 53370 -8080
rect 30770 -8245 30795 -8125
rect 30915 -8245 30960 -8125
rect 31080 -8245 31125 -8125
rect 31245 -8245 31290 -8125
rect 31410 -8245 31465 -8125
rect 31585 -8245 31630 -8125
rect 31750 -8245 31795 -8125
rect 31915 -8245 31960 -8125
rect 32080 -8245 32135 -8125
rect 32255 -8245 32300 -8125
rect 32420 -8245 32465 -8125
rect 32585 -8245 32630 -8125
rect 32750 -8245 32805 -8125
rect 32925 -8245 32970 -8125
rect 33090 -8245 33135 -8125
rect 33255 -8245 33300 -8125
rect 33420 -8245 33475 -8125
rect 33595 -8245 33640 -8125
rect 33760 -8245 33805 -8125
rect 33925 -8245 33970 -8125
rect 34090 -8245 34145 -8125
rect 34265 -8245 34310 -8125
rect 34430 -8245 34475 -8125
rect 34595 -8245 34640 -8125
rect 34760 -8245 34815 -8125
rect 34935 -8245 34980 -8125
rect 35100 -8245 35145 -8125
rect 35265 -8245 35310 -8125
rect 35430 -8245 35485 -8125
rect 35605 -8245 35650 -8125
rect 35770 -8245 35815 -8125
rect 35935 -8245 35980 -8125
rect 36100 -8245 36155 -8125
rect 36275 -8245 36485 -8125
rect 36605 -8245 36650 -8125
rect 36770 -8245 36815 -8125
rect 36935 -8245 36980 -8125
rect 37100 -8245 37155 -8125
rect 37275 -8245 37320 -8125
rect 37440 -8245 37485 -8125
rect 37605 -8245 37650 -8125
rect 37770 -8245 37825 -8125
rect 37945 -8245 37990 -8125
rect 38110 -8245 38155 -8125
rect 38275 -8245 38320 -8125
rect 38440 -8245 38495 -8125
rect 38615 -8245 38660 -8125
rect 38780 -8245 38825 -8125
rect 38945 -8245 38990 -8125
rect 39110 -8245 39165 -8125
rect 39285 -8245 39330 -8125
rect 39450 -8245 39495 -8125
rect 39615 -8245 39660 -8125
rect 39780 -8245 39835 -8125
rect 39955 -8245 40000 -8125
rect 40120 -8245 40165 -8125
rect 40285 -8245 40330 -8125
rect 40450 -8245 40505 -8125
rect 40625 -8245 40670 -8125
rect 40790 -8245 40835 -8125
rect 40955 -8245 41000 -8125
rect 41120 -8245 41175 -8125
rect 41295 -8245 41340 -8125
rect 41460 -8245 41505 -8125
rect 41625 -8245 41670 -8125
rect 41790 -8245 41845 -8125
rect 41965 -8245 42175 -8125
rect 42295 -8245 42340 -8125
rect 42460 -8245 42505 -8125
rect 42625 -8245 42670 -8125
rect 42790 -8245 42845 -8125
rect 42965 -8245 43010 -8125
rect 43130 -8245 43175 -8125
rect 43295 -8245 43340 -8125
rect 43460 -8245 43515 -8125
rect 43635 -8245 43680 -8125
rect 43800 -8245 43845 -8125
rect 43965 -8245 44010 -8125
rect 44130 -8245 44185 -8125
rect 44305 -8245 44350 -8125
rect 44470 -8245 44515 -8125
rect 44635 -8245 44680 -8125
rect 44800 -8245 44855 -8125
rect 44975 -8245 45020 -8125
rect 45140 -8245 45185 -8125
rect 45305 -8245 45350 -8125
rect 45470 -8245 45525 -8125
rect 45645 -8245 45690 -8125
rect 45810 -8245 45855 -8125
rect 45975 -8245 46020 -8125
rect 46140 -8245 46195 -8125
rect 46315 -8245 46360 -8125
rect 46480 -8245 46525 -8125
rect 46645 -8245 46690 -8125
rect 46810 -8245 46865 -8125
rect 46985 -8245 47030 -8125
rect 47150 -8245 47195 -8125
rect 47315 -8245 47360 -8125
rect 47480 -8245 47535 -8125
rect 47655 -8245 47865 -8125
rect 47985 -8245 48030 -8125
rect 48150 -8245 48195 -8125
rect 48315 -8245 48360 -8125
rect 48480 -8245 48535 -8125
rect 48655 -8245 48700 -8125
rect 48820 -8245 48865 -8125
rect 48985 -8245 49030 -8125
rect 49150 -8245 49205 -8125
rect 49325 -8245 49370 -8125
rect 49490 -8245 49535 -8125
rect 49655 -8245 49700 -8125
rect 49820 -8245 49875 -8125
rect 49995 -8245 50040 -8125
rect 50160 -8245 50205 -8125
rect 50325 -8245 50370 -8125
rect 50490 -8245 50545 -8125
rect 50665 -8245 50710 -8125
rect 50830 -8245 50875 -8125
rect 50995 -8245 51040 -8125
rect 51160 -8245 51215 -8125
rect 51335 -8245 51380 -8125
rect 51500 -8245 51545 -8125
rect 51665 -8245 51710 -8125
rect 51830 -8245 51885 -8125
rect 52005 -8245 52050 -8125
rect 52170 -8245 52215 -8125
rect 52335 -8245 52380 -8125
rect 52500 -8245 52555 -8125
rect 52675 -8245 52720 -8125
rect 52840 -8245 52885 -8125
rect 53005 -8245 53050 -8125
rect 53170 -8245 53225 -8125
rect 53345 -8245 53370 -8125
rect 30770 -8290 53370 -8245
rect 30770 -8410 30795 -8290
rect 30915 -8410 30960 -8290
rect 31080 -8410 31125 -8290
rect 31245 -8410 31290 -8290
rect 31410 -8410 31465 -8290
rect 31585 -8410 31630 -8290
rect 31750 -8410 31795 -8290
rect 31915 -8410 31960 -8290
rect 32080 -8410 32135 -8290
rect 32255 -8410 32300 -8290
rect 32420 -8410 32465 -8290
rect 32585 -8410 32630 -8290
rect 32750 -8410 32805 -8290
rect 32925 -8410 32970 -8290
rect 33090 -8410 33135 -8290
rect 33255 -8410 33300 -8290
rect 33420 -8410 33475 -8290
rect 33595 -8410 33640 -8290
rect 33760 -8410 33805 -8290
rect 33925 -8410 33970 -8290
rect 34090 -8410 34145 -8290
rect 34265 -8410 34310 -8290
rect 34430 -8410 34475 -8290
rect 34595 -8410 34640 -8290
rect 34760 -8410 34815 -8290
rect 34935 -8410 34980 -8290
rect 35100 -8410 35145 -8290
rect 35265 -8410 35310 -8290
rect 35430 -8410 35485 -8290
rect 35605 -8410 35650 -8290
rect 35770 -8410 35815 -8290
rect 35935 -8410 35980 -8290
rect 36100 -8410 36155 -8290
rect 36275 -8410 36485 -8290
rect 36605 -8410 36650 -8290
rect 36770 -8410 36815 -8290
rect 36935 -8410 36980 -8290
rect 37100 -8410 37155 -8290
rect 37275 -8410 37320 -8290
rect 37440 -8410 37485 -8290
rect 37605 -8410 37650 -8290
rect 37770 -8410 37825 -8290
rect 37945 -8410 37990 -8290
rect 38110 -8410 38155 -8290
rect 38275 -8410 38320 -8290
rect 38440 -8410 38495 -8290
rect 38615 -8410 38660 -8290
rect 38780 -8410 38825 -8290
rect 38945 -8410 38990 -8290
rect 39110 -8410 39165 -8290
rect 39285 -8410 39330 -8290
rect 39450 -8410 39495 -8290
rect 39615 -8410 39660 -8290
rect 39780 -8410 39835 -8290
rect 39955 -8410 40000 -8290
rect 40120 -8410 40165 -8290
rect 40285 -8410 40330 -8290
rect 40450 -8410 40505 -8290
rect 40625 -8410 40670 -8290
rect 40790 -8410 40835 -8290
rect 40955 -8410 41000 -8290
rect 41120 -8410 41175 -8290
rect 41295 -8410 41340 -8290
rect 41460 -8410 41505 -8290
rect 41625 -8410 41670 -8290
rect 41790 -8410 41845 -8290
rect 41965 -8410 42175 -8290
rect 42295 -8410 42340 -8290
rect 42460 -8410 42505 -8290
rect 42625 -8410 42670 -8290
rect 42790 -8410 42845 -8290
rect 42965 -8410 43010 -8290
rect 43130 -8410 43175 -8290
rect 43295 -8410 43340 -8290
rect 43460 -8410 43515 -8290
rect 43635 -8410 43680 -8290
rect 43800 -8410 43845 -8290
rect 43965 -8410 44010 -8290
rect 44130 -8410 44185 -8290
rect 44305 -8410 44350 -8290
rect 44470 -8410 44515 -8290
rect 44635 -8410 44680 -8290
rect 44800 -8410 44855 -8290
rect 44975 -8410 45020 -8290
rect 45140 -8410 45185 -8290
rect 45305 -8410 45350 -8290
rect 45470 -8410 45525 -8290
rect 45645 -8410 45690 -8290
rect 45810 -8410 45855 -8290
rect 45975 -8410 46020 -8290
rect 46140 -8410 46195 -8290
rect 46315 -8410 46360 -8290
rect 46480 -8410 46525 -8290
rect 46645 -8410 46690 -8290
rect 46810 -8410 46865 -8290
rect 46985 -8410 47030 -8290
rect 47150 -8410 47195 -8290
rect 47315 -8410 47360 -8290
rect 47480 -8410 47535 -8290
rect 47655 -8410 47865 -8290
rect 47985 -8410 48030 -8290
rect 48150 -8410 48195 -8290
rect 48315 -8410 48360 -8290
rect 48480 -8410 48535 -8290
rect 48655 -8410 48700 -8290
rect 48820 -8410 48865 -8290
rect 48985 -8410 49030 -8290
rect 49150 -8410 49205 -8290
rect 49325 -8410 49370 -8290
rect 49490 -8410 49535 -8290
rect 49655 -8410 49700 -8290
rect 49820 -8410 49875 -8290
rect 49995 -8410 50040 -8290
rect 50160 -8410 50205 -8290
rect 50325 -8410 50370 -8290
rect 50490 -8410 50545 -8290
rect 50665 -8410 50710 -8290
rect 50830 -8410 50875 -8290
rect 50995 -8410 51040 -8290
rect 51160 -8410 51215 -8290
rect 51335 -8410 51380 -8290
rect 51500 -8410 51545 -8290
rect 51665 -8410 51710 -8290
rect 51830 -8410 51885 -8290
rect 52005 -8410 52050 -8290
rect 52170 -8410 52215 -8290
rect 52335 -8410 52380 -8290
rect 52500 -8410 52555 -8290
rect 52675 -8410 52720 -8290
rect 52840 -8410 52885 -8290
rect 53005 -8410 53050 -8290
rect 53170 -8410 53225 -8290
rect 53345 -8410 53370 -8290
rect 30770 -8465 53370 -8410
rect 30770 -8585 30795 -8465
rect 30915 -8585 30960 -8465
rect 31080 -8585 31125 -8465
rect 31245 -8585 31290 -8465
rect 31410 -8585 31465 -8465
rect 31585 -8585 31630 -8465
rect 31750 -8585 31795 -8465
rect 31915 -8585 31960 -8465
rect 32080 -8585 32135 -8465
rect 32255 -8585 32300 -8465
rect 32420 -8585 32465 -8465
rect 32585 -8585 32630 -8465
rect 32750 -8585 32805 -8465
rect 32925 -8585 32970 -8465
rect 33090 -8585 33135 -8465
rect 33255 -8585 33300 -8465
rect 33420 -8585 33475 -8465
rect 33595 -8585 33640 -8465
rect 33760 -8585 33805 -8465
rect 33925 -8585 33970 -8465
rect 34090 -8585 34145 -8465
rect 34265 -8585 34310 -8465
rect 34430 -8585 34475 -8465
rect 34595 -8585 34640 -8465
rect 34760 -8585 34815 -8465
rect 34935 -8585 34980 -8465
rect 35100 -8585 35145 -8465
rect 35265 -8585 35310 -8465
rect 35430 -8585 35485 -8465
rect 35605 -8585 35650 -8465
rect 35770 -8585 35815 -8465
rect 35935 -8585 35980 -8465
rect 36100 -8585 36155 -8465
rect 36275 -8585 36485 -8465
rect 36605 -8585 36650 -8465
rect 36770 -8585 36815 -8465
rect 36935 -8585 36980 -8465
rect 37100 -8585 37155 -8465
rect 37275 -8585 37320 -8465
rect 37440 -8585 37485 -8465
rect 37605 -8585 37650 -8465
rect 37770 -8585 37825 -8465
rect 37945 -8585 37990 -8465
rect 38110 -8585 38155 -8465
rect 38275 -8585 38320 -8465
rect 38440 -8585 38495 -8465
rect 38615 -8585 38660 -8465
rect 38780 -8585 38825 -8465
rect 38945 -8585 38990 -8465
rect 39110 -8585 39165 -8465
rect 39285 -8585 39330 -8465
rect 39450 -8585 39495 -8465
rect 39615 -8585 39660 -8465
rect 39780 -8585 39835 -8465
rect 39955 -8585 40000 -8465
rect 40120 -8585 40165 -8465
rect 40285 -8585 40330 -8465
rect 40450 -8585 40505 -8465
rect 40625 -8585 40670 -8465
rect 40790 -8585 40835 -8465
rect 40955 -8585 41000 -8465
rect 41120 -8585 41175 -8465
rect 41295 -8585 41340 -8465
rect 41460 -8585 41505 -8465
rect 41625 -8585 41670 -8465
rect 41790 -8585 41845 -8465
rect 41965 -8585 42175 -8465
rect 42295 -8585 42340 -8465
rect 42460 -8585 42505 -8465
rect 42625 -8585 42670 -8465
rect 42790 -8585 42845 -8465
rect 42965 -8585 43010 -8465
rect 43130 -8585 43175 -8465
rect 43295 -8585 43340 -8465
rect 43460 -8585 43515 -8465
rect 43635 -8585 43680 -8465
rect 43800 -8585 43845 -8465
rect 43965 -8585 44010 -8465
rect 44130 -8585 44185 -8465
rect 44305 -8585 44350 -8465
rect 44470 -8585 44515 -8465
rect 44635 -8585 44680 -8465
rect 44800 -8585 44855 -8465
rect 44975 -8585 45020 -8465
rect 45140 -8585 45185 -8465
rect 45305 -8585 45350 -8465
rect 45470 -8585 45525 -8465
rect 45645 -8585 45690 -8465
rect 45810 -8585 45855 -8465
rect 45975 -8585 46020 -8465
rect 46140 -8585 46195 -8465
rect 46315 -8585 46360 -8465
rect 46480 -8585 46525 -8465
rect 46645 -8585 46690 -8465
rect 46810 -8585 46865 -8465
rect 46985 -8585 47030 -8465
rect 47150 -8585 47195 -8465
rect 47315 -8585 47360 -8465
rect 47480 -8585 47535 -8465
rect 47655 -8585 47865 -8465
rect 47985 -8585 48030 -8465
rect 48150 -8585 48195 -8465
rect 48315 -8585 48360 -8465
rect 48480 -8585 48535 -8465
rect 48655 -8585 48700 -8465
rect 48820 -8585 48865 -8465
rect 48985 -8585 49030 -8465
rect 49150 -8585 49205 -8465
rect 49325 -8585 49370 -8465
rect 49490 -8585 49535 -8465
rect 49655 -8585 49700 -8465
rect 49820 -8585 49875 -8465
rect 49995 -8585 50040 -8465
rect 50160 -8585 50205 -8465
rect 50325 -8585 50370 -8465
rect 50490 -8585 50545 -8465
rect 50665 -8585 50710 -8465
rect 50830 -8585 50875 -8465
rect 50995 -8585 51040 -8465
rect 51160 -8585 51215 -8465
rect 51335 -8585 51380 -8465
rect 51500 -8585 51545 -8465
rect 51665 -8585 51710 -8465
rect 51830 -8585 51885 -8465
rect 52005 -8585 52050 -8465
rect 52170 -8585 52215 -8465
rect 52335 -8585 52380 -8465
rect 52500 -8585 52555 -8465
rect 52675 -8585 52720 -8465
rect 52840 -8585 52885 -8465
rect 53005 -8585 53050 -8465
rect 53170 -8585 53225 -8465
rect 53345 -8585 53370 -8465
rect 30770 -8630 53370 -8585
rect 30770 -8750 30795 -8630
rect 30915 -8750 30960 -8630
rect 31080 -8750 31125 -8630
rect 31245 -8750 31290 -8630
rect 31410 -8750 31465 -8630
rect 31585 -8750 31630 -8630
rect 31750 -8750 31795 -8630
rect 31915 -8750 31960 -8630
rect 32080 -8750 32135 -8630
rect 32255 -8750 32300 -8630
rect 32420 -8750 32465 -8630
rect 32585 -8750 32630 -8630
rect 32750 -8750 32805 -8630
rect 32925 -8750 32970 -8630
rect 33090 -8750 33135 -8630
rect 33255 -8750 33300 -8630
rect 33420 -8750 33475 -8630
rect 33595 -8750 33640 -8630
rect 33760 -8750 33805 -8630
rect 33925 -8750 33970 -8630
rect 34090 -8750 34145 -8630
rect 34265 -8750 34310 -8630
rect 34430 -8750 34475 -8630
rect 34595 -8750 34640 -8630
rect 34760 -8750 34815 -8630
rect 34935 -8750 34980 -8630
rect 35100 -8750 35145 -8630
rect 35265 -8750 35310 -8630
rect 35430 -8750 35485 -8630
rect 35605 -8750 35650 -8630
rect 35770 -8750 35815 -8630
rect 35935 -8750 35980 -8630
rect 36100 -8750 36155 -8630
rect 36275 -8750 36485 -8630
rect 36605 -8750 36650 -8630
rect 36770 -8750 36815 -8630
rect 36935 -8750 36980 -8630
rect 37100 -8750 37155 -8630
rect 37275 -8750 37320 -8630
rect 37440 -8750 37485 -8630
rect 37605 -8750 37650 -8630
rect 37770 -8750 37825 -8630
rect 37945 -8750 37990 -8630
rect 38110 -8750 38155 -8630
rect 38275 -8750 38320 -8630
rect 38440 -8750 38495 -8630
rect 38615 -8750 38660 -8630
rect 38780 -8750 38825 -8630
rect 38945 -8750 38990 -8630
rect 39110 -8750 39165 -8630
rect 39285 -8750 39330 -8630
rect 39450 -8750 39495 -8630
rect 39615 -8750 39660 -8630
rect 39780 -8750 39835 -8630
rect 39955 -8750 40000 -8630
rect 40120 -8750 40165 -8630
rect 40285 -8750 40330 -8630
rect 40450 -8750 40505 -8630
rect 40625 -8750 40670 -8630
rect 40790 -8750 40835 -8630
rect 40955 -8750 41000 -8630
rect 41120 -8750 41175 -8630
rect 41295 -8750 41340 -8630
rect 41460 -8750 41505 -8630
rect 41625 -8750 41670 -8630
rect 41790 -8750 41845 -8630
rect 41965 -8750 42175 -8630
rect 42295 -8750 42340 -8630
rect 42460 -8750 42505 -8630
rect 42625 -8750 42670 -8630
rect 42790 -8750 42845 -8630
rect 42965 -8750 43010 -8630
rect 43130 -8750 43175 -8630
rect 43295 -8750 43340 -8630
rect 43460 -8750 43515 -8630
rect 43635 -8750 43680 -8630
rect 43800 -8750 43845 -8630
rect 43965 -8750 44010 -8630
rect 44130 -8750 44185 -8630
rect 44305 -8750 44350 -8630
rect 44470 -8750 44515 -8630
rect 44635 -8750 44680 -8630
rect 44800 -8750 44855 -8630
rect 44975 -8750 45020 -8630
rect 45140 -8750 45185 -8630
rect 45305 -8750 45350 -8630
rect 45470 -8750 45525 -8630
rect 45645 -8750 45690 -8630
rect 45810 -8750 45855 -8630
rect 45975 -8750 46020 -8630
rect 46140 -8750 46195 -8630
rect 46315 -8750 46360 -8630
rect 46480 -8750 46525 -8630
rect 46645 -8750 46690 -8630
rect 46810 -8750 46865 -8630
rect 46985 -8750 47030 -8630
rect 47150 -8750 47195 -8630
rect 47315 -8750 47360 -8630
rect 47480 -8750 47535 -8630
rect 47655 -8750 47865 -8630
rect 47985 -8750 48030 -8630
rect 48150 -8750 48195 -8630
rect 48315 -8750 48360 -8630
rect 48480 -8750 48535 -8630
rect 48655 -8750 48700 -8630
rect 48820 -8750 48865 -8630
rect 48985 -8750 49030 -8630
rect 49150 -8750 49205 -8630
rect 49325 -8750 49370 -8630
rect 49490 -8750 49535 -8630
rect 49655 -8750 49700 -8630
rect 49820 -8750 49875 -8630
rect 49995 -8750 50040 -8630
rect 50160 -8750 50205 -8630
rect 50325 -8750 50370 -8630
rect 50490 -8750 50545 -8630
rect 50665 -8750 50710 -8630
rect 50830 -8750 50875 -8630
rect 50995 -8750 51040 -8630
rect 51160 -8750 51215 -8630
rect 51335 -8750 51380 -8630
rect 51500 -8750 51545 -8630
rect 51665 -8750 51710 -8630
rect 51830 -8750 51885 -8630
rect 52005 -8750 52050 -8630
rect 52170 -8750 52215 -8630
rect 52335 -8750 52380 -8630
rect 52500 -8750 52555 -8630
rect 52675 -8750 52720 -8630
rect 52840 -8750 52885 -8630
rect 53005 -8750 53050 -8630
rect 53170 -8750 53225 -8630
rect 53345 -8750 53370 -8630
rect 30770 -8795 53370 -8750
rect 30770 -8915 30795 -8795
rect 30915 -8915 30960 -8795
rect 31080 -8915 31125 -8795
rect 31245 -8915 31290 -8795
rect 31410 -8915 31465 -8795
rect 31585 -8915 31630 -8795
rect 31750 -8915 31795 -8795
rect 31915 -8915 31960 -8795
rect 32080 -8915 32135 -8795
rect 32255 -8915 32300 -8795
rect 32420 -8915 32465 -8795
rect 32585 -8915 32630 -8795
rect 32750 -8915 32805 -8795
rect 32925 -8915 32970 -8795
rect 33090 -8915 33135 -8795
rect 33255 -8915 33300 -8795
rect 33420 -8915 33475 -8795
rect 33595 -8915 33640 -8795
rect 33760 -8915 33805 -8795
rect 33925 -8915 33970 -8795
rect 34090 -8915 34145 -8795
rect 34265 -8915 34310 -8795
rect 34430 -8915 34475 -8795
rect 34595 -8915 34640 -8795
rect 34760 -8915 34815 -8795
rect 34935 -8915 34980 -8795
rect 35100 -8915 35145 -8795
rect 35265 -8915 35310 -8795
rect 35430 -8915 35485 -8795
rect 35605 -8915 35650 -8795
rect 35770 -8915 35815 -8795
rect 35935 -8915 35980 -8795
rect 36100 -8915 36155 -8795
rect 36275 -8915 36485 -8795
rect 36605 -8915 36650 -8795
rect 36770 -8915 36815 -8795
rect 36935 -8915 36980 -8795
rect 37100 -8915 37155 -8795
rect 37275 -8915 37320 -8795
rect 37440 -8915 37485 -8795
rect 37605 -8915 37650 -8795
rect 37770 -8915 37825 -8795
rect 37945 -8915 37990 -8795
rect 38110 -8915 38155 -8795
rect 38275 -8915 38320 -8795
rect 38440 -8915 38495 -8795
rect 38615 -8915 38660 -8795
rect 38780 -8915 38825 -8795
rect 38945 -8915 38990 -8795
rect 39110 -8915 39165 -8795
rect 39285 -8915 39330 -8795
rect 39450 -8915 39495 -8795
rect 39615 -8915 39660 -8795
rect 39780 -8915 39835 -8795
rect 39955 -8915 40000 -8795
rect 40120 -8915 40165 -8795
rect 40285 -8915 40330 -8795
rect 40450 -8915 40505 -8795
rect 40625 -8915 40670 -8795
rect 40790 -8915 40835 -8795
rect 40955 -8915 41000 -8795
rect 41120 -8915 41175 -8795
rect 41295 -8915 41340 -8795
rect 41460 -8915 41505 -8795
rect 41625 -8915 41670 -8795
rect 41790 -8915 41845 -8795
rect 41965 -8915 42175 -8795
rect 42295 -8915 42340 -8795
rect 42460 -8915 42505 -8795
rect 42625 -8915 42670 -8795
rect 42790 -8915 42845 -8795
rect 42965 -8915 43010 -8795
rect 43130 -8915 43175 -8795
rect 43295 -8915 43340 -8795
rect 43460 -8915 43515 -8795
rect 43635 -8915 43680 -8795
rect 43800 -8915 43845 -8795
rect 43965 -8915 44010 -8795
rect 44130 -8915 44185 -8795
rect 44305 -8915 44350 -8795
rect 44470 -8915 44515 -8795
rect 44635 -8915 44680 -8795
rect 44800 -8915 44855 -8795
rect 44975 -8915 45020 -8795
rect 45140 -8915 45185 -8795
rect 45305 -8915 45350 -8795
rect 45470 -8915 45525 -8795
rect 45645 -8915 45690 -8795
rect 45810 -8915 45855 -8795
rect 45975 -8915 46020 -8795
rect 46140 -8915 46195 -8795
rect 46315 -8915 46360 -8795
rect 46480 -8915 46525 -8795
rect 46645 -8915 46690 -8795
rect 46810 -8915 46865 -8795
rect 46985 -8915 47030 -8795
rect 47150 -8915 47195 -8795
rect 47315 -8915 47360 -8795
rect 47480 -8915 47535 -8795
rect 47655 -8915 47865 -8795
rect 47985 -8915 48030 -8795
rect 48150 -8915 48195 -8795
rect 48315 -8915 48360 -8795
rect 48480 -8915 48535 -8795
rect 48655 -8915 48700 -8795
rect 48820 -8915 48865 -8795
rect 48985 -8915 49030 -8795
rect 49150 -8915 49205 -8795
rect 49325 -8915 49370 -8795
rect 49490 -8915 49535 -8795
rect 49655 -8915 49700 -8795
rect 49820 -8915 49875 -8795
rect 49995 -8915 50040 -8795
rect 50160 -8915 50205 -8795
rect 50325 -8915 50370 -8795
rect 50490 -8915 50545 -8795
rect 50665 -8915 50710 -8795
rect 50830 -8915 50875 -8795
rect 50995 -8915 51040 -8795
rect 51160 -8915 51215 -8795
rect 51335 -8915 51380 -8795
rect 51500 -8915 51545 -8795
rect 51665 -8915 51710 -8795
rect 51830 -8915 51885 -8795
rect 52005 -8915 52050 -8795
rect 52170 -8915 52215 -8795
rect 52335 -8915 52380 -8795
rect 52500 -8915 52555 -8795
rect 52675 -8915 52720 -8795
rect 52840 -8915 52885 -8795
rect 53005 -8915 53050 -8795
rect 53170 -8915 53225 -8795
rect 53345 -8915 53370 -8795
rect 30770 -8960 53370 -8915
rect 30770 -9080 30795 -8960
rect 30915 -9080 30960 -8960
rect 31080 -9080 31125 -8960
rect 31245 -9080 31290 -8960
rect 31410 -9080 31465 -8960
rect 31585 -9080 31630 -8960
rect 31750 -9080 31795 -8960
rect 31915 -9080 31960 -8960
rect 32080 -9080 32135 -8960
rect 32255 -9080 32300 -8960
rect 32420 -9080 32465 -8960
rect 32585 -9080 32630 -8960
rect 32750 -9080 32805 -8960
rect 32925 -9080 32970 -8960
rect 33090 -9080 33135 -8960
rect 33255 -9080 33300 -8960
rect 33420 -9080 33475 -8960
rect 33595 -9080 33640 -8960
rect 33760 -9080 33805 -8960
rect 33925 -9080 33970 -8960
rect 34090 -9080 34145 -8960
rect 34265 -9080 34310 -8960
rect 34430 -9080 34475 -8960
rect 34595 -9080 34640 -8960
rect 34760 -9080 34815 -8960
rect 34935 -9080 34980 -8960
rect 35100 -9080 35145 -8960
rect 35265 -9080 35310 -8960
rect 35430 -9080 35485 -8960
rect 35605 -9080 35650 -8960
rect 35770 -9080 35815 -8960
rect 35935 -9080 35980 -8960
rect 36100 -9080 36155 -8960
rect 36275 -9080 36485 -8960
rect 36605 -9080 36650 -8960
rect 36770 -9080 36815 -8960
rect 36935 -9080 36980 -8960
rect 37100 -9080 37155 -8960
rect 37275 -9080 37320 -8960
rect 37440 -9080 37485 -8960
rect 37605 -9080 37650 -8960
rect 37770 -9080 37825 -8960
rect 37945 -9080 37990 -8960
rect 38110 -9080 38155 -8960
rect 38275 -9080 38320 -8960
rect 38440 -9080 38495 -8960
rect 38615 -9080 38660 -8960
rect 38780 -9080 38825 -8960
rect 38945 -9080 38990 -8960
rect 39110 -9080 39165 -8960
rect 39285 -9080 39330 -8960
rect 39450 -9080 39495 -8960
rect 39615 -9080 39660 -8960
rect 39780 -9080 39835 -8960
rect 39955 -9080 40000 -8960
rect 40120 -9080 40165 -8960
rect 40285 -9080 40330 -8960
rect 40450 -9080 40505 -8960
rect 40625 -9080 40670 -8960
rect 40790 -9080 40835 -8960
rect 40955 -9080 41000 -8960
rect 41120 -9080 41175 -8960
rect 41295 -9080 41340 -8960
rect 41460 -9080 41505 -8960
rect 41625 -9080 41670 -8960
rect 41790 -9080 41845 -8960
rect 41965 -9080 42175 -8960
rect 42295 -9080 42340 -8960
rect 42460 -9080 42505 -8960
rect 42625 -9080 42670 -8960
rect 42790 -9080 42845 -8960
rect 42965 -9080 43010 -8960
rect 43130 -9080 43175 -8960
rect 43295 -9080 43340 -8960
rect 43460 -9080 43515 -8960
rect 43635 -9080 43680 -8960
rect 43800 -9080 43845 -8960
rect 43965 -9080 44010 -8960
rect 44130 -9080 44185 -8960
rect 44305 -9080 44350 -8960
rect 44470 -9080 44515 -8960
rect 44635 -9080 44680 -8960
rect 44800 -9080 44855 -8960
rect 44975 -9080 45020 -8960
rect 45140 -9080 45185 -8960
rect 45305 -9080 45350 -8960
rect 45470 -9080 45525 -8960
rect 45645 -9080 45690 -8960
rect 45810 -9080 45855 -8960
rect 45975 -9080 46020 -8960
rect 46140 -9080 46195 -8960
rect 46315 -9080 46360 -8960
rect 46480 -9080 46525 -8960
rect 46645 -9080 46690 -8960
rect 46810 -9080 46865 -8960
rect 46985 -9080 47030 -8960
rect 47150 -9080 47195 -8960
rect 47315 -9080 47360 -8960
rect 47480 -9080 47535 -8960
rect 47655 -9080 47865 -8960
rect 47985 -9080 48030 -8960
rect 48150 -9080 48195 -8960
rect 48315 -9080 48360 -8960
rect 48480 -9080 48535 -8960
rect 48655 -9080 48700 -8960
rect 48820 -9080 48865 -8960
rect 48985 -9080 49030 -8960
rect 49150 -9080 49205 -8960
rect 49325 -9080 49370 -8960
rect 49490 -9080 49535 -8960
rect 49655 -9080 49700 -8960
rect 49820 -9080 49875 -8960
rect 49995 -9080 50040 -8960
rect 50160 -9080 50205 -8960
rect 50325 -9080 50370 -8960
rect 50490 -9080 50545 -8960
rect 50665 -9080 50710 -8960
rect 50830 -9080 50875 -8960
rect 50995 -9080 51040 -8960
rect 51160 -9080 51215 -8960
rect 51335 -9080 51380 -8960
rect 51500 -9080 51545 -8960
rect 51665 -9080 51710 -8960
rect 51830 -9080 51885 -8960
rect 52005 -9080 52050 -8960
rect 52170 -9080 52215 -8960
rect 52335 -9080 52380 -8960
rect 52500 -9080 52555 -8960
rect 52675 -9080 52720 -8960
rect 52840 -9080 52885 -8960
rect 53005 -9080 53050 -8960
rect 53170 -9080 53225 -8960
rect 53345 -9080 53370 -8960
rect 30770 -9135 53370 -9080
rect 30770 -9255 30795 -9135
rect 30915 -9255 30960 -9135
rect 31080 -9255 31125 -9135
rect 31245 -9255 31290 -9135
rect 31410 -9255 31465 -9135
rect 31585 -9255 31630 -9135
rect 31750 -9255 31795 -9135
rect 31915 -9255 31960 -9135
rect 32080 -9255 32135 -9135
rect 32255 -9255 32300 -9135
rect 32420 -9255 32465 -9135
rect 32585 -9255 32630 -9135
rect 32750 -9255 32805 -9135
rect 32925 -9255 32970 -9135
rect 33090 -9255 33135 -9135
rect 33255 -9255 33300 -9135
rect 33420 -9255 33475 -9135
rect 33595 -9255 33640 -9135
rect 33760 -9255 33805 -9135
rect 33925 -9255 33970 -9135
rect 34090 -9255 34145 -9135
rect 34265 -9255 34310 -9135
rect 34430 -9255 34475 -9135
rect 34595 -9255 34640 -9135
rect 34760 -9255 34815 -9135
rect 34935 -9255 34980 -9135
rect 35100 -9255 35145 -9135
rect 35265 -9255 35310 -9135
rect 35430 -9255 35485 -9135
rect 35605 -9255 35650 -9135
rect 35770 -9255 35815 -9135
rect 35935 -9255 35980 -9135
rect 36100 -9255 36155 -9135
rect 36275 -9255 36485 -9135
rect 36605 -9255 36650 -9135
rect 36770 -9255 36815 -9135
rect 36935 -9255 36980 -9135
rect 37100 -9255 37155 -9135
rect 37275 -9255 37320 -9135
rect 37440 -9255 37485 -9135
rect 37605 -9255 37650 -9135
rect 37770 -9255 37825 -9135
rect 37945 -9255 37990 -9135
rect 38110 -9255 38155 -9135
rect 38275 -9255 38320 -9135
rect 38440 -9255 38495 -9135
rect 38615 -9255 38660 -9135
rect 38780 -9255 38825 -9135
rect 38945 -9255 38990 -9135
rect 39110 -9255 39165 -9135
rect 39285 -9255 39330 -9135
rect 39450 -9255 39495 -9135
rect 39615 -9255 39660 -9135
rect 39780 -9255 39835 -9135
rect 39955 -9255 40000 -9135
rect 40120 -9255 40165 -9135
rect 40285 -9255 40330 -9135
rect 40450 -9255 40505 -9135
rect 40625 -9255 40670 -9135
rect 40790 -9255 40835 -9135
rect 40955 -9255 41000 -9135
rect 41120 -9255 41175 -9135
rect 41295 -9255 41340 -9135
rect 41460 -9255 41505 -9135
rect 41625 -9255 41670 -9135
rect 41790 -9255 41845 -9135
rect 41965 -9255 42175 -9135
rect 42295 -9255 42340 -9135
rect 42460 -9255 42505 -9135
rect 42625 -9255 42670 -9135
rect 42790 -9255 42845 -9135
rect 42965 -9255 43010 -9135
rect 43130 -9255 43175 -9135
rect 43295 -9255 43340 -9135
rect 43460 -9255 43515 -9135
rect 43635 -9255 43680 -9135
rect 43800 -9255 43845 -9135
rect 43965 -9255 44010 -9135
rect 44130 -9255 44185 -9135
rect 44305 -9255 44350 -9135
rect 44470 -9255 44515 -9135
rect 44635 -9255 44680 -9135
rect 44800 -9255 44855 -9135
rect 44975 -9255 45020 -9135
rect 45140 -9255 45185 -9135
rect 45305 -9255 45350 -9135
rect 45470 -9255 45525 -9135
rect 45645 -9255 45690 -9135
rect 45810 -9255 45855 -9135
rect 45975 -9255 46020 -9135
rect 46140 -9255 46195 -9135
rect 46315 -9255 46360 -9135
rect 46480 -9255 46525 -9135
rect 46645 -9255 46690 -9135
rect 46810 -9255 46865 -9135
rect 46985 -9255 47030 -9135
rect 47150 -9255 47195 -9135
rect 47315 -9255 47360 -9135
rect 47480 -9255 47535 -9135
rect 47655 -9255 47865 -9135
rect 47985 -9255 48030 -9135
rect 48150 -9255 48195 -9135
rect 48315 -9255 48360 -9135
rect 48480 -9255 48535 -9135
rect 48655 -9255 48700 -9135
rect 48820 -9255 48865 -9135
rect 48985 -9255 49030 -9135
rect 49150 -9255 49205 -9135
rect 49325 -9255 49370 -9135
rect 49490 -9255 49535 -9135
rect 49655 -9255 49700 -9135
rect 49820 -9255 49875 -9135
rect 49995 -9255 50040 -9135
rect 50160 -9255 50205 -9135
rect 50325 -9255 50370 -9135
rect 50490 -9255 50545 -9135
rect 50665 -9255 50710 -9135
rect 50830 -9255 50875 -9135
rect 50995 -9255 51040 -9135
rect 51160 -9255 51215 -9135
rect 51335 -9255 51380 -9135
rect 51500 -9255 51545 -9135
rect 51665 -9255 51710 -9135
rect 51830 -9255 51885 -9135
rect 52005 -9255 52050 -9135
rect 52170 -9255 52215 -9135
rect 52335 -9255 52380 -9135
rect 52500 -9255 52555 -9135
rect 52675 -9255 52720 -9135
rect 52840 -9255 52885 -9135
rect 53005 -9255 53050 -9135
rect 53170 -9255 53225 -9135
rect 53345 -9255 53370 -9135
rect 30770 -9300 53370 -9255
rect 30770 -9420 30795 -9300
rect 30915 -9420 30960 -9300
rect 31080 -9420 31125 -9300
rect 31245 -9420 31290 -9300
rect 31410 -9420 31465 -9300
rect 31585 -9420 31630 -9300
rect 31750 -9420 31795 -9300
rect 31915 -9420 31960 -9300
rect 32080 -9420 32135 -9300
rect 32255 -9420 32300 -9300
rect 32420 -9420 32465 -9300
rect 32585 -9420 32630 -9300
rect 32750 -9420 32805 -9300
rect 32925 -9420 32970 -9300
rect 33090 -9420 33135 -9300
rect 33255 -9420 33300 -9300
rect 33420 -9420 33475 -9300
rect 33595 -9420 33640 -9300
rect 33760 -9420 33805 -9300
rect 33925 -9420 33970 -9300
rect 34090 -9420 34145 -9300
rect 34265 -9420 34310 -9300
rect 34430 -9420 34475 -9300
rect 34595 -9420 34640 -9300
rect 34760 -9420 34815 -9300
rect 34935 -9420 34980 -9300
rect 35100 -9420 35145 -9300
rect 35265 -9420 35310 -9300
rect 35430 -9420 35485 -9300
rect 35605 -9420 35650 -9300
rect 35770 -9420 35815 -9300
rect 35935 -9420 35980 -9300
rect 36100 -9420 36155 -9300
rect 36275 -9420 36485 -9300
rect 36605 -9420 36650 -9300
rect 36770 -9420 36815 -9300
rect 36935 -9420 36980 -9300
rect 37100 -9420 37155 -9300
rect 37275 -9420 37320 -9300
rect 37440 -9420 37485 -9300
rect 37605 -9420 37650 -9300
rect 37770 -9420 37825 -9300
rect 37945 -9420 37990 -9300
rect 38110 -9420 38155 -9300
rect 38275 -9420 38320 -9300
rect 38440 -9420 38495 -9300
rect 38615 -9420 38660 -9300
rect 38780 -9420 38825 -9300
rect 38945 -9420 38990 -9300
rect 39110 -9420 39165 -9300
rect 39285 -9420 39330 -9300
rect 39450 -9420 39495 -9300
rect 39615 -9420 39660 -9300
rect 39780 -9420 39835 -9300
rect 39955 -9420 40000 -9300
rect 40120 -9420 40165 -9300
rect 40285 -9420 40330 -9300
rect 40450 -9420 40505 -9300
rect 40625 -9420 40670 -9300
rect 40790 -9420 40835 -9300
rect 40955 -9420 41000 -9300
rect 41120 -9420 41175 -9300
rect 41295 -9420 41340 -9300
rect 41460 -9420 41505 -9300
rect 41625 -9420 41670 -9300
rect 41790 -9420 41845 -9300
rect 41965 -9420 42175 -9300
rect 42295 -9420 42340 -9300
rect 42460 -9420 42505 -9300
rect 42625 -9420 42670 -9300
rect 42790 -9420 42845 -9300
rect 42965 -9420 43010 -9300
rect 43130 -9420 43175 -9300
rect 43295 -9420 43340 -9300
rect 43460 -9420 43515 -9300
rect 43635 -9420 43680 -9300
rect 43800 -9420 43845 -9300
rect 43965 -9420 44010 -9300
rect 44130 -9420 44185 -9300
rect 44305 -9420 44350 -9300
rect 44470 -9420 44515 -9300
rect 44635 -9420 44680 -9300
rect 44800 -9420 44855 -9300
rect 44975 -9420 45020 -9300
rect 45140 -9420 45185 -9300
rect 45305 -9420 45350 -9300
rect 45470 -9420 45525 -9300
rect 45645 -9420 45690 -9300
rect 45810 -9420 45855 -9300
rect 45975 -9420 46020 -9300
rect 46140 -9420 46195 -9300
rect 46315 -9420 46360 -9300
rect 46480 -9420 46525 -9300
rect 46645 -9420 46690 -9300
rect 46810 -9420 46865 -9300
rect 46985 -9420 47030 -9300
rect 47150 -9420 47195 -9300
rect 47315 -9420 47360 -9300
rect 47480 -9420 47535 -9300
rect 47655 -9420 47865 -9300
rect 47985 -9420 48030 -9300
rect 48150 -9420 48195 -9300
rect 48315 -9420 48360 -9300
rect 48480 -9420 48535 -9300
rect 48655 -9420 48700 -9300
rect 48820 -9420 48865 -9300
rect 48985 -9420 49030 -9300
rect 49150 -9420 49205 -9300
rect 49325 -9420 49370 -9300
rect 49490 -9420 49535 -9300
rect 49655 -9420 49700 -9300
rect 49820 -9420 49875 -9300
rect 49995 -9420 50040 -9300
rect 50160 -9420 50205 -9300
rect 50325 -9420 50370 -9300
rect 50490 -9420 50545 -9300
rect 50665 -9420 50710 -9300
rect 50830 -9420 50875 -9300
rect 50995 -9420 51040 -9300
rect 51160 -9420 51215 -9300
rect 51335 -9420 51380 -9300
rect 51500 -9420 51545 -9300
rect 51665 -9420 51710 -9300
rect 51830 -9420 51885 -9300
rect 52005 -9420 52050 -9300
rect 52170 -9420 52215 -9300
rect 52335 -9420 52380 -9300
rect 52500 -9420 52555 -9300
rect 52675 -9420 52720 -9300
rect 52840 -9420 52885 -9300
rect 53005 -9420 53050 -9300
rect 53170 -9420 53225 -9300
rect 53345 -9420 53370 -9300
rect 30770 -9465 53370 -9420
rect 30770 -9585 30795 -9465
rect 30915 -9585 30960 -9465
rect 31080 -9585 31125 -9465
rect 31245 -9585 31290 -9465
rect 31410 -9585 31465 -9465
rect 31585 -9585 31630 -9465
rect 31750 -9585 31795 -9465
rect 31915 -9585 31960 -9465
rect 32080 -9585 32135 -9465
rect 32255 -9585 32300 -9465
rect 32420 -9585 32465 -9465
rect 32585 -9585 32630 -9465
rect 32750 -9585 32805 -9465
rect 32925 -9585 32970 -9465
rect 33090 -9585 33135 -9465
rect 33255 -9585 33300 -9465
rect 33420 -9585 33475 -9465
rect 33595 -9585 33640 -9465
rect 33760 -9585 33805 -9465
rect 33925 -9585 33970 -9465
rect 34090 -9585 34145 -9465
rect 34265 -9585 34310 -9465
rect 34430 -9585 34475 -9465
rect 34595 -9585 34640 -9465
rect 34760 -9585 34815 -9465
rect 34935 -9585 34980 -9465
rect 35100 -9585 35145 -9465
rect 35265 -9585 35310 -9465
rect 35430 -9585 35485 -9465
rect 35605 -9585 35650 -9465
rect 35770 -9585 35815 -9465
rect 35935 -9585 35980 -9465
rect 36100 -9585 36155 -9465
rect 36275 -9585 36485 -9465
rect 36605 -9585 36650 -9465
rect 36770 -9585 36815 -9465
rect 36935 -9585 36980 -9465
rect 37100 -9585 37155 -9465
rect 37275 -9585 37320 -9465
rect 37440 -9585 37485 -9465
rect 37605 -9585 37650 -9465
rect 37770 -9585 37825 -9465
rect 37945 -9585 37990 -9465
rect 38110 -9585 38155 -9465
rect 38275 -9585 38320 -9465
rect 38440 -9585 38495 -9465
rect 38615 -9585 38660 -9465
rect 38780 -9585 38825 -9465
rect 38945 -9585 38990 -9465
rect 39110 -9585 39165 -9465
rect 39285 -9585 39330 -9465
rect 39450 -9585 39495 -9465
rect 39615 -9585 39660 -9465
rect 39780 -9585 39835 -9465
rect 39955 -9585 40000 -9465
rect 40120 -9585 40165 -9465
rect 40285 -9585 40330 -9465
rect 40450 -9585 40505 -9465
rect 40625 -9585 40670 -9465
rect 40790 -9585 40835 -9465
rect 40955 -9585 41000 -9465
rect 41120 -9585 41175 -9465
rect 41295 -9585 41340 -9465
rect 41460 -9585 41505 -9465
rect 41625 -9585 41670 -9465
rect 41790 -9585 41845 -9465
rect 41965 -9585 42175 -9465
rect 42295 -9585 42340 -9465
rect 42460 -9585 42505 -9465
rect 42625 -9585 42670 -9465
rect 42790 -9585 42845 -9465
rect 42965 -9585 43010 -9465
rect 43130 -9585 43175 -9465
rect 43295 -9585 43340 -9465
rect 43460 -9585 43515 -9465
rect 43635 -9585 43680 -9465
rect 43800 -9585 43845 -9465
rect 43965 -9585 44010 -9465
rect 44130 -9585 44185 -9465
rect 44305 -9585 44350 -9465
rect 44470 -9585 44515 -9465
rect 44635 -9585 44680 -9465
rect 44800 -9585 44855 -9465
rect 44975 -9585 45020 -9465
rect 45140 -9585 45185 -9465
rect 45305 -9585 45350 -9465
rect 45470 -9585 45525 -9465
rect 45645 -9585 45690 -9465
rect 45810 -9585 45855 -9465
rect 45975 -9585 46020 -9465
rect 46140 -9585 46195 -9465
rect 46315 -9585 46360 -9465
rect 46480 -9585 46525 -9465
rect 46645 -9585 46690 -9465
rect 46810 -9585 46865 -9465
rect 46985 -9585 47030 -9465
rect 47150 -9585 47195 -9465
rect 47315 -9585 47360 -9465
rect 47480 -9585 47535 -9465
rect 47655 -9585 47865 -9465
rect 47985 -9585 48030 -9465
rect 48150 -9585 48195 -9465
rect 48315 -9585 48360 -9465
rect 48480 -9585 48535 -9465
rect 48655 -9585 48700 -9465
rect 48820 -9585 48865 -9465
rect 48985 -9585 49030 -9465
rect 49150 -9585 49205 -9465
rect 49325 -9585 49370 -9465
rect 49490 -9585 49535 -9465
rect 49655 -9585 49700 -9465
rect 49820 -9585 49875 -9465
rect 49995 -9585 50040 -9465
rect 50160 -9585 50205 -9465
rect 50325 -9585 50370 -9465
rect 50490 -9585 50545 -9465
rect 50665 -9585 50710 -9465
rect 50830 -9585 50875 -9465
rect 50995 -9585 51040 -9465
rect 51160 -9585 51215 -9465
rect 51335 -9585 51380 -9465
rect 51500 -9585 51545 -9465
rect 51665 -9585 51710 -9465
rect 51830 -9585 51885 -9465
rect 52005 -9585 52050 -9465
rect 52170 -9585 52215 -9465
rect 52335 -9585 52380 -9465
rect 52500 -9585 52555 -9465
rect 52675 -9585 52720 -9465
rect 52840 -9585 52885 -9465
rect 53005 -9585 53050 -9465
rect 53170 -9585 53225 -9465
rect 53345 -9585 53370 -9465
rect 30770 -9630 53370 -9585
rect 30770 -9750 30795 -9630
rect 30915 -9750 30960 -9630
rect 31080 -9750 31125 -9630
rect 31245 -9750 31290 -9630
rect 31410 -9750 31465 -9630
rect 31585 -9750 31630 -9630
rect 31750 -9750 31795 -9630
rect 31915 -9750 31960 -9630
rect 32080 -9750 32135 -9630
rect 32255 -9750 32300 -9630
rect 32420 -9750 32465 -9630
rect 32585 -9750 32630 -9630
rect 32750 -9750 32805 -9630
rect 32925 -9750 32970 -9630
rect 33090 -9750 33135 -9630
rect 33255 -9750 33300 -9630
rect 33420 -9750 33475 -9630
rect 33595 -9750 33640 -9630
rect 33760 -9750 33805 -9630
rect 33925 -9750 33970 -9630
rect 34090 -9750 34145 -9630
rect 34265 -9750 34310 -9630
rect 34430 -9750 34475 -9630
rect 34595 -9750 34640 -9630
rect 34760 -9750 34815 -9630
rect 34935 -9750 34980 -9630
rect 35100 -9750 35145 -9630
rect 35265 -9750 35310 -9630
rect 35430 -9750 35485 -9630
rect 35605 -9750 35650 -9630
rect 35770 -9750 35815 -9630
rect 35935 -9750 35980 -9630
rect 36100 -9750 36155 -9630
rect 36275 -9750 36485 -9630
rect 36605 -9750 36650 -9630
rect 36770 -9750 36815 -9630
rect 36935 -9750 36980 -9630
rect 37100 -9750 37155 -9630
rect 37275 -9750 37320 -9630
rect 37440 -9750 37485 -9630
rect 37605 -9750 37650 -9630
rect 37770 -9750 37825 -9630
rect 37945 -9750 37990 -9630
rect 38110 -9750 38155 -9630
rect 38275 -9750 38320 -9630
rect 38440 -9750 38495 -9630
rect 38615 -9750 38660 -9630
rect 38780 -9750 38825 -9630
rect 38945 -9750 38990 -9630
rect 39110 -9750 39165 -9630
rect 39285 -9750 39330 -9630
rect 39450 -9750 39495 -9630
rect 39615 -9750 39660 -9630
rect 39780 -9750 39835 -9630
rect 39955 -9750 40000 -9630
rect 40120 -9750 40165 -9630
rect 40285 -9750 40330 -9630
rect 40450 -9750 40505 -9630
rect 40625 -9750 40670 -9630
rect 40790 -9750 40835 -9630
rect 40955 -9750 41000 -9630
rect 41120 -9750 41175 -9630
rect 41295 -9750 41340 -9630
rect 41460 -9750 41505 -9630
rect 41625 -9750 41670 -9630
rect 41790 -9750 41845 -9630
rect 41965 -9750 42175 -9630
rect 42295 -9750 42340 -9630
rect 42460 -9750 42505 -9630
rect 42625 -9750 42670 -9630
rect 42790 -9750 42845 -9630
rect 42965 -9750 43010 -9630
rect 43130 -9750 43175 -9630
rect 43295 -9750 43340 -9630
rect 43460 -9750 43515 -9630
rect 43635 -9750 43680 -9630
rect 43800 -9750 43845 -9630
rect 43965 -9750 44010 -9630
rect 44130 -9750 44185 -9630
rect 44305 -9750 44350 -9630
rect 44470 -9750 44515 -9630
rect 44635 -9750 44680 -9630
rect 44800 -9750 44855 -9630
rect 44975 -9750 45020 -9630
rect 45140 -9750 45185 -9630
rect 45305 -9750 45350 -9630
rect 45470 -9750 45525 -9630
rect 45645 -9750 45690 -9630
rect 45810 -9750 45855 -9630
rect 45975 -9750 46020 -9630
rect 46140 -9750 46195 -9630
rect 46315 -9750 46360 -9630
rect 46480 -9750 46525 -9630
rect 46645 -9750 46690 -9630
rect 46810 -9750 46865 -9630
rect 46985 -9750 47030 -9630
rect 47150 -9750 47195 -9630
rect 47315 -9750 47360 -9630
rect 47480 -9750 47535 -9630
rect 47655 -9750 47865 -9630
rect 47985 -9750 48030 -9630
rect 48150 -9750 48195 -9630
rect 48315 -9750 48360 -9630
rect 48480 -9750 48535 -9630
rect 48655 -9750 48700 -9630
rect 48820 -9750 48865 -9630
rect 48985 -9750 49030 -9630
rect 49150 -9750 49205 -9630
rect 49325 -9750 49370 -9630
rect 49490 -9750 49535 -9630
rect 49655 -9750 49700 -9630
rect 49820 -9750 49875 -9630
rect 49995 -9750 50040 -9630
rect 50160 -9750 50205 -9630
rect 50325 -9750 50370 -9630
rect 50490 -9750 50545 -9630
rect 50665 -9750 50710 -9630
rect 50830 -9750 50875 -9630
rect 50995 -9750 51040 -9630
rect 51160 -9750 51215 -9630
rect 51335 -9750 51380 -9630
rect 51500 -9750 51545 -9630
rect 51665 -9750 51710 -9630
rect 51830 -9750 51885 -9630
rect 52005 -9750 52050 -9630
rect 52170 -9750 52215 -9630
rect 52335 -9750 52380 -9630
rect 52500 -9750 52555 -9630
rect 52675 -9750 52720 -9630
rect 52840 -9750 52885 -9630
rect 53005 -9750 53050 -9630
rect 53170 -9750 53225 -9630
rect 53345 -9750 53370 -9630
rect 30770 -9840 53370 -9750
rect 30770 -9960 30835 -9840
rect 30955 -9960 31000 -9840
rect 31120 -9960 31165 -9840
rect 31285 -9960 31330 -9840
rect 31450 -9960 31495 -9840
rect 31615 -9960 31660 -9840
rect 31780 -9960 31825 -9840
rect 31945 -9960 31990 -9840
rect 32110 -9960 32155 -9840
rect 32275 -9960 32320 -9840
rect 32440 -9960 32485 -9840
rect 32605 -9960 32650 -9840
rect 32770 -9960 32815 -9840
rect 32935 -9960 32980 -9840
rect 33100 -9960 33145 -9840
rect 33265 -9960 33310 -9840
rect 33430 -9960 33475 -9840
rect 33595 -9960 33640 -9840
rect 33760 -9960 33805 -9840
rect 33925 -9960 33970 -9840
rect 34090 -9960 34135 -9840
rect 34255 -9960 34300 -9840
rect 34420 -9960 34465 -9840
rect 34585 -9960 34630 -9840
rect 34750 -9960 34795 -9840
rect 34915 -9960 34960 -9840
rect 35080 -9960 35125 -9840
rect 35245 -9960 35290 -9840
rect 35410 -9960 35455 -9840
rect 35575 -9960 35620 -9840
rect 35740 -9960 35785 -9840
rect 35905 -9960 35950 -9840
rect 36070 -9960 36115 -9840
rect 36235 -9960 36525 -9840
rect 36645 -9960 36690 -9840
rect 36810 -9960 36855 -9840
rect 36975 -9960 37020 -9840
rect 37140 -9960 37185 -9840
rect 37305 -9960 37350 -9840
rect 37470 -9960 37515 -9840
rect 37635 -9960 37680 -9840
rect 37800 -9960 37845 -9840
rect 37965 -9960 38010 -9840
rect 38130 -9960 38175 -9840
rect 38295 -9960 38340 -9840
rect 38460 -9960 38505 -9840
rect 38625 -9960 38670 -9840
rect 38790 -9960 38835 -9840
rect 38955 -9960 39000 -9840
rect 39120 -9960 39165 -9840
rect 39285 -9960 39330 -9840
rect 39450 -9960 39495 -9840
rect 39615 -9960 39660 -9840
rect 39780 -9960 39825 -9840
rect 39945 -9960 39990 -9840
rect 40110 -9960 40155 -9840
rect 40275 -9960 40320 -9840
rect 40440 -9960 40485 -9840
rect 40605 -9960 40650 -9840
rect 40770 -9960 40815 -9840
rect 40935 -9960 40980 -9840
rect 41100 -9960 41145 -9840
rect 41265 -9960 41310 -9840
rect 41430 -9960 41475 -9840
rect 41595 -9960 41640 -9840
rect 41760 -9960 41805 -9840
rect 41925 -9960 42215 -9840
rect 42335 -9960 42380 -9840
rect 42500 -9960 42545 -9840
rect 42665 -9960 42710 -9840
rect 42830 -9960 42875 -9840
rect 42995 -9960 43040 -9840
rect 43160 -9960 43205 -9840
rect 43325 -9960 43370 -9840
rect 43490 -9960 43535 -9840
rect 43655 -9960 43700 -9840
rect 43820 -9960 43865 -9840
rect 43985 -9960 44030 -9840
rect 44150 -9960 44195 -9840
rect 44315 -9960 44360 -9840
rect 44480 -9960 44525 -9840
rect 44645 -9960 44690 -9840
rect 44810 -9960 44855 -9840
rect 44975 -9960 45020 -9840
rect 45140 -9960 45185 -9840
rect 45305 -9960 45350 -9840
rect 45470 -9960 45515 -9840
rect 45635 -9960 45680 -9840
rect 45800 -9960 45845 -9840
rect 45965 -9960 46010 -9840
rect 46130 -9960 46175 -9840
rect 46295 -9960 46340 -9840
rect 46460 -9960 46505 -9840
rect 46625 -9960 46670 -9840
rect 46790 -9960 46835 -9840
rect 46955 -9960 47000 -9840
rect 47120 -9960 47165 -9840
rect 47285 -9960 47330 -9840
rect 47450 -9960 47495 -9840
rect 47615 -9960 47905 -9840
rect 48025 -9960 48070 -9840
rect 48190 -9960 48235 -9840
rect 48355 -9960 48400 -9840
rect 48520 -9960 48565 -9840
rect 48685 -9960 48730 -9840
rect 48850 -9960 48895 -9840
rect 49015 -9960 49060 -9840
rect 49180 -9960 49225 -9840
rect 49345 -9960 49390 -9840
rect 49510 -9960 49555 -9840
rect 49675 -9960 49720 -9840
rect 49840 -9960 49885 -9840
rect 50005 -9960 50050 -9840
rect 50170 -9960 50215 -9840
rect 50335 -9960 50380 -9840
rect 50500 -9960 50545 -9840
rect 50665 -9960 50710 -9840
rect 50830 -9960 50875 -9840
rect 50995 -9960 51040 -9840
rect 51160 -9960 51205 -9840
rect 51325 -9960 51370 -9840
rect 51490 -9960 51535 -9840
rect 51655 -9960 51700 -9840
rect 51820 -9960 51865 -9840
rect 51985 -9960 52030 -9840
rect 52150 -9960 52195 -9840
rect 52315 -9960 52360 -9840
rect 52480 -9960 52525 -9840
rect 52645 -9960 52690 -9840
rect 52810 -9960 52855 -9840
rect 52975 -9960 53020 -9840
rect 53140 -9960 53185 -9840
rect 53305 -9960 53370 -9840
rect 30770 -10050 53370 -9960
rect 30770 -10170 30795 -10050
rect 30915 -10170 30970 -10050
rect 31090 -10170 31135 -10050
rect 31255 -10170 31300 -10050
rect 31420 -10170 31465 -10050
rect 31585 -10170 31640 -10050
rect 31760 -10170 31805 -10050
rect 31925 -10170 31970 -10050
rect 32090 -10170 32135 -10050
rect 32255 -10170 32310 -10050
rect 32430 -10170 32475 -10050
rect 32595 -10170 32640 -10050
rect 32760 -10170 32805 -10050
rect 32925 -10170 32980 -10050
rect 33100 -10170 33145 -10050
rect 33265 -10170 33310 -10050
rect 33430 -10170 33475 -10050
rect 33595 -10170 33650 -10050
rect 33770 -10170 33815 -10050
rect 33935 -10170 33980 -10050
rect 34100 -10170 34145 -10050
rect 34265 -10170 34320 -10050
rect 34440 -10170 34485 -10050
rect 34605 -10170 34650 -10050
rect 34770 -10170 34815 -10050
rect 34935 -10170 34990 -10050
rect 35110 -10170 35155 -10050
rect 35275 -10170 35320 -10050
rect 35440 -10170 35485 -10050
rect 35605 -10170 35660 -10050
rect 35780 -10170 35825 -10050
rect 35945 -10170 35990 -10050
rect 36110 -10170 36155 -10050
rect 36275 -10170 36485 -10050
rect 36605 -10170 36660 -10050
rect 36780 -10170 36825 -10050
rect 36945 -10170 36990 -10050
rect 37110 -10170 37155 -10050
rect 37275 -10170 37330 -10050
rect 37450 -10170 37495 -10050
rect 37615 -10170 37660 -10050
rect 37780 -10170 37825 -10050
rect 37945 -10170 38000 -10050
rect 38120 -10170 38165 -10050
rect 38285 -10170 38330 -10050
rect 38450 -10170 38495 -10050
rect 38615 -10170 38670 -10050
rect 38790 -10170 38835 -10050
rect 38955 -10170 39000 -10050
rect 39120 -10170 39165 -10050
rect 39285 -10170 39340 -10050
rect 39460 -10170 39505 -10050
rect 39625 -10170 39670 -10050
rect 39790 -10170 39835 -10050
rect 39955 -10170 40010 -10050
rect 40130 -10170 40175 -10050
rect 40295 -10170 40340 -10050
rect 40460 -10170 40505 -10050
rect 40625 -10170 40680 -10050
rect 40800 -10170 40845 -10050
rect 40965 -10170 41010 -10050
rect 41130 -10170 41175 -10050
rect 41295 -10170 41350 -10050
rect 41470 -10170 41515 -10050
rect 41635 -10170 41680 -10050
rect 41800 -10170 41845 -10050
rect 41965 -10170 42175 -10050
rect 42295 -10170 42350 -10050
rect 42470 -10170 42515 -10050
rect 42635 -10170 42680 -10050
rect 42800 -10170 42845 -10050
rect 42965 -10170 43020 -10050
rect 43140 -10170 43185 -10050
rect 43305 -10170 43350 -10050
rect 43470 -10170 43515 -10050
rect 43635 -10170 43690 -10050
rect 43810 -10170 43855 -10050
rect 43975 -10170 44020 -10050
rect 44140 -10170 44185 -10050
rect 44305 -10170 44360 -10050
rect 44480 -10170 44525 -10050
rect 44645 -10170 44690 -10050
rect 44810 -10170 44855 -10050
rect 44975 -10170 45030 -10050
rect 45150 -10170 45195 -10050
rect 45315 -10170 45360 -10050
rect 45480 -10170 45525 -10050
rect 45645 -10170 45700 -10050
rect 45820 -10170 45865 -10050
rect 45985 -10170 46030 -10050
rect 46150 -10170 46195 -10050
rect 46315 -10170 46370 -10050
rect 46490 -10170 46535 -10050
rect 46655 -10170 46700 -10050
rect 46820 -10170 46865 -10050
rect 46985 -10170 47040 -10050
rect 47160 -10170 47205 -10050
rect 47325 -10170 47370 -10050
rect 47490 -10170 47535 -10050
rect 47655 -10170 47865 -10050
rect 47985 -10170 48040 -10050
rect 48160 -10170 48205 -10050
rect 48325 -10170 48370 -10050
rect 48490 -10170 48535 -10050
rect 48655 -10170 48710 -10050
rect 48830 -10170 48875 -10050
rect 48995 -10170 49040 -10050
rect 49160 -10170 49205 -10050
rect 49325 -10170 49380 -10050
rect 49500 -10170 49545 -10050
rect 49665 -10170 49710 -10050
rect 49830 -10170 49875 -10050
rect 49995 -10170 50050 -10050
rect 50170 -10170 50215 -10050
rect 50335 -10170 50380 -10050
rect 50500 -10170 50545 -10050
rect 50665 -10170 50720 -10050
rect 50840 -10170 50885 -10050
rect 51005 -10170 51050 -10050
rect 51170 -10170 51215 -10050
rect 51335 -10170 51390 -10050
rect 51510 -10170 51555 -10050
rect 51675 -10170 51720 -10050
rect 51840 -10170 51885 -10050
rect 52005 -10170 52060 -10050
rect 52180 -10170 52225 -10050
rect 52345 -10170 52390 -10050
rect 52510 -10170 52555 -10050
rect 52675 -10170 52730 -10050
rect 52850 -10170 52895 -10050
rect 53015 -10170 53060 -10050
rect 53180 -10170 53225 -10050
rect 53345 -10170 53370 -10050
rect 30770 -10215 53370 -10170
rect 30770 -10335 30795 -10215
rect 30915 -10335 30970 -10215
rect 31090 -10335 31135 -10215
rect 31255 -10335 31300 -10215
rect 31420 -10335 31465 -10215
rect 31585 -10335 31640 -10215
rect 31760 -10335 31805 -10215
rect 31925 -10335 31970 -10215
rect 32090 -10335 32135 -10215
rect 32255 -10335 32310 -10215
rect 32430 -10335 32475 -10215
rect 32595 -10335 32640 -10215
rect 32760 -10335 32805 -10215
rect 32925 -10335 32980 -10215
rect 33100 -10335 33145 -10215
rect 33265 -10335 33310 -10215
rect 33430 -10335 33475 -10215
rect 33595 -10335 33650 -10215
rect 33770 -10335 33815 -10215
rect 33935 -10335 33980 -10215
rect 34100 -10335 34145 -10215
rect 34265 -10335 34320 -10215
rect 34440 -10335 34485 -10215
rect 34605 -10335 34650 -10215
rect 34770 -10335 34815 -10215
rect 34935 -10335 34990 -10215
rect 35110 -10335 35155 -10215
rect 35275 -10335 35320 -10215
rect 35440 -10335 35485 -10215
rect 35605 -10335 35660 -10215
rect 35780 -10335 35825 -10215
rect 35945 -10335 35990 -10215
rect 36110 -10335 36155 -10215
rect 36275 -10335 36485 -10215
rect 36605 -10335 36660 -10215
rect 36780 -10335 36825 -10215
rect 36945 -10335 36990 -10215
rect 37110 -10335 37155 -10215
rect 37275 -10335 37330 -10215
rect 37450 -10335 37495 -10215
rect 37615 -10335 37660 -10215
rect 37780 -10335 37825 -10215
rect 37945 -10335 38000 -10215
rect 38120 -10335 38165 -10215
rect 38285 -10335 38330 -10215
rect 38450 -10335 38495 -10215
rect 38615 -10335 38670 -10215
rect 38790 -10335 38835 -10215
rect 38955 -10335 39000 -10215
rect 39120 -10335 39165 -10215
rect 39285 -10335 39340 -10215
rect 39460 -10335 39505 -10215
rect 39625 -10335 39670 -10215
rect 39790 -10335 39835 -10215
rect 39955 -10335 40010 -10215
rect 40130 -10335 40175 -10215
rect 40295 -10335 40340 -10215
rect 40460 -10335 40505 -10215
rect 40625 -10335 40680 -10215
rect 40800 -10335 40845 -10215
rect 40965 -10335 41010 -10215
rect 41130 -10335 41175 -10215
rect 41295 -10335 41350 -10215
rect 41470 -10335 41515 -10215
rect 41635 -10335 41680 -10215
rect 41800 -10335 41845 -10215
rect 41965 -10335 42175 -10215
rect 42295 -10335 42350 -10215
rect 42470 -10335 42515 -10215
rect 42635 -10335 42680 -10215
rect 42800 -10335 42845 -10215
rect 42965 -10335 43020 -10215
rect 43140 -10335 43185 -10215
rect 43305 -10335 43350 -10215
rect 43470 -10335 43515 -10215
rect 43635 -10335 43690 -10215
rect 43810 -10335 43855 -10215
rect 43975 -10335 44020 -10215
rect 44140 -10335 44185 -10215
rect 44305 -10335 44360 -10215
rect 44480 -10335 44525 -10215
rect 44645 -10335 44690 -10215
rect 44810 -10335 44855 -10215
rect 44975 -10335 45030 -10215
rect 45150 -10335 45195 -10215
rect 45315 -10335 45360 -10215
rect 45480 -10335 45525 -10215
rect 45645 -10335 45700 -10215
rect 45820 -10335 45865 -10215
rect 45985 -10335 46030 -10215
rect 46150 -10335 46195 -10215
rect 46315 -10335 46370 -10215
rect 46490 -10335 46535 -10215
rect 46655 -10335 46700 -10215
rect 46820 -10335 46865 -10215
rect 46985 -10335 47040 -10215
rect 47160 -10335 47205 -10215
rect 47325 -10335 47370 -10215
rect 47490 -10335 47535 -10215
rect 47655 -10335 47865 -10215
rect 47985 -10335 48040 -10215
rect 48160 -10335 48205 -10215
rect 48325 -10335 48370 -10215
rect 48490 -10335 48535 -10215
rect 48655 -10335 48710 -10215
rect 48830 -10335 48875 -10215
rect 48995 -10335 49040 -10215
rect 49160 -10335 49205 -10215
rect 49325 -10335 49380 -10215
rect 49500 -10335 49545 -10215
rect 49665 -10335 49710 -10215
rect 49830 -10335 49875 -10215
rect 49995 -10335 50050 -10215
rect 50170 -10335 50215 -10215
rect 50335 -10335 50380 -10215
rect 50500 -10335 50545 -10215
rect 50665 -10335 50720 -10215
rect 50840 -10335 50885 -10215
rect 51005 -10335 51050 -10215
rect 51170 -10335 51215 -10215
rect 51335 -10335 51390 -10215
rect 51510 -10335 51555 -10215
rect 51675 -10335 51720 -10215
rect 51840 -10335 51885 -10215
rect 52005 -10335 52060 -10215
rect 52180 -10335 52225 -10215
rect 52345 -10335 52390 -10215
rect 52510 -10335 52555 -10215
rect 52675 -10335 52730 -10215
rect 52850 -10335 52895 -10215
rect 53015 -10335 53060 -10215
rect 53180 -10335 53225 -10215
rect 53345 -10335 53370 -10215
rect 30770 -10380 53370 -10335
rect 30770 -10459 30795 -10380
rect 30365 -10500 30795 -10459
rect 30915 -10500 30970 -10380
rect 31090 -10500 31135 -10380
rect 31255 -10500 31300 -10380
rect 31420 -10500 31465 -10380
rect 31585 -10500 31640 -10380
rect 31760 -10500 31805 -10380
rect 31925 -10500 31970 -10380
rect 32090 -10500 32135 -10380
rect 32255 -10500 32310 -10380
rect 32430 -10500 32475 -10380
rect 32595 -10500 32640 -10380
rect 32760 -10500 32805 -10380
rect 32925 -10500 32980 -10380
rect 33100 -10500 33145 -10380
rect 33265 -10500 33310 -10380
rect 33430 -10500 33475 -10380
rect 33595 -10500 33650 -10380
rect 33770 -10500 33815 -10380
rect 33935 -10500 33980 -10380
rect 34100 -10500 34145 -10380
rect 34265 -10500 34320 -10380
rect 34440 -10500 34485 -10380
rect 34605 -10500 34650 -10380
rect 34770 -10500 34815 -10380
rect 34935 -10500 34990 -10380
rect 35110 -10500 35155 -10380
rect 35275 -10500 35320 -10380
rect 35440 -10500 35485 -10380
rect 35605 -10500 35660 -10380
rect 35780 -10500 35825 -10380
rect 35945 -10500 35990 -10380
rect 36110 -10500 36155 -10380
rect 36275 -10500 36485 -10380
rect 36605 -10500 36660 -10380
rect 36780 -10500 36825 -10380
rect 36945 -10500 36990 -10380
rect 37110 -10500 37155 -10380
rect 37275 -10500 37330 -10380
rect 37450 -10500 37495 -10380
rect 37615 -10500 37660 -10380
rect 37780 -10500 37825 -10380
rect 37945 -10500 38000 -10380
rect 38120 -10500 38165 -10380
rect 38285 -10500 38330 -10380
rect 38450 -10500 38495 -10380
rect 38615 -10500 38670 -10380
rect 38790 -10500 38835 -10380
rect 38955 -10500 39000 -10380
rect 39120 -10500 39165 -10380
rect 39285 -10500 39340 -10380
rect 39460 -10500 39505 -10380
rect 39625 -10500 39670 -10380
rect 39790 -10500 39835 -10380
rect 39955 -10500 40010 -10380
rect 40130 -10500 40175 -10380
rect 40295 -10500 40340 -10380
rect 40460 -10500 40505 -10380
rect 40625 -10500 40680 -10380
rect 40800 -10500 40845 -10380
rect 40965 -10500 41010 -10380
rect 41130 -10500 41175 -10380
rect 41295 -10500 41350 -10380
rect 41470 -10500 41515 -10380
rect 41635 -10500 41680 -10380
rect 41800 -10500 41845 -10380
rect 41965 -10500 42175 -10380
rect 42295 -10500 42350 -10380
rect 42470 -10500 42515 -10380
rect 42635 -10500 42680 -10380
rect 42800 -10500 42845 -10380
rect 42965 -10500 43020 -10380
rect 43140 -10500 43185 -10380
rect 43305 -10500 43350 -10380
rect 43470 -10500 43515 -10380
rect 43635 -10500 43690 -10380
rect 43810 -10500 43855 -10380
rect 43975 -10500 44020 -10380
rect 44140 -10500 44185 -10380
rect 44305 -10500 44360 -10380
rect 44480 -10500 44525 -10380
rect 44645 -10500 44690 -10380
rect 44810 -10500 44855 -10380
rect 44975 -10500 45030 -10380
rect 45150 -10500 45195 -10380
rect 45315 -10500 45360 -10380
rect 45480 -10500 45525 -10380
rect 45645 -10500 45700 -10380
rect 45820 -10500 45865 -10380
rect 45985 -10500 46030 -10380
rect 46150 -10500 46195 -10380
rect 46315 -10500 46370 -10380
rect 46490 -10500 46535 -10380
rect 46655 -10500 46700 -10380
rect 46820 -10500 46865 -10380
rect 46985 -10500 47040 -10380
rect 47160 -10500 47205 -10380
rect 47325 -10500 47370 -10380
rect 47490 -10500 47535 -10380
rect 47655 -10500 47865 -10380
rect 47985 -10500 48040 -10380
rect 48160 -10500 48205 -10380
rect 48325 -10500 48370 -10380
rect 48490 -10500 48535 -10380
rect 48655 -10500 48710 -10380
rect 48830 -10500 48875 -10380
rect 48995 -10500 49040 -10380
rect 49160 -10500 49205 -10380
rect 49325 -10500 49380 -10380
rect 49500 -10500 49545 -10380
rect 49665 -10500 49710 -10380
rect 49830 -10500 49875 -10380
rect 49995 -10500 50050 -10380
rect 50170 -10500 50215 -10380
rect 50335 -10500 50380 -10380
rect 50500 -10500 50545 -10380
rect 50665 -10500 50720 -10380
rect 50840 -10500 50885 -10380
rect 51005 -10500 51050 -10380
rect 51170 -10500 51215 -10380
rect 51335 -10500 51390 -10380
rect 51510 -10500 51555 -10380
rect 51675 -10500 51720 -10380
rect 51840 -10500 51885 -10380
rect 52005 -10500 52060 -10380
rect 52180 -10500 52225 -10380
rect 52345 -10500 52390 -10380
rect 52510 -10500 52555 -10380
rect 52675 -10500 52730 -10380
rect 52850 -10500 52895 -10380
rect 53015 -10500 53060 -10380
rect 53180 -10500 53225 -10380
rect 53345 -10500 53370 -10380
rect 30365 -10545 53370 -10500
rect 30365 -10665 30795 -10545
rect 30915 -10665 30970 -10545
rect 31090 -10665 31135 -10545
rect 31255 -10665 31300 -10545
rect 31420 -10665 31465 -10545
rect 31585 -10665 31640 -10545
rect 31760 -10665 31805 -10545
rect 31925 -10665 31970 -10545
rect 32090 -10665 32135 -10545
rect 32255 -10665 32310 -10545
rect 32430 -10665 32475 -10545
rect 32595 -10665 32640 -10545
rect 32760 -10665 32805 -10545
rect 32925 -10665 32980 -10545
rect 33100 -10665 33145 -10545
rect 33265 -10665 33310 -10545
rect 33430 -10665 33475 -10545
rect 33595 -10665 33650 -10545
rect 33770 -10665 33815 -10545
rect 33935 -10665 33980 -10545
rect 34100 -10665 34145 -10545
rect 34265 -10665 34320 -10545
rect 34440 -10665 34485 -10545
rect 34605 -10665 34650 -10545
rect 34770 -10665 34815 -10545
rect 34935 -10665 34990 -10545
rect 35110 -10665 35155 -10545
rect 35275 -10665 35320 -10545
rect 35440 -10665 35485 -10545
rect 35605 -10665 35660 -10545
rect 35780 -10665 35825 -10545
rect 35945 -10665 35990 -10545
rect 36110 -10665 36155 -10545
rect 36275 -10665 36485 -10545
rect 36605 -10665 36660 -10545
rect 36780 -10665 36825 -10545
rect 36945 -10665 36990 -10545
rect 37110 -10665 37155 -10545
rect 37275 -10665 37330 -10545
rect 37450 -10665 37495 -10545
rect 37615 -10665 37660 -10545
rect 37780 -10665 37825 -10545
rect 37945 -10665 38000 -10545
rect 38120 -10665 38165 -10545
rect 38285 -10665 38330 -10545
rect 38450 -10665 38495 -10545
rect 38615 -10665 38670 -10545
rect 38790 -10665 38835 -10545
rect 38955 -10665 39000 -10545
rect 39120 -10665 39165 -10545
rect 39285 -10665 39340 -10545
rect 39460 -10665 39505 -10545
rect 39625 -10665 39670 -10545
rect 39790 -10665 39835 -10545
rect 39955 -10665 40010 -10545
rect 40130 -10665 40175 -10545
rect 40295 -10665 40340 -10545
rect 40460 -10665 40505 -10545
rect 40625 -10665 40680 -10545
rect 40800 -10665 40845 -10545
rect 40965 -10665 41010 -10545
rect 41130 -10665 41175 -10545
rect 41295 -10665 41350 -10545
rect 41470 -10665 41515 -10545
rect 41635 -10665 41680 -10545
rect 41800 -10665 41845 -10545
rect 41965 -10665 42175 -10545
rect 42295 -10665 42350 -10545
rect 42470 -10665 42515 -10545
rect 42635 -10665 42680 -10545
rect 42800 -10665 42845 -10545
rect 42965 -10665 43020 -10545
rect 43140 -10665 43185 -10545
rect 43305 -10665 43350 -10545
rect 43470 -10665 43515 -10545
rect 43635 -10665 43690 -10545
rect 43810 -10665 43855 -10545
rect 43975 -10665 44020 -10545
rect 44140 -10665 44185 -10545
rect 44305 -10665 44360 -10545
rect 44480 -10665 44525 -10545
rect 44645 -10665 44690 -10545
rect 44810 -10665 44855 -10545
rect 44975 -10665 45030 -10545
rect 45150 -10665 45195 -10545
rect 45315 -10665 45360 -10545
rect 45480 -10665 45525 -10545
rect 45645 -10665 45700 -10545
rect 45820 -10665 45865 -10545
rect 45985 -10665 46030 -10545
rect 46150 -10665 46195 -10545
rect 46315 -10665 46370 -10545
rect 46490 -10665 46535 -10545
rect 46655 -10665 46700 -10545
rect 46820 -10665 46865 -10545
rect 46985 -10665 47040 -10545
rect 47160 -10665 47205 -10545
rect 47325 -10665 47370 -10545
rect 47490 -10665 47535 -10545
rect 47655 -10665 47865 -10545
rect 47985 -10665 48040 -10545
rect 48160 -10665 48205 -10545
rect 48325 -10665 48370 -10545
rect 48490 -10665 48535 -10545
rect 48655 -10665 48710 -10545
rect 48830 -10665 48875 -10545
rect 48995 -10665 49040 -10545
rect 49160 -10665 49205 -10545
rect 49325 -10665 49380 -10545
rect 49500 -10665 49545 -10545
rect 49665 -10665 49710 -10545
rect 49830 -10665 49875 -10545
rect 49995 -10665 50050 -10545
rect 50170 -10665 50215 -10545
rect 50335 -10665 50380 -10545
rect 50500 -10665 50545 -10545
rect 50665 -10665 50720 -10545
rect 50840 -10665 50885 -10545
rect 51005 -10665 51050 -10545
rect 51170 -10665 51215 -10545
rect 51335 -10665 51390 -10545
rect 51510 -10665 51555 -10545
rect 51675 -10665 51720 -10545
rect 51840 -10665 51885 -10545
rect 52005 -10665 52060 -10545
rect 52180 -10665 52225 -10545
rect 52345 -10665 52390 -10545
rect 52510 -10665 52555 -10545
rect 52675 -10665 52730 -10545
rect 52850 -10665 52895 -10545
rect 53015 -10665 53060 -10545
rect 53180 -10665 53225 -10545
rect 53345 -10665 53370 -10545
rect 30365 -10720 53370 -10665
rect 30365 -10840 30795 -10720
rect 30915 -10840 30970 -10720
rect 31090 -10840 31135 -10720
rect 31255 -10840 31300 -10720
rect 31420 -10840 31465 -10720
rect 31585 -10840 31640 -10720
rect 31760 -10840 31805 -10720
rect 31925 -10840 31970 -10720
rect 32090 -10840 32135 -10720
rect 32255 -10840 32310 -10720
rect 32430 -10840 32475 -10720
rect 32595 -10840 32640 -10720
rect 32760 -10840 32805 -10720
rect 32925 -10840 32980 -10720
rect 33100 -10840 33145 -10720
rect 33265 -10840 33310 -10720
rect 33430 -10840 33475 -10720
rect 33595 -10840 33650 -10720
rect 33770 -10840 33815 -10720
rect 33935 -10840 33980 -10720
rect 34100 -10840 34145 -10720
rect 34265 -10840 34320 -10720
rect 34440 -10840 34485 -10720
rect 34605 -10840 34650 -10720
rect 34770 -10840 34815 -10720
rect 34935 -10840 34990 -10720
rect 35110 -10840 35155 -10720
rect 35275 -10840 35320 -10720
rect 35440 -10840 35485 -10720
rect 35605 -10840 35660 -10720
rect 35780 -10840 35825 -10720
rect 35945 -10840 35990 -10720
rect 36110 -10840 36155 -10720
rect 36275 -10840 36485 -10720
rect 36605 -10840 36660 -10720
rect 36780 -10840 36825 -10720
rect 36945 -10840 36990 -10720
rect 37110 -10840 37155 -10720
rect 37275 -10840 37330 -10720
rect 37450 -10840 37495 -10720
rect 37615 -10840 37660 -10720
rect 37780 -10840 37825 -10720
rect 37945 -10840 38000 -10720
rect 38120 -10840 38165 -10720
rect 38285 -10840 38330 -10720
rect 38450 -10840 38495 -10720
rect 38615 -10840 38670 -10720
rect 38790 -10840 38835 -10720
rect 38955 -10840 39000 -10720
rect 39120 -10840 39165 -10720
rect 39285 -10840 39340 -10720
rect 39460 -10840 39505 -10720
rect 39625 -10840 39670 -10720
rect 39790 -10840 39835 -10720
rect 39955 -10840 40010 -10720
rect 40130 -10840 40175 -10720
rect 40295 -10840 40340 -10720
rect 40460 -10840 40505 -10720
rect 40625 -10840 40680 -10720
rect 40800 -10840 40845 -10720
rect 40965 -10840 41010 -10720
rect 41130 -10840 41175 -10720
rect 41295 -10840 41350 -10720
rect 41470 -10840 41515 -10720
rect 41635 -10840 41680 -10720
rect 41800 -10840 41845 -10720
rect 41965 -10840 42175 -10720
rect 42295 -10840 42350 -10720
rect 42470 -10840 42515 -10720
rect 42635 -10840 42680 -10720
rect 42800 -10840 42845 -10720
rect 42965 -10840 43020 -10720
rect 43140 -10840 43185 -10720
rect 43305 -10840 43350 -10720
rect 43470 -10840 43515 -10720
rect 43635 -10840 43690 -10720
rect 43810 -10840 43855 -10720
rect 43975 -10840 44020 -10720
rect 44140 -10840 44185 -10720
rect 44305 -10840 44360 -10720
rect 44480 -10840 44525 -10720
rect 44645 -10840 44690 -10720
rect 44810 -10840 44855 -10720
rect 44975 -10840 45030 -10720
rect 45150 -10840 45195 -10720
rect 45315 -10840 45360 -10720
rect 45480 -10840 45525 -10720
rect 45645 -10840 45700 -10720
rect 45820 -10840 45865 -10720
rect 45985 -10840 46030 -10720
rect 46150 -10840 46195 -10720
rect 46315 -10840 46370 -10720
rect 46490 -10840 46535 -10720
rect 46655 -10840 46700 -10720
rect 46820 -10840 46865 -10720
rect 46985 -10840 47040 -10720
rect 47160 -10840 47205 -10720
rect 47325 -10840 47370 -10720
rect 47490 -10840 47535 -10720
rect 47655 -10840 47865 -10720
rect 47985 -10840 48040 -10720
rect 48160 -10840 48205 -10720
rect 48325 -10840 48370 -10720
rect 48490 -10840 48535 -10720
rect 48655 -10840 48710 -10720
rect 48830 -10840 48875 -10720
rect 48995 -10840 49040 -10720
rect 49160 -10840 49205 -10720
rect 49325 -10840 49380 -10720
rect 49500 -10840 49545 -10720
rect 49665 -10840 49710 -10720
rect 49830 -10840 49875 -10720
rect 49995 -10840 50050 -10720
rect 50170 -10840 50215 -10720
rect 50335 -10840 50380 -10720
rect 50500 -10840 50545 -10720
rect 50665 -10840 50720 -10720
rect 50840 -10840 50885 -10720
rect 51005 -10840 51050 -10720
rect 51170 -10840 51215 -10720
rect 51335 -10840 51390 -10720
rect 51510 -10840 51555 -10720
rect 51675 -10840 51720 -10720
rect 51840 -10840 51885 -10720
rect 52005 -10840 52060 -10720
rect 52180 -10840 52225 -10720
rect 52345 -10840 52390 -10720
rect 52510 -10840 52555 -10720
rect 52675 -10840 52730 -10720
rect 52850 -10840 52895 -10720
rect 53015 -10840 53060 -10720
rect 53180 -10840 53225 -10720
rect 53345 -10840 53370 -10720
rect 30365 -10844 53370 -10840
rect 30770 -10885 53370 -10844
rect 30770 -11005 30795 -10885
rect 30915 -11005 30970 -10885
rect 31090 -11005 31135 -10885
rect 31255 -11005 31300 -10885
rect 31420 -11005 31465 -10885
rect 31585 -11005 31640 -10885
rect 31760 -11005 31805 -10885
rect 31925 -11005 31970 -10885
rect 32090 -11005 32135 -10885
rect 32255 -11005 32310 -10885
rect 32430 -11005 32475 -10885
rect 32595 -11005 32640 -10885
rect 32760 -11005 32805 -10885
rect 32925 -11005 32980 -10885
rect 33100 -11005 33145 -10885
rect 33265 -11005 33310 -10885
rect 33430 -11005 33475 -10885
rect 33595 -11005 33650 -10885
rect 33770 -11005 33815 -10885
rect 33935 -11005 33980 -10885
rect 34100 -11005 34145 -10885
rect 34265 -11005 34320 -10885
rect 34440 -11005 34485 -10885
rect 34605 -11005 34650 -10885
rect 34770 -11005 34815 -10885
rect 34935 -11005 34990 -10885
rect 35110 -11005 35155 -10885
rect 35275 -11005 35320 -10885
rect 35440 -11005 35485 -10885
rect 35605 -11005 35660 -10885
rect 35780 -11005 35825 -10885
rect 35945 -11005 35990 -10885
rect 36110 -11005 36155 -10885
rect 36275 -11005 36485 -10885
rect 36605 -11005 36660 -10885
rect 36780 -11005 36825 -10885
rect 36945 -11005 36990 -10885
rect 37110 -11005 37155 -10885
rect 37275 -11005 37330 -10885
rect 37450 -11005 37495 -10885
rect 37615 -11005 37660 -10885
rect 37780 -11005 37825 -10885
rect 37945 -11005 38000 -10885
rect 38120 -11005 38165 -10885
rect 38285 -11005 38330 -10885
rect 38450 -11005 38495 -10885
rect 38615 -11005 38670 -10885
rect 38790 -11005 38835 -10885
rect 38955 -11005 39000 -10885
rect 39120 -11005 39165 -10885
rect 39285 -11005 39340 -10885
rect 39460 -11005 39505 -10885
rect 39625 -11005 39670 -10885
rect 39790 -11005 39835 -10885
rect 39955 -11005 40010 -10885
rect 40130 -11005 40175 -10885
rect 40295 -11005 40340 -10885
rect 40460 -11005 40505 -10885
rect 40625 -11005 40680 -10885
rect 40800 -11005 40845 -10885
rect 40965 -11005 41010 -10885
rect 41130 -11005 41175 -10885
rect 41295 -11005 41350 -10885
rect 41470 -11005 41515 -10885
rect 41635 -11005 41680 -10885
rect 41800 -11005 41845 -10885
rect 41965 -11005 42175 -10885
rect 42295 -11005 42350 -10885
rect 42470 -11005 42515 -10885
rect 42635 -11005 42680 -10885
rect 42800 -11005 42845 -10885
rect 42965 -11005 43020 -10885
rect 43140 -11005 43185 -10885
rect 43305 -11005 43350 -10885
rect 43470 -11005 43515 -10885
rect 43635 -11005 43690 -10885
rect 43810 -11005 43855 -10885
rect 43975 -11005 44020 -10885
rect 44140 -11005 44185 -10885
rect 44305 -11005 44360 -10885
rect 44480 -11005 44525 -10885
rect 44645 -11005 44690 -10885
rect 44810 -11005 44855 -10885
rect 44975 -11005 45030 -10885
rect 45150 -11005 45195 -10885
rect 45315 -11005 45360 -10885
rect 45480 -11005 45525 -10885
rect 45645 -11005 45700 -10885
rect 45820 -11005 45865 -10885
rect 45985 -11005 46030 -10885
rect 46150 -11005 46195 -10885
rect 46315 -11005 46370 -10885
rect 46490 -11005 46535 -10885
rect 46655 -11005 46700 -10885
rect 46820 -11005 46865 -10885
rect 46985 -11005 47040 -10885
rect 47160 -11005 47205 -10885
rect 47325 -11005 47370 -10885
rect 47490 -11005 47535 -10885
rect 47655 -11005 47865 -10885
rect 47985 -11005 48040 -10885
rect 48160 -11005 48205 -10885
rect 48325 -11005 48370 -10885
rect 48490 -11005 48535 -10885
rect 48655 -11005 48710 -10885
rect 48830 -11005 48875 -10885
rect 48995 -11005 49040 -10885
rect 49160 -11005 49205 -10885
rect 49325 -11005 49380 -10885
rect 49500 -11005 49545 -10885
rect 49665 -11005 49710 -10885
rect 49830 -11005 49875 -10885
rect 49995 -11005 50050 -10885
rect 50170 -11005 50215 -10885
rect 50335 -11005 50380 -10885
rect 50500 -11005 50545 -10885
rect 50665 -11005 50720 -10885
rect 50840 -11005 50885 -10885
rect 51005 -11005 51050 -10885
rect 51170 -11005 51215 -10885
rect 51335 -11005 51390 -10885
rect 51510 -11005 51555 -10885
rect 51675 -11005 51720 -10885
rect 51840 -11005 51885 -10885
rect 52005 -11005 52060 -10885
rect 52180 -11005 52225 -10885
rect 52345 -11005 52390 -10885
rect 52510 -11005 52555 -10885
rect 52675 -11005 52730 -10885
rect 52850 -11005 52895 -10885
rect 53015 -11005 53060 -10885
rect 53180 -11005 53225 -10885
rect 53345 -11005 53370 -10885
rect 30770 -11050 53370 -11005
rect 30770 -11170 30795 -11050
rect 30915 -11170 30970 -11050
rect 31090 -11170 31135 -11050
rect 31255 -11170 31300 -11050
rect 31420 -11170 31465 -11050
rect 31585 -11170 31640 -11050
rect 31760 -11170 31805 -11050
rect 31925 -11170 31970 -11050
rect 32090 -11170 32135 -11050
rect 32255 -11170 32310 -11050
rect 32430 -11170 32475 -11050
rect 32595 -11170 32640 -11050
rect 32760 -11170 32805 -11050
rect 32925 -11170 32980 -11050
rect 33100 -11170 33145 -11050
rect 33265 -11170 33310 -11050
rect 33430 -11170 33475 -11050
rect 33595 -11170 33650 -11050
rect 33770 -11170 33815 -11050
rect 33935 -11170 33980 -11050
rect 34100 -11170 34145 -11050
rect 34265 -11170 34320 -11050
rect 34440 -11170 34485 -11050
rect 34605 -11170 34650 -11050
rect 34770 -11170 34815 -11050
rect 34935 -11170 34990 -11050
rect 35110 -11170 35155 -11050
rect 35275 -11170 35320 -11050
rect 35440 -11170 35485 -11050
rect 35605 -11170 35660 -11050
rect 35780 -11170 35825 -11050
rect 35945 -11170 35990 -11050
rect 36110 -11170 36155 -11050
rect 36275 -11170 36485 -11050
rect 36605 -11170 36660 -11050
rect 36780 -11170 36825 -11050
rect 36945 -11170 36990 -11050
rect 37110 -11170 37155 -11050
rect 37275 -11170 37330 -11050
rect 37450 -11170 37495 -11050
rect 37615 -11170 37660 -11050
rect 37780 -11170 37825 -11050
rect 37945 -11170 38000 -11050
rect 38120 -11170 38165 -11050
rect 38285 -11170 38330 -11050
rect 38450 -11170 38495 -11050
rect 38615 -11170 38670 -11050
rect 38790 -11170 38835 -11050
rect 38955 -11170 39000 -11050
rect 39120 -11170 39165 -11050
rect 39285 -11170 39340 -11050
rect 39460 -11170 39505 -11050
rect 39625 -11170 39670 -11050
rect 39790 -11170 39835 -11050
rect 39955 -11170 40010 -11050
rect 40130 -11170 40175 -11050
rect 40295 -11170 40340 -11050
rect 40460 -11170 40505 -11050
rect 40625 -11170 40680 -11050
rect 40800 -11170 40845 -11050
rect 40965 -11170 41010 -11050
rect 41130 -11170 41175 -11050
rect 41295 -11170 41350 -11050
rect 41470 -11170 41515 -11050
rect 41635 -11170 41680 -11050
rect 41800 -11170 41845 -11050
rect 41965 -11170 42175 -11050
rect 42295 -11170 42350 -11050
rect 42470 -11170 42515 -11050
rect 42635 -11170 42680 -11050
rect 42800 -11170 42845 -11050
rect 42965 -11170 43020 -11050
rect 43140 -11170 43185 -11050
rect 43305 -11170 43350 -11050
rect 43470 -11170 43515 -11050
rect 43635 -11170 43690 -11050
rect 43810 -11170 43855 -11050
rect 43975 -11170 44020 -11050
rect 44140 -11170 44185 -11050
rect 44305 -11170 44360 -11050
rect 44480 -11170 44525 -11050
rect 44645 -11170 44690 -11050
rect 44810 -11170 44855 -11050
rect 44975 -11170 45030 -11050
rect 45150 -11170 45195 -11050
rect 45315 -11170 45360 -11050
rect 45480 -11170 45525 -11050
rect 45645 -11170 45700 -11050
rect 45820 -11170 45865 -11050
rect 45985 -11170 46030 -11050
rect 46150 -11170 46195 -11050
rect 46315 -11170 46370 -11050
rect 46490 -11170 46535 -11050
rect 46655 -11170 46700 -11050
rect 46820 -11170 46865 -11050
rect 46985 -11170 47040 -11050
rect 47160 -11170 47205 -11050
rect 47325 -11170 47370 -11050
rect 47490 -11170 47535 -11050
rect 47655 -11170 47865 -11050
rect 47985 -11170 48040 -11050
rect 48160 -11170 48205 -11050
rect 48325 -11170 48370 -11050
rect 48490 -11170 48535 -11050
rect 48655 -11170 48710 -11050
rect 48830 -11170 48875 -11050
rect 48995 -11170 49040 -11050
rect 49160 -11170 49205 -11050
rect 49325 -11170 49380 -11050
rect 49500 -11170 49545 -11050
rect 49665 -11170 49710 -11050
rect 49830 -11170 49875 -11050
rect 49995 -11170 50050 -11050
rect 50170 -11170 50215 -11050
rect 50335 -11170 50380 -11050
rect 50500 -11170 50545 -11050
rect 50665 -11170 50720 -11050
rect 50840 -11170 50885 -11050
rect 51005 -11170 51050 -11050
rect 51170 -11170 51215 -11050
rect 51335 -11170 51390 -11050
rect 51510 -11170 51555 -11050
rect 51675 -11170 51720 -11050
rect 51840 -11170 51885 -11050
rect 52005 -11170 52060 -11050
rect 52180 -11170 52225 -11050
rect 52345 -11170 52390 -11050
rect 52510 -11170 52555 -11050
rect 52675 -11170 52730 -11050
rect 52850 -11170 52895 -11050
rect 53015 -11170 53060 -11050
rect 53180 -11170 53225 -11050
rect 53345 -11170 53370 -11050
rect 30770 -11215 53370 -11170
rect 30770 -11335 30795 -11215
rect 30915 -11335 30970 -11215
rect 31090 -11335 31135 -11215
rect 31255 -11335 31300 -11215
rect 31420 -11335 31465 -11215
rect 31585 -11335 31640 -11215
rect 31760 -11335 31805 -11215
rect 31925 -11335 31970 -11215
rect 32090 -11335 32135 -11215
rect 32255 -11335 32310 -11215
rect 32430 -11335 32475 -11215
rect 32595 -11335 32640 -11215
rect 32760 -11335 32805 -11215
rect 32925 -11335 32980 -11215
rect 33100 -11335 33145 -11215
rect 33265 -11335 33310 -11215
rect 33430 -11335 33475 -11215
rect 33595 -11335 33650 -11215
rect 33770 -11335 33815 -11215
rect 33935 -11335 33980 -11215
rect 34100 -11335 34145 -11215
rect 34265 -11335 34320 -11215
rect 34440 -11335 34485 -11215
rect 34605 -11335 34650 -11215
rect 34770 -11335 34815 -11215
rect 34935 -11335 34990 -11215
rect 35110 -11335 35155 -11215
rect 35275 -11335 35320 -11215
rect 35440 -11335 35485 -11215
rect 35605 -11335 35660 -11215
rect 35780 -11335 35825 -11215
rect 35945 -11335 35990 -11215
rect 36110 -11335 36155 -11215
rect 36275 -11335 36485 -11215
rect 36605 -11335 36660 -11215
rect 36780 -11335 36825 -11215
rect 36945 -11335 36990 -11215
rect 37110 -11335 37155 -11215
rect 37275 -11335 37330 -11215
rect 37450 -11335 37495 -11215
rect 37615 -11335 37660 -11215
rect 37780 -11335 37825 -11215
rect 37945 -11335 38000 -11215
rect 38120 -11335 38165 -11215
rect 38285 -11335 38330 -11215
rect 38450 -11335 38495 -11215
rect 38615 -11335 38670 -11215
rect 38790 -11335 38835 -11215
rect 38955 -11335 39000 -11215
rect 39120 -11335 39165 -11215
rect 39285 -11335 39340 -11215
rect 39460 -11335 39505 -11215
rect 39625 -11335 39670 -11215
rect 39790 -11335 39835 -11215
rect 39955 -11335 40010 -11215
rect 40130 -11335 40175 -11215
rect 40295 -11335 40340 -11215
rect 40460 -11335 40505 -11215
rect 40625 -11335 40680 -11215
rect 40800 -11335 40845 -11215
rect 40965 -11335 41010 -11215
rect 41130 -11335 41175 -11215
rect 41295 -11335 41350 -11215
rect 41470 -11335 41515 -11215
rect 41635 -11335 41680 -11215
rect 41800 -11335 41845 -11215
rect 41965 -11335 42175 -11215
rect 42295 -11335 42350 -11215
rect 42470 -11335 42515 -11215
rect 42635 -11335 42680 -11215
rect 42800 -11335 42845 -11215
rect 42965 -11335 43020 -11215
rect 43140 -11335 43185 -11215
rect 43305 -11335 43350 -11215
rect 43470 -11335 43515 -11215
rect 43635 -11335 43690 -11215
rect 43810 -11335 43855 -11215
rect 43975 -11335 44020 -11215
rect 44140 -11335 44185 -11215
rect 44305 -11335 44360 -11215
rect 44480 -11335 44525 -11215
rect 44645 -11335 44690 -11215
rect 44810 -11335 44855 -11215
rect 44975 -11335 45030 -11215
rect 45150 -11335 45195 -11215
rect 45315 -11335 45360 -11215
rect 45480 -11335 45525 -11215
rect 45645 -11335 45700 -11215
rect 45820 -11335 45865 -11215
rect 45985 -11335 46030 -11215
rect 46150 -11335 46195 -11215
rect 46315 -11335 46370 -11215
rect 46490 -11335 46535 -11215
rect 46655 -11335 46700 -11215
rect 46820 -11335 46865 -11215
rect 46985 -11335 47040 -11215
rect 47160 -11335 47205 -11215
rect 47325 -11335 47370 -11215
rect 47490 -11335 47535 -11215
rect 47655 -11335 47865 -11215
rect 47985 -11335 48040 -11215
rect 48160 -11335 48205 -11215
rect 48325 -11335 48370 -11215
rect 48490 -11335 48535 -11215
rect 48655 -11335 48710 -11215
rect 48830 -11335 48875 -11215
rect 48995 -11335 49040 -11215
rect 49160 -11335 49205 -11215
rect 49325 -11335 49380 -11215
rect 49500 -11335 49545 -11215
rect 49665 -11335 49710 -11215
rect 49830 -11335 49875 -11215
rect 49995 -11335 50050 -11215
rect 50170 -11335 50215 -11215
rect 50335 -11335 50380 -11215
rect 50500 -11335 50545 -11215
rect 50665 -11335 50720 -11215
rect 50840 -11335 50885 -11215
rect 51005 -11335 51050 -11215
rect 51170 -11335 51215 -11215
rect 51335 -11335 51390 -11215
rect 51510 -11335 51555 -11215
rect 51675 -11335 51720 -11215
rect 51840 -11335 51885 -11215
rect 52005 -11335 52060 -11215
rect 52180 -11335 52225 -11215
rect 52345 -11335 52390 -11215
rect 52510 -11335 52555 -11215
rect 52675 -11335 52730 -11215
rect 52850 -11335 52895 -11215
rect 53015 -11335 53060 -11215
rect 53180 -11335 53225 -11215
rect 53345 -11335 53370 -11215
rect 30770 -11390 53370 -11335
rect 30770 -11510 30795 -11390
rect 30915 -11510 30970 -11390
rect 31090 -11510 31135 -11390
rect 31255 -11510 31300 -11390
rect 31420 -11510 31465 -11390
rect 31585 -11510 31640 -11390
rect 31760 -11510 31805 -11390
rect 31925 -11510 31970 -11390
rect 32090 -11510 32135 -11390
rect 32255 -11510 32310 -11390
rect 32430 -11510 32475 -11390
rect 32595 -11510 32640 -11390
rect 32760 -11510 32805 -11390
rect 32925 -11510 32980 -11390
rect 33100 -11510 33145 -11390
rect 33265 -11510 33310 -11390
rect 33430 -11510 33475 -11390
rect 33595 -11510 33650 -11390
rect 33770 -11510 33815 -11390
rect 33935 -11510 33980 -11390
rect 34100 -11510 34145 -11390
rect 34265 -11510 34320 -11390
rect 34440 -11510 34485 -11390
rect 34605 -11510 34650 -11390
rect 34770 -11510 34815 -11390
rect 34935 -11510 34990 -11390
rect 35110 -11510 35155 -11390
rect 35275 -11510 35320 -11390
rect 35440 -11510 35485 -11390
rect 35605 -11510 35660 -11390
rect 35780 -11510 35825 -11390
rect 35945 -11510 35990 -11390
rect 36110 -11510 36155 -11390
rect 36275 -11510 36485 -11390
rect 36605 -11510 36660 -11390
rect 36780 -11510 36825 -11390
rect 36945 -11510 36990 -11390
rect 37110 -11510 37155 -11390
rect 37275 -11510 37330 -11390
rect 37450 -11510 37495 -11390
rect 37615 -11510 37660 -11390
rect 37780 -11510 37825 -11390
rect 37945 -11510 38000 -11390
rect 38120 -11510 38165 -11390
rect 38285 -11510 38330 -11390
rect 38450 -11510 38495 -11390
rect 38615 -11510 38670 -11390
rect 38790 -11510 38835 -11390
rect 38955 -11510 39000 -11390
rect 39120 -11510 39165 -11390
rect 39285 -11510 39340 -11390
rect 39460 -11510 39505 -11390
rect 39625 -11510 39670 -11390
rect 39790 -11510 39835 -11390
rect 39955 -11510 40010 -11390
rect 40130 -11510 40175 -11390
rect 40295 -11510 40340 -11390
rect 40460 -11510 40505 -11390
rect 40625 -11510 40680 -11390
rect 40800 -11510 40845 -11390
rect 40965 -11510 41010 -11390
rect 41130 -11510 41175 -11390
rect 41295 -11510 41350 -11390
rect 41470 -11510 41515 -11390
rect 41635 -11510 41680 -11390
rect 41800 -11510 41845 -11390
rect 41965 -11510 42175 -11390
rect 42295 -11510 42350 -11390
rect 42470 -11510 42515 -11390
rect 42635 -11510 42680 -11390
rect 42800 -11510 42845 -11390
rect 42965 -11510 43020 -11390
rect 43140 -11510 43185 -11390
rect 43305 -11510 43350 -11390
rect 43470 -11510 43515 -11390
rect 43635 -11510 43690 -11390
rect 43810 -11510 43855 -11390
rect 43975 -11510 44020 -11390
rect 44140 -11510 44185 -11390
rect 44305 -11510 44360 -11390
rect 44480 -11510 44525 -11390
rect 44645 -11510 44690 -11390
rect 44810 -11510 44855 -11390
rect 44975 -11510 45030 -11390
rect 45150 -11510 45195 -11390
rect 45315 -11510 45360 -11390
rect 45480 -11510 45525 -11390
rect 45645 -11510 45700 -11390
rect 45820 -11510 45865 -11390
rect 45985 -11510 46030 -11390
rect 46150 -11510 46195 -11390
rect 46315 -11510 46370 -11390
rect 46490 -11510 46535 -11390
rect 46655 -11510 46700 -11390
rect 46820 -11510 46865 -11390
rect 46985 -11510 47040 -11390
rect 47160 -11510 47205 -11390
rect 47325 -11510 47370 -11390
rect 47490 -11510 47535 -11390
rect 47655 -11510 47865 -11390
rect 47985 -11510 48040 -11390
rect 48160 -11510 48205 -11390
rect 48325 -11510 48370 -11390
rect 48490 -11510 48535 -11390
rect 48655 -11510 48710 -11390
rect 48830 -11510 48875 -11390
rect 48995 -11510 49040 -11390
rect 49160 -11510 49205 -11390
rect 49325 -11510 49380 -11390
rect 49500 -11510 49545 -11390
rect 49665 -11510 49710 -11390
rect 49830 -11510 49875 -11390
rect 49995 -11510 50050 -11390
rect 50170 -11510 50215 -11390
rect 50335 -11510 50380 -11390
rect 50500 -11510 50545 -11390
rect 50665 -11510 50720 -11390
rect 50840 -11510 50885 -11390
rect 51005 -11510 51050 -11390
rect 51170 -11510 51215 -11390
rect 51335 -11510 51390 -11390
rect 51510 -11510 51555 -11390
rect 51675 -11510 51720 -11390
rect 51840 -11510 51885 -11390
rect 52005 -11510 52060 -11390
rect 52180 -11510 52225 -11390
rect 52345 -11510 52390 -11390
rect 52510 -11510 52555 -11390
rect 52675 -11510 52730 -11390
rect 52850 -11510 52895 -11390
rect 53015 -11510 53060 -11390
rect 53180 -11510 53225 -11390
rect 53345 -11510 53370 -11390
rect 30770 -11555 53370 -11510
rect 30770 -11675 30795 -11555
rect 30915 -11675 30970 -11555
rect 31090 -11675 31135 -11555
rect 31255 -11675 31300 -11555
rect 31420 -11675 31465 -11555
rect 31585 -11675 31640 -11555
rect 31760 -11675 31805 -11555
rect 31925 -11675 31970 -11555
rect 32090 -11675 32135 -11555
rect 32255 -11675 32310 -11555
rect 32430 -11675 32475 -11555
rect 32595 -11675 32640 -11555
rect 32760 -11675 32805 -11555
rect 32925 -11675 32980 -11555
rect 33100 -11675 33145 -11555
rect 33265 -11675 33310 -11555
rect 33430 -11675 33475 -11555
rect 33595 -11675 33650 -11555
rect 33770 -11675 33815 -11555
rect 33935 -11675 33980 -11555
rect 34100 -11675 34145 -11555
rect 34265 -11675 34320 -11555
rect 34440 -11675 34485 -11555
rect 34605 -11675 34650 -11555
rect 34770 -11675 34815 -11555
rect 34935 -11675 34990 -11555
rect 35110 -11675 35155 -11555
rect 35275 -11675 35320 -11555
rect 35440 -11675 35485 -11555
rect 35605 -11675 35660 -11555
rect 35780 -11675 35825 -11555
rect 35945 -11675 35990 -11555
rect 36110 -11675 36155 -11555
rect 36275 -11675 36485 -11555
rect 36605 -11675 36660 -11555
rect 36780 -11675 36825 -11555
rect 36945 -11675 36990 -11555
rect 37110 -11675 37155 -11555
rect 37275 -11675 37330 -11555
rect 37450 -11675 37495 -11555
rect 37615 -11675 37660 -11555
rect 37780 -11675 37825 -11555
rect 37945 -11675 38000 -11555
rect 38120 -11675 38165 -11555
rect 38285 -11675 38330 -11555
rect 38450 -11675 38495 -11555
rect 38615 -11675 38670 -11555
rect 38790 -11675 38835 -11555
rect 38955 -11675 39000 -11555
rect 39120 -11675 39165 -11555
rect 39285 -11675 39340 -11555
rect 39460 -11675 39505 -11555
rect 39625 -11675 39670 -11555
rect 39790 -11675 39835 -11555
rect 39955 -11675 40010 -11555
rect 40130 -11675 40175 -11555
rect 40295 -11675 40340 -11555
rect 40460 -11675 40505 -11555
rect 40625 -11675 40680 -11555
rect 40800 -11675 40845 -11555
rect 40965 -11675 41010 -11555
rect 41130 -11675 41175 -11555
rect 41295 -11675 41350 -11555
rect 41470 -11675 41515 -11555
rect 41635 -11675 41680 -11555
rect 41800 -11675 41845 -11555
rect 41965 -11675 42175 -11555
rect 42295 -11675 42350 -11555
rect 42470 -11675 42515 -11555
rect 42635 -11675 42680 -11555
rect 42800 -11675 42845 -11555
rect 42965 -11675 43020 -11555
rect 43140 -11675 43185 -11555
rect 43305 -11675 43350 -11555
rect 43470 -11675 43515 -11555
rect 43635 -11675 43690 -11555
rect 43810 -11675 43855 -11555
rect 43975 -11675 44020 -11555
rect 44140 -11675 44185 -11555
rect 44305 -11675 44360 -11555
rect 44480 -11675 44525 -11555
rect 44645 -11675 44690 -11555
rect 44810 -11675 44855 -11555
rect 44975 -11675 45030 -11555
rect 45150 -11675 45195 -11555
rect 45315 -11675 45360 -11555
rect 45480 -11675 45525 -11555
rect 45645 -11675 45700 -11555
rect 45820 -11675 45865 -11555
rect 45985 -11675 46030 -11555
rect 46150 -11675 46195 -11555
rect 46315 -11675 46370 -11555
rect 46490 -11675 46535 -11555
rect 46655 -11675 46700 -11555
rect 46820 -11675 46865 -11555
rect 46985 -11675 47040 -11555
rect 47160 -11675 47205 -11555
rect 47325 -11675 47370 -11555
rect 47490 -11675 47535 -11555
rect 47655 -11675 47865 -11555
rect 47985 -11675 48040 -11555
rect 48160 -11675 48205 -11555
rect 48325 -11675 48370 -11555
rect 48490 -11675 48535 -11555
rect 48655 -11675 48710 -11555
rect 48830 -11675 48875 -11555
rect 48995 -11675 49040 -11555
rect 49160 -11675 49205 -11555
rect 49325 -11675 49380 -11555
rect 49500 -11675 49545 -11555
rect 49665 -11675 49710 -11555
rect 49830 -11675 49875 -11555
rect 49995 -11675 50050 -11555
rect 50170 -11675 50215 -11555
rect 50335 -11675 50380 -11555
rect 50500 -11675 50545 -11555
rect 50665 -11675 50720 -11555
rect 50840 -11675 50885 -11555
rect 51005 -11675 51050 -11555
rect 51170 -11675 51215 -11555
rect 51335 -11675 51390 -11555
rect 51510 -11675 51555 -11555
rect 51675 -11675 51720 -11555
rect 51840 -11675 51885 -11555
rect 52005 -11675 52060 -11555
rect 52180 -11675 52225 -11555
rect 52345 -11675 52390 -11555
rect 52510 -11675 52555 -11555
rect 52675 -11675 52730 -11555
rect 52850 -11675 52895 -11555
rect 53015 -11675 53060 -11555
rect 53180 -11675 53225 -11555
rect 53345 -11675 53370 -11555
rect 30770 -11720 53370 -11675
rect 30770 -11840 30795 -11720
rect 30915 -11840 30970 -11720
rect 31090 -11840 31135 -11720
rect 31255 -11840 31300 -11720
rect 31420 -11840 31465 -11720
rect 31585 -11840 31640 -11720
rect 31760 -11840 31805 -11720
rect 31925 -11840 31970 -11720
rect 32090 -11840 32135 -11720
rect 32255 -11840 32310 -11720
rect 32430 -11840 32475 -11720
rect 32595 -11840 32640 -11720
rect 32760 -11840 32805 -11720
rect 32925 -11840 32980 -11720
rect 33100 -11840 33145 -11720
rect 33265 -11840 33310 -11720
rect 33430 -11840 33475 -11720
rect 33595 -11840 33650 -11720
rect 33770 -11840 33815 -11720
rect 33935 -11840 33980 -11720
rect 34100 -11840 34145 -11720
rect 34265 -11840 34320 -11720
rect 34440 -11840 34485 -11720
rect 34605 -11840 34650 -11720
rect 34770 -11840 34815 -11720
rect 34935 -11840 34990 -11720
rect 35110 -11840 35155 -11720
rect 35275 -11840 35320 -11720
rect 35440 -11840 35485 -11720
rect 35605 -11840 35660 -11720
rect 35780 -11840 35825 -11720
rect 35945 -11840 35990 -11720
rect 36110 -11840 36155 -11720
rect 36275 -11840 36485 -11720
rect 36605 -11840 36660 -11720
rect 36780 -11840 36825 -11720
rect 36945 -11840 36990 -11720
rect 37110 -11840 37155 -11720
rect 37275 -11840 37330 -11720
rect 37450 -11840 37495 -11720
rect 37615 -11840 37660 -11720
rect 37780 -11840 37825 -11720
rect 37945 -11840 38000 -11720
rect 38120 -11840 38165 -11720
rect 38285 -11840 38330 -11720
rect 38450 -11840 38495 -11720
rect 38615 -11840 38670 -11720
rect 38790 -11840 38835 -11720
rect 38955 -11840 39000 -11720
rect 39120 -11840 39165 -11720
rect 39285 -11840 39340 -11720
rect 39460 -11840 39505 -11720
rect 39625 -11840 39670 -11720
rect 39790 -11840 39835 -11720
rect 39955 -11840 40010 -11720
rect 40130 -11840 40175 -11720
rect 40295 -11840 40340 -11720
rect 40460 -11840 40505 -11720
rect 40625 -11840 40680 -11720
rect 40800 -11840 40845 -11720
rect 40965 -11840 41010 -11720
rect 41130 -11840 41175 -11720
rect 41295 -11840 41350 -11720
rect 41470 -11840 41515 -11720
rect 41635 -11840 41680 -11720
rect 41800 -11840 41845 -11720
rect 41965 -11840 42175 -11720
rect 42295 -11840 42350 -11720
rect 42470 -11840 42515 -11720
rect 42635 -11840 42680 -11720
rect 42800 -11840 42845 -11720
rect 42965 -11840 43020 -11720
rect 43140 -11840 43185 -11720
rect 43305 -11840 43350 -11720
rect 43470 -11840 43515 -11720
rect 43635 -11840 43690 -11720
rect 43810 -11840 43855 -11720
rect 43975 -11840 44020 -11720
rect 44140 -11840 44185 -11720
rect 44305 -11840 44360 -11720
rect 44480 -11840 44525 -11720
rect 44645 -11840 44690 -11720
rect 44810 -11840 44855 -11720
rect 44975 -11840 45030 -11720
rect 45150 -11840 45195 -11720
rect 45315 -11840 45360 -11720
rect 45480 -11840 45525 -11720
rect 45645 -11840 45700 -11720
rect 45820 -11840 45865 -11720
rect 45985 -11840 46030 -11720
rect 46150 -11840 46195 -11720
rect 46315 -11840 46370 -11720
rect 46490 -11840 46535 -11720
rect 46655 -11840 46700 -11720
rect 46820 -11840 46865 -11720
rect 46985 -11840 47040 -11720
rect 47160 -11840 47205 -11720
rect 47325 -11840 47370 -11720
rect 47490 -11840 47535 -11720
rect 47655 -11840 47865 -11720
rect 47985 -11840 48040 -11720
rect 48160 -11840 48205 -11720
rect 48325 -11840 48370 -11720
rect 48490 -11840 48535 -11720
rect 48655 -11840 48710 -11720
rect 48830 -11840 48875 -11720
rect 48995 -11840 49040 -11720
rect 49160 -11840 49205 -11720
rect 49325 -11840 49380 -11720
rect 49500 -11840 49545 -11720
rect 49665 -11840 49710 -11720
rect 49830 -11840 49875 -11720
rect 49995 -11840 50050 -11720
rect 50170 -11840 50215 -11720
rect 50335 -11840 50380 -11720
rect 50500 -11840 50545 -11720
rect 50665 -11840 50720 -11720
rect 50840 -11840 50885 -11720
rect 51005 -11840 51050 -11720
rect 51170 -11840 51215 -11720
rect 51335 -11840 51390 -11720
rect 51510 -11840 51555 -11720
rect 51675 -11840 51720 -11720
rect 51840 -11840 51885 -11720
rect 52005 -11840 52060 -11720
rect 52180 -11840 52225 -11720
rect 52345 -11840 52390 -11720
rect 52510 -11840 52555 -11720
rect 52675 -11840 52730 -11720
rect 52850 -11840 52895 -11720
rect 53015 -11840 53060 -11720
rect 53180 -11840 53225 -11720
rect 53345 -11840 53370 -11720
rect 30770 -11885 53370 -11840
rect 30770 -12005 30795 -11885
rect 30915 -12005 30970 -11885
rect 31090 -12005 31135 -11885
rect 31255 -12005 31300 -11885
rect 31420 -12005 31465 -11885
rect 31585 -12005 31640 -11885
rect 31760 -12005 31805 -11885
rect 31925 -12005 31970 -11885
rect 32090 -12005 32135 -11885
rect 32255 -12005 32310 -11885
rect 32430 -12005 32475 -11885
rect 32595 -12005 32640 -11885
rect 32760 -12005 32805 -11885
rect 32925 -12005 32980 -11885
rect 33100 -12005 33145 -11885
rect 33265 -12005 33310 -11885
rect 33430 -12005 33475 -11885
rect 33595 -12005 33650 -11885
rect 33770 -12005 33815 -11885
rect 33935 -12005 33980 -11885
rect 34100 -12005 34145 -11885
rect 34265 -12005 34320 -11885
rect 34440 -12005 34485 -11885
rect 34605 -12005 34650 -11885
rect 34770 -12005 34815 -11885
rect 34935 -12005 34990 -11885
rect 35110 -12005 35155 -11885
rect 35275 -12005 35320 -11885
rect 35440 -12005 35485 -11885
rect 35605 -12005 35660 -11885
rect 35780 -12005 35825 -11885
rect 35945 -12005 35990 -11885
rect 36110 -12005 36155 -11885
rect 36275 -12005 36485 -11885
rect 36605 -12005 36660 -11885
rect 36780 -12005 36825 -11885
rect 36945 -12005 36990 -11885
rect 37110 -12005 37155 -11885
rect 37275 -12005 37330 -11885
rect 37450 -12005 37495 -11885
rect 37615 -12005 37660 -11885
rect 37780 -12005 37825 -11885
rect 37945 -12005 38000 -11885
rect 38120 -12005 38165 -11885
rect 38285 -12005 38330 -11885
rect 38450 -12005 38495 -11885
rect 38615 -12005 38670 -11885
rect 38790 -12005 38835 -11885
rect 38955 -12005 39000 -11885
rect 39120 -12005 39165 -11885
rect 39285 -12005 39340 -11885
rect 39460 -12005 39505 -11885
rect 39625 -12005 39670 -11885
rect 39790 -12005 39835 -11885
rect 39955 -12005 40010 -11885
rect 40130 -12005 40175 -11885
rect 40295 -12005 40340 -11885
rect 40460 -12005 40505 -11885
rect 40625 -12005 40680 -11885
rect 40800 -12005 40845 -11885
rect 40965 -12005 41010 -11885
rect 41130 -12005 41175 -11885
rect 41295 -12005 41350 -11885
rect 41470 -12005 41515 -11885
rect 41635 -12005 41680 -11885
rect 41800 -12005 41845 -11885
rect 41965 -12005 42175 -11885
rect 42295 -12005 42350 -11885
rect 42470 -12005 42515 -11885
rect 42635 -12005 42680 -11885
rect 42800 -12005 42845 -11885
rect 42965 -12005 43020 -11885
rect 43140 -12005 43185 -11885
rect 43305 -12005 43350 -11885
rect 43470 -12005 43515 -11885
rect 43635 -12005 43690 -11885
rect 43810 -12005 43855 -11885
rect 43975 -12005 44020 -11885
rect 44140 -12005 44185 -11885
rect 44305 -12005 44360 -11885
rect 44480 -12005 44525 -11885
rect 44645 -12005 44690 -11885
rect 44810 -12005 44855 -11885
rect 44975 -12005 45030 -11885
rect 45150 -12005 45195 -11885
rect 45315 -12005 45360 -11885
rect 45480 -12005 45525 -11885
rect 45645 -12005 45700 -11885
rect 45820 -12005 45865 -11885
rect 45985 -12005 46030 -11885
rect 46150 -12005 46195 -11885
rect 46315 -12005 46370 -11885
rect 46490 -12005 46535 -11885
rect 46655 -12005 46700 -11885
rect 46820 -12005 46865 -11885
rect 46985 -12005 47040 -11885
rect 47160 -12005 47205 -11885
rect 47325 -12005 47370 -11885
rect 47490 -12005 47535 -11885
rect 47655 -12005 47865 -11885
rect 47985 -12005 48040 -11885
rect 48160 -12005 48205 -11885
rect 48325 -12005 48370 -11885
rect 48490 -12005 48535 -11885
rect 48655 -12005 48710 -11885
rect 48830 -12005 48875 -11885
rect 48995 -12005 49040 -11885
rect 49160 -12005 49205 -11885
rect 49325 -12005 49380 -11885
rect 49500 -12005 49545 -11885
rect 49665 -12005 49710 -11885
rect 49830 -12005 49875 -11885
rect 49995 -12005 50050 -11885
rect 50170 -12005 50215 -11885
rect 50335 -12005 50380 -11885
rect 50500 -12005 50545 -11885
rect 50665 -12005 50720 -11885
rect 50840 -12005 50885 -11885
rect 51005 -12005 51050 -11885
rect 51170 -12005 51215 -11885
rect 51335 -12005 51390 -11885
rect 51510 -12005 51555 -11885
rect 51675 -12005 51720 -11885
rect 51840 -12005 51885 -11885
rect 52005 -12005 52060 -11885
rect 52180 -12005 52225 -11885
rect 52345 -12005 52390 -11885
rect 52510 -12005 52555 -11885
rect 52675 -12005 52730 -11885
rect 52850 -12005 52895 -11885
rect 53015 -12005 53060 -11885
rect 53180 -12005 53225 -11885
rect 53345 -12005 53370 -11885
rect 30770 -12060 53370 -12005
rect 30770 -12180 30795 -12060
rect 30915 -12180 30970 -12060
rect 31090 -12180 31135 -12060
rect 31255 -12180 31300 -12060
rect 31420 -12180 31465 -12060
rect 31585 -12180 31640 -12060
rect 31760 -12180 31805 -12060
rect 31925 -12180 31970 -12060
rect 32090 -12180 32135 -12060
rect 32255 -12180 32310 -12060
rect 32430 -12180 32475 -12060
rect 32595 -12180 32640 -12060
rect 32760 -12180 32805 -12060
rect 32925 -12180 32980 -12060
rect 33100 -12180 33145 -12060
rect 33265 -12180 33310 -12060
rect 33430 -12180 33475 -12060
rect 33595 -12180 33650 -12060
rect 33770 -12180 33815 -12060
rect 33935 -12180 33980 -12060
rect 34100 -12180 34145 -12060
rect 34265 -12180 34320 -12060
rect 34440 -12180 34485 -12060
rect 34605 -12180 34650 -12060
rect 34770 -12180 34815 -12060
rect 34935 -12180 34990 -12060
rect 35110 -12180 35155 -12060
rect 35275 -12180 35320 -12060
rect 35440 -12180 35485 -12060
rect 35605 -12180 35660 -12060
rect 35780 -12180 35825 -12060
rect 35945 -12180 35990 -12060
rect 36110 -12180 36155 -12060
rect 36275 -12180 36485 -12060
rect 36605 -12180 36660 -12060
rect 36780 -12180 36825 -12060
rect 36945 -12180 36990 -12060
rect 37110 -12180 37155 -12060
rect 37275 -12180 37330 -12060
rect 37450 -12180 37495 -12060
rect 37615 -12180 37660 -12060
rect 37780 -12180 37825 -12060
rect 37945 -12180 38000 -12060
rect 38120 -12180 38165 -12060
rect 38285 -12180 38330 -12060
rect 38450 -12180 38495 -12060
rect 38615 -12180 38670 -12060
rect 38790 -12180 38835 -12060
rect 38955 -12180 39000 -12060
rect 39120 -12180 39165 -12060
rect 39285 -12180 39340 -12060
rect 39460 -12180 39505 -12060
rect 39625 -12180 39670 -12060
rect 39790 -12180 39835 -12060
rect 39955 -12180 40010 -12060
rect 40130 -12180 40175 -12060
rect 40295 -12180 40340 -12060
rect 40460 -12180 40505 -12060
rect 40625 -12180 40680 -12060
rect 40800 -12180 40845 -12060
rect 40965 -12180 41010 -12060
rect 41130 -12180 41175 -12060
rect 41295 -12180 41350 -12060
rect 41470 -12180 41515 -12060
rect 41635 -12180 41680 -12060
rect 41800 -12180 41845 -12060
rect 41965 -12180 42175 -12060
rect 42295 -12180 42350 -12060
rect 42470 -12180 42515 -12060
rect 42635 -12180 42680 -12060
rect 42800 -12180 42845 -12060
rect 42965 -12180 43020 -12060
rect 43140 -12180 43185 -12060
rect 43305 -12180 43350 -12060
rect 43470 -12180 43515 -12060
rect 43635 -12180 43690 -12060
rect 43810 -12180 43855 -12060
rect 43975 -12180 44020 -12060
rect 44140 -12180 44185 -12060
rect 44305 -12180 44360 -12060
rect 44480 -12180 44525 -12060
rect 44645 -12180 44690 -12060
rect 44810 -12180 44855 -12060
rect 44975 -12180 45030 -12060
rect 45150 -12180 45195 -12060
rect 45315 -12180 45360 -12060
rect 45480 -12180 45525 -12060
rect 45645 -12180 45700 -12060
rect 45820 -12180 45865 -12060
rect 45985 -12180 46030 -12060
rect 46150 -12180 46195 -12060
rect 46315 -12180 46370 -12060
rect 46490 -12180 46535 -12060
rect 46655 -12180 46700 -12060
rect 46820 -12180 46865 -12060
rect 46985 -12180 47040 -12060
rect 47160 -12180 47205 -12060
rect 47325 -12180 47370 -12060
rect 47490 -12180 47535 -12060
rect 47655 -12180 47865 -12060
rect 47985 -12180 48040 -12060
rect 48160 -12180 48205 -12060
rect 48325 -12180 48370 -12060
rect 48490 -12180 48535 -12060
rect 48655 -12180 48710 -12060
rect 48830 -12180 48875 -12060
rect 48995 -12180 49040 -12060
rect 49160 -12180 49205 -12060
rect 49325 -12180 49380 -12060
rect 49500 -12180 49545 -12060
rect 49665 -12180 49710 -12060
rect 49830 -12180 49875 -12060
rect 49995 -12180 50050 -12060
rect 50170 -12180 50215 -12060
rect 50335 -12180 50380 -12060
rect 50500 -12180 50545 -12060
rect 50665 -12180 50720 -12060
rect 50840 -12180 50885 -12060
rect 51005 -12180 51050 -12060
rect 51170 -12180 51215 -12060
rect 51335 -12180 51390 -12060
rect 51510 -12180 51555 -12060
rect 51675 -12180 51720 -12060
rect 51840 -12180 51885 -12060
rect 52005 -12180 52060 -12060
rect 52180 -12180 52225 -12060
rect 52345 -12180 52390 -12060
rect 52510 -12180 52555 -12060
rect 52675 -12180 52730 -12060
rect 52850 -12180 52895 -12060
rect 53015 -12180 53060 -12060
rect 53180 -12180 53225 -12060
rect 53345 -12180 53370 -12060
rect 30770 -12225 53370 -12180
rect 30770 -12345 30795 -12225
rect 30915 -12345 30970 -12225
rect 31090 -12345 31135 -12225
rect 31255 -12345 31300 -12225
rect 31420 -12345 31465 -12225
rect 31585 -12345 31640 -12225
rect 31760 -12345 31805 -12225
rect 31925 -12345 31970 -12225
rect 32090 -12345 32135 -12225
rect 32255 -12345 32310 -12225
rect 32430 -12345 32475 -12225
rect 32595 -12345 32640 -12225
rect 32760 -12345 32805 -12225
rect 32925 -12345 32980 -12225
rect 33100 -12345 33145 -12225
rect 33265 -12345 33310 -12225
rect 33430 -12345 33475 -12225
rect 33595 -12345 33650 -12225
rect 33770 -12345 33815 -12225
rect 33935 -12345 33980 -12225
rect 34100 -12345 34145 -12225
rect 34265 -12345 34320 -12225
rect 34440 -12345 34485 -12225
rect 34605 -12345 34650 -12225
rect 34770 -12345 34815 -12225
rect 34935 -12345 34990 -12225
rect 35110 -12345 35155 -12225
rect 35275 -12345 35320 -12225
rect 35440 -12345 35485 -12225
rect 35605 -12345 35660 -12225
rect 35780 -12345 35825 -12225
rect 35945 -12345 35990 -12225
rect 36110 -12345 36155 -12225
rect 36275 -12345 36485 -12225
rect 36605 -12345 36660 -12225
rect 36780 -12345 36825 -12225
rect 36945 -12345 36990 -12225
rect 37110 -12345 37155 -12225
rect 37275 -12345 37330 -12225
rect 37450 -12345 37495 -12225
rect 37615 -12345 37660 -12225
rect 37780 -12345 37825 -12225
rect 37945 -12345 38000 -12225
rect 38120 -12345 38165 -12225
rect 38285 -12345 38330 -12225
rect 38450 -12345 38495 -12225
rect 38615 -12345 38670 -12225
rect 38790 -12345 38835 -12225
rect 38955 -12345 39000 -12225
rect 39120 -12345 39165 -12225
rect 39285 -12345 39340 -12225
rect 39460 -12345 39505 -12225
rect 39625 -12345 39670 -12225
rect 39790 -12345 39835 -12225
rect 39955 -12345 40010 -12225
rect 40130 -12345 40175 -12225
rect 40295 -12345 40340 -12225
rect 40460 -12345 40505 -12225
rect 40625 -12345 40680 -12225
rect 40800 -12345 40845 -12225
rect 40965 -12345 41010 -12225
rect 41130 -12345 41175 -12225
rect 41295 -12345 41350 -12225
rect 41470 -12345 41515 -12225
rect 41635 -12345 41680 -12225
rect 41800 -12345 41845 -12225
rect 41965 -12345 42175 -12225
rect 42295 -12345 42350 -12225
rect 42470 -12345 42515 -12225
rect 42635 -12345 42680 -12225
rect 42800 -12345 42845 -12225
rect 42965 -12345 43020 -12225
rect 43140 -12345 43185 -12225
rect 43305 -12345 43350 -12225
rect 43470 -12345 43515 -12225
rect 43635 -12345 43690 -12225
rect 43810 -12345 43855 -12225
rect 43975 -12345 44020 -12225
rect 44140 -12345 44185 -12225
rect 44305 -12345 44360 -12225
rect 44480 -12345 44525 -12225
rect 44645 -12345 44690 -12225
rect 44810 -12345 44855 -12225
rect 44975 -12345 45030 -12225
rect 45150 -12345 45195 -12225
rect 45315 -12345 45360 -12225
rect 45480 -12345 45525 -12225
rect 45645 -12345 45700 -12225
rect 45820 -12345 45865 -12225
rect 45985 -12345 46030 -12225
rect 46150 -12345 46195 -12225
rect 46315 -12345 46370 -12225
rect 46490 -12345 46535 -12225
rect 46655 -12345 46700 -12225
rect 46820 -12345 46865 -12225
rect 46985 -12345 47040 -12225
rect 47160 -12345 47205 -12225
rect 47325 -12345 47370 -12225
rect 47490 -12345 47535 -12225
rect 47655 -12345 47865 -12225
rect 47985 -12345 48040 -12225
rect 48160 -12345 48205 -12225
rect 48325 -12345 48370 -12225
rect 48490 -12345 48535 -12225
rect 48655 -12345 48710 -12225
rect 48830 -12345 48875 -12225
rect 48995 -12345 49040 -12225
rect 49160 -12345 49205 -12225
rect 49325 -12345 49380 -12225
rect 49500 -12345 49545 -12225
rect 49665 -12345 49710 -12225
rect 49830 -12345 49875 -12225
rect 49995 -12345 50050 -12225
rect 50170 -12345 50215 -12225
rect 50335 -12345 50380 -12225
rect 50500 -12345 50545 -12225
rect 50665 -12345 50720 -12225
rect 50840 -12345 50885 -12225
rect 51005 -12345 51050 -12225
rect 51170 -12345 51215 -12225
rect 51335 -12345 51390 -12225
rect 51510 -12345 51555 -12225
rect 51675 -12345 51720 -12225
rect 51840 -12345 51885 -12225
rect 52005 -12345 52060 -12225
rect 52180 -12345 52225 -12225
rect 52345 -12345 52390 -12225
rect 52510 -12345 52555 -12225
rect 52675 -12345 52730 -12225
rect 52850 -12345 52895 -12225
rect 53015 -12345 53060 -12225
rect 53180 -12345 53225 -12225
rect 53345 -12345 53370 -12225
rect 30770 -12390 53370 -12345
rect 30770 -12510 30795 -12390
rect 30915 -12510 30970 -12390
rect 31090 -12510 31135 -12390
rect 31255 -12510 31300 -12390
rect 31420 -12510 31465 -12390
rect 31585 -12510 31640 -12390
rect 31760 -12510 31805 -12390
rect 31925 -12510 31970 -12390
rect 32090 -12510 32135 -12390
rect 32255 -12510 32310 -12390
rect 32430 -12510 32475 -12390
rect 32595 -12510 32640 -12390
rect 32760 -12510 32805 -12390
rect 32925 -12510 32980 -12390
rect 33100 -12510 33145 -12390
rect 33265 -12510 33310 -12390
rect 33430 -12510 33475 -12390
rect 33595 -12510 33650 -12390
rect 33770 -12510 33815 -12390
rect 33935 -12510 33980 -12390
rect 34100 -12510 34145 -12390
rect 34265 -12510 34320 -12390
rect 34440 -12510 34485 -12390
rect 34605 -12510 34650 -12390
rect 34770 -12510 34815 -12390
rect 34935 -12510 34990 -12390
rect 35110 -12510 35155 -12390
rect 35275 -12510 35320 -12390
rect 35440 -12510 35485 -12390
rect 35605 -12510 35660 -12390
rect 35780 -12510 35825 -12390
rect 35945 -12510 35990 -12390
rect 36110 -12510 36155 -12390
rect 36275 -12510 36485 -12390
rect 36605 -12510 36660 -12390
rect 36780 -12510 36825 -12390
rect 36945 -12510 36990 -12390
rect 37110 -12510 37155 -12390
rect 37275 -12510 37330 -12390
rect 37450 -12510 37495 -12390
rect 37615 -12510 37660 -12390
rect 37780 -12510 37825 -12390
rect 37945 -12510 38000 -12390
rect 38120 -12510 38165 -12390
rect 38285 -12510 38330 -12390
rect 38450 -12510 38495 -12390
rect 38615 -12510 38670 -12390
rect 38790 -12510 38835 -12390
rect 38955 -12510 39000 -12390
rect 39120 -12510 39165 -12390
rect 39285 -12510 39340 -12390
rect 39460 -12510 39505 -12390
rect 39625 -12510 39670 -12390
rect 39790 -12510 39835 -12390
rect 39955 -12510 40010 -12390
rect 40130 -12510 40175 -12390
rect 40295 -12510 40340 -12390
rect 40460 -12510 40505 -12390
rect 40625 -12510 40680 -12390
rect 40800 -12510 40845 -12390
rect 40965 -12510 41010 -12390
rect 41130 -12510 41175 -12390
rect 41295 -12510 41350 -12390
rect 41470 -12510 41515 -12390
rect 41635 -12510 41680 -12390
rect 41800 -12510 41845 -12390
rect 41965 -12510 42175 -12390
rect 42295 -12510 42350 -12390
rect 42470 -12510 42515 -12390
rect 42635 -12510 42680 -12390
rect 42800 -12510 42845 -12390
rect 42965 -12510 43020 -12390
rect 43140 -12510 43185 -12390
rect 43305 -12510 43350 -12390
rect 43470 -12510 43515 -12390
rect 43635 -12510 43690 -12390
rect 43810 -12510 43855 -12390
rect 43975 -12510 44020 -12390
rect 44140 -12510 44185 -12390
rect 44305 -12510 44360 -12390
rect 44480 -12510 44525 -12390
rect 44645 -12510 44690 -12390
rect 44810 -12510 44855 -12390
rect 44975 -12510 45030 -12390
rect 45150 -12510 45195 -12390
rect 45315 -12510 45360 -12390
rect 45480 -12510 45525 -12390
rect 45645 -12510 45700 -12390
rect 45820 -12510 45865 -12390
rect 45985 -12510 46030 -12390
rect 46150 -12510 46195 -12390
rect 46315 -12510 46370 -12390
rect 46490 -12510 46535 -12390
rect 46655 -12510 46700 -12390
rect 46820 -12510 46865 -12390
rect 46985 -12510 47040 -12390
rect 47160 -12510 47205 -12390
rect 47325 -12510 47370 -12390
rect 47490 -12510 47535 -12390
rect 47655 -12510 47865 -12390
rect 47985 -12510 48040 -12390
rect 48160 -12510 48205 -12390
rect 48325 -12510 48370 -12390
rect 48490 -12510 48535 -12390
rect 48655 -12510 48710 -12390
rect 48830 -12510 48875 -12390
rect 48995 -12510 49040 -12390
rect 49160 -12510 49205 -12390
rect 49325 -12510 49380 -12390
rect 49500 -12510 49545 -12390
rect 49665 -12510 49710 -12390
rect 49830 -12510 49875 -12390
rect 49995 -12510 50050 -12390
rect 50170 -12510 50215 -12390
rect 50335 -12510 50380 -12390
rect 50500 -12510 50545 -12390
rect 50665 -12510 50720 -12390
rect 50840 -12510 50885 -12390
rect 51005 -12510 51050 -12390
rect 51170 -12510 51215 -12390
rect 51335 -12510 51390 -12390
rect 51510 -12510 51555 -12390
rect 51675 -12510 51720 -12390
rect 51840 -12510 51885 -12390
rect 52005 -12510 52060 -12390
rect 52180 -12510 52225 -12390
rect 52345 -12510 52390 -12390
rect 52510 -12510 52555 -12390
rect 52675 -12510 52730 -12390
rect 52850 -12510 52895 -12390
rect 53015 -12510 53060 -12390
rect 53180 -12510 53225 -12390
rect 53345 -12510 53370 -12390
rect 30770 -12555 53370 -12510
rect 30770 -12675 30795 -12555
rect 30915 -12675 30970 -12555
rect 31090 -12675 31135 -12555
rect 31255 -12675 31300 -12555
rect 31420 -12675 31465 -12555
rect 31585 -12675 31640 -12555
rect 31760 -12675 31805 -12555
rect 31925 -12675 31970 -12555
rect 32090 -12675 32135 -12555
rect 32255 -12675 32310 -12555
rect 32430 -12675 32475 -12555
rect 32595 -12675 32640 -12555
rect 32760 -12675 32805 -12555
rect 32925 -12675 32980 -12555
rect 33100 -12675 33145 -12555
rect 33265 -12675 33310 -12555
rect 33430 -12675 33475 -12555
rect 33595 -12675 33650 -12555
rect 33770 -12675 33815 -12555
rect 33935 -12675 33980 -12555
rect 34100 -12675 34145 -12555
rect 34265 -12675 34320 -12555
rect 34440 -12675 34485 -12555
rect 34605 -12675 34650 -12555
rect 34770 -12675 34815 -12555
rect 34935 -12675 34990 -12555
rect 35110 -12675 35155 -12555
rect 35275 -12675 35320 -12555
rect 35440 -12675 35485 -12555
rect 35605 -12675 35660 -12555
rect 35780 -12675 35825 -12555
rect 35945 -12675 35990 -12555
rect 36110 -12675 36155 -12555
rect 36275 -12675 36485 -12555
rect 36605 -12675 36660 -12555
rect 36780 -12675 36825 -12555
rect 36945 -12675 36990 -12555
rect 37110 -12675 37155 -12555
rect 37275 -12675 37330 -12555
rect 37450 -12675 37495 -12555
rect 37615 -12675 37660 -12555
rect 37780 -12675 37825 -12555
rect 37945 -12675 38000 -12555
rect 38120 -12675 38165 -12555
rect 38285 -12675 38330 -12555
rect 38450 -12675 38495 -12555
rect 38615 -12675 38670 -12555
rect 38790 -12675 38835 -12555
rect 38955 -12675 39000 -12555
rect 39120 -12675 39165 -12555
rect 39285 -12675 39340 -12555
rect 39460 -12675 39505 -12555
rect 39625 -12675 39670 -12555
rect 39790 -12675 39835 -12555
rect 39955 -12675 40010 -12555
rect 40130 -12675 40175 -12555
rect 40295 -12675 40340 -12555
rect 40460 -12675 40505 -12555
rect 40625 -12675 40680 -12555
rect 40800 -12675 40845 -12555
rect 40965 -12675 41010 -12555
rect 41130 -12675 41175 -12555
rect 41295 -12675 41350 -12555
rect 41470 -12675 41515 -12555
rect 41635 -12675 41680 -12555
rect 41800 -12675 41845 -12555
rect 41965 -12675 42175 -12555
rect 42295 -12675 42350 -12555
rect 42470 -12675 42515 -12555
rect 42635 -12675 42680 -12555
rect 42800 -12675 42845 -12555
rect 42965 -12675 43020 -12555
rect 43140 -12675 43185 -12555
rect 43305 -12675 43350 -12555
rect 43470 -12675 43515 -12555
rect 43635 -12675 43690 -12555
rect 43810 -12675 43855 -12555
rect 43975 -12675 44020 -12555
rect 44140 -12675 44185 -12555
rect 44305 -12675 44360 -12555
rect 44480 -12675 44525 -12555
rect 44645 -12675 44690 -12555
rect 44810 -12675 44855 -12555
rect 44975 -12675 45030 -12555
rect 45150 -12675 45195 -12555
rect 45315 -12675 45360 -12555
rect 45480 -12675 45525 -12555
rect 45645 -12675 45700 -12555
rect 45820 -12675 45865 -12555
rect 45985 -12675 46030 -12555
rect 46150 -12675 46195 -12555
rect 46315 -12675 46370 -12555
rect 46490 -12675 46535 -12555
rect 46655 -12675 46700 -12555
rect 46820 -12675 46865 -12555
rect 46985 -12675 47040 -12555
rect 47160 -12675 47205 -12555
rect 47325 -12675 47370 -12555
rect 47490 -12675 47535 -12555
rect 47655 -12675 47865 -12555
rect 47985 -12675 48040 -12555
rect 48160 -12675 48205 -12555
rect 48325 -12675 48370 -12555
rect 48490 -12675 48535 -12555
rect 48655 -12675 48710 -12555
rect 48830 -12675 48875 -12555
rect 48995 -12675 49040 -12555
rect 49160 -12675 49205 -12555
rect 49325 -12675 49380 -12555
rect 49500 -12675 49545 -12555
rect 49665 -12675 49710 -12555
rect 49830 -12675 49875 -12555
rect 49995 -12675 50050 -12555
rect 50170 -12675 50215 -12555
rect 50335 -12675 50380 -12555
rect 50500 -12675 50545 -12555
rect 50665 -12675 50720 -12555
rect 50840 -12675 50885 -12555
rect 51005 -12675 51050 -12555
rect 51170 -12675 51215 -12555
rect 51335 -12675 51390 -12555
rect 51510 -12675 51555 -12555
rect 51675 -12675 51720 -12555
rect 51840 -12675 51885 -12555
rect 52005 -12675 52060 -12555
rect 52180 -12675 52225 -12555
rect 52345 -12675 52390 -12555
rect 52510 -12675 52555 -12555
rect 52675 -12675 52730 -12555
rect 52850 -12675 52895 -12555
rect 53015 -12675 53060 -12555
rect 53180 -12675 53225 -12555
rect 53345 -12675 53370 -12555
rect 30770 -12730 53370 -12675
rect 30770 -12850 30795 -12730
rect 30915 -12850 30970 -12730
rect 31090 -12850 31135 -12730
rect 31255 -12850 31300 -12730
rect 31420 -12850 31465 -12730
rect 31585 -12850 31640 -12730
rect 31760 -12850 31805 -12730
rect 31925 -12850 31970 -12730
rect 32090 -12850 32135 -12730
rect 32255 -12850 32310 -12730
rect 32430 -12850 32475 -12730
rect 32595 -12850 32640 -12730
rect 32760 -12850 32805 -12730
rect 32925 -12850 32980 -12730
rect 33100 -12850 33145 -12730
rect 33265 -12850 33310 -12730
rect 33430 -12850 33475 -12730
rect 33595 -12850 33650 -12730
rect 33770 -12850 33815 -12730
rect 33935 -12850 33980 -12730
rect 34100 -12850 34145 -12730
rect 34265 -12850 34320 -12730
rect 34440 -12850 34485 -12730
rect 34605 -12850 34650 -12730
rect 34770 -12850 34815 -12730
rect 34935 -12850 34990 -12730
rect 35110 -12850 35155 -12730
rect 35275 -12850 35320 -12730
rect 35440 -12850 35485 -12730
rect 35605 -12850 35660 -12730
rect 35780 -12850 35825 -12730
rect 35945 -12850 35990 -12730
rect 36110 -12850 36155 -12730
rect 36275 -12850 36485 -12730
rect 36605 -12850 36660 -12730
rect 36780 -12850 36825 -12730
rect 36945 -12850 36990 -12730
rect 37110 -12850 37155 -12730
rect 37275 -12850 37330 -12730
rect 37450 -12850 37495 -12730
rect 37615 -12850 37660 -12730
rect 37780 -12850 37825 -12730
rect 37945 -12850 38000 -12730
rect 38120 -12850 38165 -12730
rect 38285 -12850 38330 -12730
rect 38450 -12850 38495 -12730
rect 38615 -12850 38670 -12730
rect 38790 -12850 38835 -12730
rect 38955 -12850 39000 -12730
rect 39120 -12850 39165 -12730
rect 39285 -12850 39340 -12730
rect 39460 -12850 39505 -12730
rect 39625 -12850 39670 -12730
rect 39790 -12850 39835 -12730
rect 39955 -12850 40010 -12730
rect 40130 -12850 40175 -12730
rect 40295 -12850 40340 -12730
rect 40460 -12850 40505 -12730
rect 40625 -12850 40680 -12730
rect 40800 -12850 40845 -12730
rect 40965 -12850 41010 -12730
rect 41130 -12850 41175 -12730
rect 41295 -12850 41350 -12730
rect 41470 -12850 41515 -12730
rect 41635 -12850 41680 -12730
rect 41800 -12850 41845 -12730
rect 41965 -12850 42175 -12730
rect 42295 -12850 42350 -12730
rect 42470 -12850 42515 -12730
rect 42635 -12850 42680 -12730
rect 42800 -12850 42845 -12730
rect 42965 -12850 43020 -12730
rect 43140 -12850 43185 -12730
rect 43305 -12850 43350 -12730
rect 43470 -12850 43515 -12730
rect 43635 -12850 43690 -12730
rect 43810 -12850 43855 -12730
rect 43975 -12850 44020 -12730
rect 44140 -12850 44185 -12730
rect 44305 -12850 44360 -12730
rect 44480 -12850 44525 -12730
rect 44645 -12850 44690 -12730
rect 44810 -12850 44855 -12730
rect 44975 -12850 45030 -12730
rect 45150 -12850 45195 -12730
rect 45315 -12850 45360 -12730
rect 45480 -12850 45525 -12730
rect 45645 -12850 45700 -12730
rect 45820 -12850 45865 -12730
rect 45985 -12850 46030 -12730
rect 46150 -12850 46195 -12730
rect 46315 -12850 46370 -12730
rect 46490 -12850 46535 -12730
rect 46655 -12850 46700 -12730
rect 46820 -12850 46865 -12730
rect 46985 -12850 47040 -12730
rect 47160 -12850 47205 -12730
rect 47325 -12850 47370 -12730
rect 47490 -12850 47535 -12730
rect 47655 -12850 47865 -12730
rect 47985 -12850 48040 -12730
rect 48160 -12850 48205 -12730
rect 48325 -12850 48370 -12730
rect 48490 -12850 48535 -12730
rect 48655 -12850 48710 -12730
rect 48830 -12850 48875 -12730
rect 48995 -12850 49040 -12730
rect 49160 -12850 49205 -12730
rect 49325 -12850 49380 -12730
rect 49500 -12850 49545 -12730
rect 49665 -12850 49710 -12730
rect 49830 -12850 49875 -12730
rect 49995 -12850 50050 -12730
rect 50170 -12850 50215 -12730
rect 50335 -12850 50380 -12730
rect 50500 -12850 50545 -12730
rect 50665 -12850 50720 -12730
rect 50840 -12850 50885 -12730
rect 51005 -12850 51050 -12730
rect 51170 -12850 51215 -12730
rect 51335 -12850 51390 -12730
rect 51510 -12850 51555 -12730
rect 51675 -12850 51720 -12730
rect 51840 -12850 51885 -12730
rect 52005 -12850 52060 -12730
rect 52180 -12850 52225 -12730
rect 52345 -12850 52390 -12730
rect 52510 -12850 52555 -12730
rect 52675 -12850 52730 -12730
rect 52850 -12850 52895 -12730
rect 53015 -12850 53060 -12730
rect 53180 -12850 53225 -12730
rect 53345 -12850 53370 -12730
rect 30770 -12895 53370 -12850
rect 30770 -13015 30795 -12895
rect 30915 -13015 30970 -12895
rect 31090 -13015 31135 -12895
rect 31255 -13015 31300 -12895
rect 31420 -13015 31465 -12895
rect 31585 -13015 31640 -12895
rect 31760 -13015 31805 -12895
rect 31925 -13015 31970 -12895
rect 32090 -13015 32135 -12895
rect 32255 -13015 32310 -12895
rect 32430 -13015 32475 -12895
rect 32595 -13015 32640 -12895
rect 32760 -13015 32805 -12895
rect 32925 -13015 32980 -12895
rect 33100 -13015 33145 -12895
rect 33265 -13015 33310 -12895
rect 33430 -13015 33475 -12895
rect 33595 -13015 33650 -12895
rect 33770 -13015 33815 -12895
rect 33935 -13015 33980 -12895
rect 34100 -13015 34145 -12895
rect 34265 -13015 34320 -12895
rect 34440 -13015 34485 -12895
rect 34605 -13015 34650 -12895
rect 34770 -13015 34815 -12895
rect 34935 -13015 34990 -12895
rect 35110 -13015 35155 -12895
rect 35275 -13015 35320 -12895
rect 35440 -13015 35485 -12895
rect 35605 -13015 35660 -12895
rect 35780 -13015 35825 -12895
rect 35945 -13015 35990 -12895
rect 36110 -13015 36155 -12895
rect 36275 -13015 36485 -12895
rect 36605 -13015 36660 -12895
rect 36780 -13015 36825 -12895
rect 36945 -13015 36990 -12895
rect 37110 -13015 37155 -12895
rect 37275 -13015 37330 -12895
rect 37450 -13015 37495 -12895
rect 37615 -13015 37660 -12895
rect 37780 -13015 37825 -12895
rect 37945 -13015 38000 -12895
rect 38120 -13015 38165 -12895
rect 38285 -13015 38330 -12895
rect 38450 -13015 38495 -12895
rect 38615 -13015 38670 -12895
rect 38790 -13015 38835 -12895
rect 38955 -13015 39000 -12895
rect 39120 -13015 39165 -12895
rect 39285 -13015 39340 -12895
rect 39460 -13015 39505 -12895
rect 39625 -13015 39670 -12895
rect 39790 -13015 39835 -12895
rect 39955 -13015 40010 -12895
rect 40130 -13015 40175 -12895
rect 40295 -13015 40340 -12895
rect 40460 -13015 40505 -12895
rect 40625 -13015 40680 -12895
rect 40800 -13015 40845 -12895
rect 40965 -13015 41010 -12895
rect 41130 -13015 41175 -12895
rect 41295 -13015 41350 -12895
rect 41470 -13015 41515 -12895
rect 41635 -13015 41680 -12895
rect 41800 -13015 41845 -12895
rect 41965 -13015 42175 -12895
rect 42295 -13015 42350 -12895
rect 42470 -13015 42515 -12895
rect 42635 -13015 42680 -12895
rect 42800 -13015 42845 -12895
rect 42965 -13015 43020 -12895
rect 43140 -13015 43185 -12895
rect 43305 -13015 43350 -12895
rect 43470 -13015 43515 -12895
rect 43635 -13015 43690 -12895
rect 43810 -13015 43855 -12895
rect 43975 -13015 44020 -12895
rect 44140 -13015 44185 -12895
rect 44305 -13015 44360 -12895
rect 44480 -13015 44525 -12895
rect 44645 -13015 44690 -12895
rect 44810 -13015 44855 -12895
rect 44975 -13015 45030 -12895
rect 45150 -13015 45195 -12895
rect 45315 -13015 45360 -12895
rect 45480 -13015 45525 -12895
rect 45645 -13015 45700 -12895
rect 45820 -13015 45865 -12895
rect 45985 -13015 46030 -12895
rect 46150 -13015 46195 -12895
rect 46315 -13015 46370 -12895
rect 46490 -13015 46535 -12895
rect 46655 -13015 46700 -12895
rect 46820 -13015 46865 -12895
rect 46985 -13015 47040 -12895
rect 47160 -13015 47205 -12895
rect 47325 -13015 47370 -12895
rect 47490 -13015 47535 -12895
rect 47655 -13015 47865 -12895
rect 47985 -13015 48040 -12895
rect 48160 -13015 48205 -12895
rect 48325 -13015 48370 -12895
rect 48490 -13015 48535 -12895
rect 48655 -13015 48710 -12895
rect 48830 -13015 48875 -12895
rect 48995 -13015 49040 -12895
rect 49160 -13015 49205 -12895
rect 49325 -13015 49380 -12895
rect 49500 -13015 49545 -12895
rect 49665 -13015 49710 -12895
rect 49830 -13015 49875 -12895
rect 49995 -13015 50050 -12895
rect 50170 -13015 50215 -12895
rect 50335 -13015 50380 -12895
rect 50500 -13015 50545 -12895
rect 50665 -13015 50720 -12895
rect 50840 -13015 50885 -12895
rect 51005 -13015 51050 -12895
rect 51170 -13015 51215 -12895
rect 51335 -13015 51390 -12895
rect 51510 -13015 51555 -12895
rect 51675 -13015 51720 -12895
rect 51840 -13015 51885 -12895
rect 52005 -13015 52060 -12895
rect 52180 -13015 52225 -12895
rect 52345 -13015 52390 -12895
rect 52510 -13015 52555 -12895
rect 52675 -13015 52730 -12895
rect 52850 -13015 52895 -12895
rect 53015 -13015 53060 -12895
rect 53180 -13015 53225 -12895
rect 53345 -13015 53370 -12895
rect 30770 -13060 53370 -13015
rect 30770 -13180 30795 -13060
rect 30915 -13180 30970 -13060
rect 31090 -13180 31135 -13060
rect 31255 -13180 31300 -13060
rect 31420 -13180 31465 -13060
rect 31585 -13180 31640 -13060
rect 31760 -13180 31805 -13060
rect 31925 -13180 31970 -13060
rect 32090 -13180 32135 -13060
rect 32255 -13180 32310 -13060
rect 32430 -13180 32475 -13060
rect 32595 -13180 32640 -13060
rect 32760 -13180 32805 -13060
rect 32925 -13180 32980 -13060
rect 33100 -13180 33145 -13060
rect 33265 -13180 33310 -13060
rect 33430 -13180 33475 -13060
rect 33595 -13180 33650 -13060
rect 33770 -13180 33815 -13060
rect 33935 -13180 33980 -13060
rect 34100 -13180 34145 -13060
rect 34265 -13180 34320 -13060
rect 34440 -13180 34485 -13060
rect 34605 -13180 34650 -13060
rect 34770 -13180 34815 -13060
rect 34935 -13180 34990 -13060
rect 35110 -13180 35155 -13060
rect 35275 -13180 35320 -13060
rect 35440 -13180 35485 -13060
rect 35605 -13180 35660 -13060
rect 35780 -13180 35825 -13060
rect 35945 -13180 35990 -13060
rect 36110 -13180 36155 -13060
rect 36275 -13180 36485 -13060
rect 36605 -13180 36660 -13060
rect 36780 -13180 36825 -13060
rect 36945 -13180 36990 -13060
rect 37110 -13180 37155 -13060
rect 37275 -13180 37330 -13060
rect 37450 -13180 37495 -13060
rect 37615 -13180 37660 -13060
rect 37780 -13180 37825 -13060
rect 37945 -13180 38000 -13060
rect 38120 -13180 38165 -13060
rect 38285 -13180 38330 -13060
rect 38450 -13180 38495 -13060
rect 38615 -13180 38670 -13060
rect 38790 -13180 38835 -13060
rect 38955 -13180 39000 -13060
rect 39120 -13180 39165 -13060
rect 39285 -13180 39340 -13060
rect 39460 -13180 39505 -13060
rect 39625 -13180 39670 -13060
rect 39790 -13180 39835 -13060
rect 39955 -13180 40010 -13060
rect 40130 -13180 40175 -13060
rect 40295 -13180 40340 -13060
rect 40460 -13180 40505 -13060
rect 40625 -13180 40680 -13060
rect 40800 -13180 40845 -13060
rect 40965 -13180 41010 -13060
rect 41130 -13180 41175 -13060
rect 41295 -13180 41350 -13060
rect 41470 -13180 41515 -13060
rect 41635 -13180 41680 -13060
rect 41800 -13180 41845 -13060
rect 41965 -13180 42175 -13060
rect 42295 -13180 42350 -13060
rect 42470 -13180 42515 -13060
rect 42635 -13180 42680 -13060
rect 42800 -13180 42845 -13060
rect 42965 -13180 43020 -13060
rect 43140 -13180 43185 -13060
rect 43305 -13180 43350 -13060
rect 43470 -13180 43515 -13060
rect 43635 -13180 43690 -13060
rect 43810 -13180 43855 -13060
rect 43975 -13180 44020 -13060
rect 44140 -13180 44185 -13060
rect 44305 -13180 44360 -13060
rect 44480 -13180 44525 -13060
rect 44645 -13180 44690 -13060
rect 44810 -13180 44855 -13060
rect 44975 -13180 45030 -13060
rect 45150 -13180 45195 -13060
rect 45315 -13180 45360 -13060
rect 45480 -13180 45525 -13060
rect 45645 -13180 45700 -13060
rect 45820 -13180 45865 -13060
rect 45985 -13180 46030 -13060
rect 46150 -13180 46195 -13060
rect 46315 -13180 46370 -13060
rect 46490 -13180 46535 -13060
rect 46655 -13180 46700 -13060
rect 46820 -13180 46865 -13060
rect 46985 -13180 47040 -13060
rect 47160 -13180 47205 -13060
rect 47325 -13180 47370 -13060
rect 47490 -13180 47535 -13060
rect 47655 -13180 47865 -13060
rect 47985 -13180 48040 -13060
rect 48160 -13180 48205 -13060
rect 48325 -13180 48370 -13060
rect 48490 -13180 48535 -13060
rect 48655 -13180 48710 -13060
rect 48830 -13180 48875 -13060
rect 48995 -13180 49040 -13060
rect 49160 -13180 49205 -13060
rect 49325 -13180 49380 -13060
rect 49500 -13180 49545 -13060
rect 49665 -13180 49710 -13060
rect 49830 -13180 49875 -13060
rect 49995 -13180 50050 -13060
rect 50170 -13180 50215 -13060
rect 50335 -13180 50380 -13060
rect 50500 -13180 50545 -13060
rect 50665 -13180 50720 -13060
rect 50840 -13180 50885 -13060
rect 51005 -13180 51050 -13060
rect 51170 -13180 51215 -13060
rect 51335 -13180 51390 -13060
rect 51510 -13180 51555 -13060
rect 51675 -13180 51720 -13060
rect 51840 -13180 51885 -13060
rect 52005 -13180 52060 -13060
rect 52180 -13180 52225 -13060
rect 52345 -13180 52390 -13060
rect 52510 -13180 52555 -13060
rect 52675 -13180 52730 -13060
rect 52850 -13180 52895 -13060
rect 53015 -13180 53060 -13060
rect 53180 -13180 53225 -13060
rect 53345 -13180 53370 -13060
rect 30770 -13225 53370 -13180
rect 30770 -13345 30795 -13225
rect 30915 -13345 30970 -13225
rect 31090 -13345 31135 -13225
rect 31255 -13345 31300 -13225
rect 31420 -13345 31465 -13225
rect 31585 -13345 31640 -13225
rect 31760 -13345 31805 -13225
rect 31925 -13345 31970 -13225
rect 32090 -13345 32135 -13225
rect 32255 -13345 32310 -13225
rect 32430 -13345 32475 -13225
rect 32595 -13345 32640 -13225
rect 32760 -13345 32805 -13225
rect 32925 -13345 32980 -13225
rect 33100 -13345 33145 -13225
rect 33265 -13345 33310 -13225
rect 33430 -13345 33475 -13225
rect 33595 -13345 33650 -13225
rect 33770 -13345 33815 -13225
rect 33935 -13345 33980 -13225
rect 34100 -13345 34145 -13225
rect 34265 -13345 34320 -13225
rect 34440 -13345 34485 -13225
rect 34605 -13345 34650 -13225
rect 34770 -13345 34815 -13225
rect 34935 -13345 34990 -13225
rect 35110 -13345 35155 -13225
rect 35275 -13345 35320 -13225
rect 35440 -13345 35485 -13225
rect 35605 -13345 35660 -13225
rect 35780 -13345 35825 -13225
rect 35945 -13345 35990 -13225
rect 36110 -13345 36155 -13225
rect 36275 -13345 36485 -13225
rect 36605 -13345 36660 -13225
rect 36780 -13345 36825 -13225
rect 36945 -13345 36990 -13225
rect 37110 -13345 37155 -13225
rect 37275 -13345 37330 -13225
rect 37450 -13345 37495 -13225
rect 37615 -13345 37660 -13225
rect 37780 -13345 37825 -13225
rect 37945 -13345 38000 -13225
rect 38120 -13345 38165 -13225
rect 38285 -13345 38330 -13225
rect 38450 -13345 38495 -13225
rect 38615 -13345 38670 -13225
rect 38790 -13345 38835 -13225
rect 38955 -13345 39000 -13225
rect 39120 -13345 39165 -13225
rect 39285 -13345 39340 -13225
rect 39460 -13345 39505 -13225
rect 39625 -13345 39670 -13225
rect 39790 -13345 39835 -13225
rect 39955 -13345 40010 -13225
rect 40130 -13345 40175 -13225
rect 40295 -13345 40340 -13225
rect 40460 -13345 40505 -13225
rect 40625 -13345 40680 -13225
rect 40800 -13345 40845 -13225
rect 40965 -13345 41010 -13225
rect 41130 -13345 41175 -13225
rect 41295 -13345 41350 -13225
rect 41470 -13345 41515 -13225
rect 41635 -13345 41680 -13225
rect 41800 -13345 41845 -13225
rect 41965 -13345 42175 -13225
rect 42295 -13345 42350 -13225
rect 42470 -13345 42515 -13225
rect 42635 -13345 42680 -13225
rect 42800 -13345 42845 -13225
rect 42965 -13345 43020 -13225
rect 43140 -13345 43185 -13225
rect 43305 -13345 43350 -13225
rect 43470 -13345 43515 -13225
rect 43635 -13345 43690 -13225
rect 43810 -13345 43855 -13225
rect 43975 -13345 44020 -13225
rect 44140 -13345 44185 -13225
rect 44305 -13345 44360 -13225
rect 44480 -13345 44525 -13225
rect 44645 -13345 44690 -13225
rect 44810 -13345 44855 -13225
rect 44975 -13345 45030 -13225
rect 45150 -13345 45195 -13225
rect 45315 -13345 45360 -13225
rect 45480 -13345 45525 -13225
rect 45645 -13345 45700 -13225
rect 45820 -13345 45865 -13225
rect 45985 -13345 46030 -13225
rect 46150 -13345 46195 -13225
rect 46315 -13345 46370 -13225
rect 46490 -13345 46535 -13225
rect 46655 -13345 46700 -13225
rect 46820 -13345 46865 -13225
rect 46985 -13345 47040 -13225
rect 47160 -13345 47205 -13225
rect 47325 -13345 47370 -13225
rect 47490 -13345 47535 -13225
rect 47655 -13345 47865 -13225
rect 47985 -13345 48040 -13225
rect 48160 -13345 48205 -13225
rect 48325 -13345 48370 -13225
rect 48490 -13345 48535 -13225
rect 48655 -13345 48710 -13225
rect 48830 -13345 48875 -13225
rect 48995 -13345 49040 -13225
rect 49160 -13345 49205 -13225
rect 49325 -13345 49380 -13225
rect 49500 -13345 49545 -13225
rect 49665 -13345 49710 -13225
rect 49830 -13345 49875 -13225
rect 49995 -13345 50050 -13225
rect 50170 -13345 50215 -13225
rect 50335 -13345 50380 -13225
rect 50500 -13345 50545 -13225
rect 50665 -13345 50720 -13225
rect 50840 -13345 50885 -13225
rect 51005 -13345 51050 -13225
rect 51170 -13345 51215 -13225
rect 51335 -13345 51390 -13225
rect 51510 -13345 51555 -13225
rect 51675 -13345 51720 -13225
rect 51840 -13345 51885 -13225
rect 52005 -13345 52060 -13225
rect 52180 -13345 52225 -13225
rect 52345 -13345 52390 -13225
rect 52510 -13345 52555 -13225
rect 52675 -13345 52730 -13225
rect 52850 -13345 52895 -13225
rect 53015 -13345 53060 -13225
rect 53180 -13345 53225 -13225
rect 53345 -13345 53370 -13225
rect 30770 -13400 53370 -13345
rect 30770 -13520 30795 -13400
rect 30915 -13520 30970 -13400
rect 31090 -13520 31135 -13400
rect 31255 -13520 31300 -13400
rect 31420 -13520 31465 -13400
rect 31585 -13520 31640 -13400
rect 31760 -13520 31805 -13400
rect 31925 -13520 31970 -13400
rect 32090 -13520 32135 -13400
rect 32255 -13520 32310 -13400
rect 32430 -13520 32475 -13400
rect 32595 -13520 32640 -13400
rect 32760 -13520 32805 -13400
rect 32925 -13520 32980 -13400
rect 33100 -13520 33145 -13400
rect 33265 -13520 33310 -13400
rect 33430 -13520 33475 -13400
rect 33595 -13520 33650 -13400
rect 33770 -13520 33815 -13400
rect 33935 -13520 33980 -13400
rect 34100 -13520 34145 -13400
rect 34265 -13520 34320 -13400
rect 34440 -13520 34485 -13400
rect 34605 -13520 34650 -13400
rect 34770 -13520 34815 -13400
rect 34935 -13520 34990 -13400
rect 35110 -13520 35155 -13400
rect 35275 -13520 35320 -13400
rect 35440 -13520 35485 -13400
rect 35605 -13520 35660 -13400
rect 35780 -13520 35825 -13400
rect 35945 -13520 35990 -13400
rect 36110 -13520 36155 -13400
rect 36275 -13520 36485 -13400
rect 36605 -13520 36660 -13400
rect 36780 -13520 36825 -13400
rect 36945 -13520 36990 -13400
rect 37110 -13520 37155 -13400
rect 37275 -13520 37330 -13400
rect 37450 -13520 37495 -13400
rect 37615 -13520 37660 -13400
rect 37780 -13520 37825 -13400
rect 37945 -13520 38000 -13400
rect 38120 -13520 38165 -13400
rect 38285 -13520 38330 -13400
rect 38450 -13520 38495 -13400
rect 38615 -13520 38670 -13400
rect 38790 -13520 38835 -13400
rect 38955 -13520 39000 -13400
rect 39120 -13520 39165 -13400
rect 39285 -13520 39340 -13400
rect 39460 -13520 39505 -13400
rect 39625 -13520 39670 -13400
rect 39790 -13520 39835 -13400
rect 39955 -13520 40010 -13400
rect 40130 -13520 40175 -13400
rect 40295 -13520 40340 -13400
rect 40460 -13520 40505 -13400
rect 40625 -13520 40680 -13400
rect 40800 -13520 40845 -13400
rect 40965 -13520 41010 -13400
rect 41130 -13520 41175 -13400
rect 41295 -13520 41350 -13400
rect 41470 -13520 41515 -13400
rect 41635 -13520 41680 -13400
rect 41800 -13520 41845 -13400
rect 41965 -13520 42175 -13400
rect 42295 -13520 42350 -13400
rect 42470 -13520 42515 -13400
rect 42635 -13520 42680 -13400
rect 42800 -13520 42845 -13400
rect 42965 -13520 43020 -13400
rect 43140 -13520 43185 -13400
rect 43305 -13520 43350 -13400
rect 43470 -13520 43515 -13400
rect 43635 -13520 43690 -13400
rect 43810 -13520 43855 -13400
rect 43975 -13520 44020 -13400
rect 44140 -13520 44185 -13400
rect 44305 -13520 44360 -13400
rect 44480 -13520 44525 -13400
rect 44645 -13520 44690 -13400
rect 44810 -13520 44855 -13400
rect 44975 -13520 45030 -13400
rect 45150 -13520 45195 -13400
rect 45315 -13520 45360 -13400
rect 45480 -13520 45525 -13400
rect 45645 -13520 45700 -13400
rect 45820 -13520 45865 -13400
rect 45985 -13520 46030 -13400
rect 46150 -13520 46195 -13400
rect 46315 -13520 46370 -13400
rect 46490 -13520 46535 -13400
rect 46655 -13520 46700 -13400
rect 46820 -13520 46865 -13400
rect 46985 -13520 47040 -13400
rect 47160 -13520 47205 -13400
rect 47325 -13520 47370 -13400
rect 47490 -13520 47535 -13400
rect 47655 -13520 47865 -13400
rect 47985 -13520 48040 -13400
rect 48160 -13520 48205 -13400
rect 48325 -13520 48370 -13400
rect 48490 -13520 48535 -13400
rect 48655 -13520 48710 -13400
rect 48830 -13520 48875 -13400
rect 48995 -13520 49040 -13400
rect 49160 -13520 49205 -13400
rect 49325 -13520 49380 -13400
rect 49500 -13520 49545 -13400
rect 49665 -13520 49710 -13400
rect 49830 -13520 49875 -13400
rect 49995 -13520 50050 -13400
rect 50170 -13520 50215 -13400
rect 50335 -13520 50380 -13400
rect 50500 -13520 50545 -13400
rect 50665 -13520 50720 -13400
rect 50840 -13520 50885 -13400
rect 51005 -13520 51050 -13400
rect 51170 -13520 51215 -13400
rect 51335 -13520 51390 -13400
rect 51510 -13520 51555 -13400
rect 51675 -13520 51720 -13400
rect 51840 -13520 51885 -13400
rect 52005 -13520 52060 -13400
rect 52180 -13520 52225 -13400
rect 52345 -13520 52390 -13400
rect 52510 -13520 52555 -13400
rect 52675 -13520 52730 -13400
rect 52850 -13520 52895 -13400
rect 53015 -13520 53060 -13400
rect 53180 -13520 53225 -13400
rect 53345 -13520 53370 -13400
rect 30770 -13565 53370 -13520
rect 30770 -13685 30795 -13565
rect 30915 -13685 30970 -13565
rect 31090 -13685 31135 -13565
rect 31255 -13685 31300 -13565
rect 31420 -13685 31465 -13565
rect 31585 -13685 31640 -13565
rect 31760 -13685 31805 -13565
rect 31925 -13685 31970 -13565
rect 32090 -13685 32135 -13565
rect 32255 -13685 32310 -13565
rect 32430 -13685 32475 -13565
rect 32595 -13685 32640 -13565
rect 32760 -13685 32805 -13565
rect 32925 -13685 32980 -13565
rect 33100 -13685 33145 -13565
rect 33265 -13685 33310 -13565
rect 33430 -13685 33475 -13565
rect 33595 -13685 33650 -13565
rect 33770 -13685 33815 -13565
rect 33935 -13685 33980 -13565
rect 34100 -13685 34145 -13565
rect 34265 -13685 34320 -13565
rect 34440 -13685 34485 -13565
rect 34605 -13685 34650 -13565
rect 34770 -13685 34815 -13565
rect 34935 -13685 34990 -13565
rect 35110 -13685 35155 -13565
rect 35275 -13685 35320 -13565
rect 35440 -13685 35485 -13565
rect 35605 -13685 35660 -13565
rect 35780 -13685 35825 -13565
rect 35945 -13685 35990 -13565
rect 36110 -13685 36155 -13565
rect 36275 -13685 36485 -13565
rect 36605 -13685 36660 -13565
rect 36780 -13685 36825 -13565
rect 36945 -13685 36990 -13565
rect 37110 -13685 37155 -13565
rect 37275 -13685 37330 -13565
rect 37450 -13685 37495 -13565
rect 37615 -13685 37660 -13565
rect 37780 -13685 37825 -13565
rect 37945 -13685 38000 -13565
rect 38120 -13685 38165 -13565
rect 38285 -13685 38330 -13565
rect 38450 -13685 38495 -13565
rect 38615 -13685 38670 -13565
rect 38790 -13685 38835 -13565
rect 38955 -13685 39000 -13565
rect 39120 -13685 39165 -13565
rect 39285 -13685 39340 -13565
rect 39460 -13685 39505 -13565
rect 39625 -13685 39670 -13565
rect 39790 -13685 39835 -13565
rect 39955 -13685 40010 -13565
rect 40130 -13685 40175 -13565
rect 40295 -13685 40340 -13565
rect 40460 -13685 40505 -13565
rect 40625 -13685 40680 -13565
rect 40800 -13685 40845 -13565
rect 40965 -13685 41010 -13565
rect 41130 -13685 41175 -13565
rect 41295 -13685 41350 -13565
rect 41470 -13685 41515 -13565
rect 41635 -13685 41680 -13565
rect 41800 -13685 41845 -13565
rect 41965 -13685 42175 -13565
rect 42295 -13685 42350 -13565
rect 42470 -13685 42515 -13565
rect 42635 -13685 42680 -13565
rect 42800 -13685 42845 -13565
rect 42965 -13685 43020 -13565
rect 43140 -13685 43185 -13565
rect 43305 -13685 43350 -13565
rect 43470 -13685 43515 -13565
rect 43635 -13685 43690 -13565
rect 43810 -13685 43855 -13565
rect 43975 -13685 44020 -13565
rect 44140 -13685 44185 -13565
rect 44305 -13685 44360 -13565
rect 44480 -13685 44525 -13565
rect 44645 -13685 44690 -13565
rect 44810 -13685 44855 -13565
rect 44975 -13685 45030 -13565
rect 45150 -13685 45195 -13565
rect 45315 -13685 45360 -13565
rect 45480 -13685 45525 -13565
rect 45645 -13685 45700 -13565
rect 45820 -13685 45865 -13565
rect 45985 -13685 46030 -13565
rect 46150 -13685 46195 -13565
rect 46315 -13685 46370 -13565
rect 46490 -13685 46535 -13565
rect 46655 -13685 46700 -13565
rect 46820 -13685 46865 -13565
rect 46985 -13685 47040 -13565
rect 47160 -13685 47205 -13565
rect 47325 -13685 47370 -13565
rect 47490 -13685 47535 -13565
rect 47655 -13685 47865 -13565
rect 47985 -13685 48040 -13565
rect 48160 -13685 48205 -13565
rect 48325 -13685 48370 -13565
rect 48490 -13685 48535 -13565
rect 48655 -13685 48710 -13565
rect 48830 -13685 48875 -13565
rect 48995 -13685 49040 -13565
rect 49160 -13685 49205 -13565
rect 49325 -13685 49380 -13565
rect 49500 -13685 49545 -13565
rect 49665 -13685 49710 -13565
rect 49830 -13685 49875 -13565
rect 49995 -13685 50050 -13565
rect 50170 -13685 50215 -13565
rect 50335 -13685 50380 -13565
rect 50500 -13685 50545 -13565
rect 50665 -13685 50720 -13565
rect 50840 -13685 50885 -13565
rect 51005 -13685 51050 -13565
rect 51170 -13685 51215 -13565
rect 51335 -13685 51390 -13565
rect 51510 -13685 51555 -13565
rect 51675 -13685 51720 -13565
rect 51840 -13685 51885 -13565
rect 52005 -13685 52060 -13565
rect 52180 -13685 52225 -13565
rect 52345 -13685 52390 -13565
rect 52510 -13685 52555 -13565
rect 52675 -13685 52730 -13565
rect 52850 -13685 52895 -13565
rect 53015 -13685 53060 -13565
rect 53180 -13685 53225 -13565
rect 53345 -13685 53370 -13565
rect 30770 -13730 53370 -13685
rect 30770 -13850 30795 -13730
rect 30915 -13850 30970 -13730
rect 31090 -13850 31135 -13730
rect 31255 -13850 31300 -13730
rect 31420 -13850 31465 -13730
rect 31585 -13850 31640 -13730
rect 31760 -13850 31805 -13730
rect 31925 -13850 31970 -13730
rect 32090 -13850 32135 -13730
rect 32255 -13850 32310 -13730
rect 32430 -13850 32475 -13730
rect 32595 -13850 32640 -13730
rect 32760 -13850 32805 -13730
rect 32925 -13850 32980 -13730
rect 33100 -13850 33145 -13730
rect 33265 -13850 33310 -13730
rect 33430 -13850 33475 -13730
rect 33595 -13850 33650 -13730
rect 33770 -13850 33815 -13730
rect 33935 -13850 33980 -13730
rect 34100 -13850 34145 -13730
rect 34265 -13850 34320 -13730
rect 34440 -13850 34485 -13730
rect 34605 -13850 34650 -13730
rect 34770 -13850 34815 -13730
rect 34935 -13850 34990 -13730
rect 35110 -13850 35155 -13730
rect 35275 -13850 35320 -13730
rect 35440 -13850 35485 -13730
rect 35605 -13850 35660 -13730
rect 35780 -13850 35825 -13730
rect 35945 -13850 35990 -13730
rect 36110 -13850 36155 -13730
rect 36275 -13850 36485 -13730
rect 36605 -13850 36660 -13730
rect 36780 -13850 36825 -13730
rect 36945 -13850 36990 -13730
rect 37110 -13850 37155 -13730
rect 37275 -13850 37330 -13730
rect 37450 -13850 37495 -13730
rect 37615 -13850 37660 -13730
rect 37780 -13850 37825 -13730
rect 37945 -13850 38000 -13730
rect 38120 -13850 38165 -13730
rect 38285 -13850 38330 -13730
rect 38450 -13850 38495 -13730
rect 38615 -13850 38670 -13730
rect 38790 -13850 38835 -13730
rect 38955 -13850 39000 -13730
rect 39120 -13850 39165 -13730
rect 39285 -13850 39340 -13730
rect 39460 -13850 39505 -13730
rect 39625 -13850 39670 -13730
rect 39790 -13850 39835 -13730
rect 39955 -13850 40010 -13730
rect 40130 -13850 40175 -13730
rect 40295 -13850 40340 -13730
rect 40460 -13850 40505 -13730
rect 40625 -13850 40680 -13730
rect 40800 -13850 40845 -13730
rect 40965 -13850 41010 -13730
rect 41130 -13850 41175 -13730
rect 41295 -13850 41350 -13730
rect 41470 -13850 41515 -13730
rect 41635 -13850 41680 -13730
rect 41800 -13850 41845 -13730
rect 41965 -13850 42175 -13730
rect 42295 -13850 42350 -13730
rect 42470 -13850 42515 -13730
rect 42635 -13850 42680 -13730
rect 42800 -13850 42845 -13730
rect 42965 -13850 43020 -13730
rect 43140 -13850 43185 -13730
rect 43305 -13850 43350 -13730
rect 43470 -13850 43515 -13730
rect 43635 -13850 43690 -13730
rect 43810 -13850 43855 -13730
rect 43975 -13850 44020 -13730
rect 44140 -13850 44185 -13730
rect 44305 -13850 44360 -13730
rect 44480 -13850 44525 -13730
rect 44645 -13850 44690 -13730
rect 44810 -13850 44855 -13730
rect 44975 -13850 45030 -13730
rect 45150 -13850 45195 -13730
rect 45315 -13850 45360 -13730
rect 45480 -13850 45525 -13730
rect 45645 -13850 45700 -13730
rect 45820 -13850 45865 -13730
rect 45985 -13850 46030 -13730
rect 46150 -13850 46195 -13730
rect 46315 -13850 46370 -13730
rect 46490 -13850 46535 -13730
rect 46655 -13850 46700 -13730
rect 46820 -13850 46865 -13730
rect 46985 -13850 47040 -13730
rect 47160 -13850 47205 -13730
rect 47325 -13850 47370 -13730
rect 47490 -13850 47535 -13730
rect 47655 -13850 47865 -13730
rect 47985 -13850 48040 -13730
rect 48160 -13850 48205 -13730
rect 48325 -13850 48370 -13730
rect 48490 -13850 48535 -13730
rect 48655 -13850 48710 -13730
rect 48830 -13850 48875 -13730
rect 48995 -13850 49040 -13730
rect 49160 -13850 49205 -13730
rect 49325 -13850 49380 -13730
rect 49500 -13850 49545 -13730
rect 49665 -13850 49710 -13730
rect 49830 -13850 49875 -13730
rect 49995 -13850 50050 -13730
rect 50170 -13850 50215 -13730
rect 50335 -13850 50380 -13730
rect 50500 -13850 50545 -13730
rect 50665 -13850 50720 -13730
rect 50840 -13850 50885 -13730
rect 51005 -13850 51050 -13730
rect 51170 -13850 51215 -13730
rect 51335 -13850 51390 -13730
rect 51510 -13850 51555 -13730
rect 51675 -13850 51720 -13730
rect 51840 -13850 51885 -13730
rect 52005 -13850 52060 -13730
rect 52180 -13850 52225 -13730
rect 52345 -13850 52390 -13730
rect 52510 -13850 52555 -13730
rect 52675 -13850 52730 -13730
rect 52850 -13850 52895 -13730
rect 53015 -13850 53060 -13730
rect 53180 -13850 53225 -13730
rect 53345 -13850 53370 -13730
rect 30770 -13895 53370 -13850
rect 30770 -14015 30795 -13895
rect 30915 -14015 30970 -13895
rect 31090 -14015 31135 -13895
rect 31255 -14015 31300 -13895
rect 31420 -14015 31465 -13895
rect 31585 -14015 31640 -13895
rect 31760 -14015 31805 -13895
rect 31925 -14015 31970 -13895
rect 32090 -14015 32135 -13895
rect 32255 -14015 32310 -13895
rect 32430 -14015 32475 -13895
rect 32595 -14015 32640 -13895
rect 32760 -14015 32805 -13895
rect 32925 -14015 32980 -13895
rect 33100 -14015 33145 -13895
rect 33265 -14015 33310 -13895
rect 33430 -14015 33475 -13895
rect 33595 -14015 33650 -13895
rect 33770 -14015 33815 -13895
rect 33935 -14015 33980 -13895
rect 34100 -14015 34145 -13895
rect 34265 -14015 34320 -13895
rect 34440 -14015 34485 -13895
rect 34605 -14015 34650 -13895
rect 34770 -14015 34815 -13895
rect 34935 -14015 34990 -13895
rect 35110 -14015 35155 -13895
rect 35275 -14015 35320 -13895
rect 35440 -14015 35485 -13895
rect 35605 -14015 35660 -13895
rect 35780 -14015 35825 -13895
rect 35945 -14015 35990 -13895
rect 36110 -14015 36155 -13895
rect 36275 -14015 36485 -13895
rect 36605 -14015 36660 -13895
rect 36780 -14015 36825 -13895
rect 36945 -14015 36990 -13895
rect 37110 -14015 37155 -13895
rect 37275 -14015 37330 -13895
rect 37450 -14015 37495 -13895
rect 37615 -14015 37660 -13895
rect 37780 -14015 37825 -13895
rect 37945 -14015 38000 -13895
rect 38120 -14015 38165 -13895
rect 38285 -14015 38330 -13895
rect 38450 -14015 38495 -13895
rect 38615 -14015 38670 -13895
rect 38790 -14015 38835 -13895
rect 38955 -14015 39000 -13895
rect 39120 -14015 39165 -13895
rect 39285 -14015 39340 -13895
rect 39460 -14015 39505 -13895
rect 39625 -14015 39670 -13895
rect 39790 -14015 39835 -13895
rect 39955 -14015 40010 -13895
rect 40130 -14015 40175 -13895
rect 40295 -14015 40340 -13895
rect 40460 -14015 40505 -13895
rect 40625 -14015 40680 -13895
rect 40800 -14015 40845 -13895
rect 40965 -14015 41010 -13895
rect 41130 -14015 41175 -13895
rect 41295 -14015 41350 -13895
rect 41470 -14015 41515 -13895
rect 41635 -14015 41680 -13895
rect 41800 -14015 41845 -13895
rect 41965 -14015 42175 -13895
rect 42295 -14015 42350 -13895
rect 42470 -14015 42515 -13895
rect 42635 -14015 42680 -13895
rect 42800 -14015 42845 -13895
rect 42965 -14015 43020 -13895
rect 43140 -14015 43185 -13895
rect 43305 -14015 43350 -13895
rect 43470 -14015 43515 -13895
rect 43635 -14015 43690 -13895
rect 43810 -14015 43855 -13895
rect 43975 -14015 44020 -13895
rect 44140 -14015 44185 -13895
rect 44305 -14015 44360 -13895
rect 44480 -14015 44525 -13895
rect 44645 -14015 44690 -13895
rect 44810 -14015 44855 -13895
rect 44975 -14015 45030 -13895
rect 45150 -14015 45195 -13895
rect 45315 -14015 45360 -13895
rect 45480 -14015 45525 -13895
rect 45645 -14015 45700 -13895
rect 45820 -14015 45865 -13895
rect 45985 -14015 46030 -13895
rect 46150 -14015 46195 -13895
rect 46315 -14015 46370 -13895
rect 46490 -14015 46535 -13895
rect 46655 -14015 46700 -13895
rect 46820 -14015 46865 -13895
rect 46985 -14015 47040 -13895
rect 47160 -14015 47205 -13895
rect 47325 -14015 47370 -13895
rect 47490 -14015 47535 -13895
rect 47655 -14015 47865 -13895
rect 47985 -14015 48040 -13895
rect 48160 -14015 48205 -13895
rect 48325 -14015 48370 -13895
rect 48490 -14015 48535 -13895
rect 48655 -14015 48710 -13895
rect 48830 -14015 48875 -13895
rect 48995 -14015 49040 -13895
rect 49160 -14015 49205 -13895
rect 49325 -14015 49380 -13895
rect 49500 -14015 49545 -13895
rect 49665 -14015 49710 -13895
rect 49830 -14015 49875 -13895
rect 49995 -14015 50050 -13895
rect 50170 -14015 50215 -13895
rect 50335 -14015 50380 -13895
rect 50500 -14015 50545 -13895
rect 50665 -14015 50720 -13895
rect 50840 -14015 50885 -13895
rect 51005 -14015 51050 -13895
rect 51170 -14015 51215 -13895
rect 51335 -14015 51390 -13895
rect 51510 -14015 51555 -13895
rect 51675 -14015 51720 -13895
rect 51840 -14015 51885 -13895
rect 52005 -14015 52060 -13895
rect 52180 -14015 52225 -13895
rect 52345 -14015 52390 -13895
rect 52510 -14015 52555 -13895
rect 52675 -14015 52730 -13895
rect 52850 -14015 52895 -13895
rect 53015 -14015 53060 -13895
rect 53180 -14015 53225 -13895
rect 53345 -14015 53370 -13895
rect 30770 -14070 53370 -14015
rect 30770 -14190 30795 -14070
rect 30915 -14190 30970 -14070
rect 31090 -14190 31135 -14070
rect 31255 -14190 31300 -14070
rect 31420 -14190 31465 -14070
rect 31585 -14190 31640 -14070
rect 31760 -14190 31805 -14070
rect 31925 -14190 31970 -14070
rect 32090 -14190 32135 -14070
rect 32255 -14190 32310 -14070
rect 32430 -14190 32475 -14070
rect 32595 -14190 32640 -14070
rect 32760 -14190 32805 -14070
rect 32925 -14190 32980 -14070
rect 33100 -14190 33145 -14070
rect 33265 -14190 33310 -14070
rect 33430 -14190 33475 -14070
rect 33595 -14190 33650 -14070
rect 33770 -14190 33815 -14070
rect 33935 -14190 33980 -14070
rect 34100 -14190 34145 -14070
rect 34265 -14190 34320 -14070
rect 34440 -14190 34485 -14070
rect 34605 -14190 34650 -14070
rect 34770 -14190 34815 -14070
rect 34935 -14190 34990 -14070
rect 35110 -14190 35155 -14070
rect 35275 -14190 35320 -14070
rect 35440 -14190 35485 -14070
rect 35605 -14190 35660 -14070
rect 35780 -14190 35825 -14070
rect 35945 -14190 35990 -14070
rect 36110 -14190 36155 -14070
rect 36275 -14190 36485 -14070
rect 36605 -14190 36660 -14070
rect 36780 -14190 36825 -14070
rect 36945 -14190 36990 -14070
rect 37110 -14190 37155 -14070
rect 37275 -14190 37330 -14070
rect 37450 -14190 37495 -14070
rect 37615 -14190 37660 -14070
rect 37780 -14190 37825 -14070
rect 37945 -14190 38000 -14070
rect 38120 -14190 38165 -14070
rect 38285 -14190 38330 -14070
rect 38450 -14190 38495 -14070
rect 38615 -14190 38670 -14070
rect 38790 -14190 38835 -14070
rect 38955 -14190 39000 -14070
rect 39120 -14190 39165 -14070
rect 39285 -14190 39340 -14070
rect 39460 -14190 39505 -14070
rect 39625 -14190 39670 -14070
rect 39790 -14190 39835 -14070
rect 39955 -14190 40010 -14070
rect 40130 -14190 40175 -14070
rect 40295 -14190 40340 -14070
rect 40460 -14190 40505 -14070
rect 40625 -14190 40680 -14070
rect 40800 -14190 40845 -14070
rect 40965 -14190 41010 -14070
rect 41130 -14190 41175 -14070
rect 41295 -14190 41350 -14070
rect 41470 -14190 41515 -14070
rect 41635 -14190 41680 -14070
rect 41800 -14190 41845 -14070
rect 41965 -14190 42175 -14070
rect 42295 -14190 42350 -14070
rect 42470 -14190 42515 -14070
rect 42635 -14190 42680 -14070
rect 42800 -14190 42845 -14070
rect 42965 -14190 43020 -14070
rect 43140 -14190 43185 -14070
rect 43305 -14190 43350 -14070
rect 43470 -14190 43515 -14070
rect 43635 -14190 43690 -14070
rect 43810 -14190 43855 -14070
rect 43975 -14190 44020 -14070
rect 44140 -14190 44185 -14070
rect 44305 -14190 44360 -14070
rect 44480 -14190 44525 -14070
rect 44645 -14190 44690 -14070
rect 44810 -14190 44855 -14070
rect 44975 -14190 45030 -14070
rect 45150 -14190 45195 -14070
rect 45315 -14190 45360 -14070
rect 45480 -14190 45525 -14070
rect 45645 -14190 45700 -14070
rect 45820 -14190 45865 -14070
rect 45985 -14190 46030 -14070
rect 46150 -14190 46195 -14070
rect 46315 -14190 46370 -14070
rect 46490 -14190 46535 -14070
rect 46655 -14190 46700 -14070
rect 46820 -14190 46865 -14070
rect 46985 -14190 47040 -14070
rect 47160 -14190 47205 -14070
rect 47325 -14190 47370 -14070
rect 47490 -14190 47535 -14070
rect 47655 -14190 47865 -14070
rect 47985 -14190 48040 -14070
rect 48160 -14190 48205 -14070
rect 48325 -14190 48370 -14070
rect 48490 -14190 48535 -14070
rect 48655 -14190 48710 -14070
rect 48830 -14190 48875 -14070
rect 48995 -14190 49040 -14070
rect 49160 -14190 49205 -14070
rect 49325 -14190 49380 -14070
rect 49500 -14190 49545 -14070
rect 49665 -14190 49710 -14070
rect 49830 -14190 49875 -14070
rect 49995 -14190 50050 -14070
rect 50170 -14190 50215 -14070
rect 50335 -14190 50380 -14070
rect 50500 -14190 50545 -14070
rect 50665 -14190 50720 -14070
rect 50840 -14190 50885 -14070
rect 51005 -14190 51050 -14070
rect 51170 -14190 51215 -14070
rect 51335 -14190 51390 -14070
rect 51510 -14190 51555 -14070
rect 51675 -14190 51720 -14070
rect 51840 -14190 51885 -14070
rect 52005 -14190 52060 -14070
rect 52180 -14190 52225 -14070
rect 52345 -14190 52390 -14070
rect 52510 -14190 52555 -14070
rect 52675 -14190 52730 -14070
rect 52850 -14190 52895 -14070
rect 53015 -14190 53060 -14070
rect 53180 -14190 53225 -14070
rect 53345 -14190 53370 -14070
rect 30770 -14235 53370 -14190
rect 30770 -14355 30795 -14235
rect 30915 -14355 30970 -14235
rect 31090 -14355 31135 -14235
rect 31255 -14355 31300 -14235
rect 31420 -14355 31465 -14235
rect 31585 -14355 31640 -14235
rect 31760 -14355 31805 -14235
rect 31925 -14355 31970 -14235
rect 32090 -14355 32135 -14235
rect 32255 -14355 32310 -14235
rect 32430 -14355 32475 -14235
rect 32595 -14355 32640 -14235
rect 32760 -14355 32805 -14235
rect 32925 -14355 32980 -14235
rect 33100 -14355 33145 -14235
rect 33265 -14355 33310 -14235
rect 33430 -14355 33475 -14235
rect 33595 -14355 33650 -14235
rect 33770 -14355 33815 -14235
rect 33935 -14355 33980 -14235
rect 34100 -14355 34145 -14235
rect 34265 -14355 34320 -14235
rect 34440 -14355 34485 -14235
rect 34605 -14355 34650 -14235
rect 34770 -14355 34815 -14235
rect 34935 -14355 34990 -14235
rect 35110 -14355 35155 -14235
rect 35275 -14355 35320 -14235
rect 35440 -14355 35485 -14235
rect 35605 -14355 35660 -14235
rect 35780 -14355 35825 -14235
rect 35945 -14355 35990 -14235
rect 36110 -14355 36155 -14235
rect 36275 -14355 36485 -14235
rect 36605 -14355 36660 -14235
rect 36780 -14355 36825 -14235
rect 36945 -14355 36990 -14235
rect 37110 -14355 37155 -14235
rect 37275 -14355 37330 -14235
rect 37450 -14355 37495 -14235
rect 37615 -14355 37660 -14235
rect 37780 -14355 37825 -14235
rect 37945 -14355 38000 -14235
rect 38120 -14355 38165 -14235
rect 38285 -14355 38330 -14235
rect 38450 -14355 38495 -14235
rect 38615 -14355 38670 -14235
rect 38790 -14355 38835 -14235
rect 38955 -14355 39000 -14235
rect 39120 -14355 39165 -14235
rect 39285 -14355 39340 -14235
rect 39460 -14355 39505 -14235
rect 39625 -14355 39670 -14235
rect 39790 -14355 39835 -14235
rect 39955 -14355 40010 -14235
rect 40130 -14355 40175 -14235
rect 40295 -14355 40340 -14235
rect 40460 -14355 40505 -14235
rect 40625 -14355 40680 -14235
rect 40800 -14355 40845 -14235
rect 40965 -14355 41010 -14235
rect 41130 -14355 41175 -14235
rect 41295 -14355 41350 -14235
rect 41470 -14355 41515 -14235
rect 41635 -14355 41680 -14235
rect 41800 -14355 41845 -14235
rect 41965 -14355 42175 -14235
rect 42295 -14355 42350 -14235
rect 42470 -14355 42515 -14235
rect 42635 -14355 42680 -14235
rect 42800 -14355 42845 -14235
rect 42965 -14355 43020 -14235
rect 43140 -14355 43185 -14235
rect 43305 -14355 43350 -14235
rect 43470 -14355 43515 -14235
rect 43635 -14355 43690 -14235
rect 43810 -14355 43855 -14235
rect 43975 -14355 44020 -14235
rect 44140 -14355 44185 -14235
rect 44305 -14355 44360 -14235
rect 44480 -14355 44525 -14235
rect 44645 -14355 44690 -14235
rect 44810 -14355 44855 -14235
rect 44975 -14355 45030 -14235
rect 45150 -14355 45195 -14235
rect 45315 -14355 45360 -14235
rect 45480 -14355 45525 -14235
rect 45645 -14355 45700 -14235
rect 45820 -14355 45865 -14235
rect 45985 -14355 46030 -14235
rect 46150 -14355 46195 -14235
rect 46315 -14355 46370 -14235
rect 46490 -14355 46535 -14235
rect 46655 -14355 46700 -14235
rect 46820 -14355 46865 -14235
rect 46985 -14355 47040 -14235
rect 47160 -14355 47205 -14235
rect 47325 -14355 47370 -14235
rect 47490 -14355 47535 -14235
rect 47655 -14355 47865 -14235
rect 47985 -14355 48040 -14235
rect 48160 -14355 48205 -14235
rect 48325 -14355 48370 -14235
rect 48490 -14355 48535 -14235
rect 48655 -14355 48710 -14235
rect 48830 -14355 48875 -14235
rect 48995 -14355 49040 -14235
rect 49160 -14355 49205 -14235
rect 49325 -14355 49380 -14235
rect 49500 -14355 49545 -14235
rect 49665 -14355 49710 -14235
rect 49830 -14355 49875 -14235
rect 49995 -14355 50050 -14235
rect 50170 -14355 50215 -14235
rect 50335 -14355 50380 -14235
rect 50500 -14355 50545 -14235
rect 50665 -14355 50720 -14235
rect 50840 -14355 50885 -14235
rect 51005 -14355 51050 -14235
rect 51170 -14355 51215 -14235
rect 51335 -14355 51390 -14235
rect 51510 -14355 51555 -14235
rect 51675 -14355 51720 -14235
rect 51840 -14355 51885 -14235
rect 52005 -14355 52060 -14235
rect 52180 -14355 52225 -14235
rect 52345 -14355 52390 -14235
rect 52510 -14355 52555 -14235
rect 52675 -14355 52730 -14235
rect 52850 -14355 52895 -14235
rect 53015 -14355 53060 -14235
rect 53180 -14355 53225 -14235
rect 53345 -14355 53370 -14235
rect 30770 -14400 53370 -14355
rect 30770 -14520 30795 -14400
rect 30915 -14520 30970 -14400
rect 31090 -14520 31135 -14400
rect 31255 -14520 31300 -14400
rect 31420 -14520 31465 -14400
rect 31585 -14520 31640 -14400
rect 31760 -14520 31805 -14400
rect 31925 -14520 31970 -14400
rect 32090 -14520 32135 -14400
rect 32255 -14520 32310 -14400
rect 32430 -14520 32475 -14400
rect 32595 -14520 32640 -14400
rect 32760 -14520 32805 -14400
rect 32925 -14520 32980 -14400
rect 33100 -14520 33145 -14400
rect 33265 -14520 33310 -14400
rect 33430 -14520 33475 -14400
rect 33595 -14520 33650 -14400
rect 33770 -14520 33815 -14400
rect 33935 -14520 33980 -14400
rect 34100 -14520 34145 -14400
rect 34265 -14520 34320 -14400
rect 34440 -14520 34485 -14400
rect 34605 -14520 34650 -14400
rect 34770 -14520 34815 -14400
rect 34935 -14520 34990 -14400
rect 35110 -14520 35155 -14400
rect 35275 -14520 35320 -14400
rect 35440 -14520 35485 -14400
rect 35605 -14520 35660 -14400
rect 35780 -14520 35825 -14400
rect 35945 -14520 35990 -14400
rect 36110 -14520 36155 -14400
rect 36275 -14520 36485 -14400
rect 36605 -14520 36660 -14400
rect 36780 -14520 36825 -14400
rect 36945 -14520 36990 -14400
rect 37110 -14520 37155 -14400
rect 37275 -14520 37330 -14400
rect 37450 -14520 37495 -14400
rect 37615 -14520 37660 -14400
rect 37780 -14520 37825 -14400
rect 37945 -14520 38000 -14400
rect 38120 -14520 38165 -14400
rect 38285 -14520 38330 -14400
rect 38450 -14520 38495 -14400
rect 38615 -14520 38670 -14400
rect 38790 -14520 38835 -14400
rect 38955 -14520 39000 -14400
rect 39120 -14520 39165 -14400
rect 39285 -14520 39340 -14400
rect 39460 -14520 39505 -14400
rect 39625 -14520 39670 -14400
rect 39790 -14520 39835 -14400
rect 39955 -14520 40010 -14400
rect 40130 -14520 40175 -14400
rect 40295 -14520 40340 -14400
rect 40460 -14520 40505 -14400
rect 40625 -14520 40680 -14400
rect 40800 -14520 40845 -14400
rect 40965 -14520 41010 -14400
rect 41130 -14520 41175 -14400
rect 41295 -14520 41350 -14400
rect 41470 -14520 41515 -14400
rect 41635 -14520 41680 -14400
rect 41800 -14520 41845 -14400
rect 41965 -14520 42175 -14400
rect 42295 -14520 42350 -14400
rect 42470 -14520 42515 -14400
rect 42635 -14520 42680 -14400
rect 42800 -14520 42845 -14400
rect 42965 -14520 43020 -14400
rect 43140 -14520 43185 -14400
rect 43305 -14520 43350 -14400
rect 43470 -14520 43515 -14400
rect 43635 -14520 43690 -14400
rect 43810 -14520 43855 -14400
rect 43975 -14520 44020 -14400
rect 44140 -14520 44185 -14400
rect 44305 -14520 44360 -14400
rect 44480 -14520 44525 -14400
rect 44645 -14520 44690 -14400
rect 44810 -14520 44855 -14400
rect 44975 -14520 45030 -14400
rect 45150 -14520 45195 -14400
rect 45315 -14520 45360 -14400
rect 45480 -14520 45525 -14400
rect 45645 -14520 45700 -14400
rect 45820 -14520 45865 -14400
rect 45985 -14520 46030 -14400
rect 46150 -14520 46195 -14400
rect 46315 -14520 46370 -14400
rect 46490 -14520 46535 -14400
rect 46655 -14520 46700 -14400
rect 46820 -14520 46865 -14400
rect 46985 -14520 47040 -14400
rect 47160 -14520 47205 -14400
rect 47325 -14520 47370 -14400
rect 47490 -14520 47535 -14400
rect 47655 -14520 47865 -14400
rect 47985 -14520 48040 -14400
rect 48160 -14520 48205 -14400
rect 48325 -14520 48370 -14400
rect 48490 -14520 48535 -14400
rect 48655 -14520 48710 -14400
rect 48830 -14520 48875 -14400
rect 48995 -14520 49040 -14400
rect 49160 -14520 49205 -14400
rect 49325 -14520 49380 -14400
rect 49500 -14520 49545 -14400
rect 49665 -14520 49710 -14400
rect 49830 -14520 49875 -14400
rect 49995 -14520 50050 -14400
rect 50170 -14520 50215 -14400
rect 50335 -14520 50380 -14400
rect 50500 -14520 50545 -14400
rect 50665 -14520 50720 -14400
rect 50840 -14520 50885 -14400
rect 51005 -14520 51050 -14400
rect 51170 -14520 51215 -14400
rect 51335 -14520 51390 -14400
rect 51510 -14520 51555 -14400
rect 51675 -14520 51720 -14400
rect 51840 -14520 51885 -14400
rect 52005 -14520 52060 -14400
rect 52180 -14520 52225 -14400
rect 52345 -14520 52390 -14400
rect 52510 -14520 52555 -14400
rect 52675 -14520 52730 -14400
rect 52850 -14520 52895 -14400
rect 53015 -14520 53060 -14400
rect 53180 -14520 53225 -14400
rect 53345 -14520 53370 -14400
rect 30770 -14565 53370 -14520
rect 30770 -14685 30795 -14565
rect 30915 -14685 30970 -14565
rect 31090 -14685 31135 -14565
rect 31255 -14685 31300 -14565
rect 31420 -14685 31465 -14565
rect 31585 -14685 31640 -14565
rect 31760 -14685 31805 -14565
rect 31925 -14685 31970 -14565
rect 32090 -14685 32135 -14565
rect 32255 -14685 32310 -14565
rect 32430 -14685 32475 -14565
rect 32595 -14685 32640 -14565
rect 32760 -14685 32805 -14565
rect 32925 -14685 32980 -14565
rect 33100 -14685 33145 -14565
rect 33265 -14685 33310 -14565
rect 33430 -14685 33475 -14565
rect 33595 -14685 33650 -14565
rect 33770 -14685 33815 -14565
rect 33935 -14685 33980 -14565
rect 34100 -14685 34145 -14565
rect 34265 -14685 34320 -14565
rect 34440 -14685 34485 -14565
rect 34605 -14685 34650 -14565
rect 34770 -14685 34815 -14565
rect 34935 -14685 34990 -14565
rect 35110 -14685 35155 -14565
rect 35275 -14685 35320 -14565
rect 35440 -14685 35485 -14565
rect 35605 -14685 35660 -14565
rect 35780 -14685 35825 -14565
rect 35945 -14685 35990 -14565
rect 36110 -14685 36155 -14565
rect 36275 -14685 36485 -14565
rect 36605 -14685 36660 -14565
rect 36780 -14685 36825 -14565
rect 36945 -14685 36990 -14565
rect 37110 -14685 37155 -14565
rect 37275 -14685 37330 -14565
rect 37450 -14685 37495 -14565
rect 37615 -14685 37660 -14565
rect 37780 -14685 37825 -14565
rect 37945 -14685 38000 -14565
rect 38120 -14685 38165 -14565
rect 38285 -14685 38330 -14565
rect 38450 -14685 38495 -14565
rect 38615 -14685 38670 -14565
rect 38790 -14685 38835 -14565
rect 38955 -14685 39000 -14565
rect 39120 -14685 39165 -14565
rect 39285 -14685 39340 -14565
rect 39460 -14685 39505 -14565
rect 39625 -14685 39670 -14565
rect 39790 -14685 39835 -14565
rect 39955 -14685 40010 -14565
rect 40130 -14685 40175 -14565
rect 40295 -14685 40340 -14565
rect 40460 -14685 40505 -14565
rect 40625 -14685 40680 -14565
rect 40800 -14685 40845 -14565
rect 40965 -14685 41010 -14565
rect 41130 -14685 41175 -14565
rect 41295 -14685 41350 -14565
rect 41470 -14685 41515 -14565
rect 41635 -14685 41680 -14565
rect 41800 -14685 41845 -14565
rect 41965 -14685 42175 -14565
rect 42295 -14685 42350 -14565
rect 42470 -14685 42515 -14565
rect 42635 -14685 42680 -14565
rect 42800 -14685 42845 -14565
rect 42965 -14685 43020 -14565
rect 43140 -14685 43185 -14565
rect 43305 -14685 43350 -14565
rect 43470 -14685 43515 -14565
rect 43635 -14685 43690 -14565
rect 43810 -14685 43855 -14565
rect 43975 -14685 44020 -14565
rect 44140 -14685 44185 -14565
rect 44305 -14685 44360 -14565
rect 44480 -14685 44525 -14565
rect 44645 -14685 44690 -14565
rect 44810 -14685 44855 -14565
rect 44975 -14685 45030 -14565
rect 45150 -14685 45195 -14565
rect 45315 -14685 45360 -14565
rect 45480 -14685 45525 -14565
rect 45645 -14685 45700 -14565
rect 45820 -14685 45865 -14565
rect 45985 -14685 46030 -14565
rect 46150 -14685 46195 -14565
rect 46315 -14685 46370 -14565
rect 46490 -14685 46535 -14565
rect 46655 -14685 46700 -14565
rect 46820 -14685 46865 -14565
rect 46985 -14685 47040 -14565
rect 47160 -14685 47205 -14565
rect 47325 -14685 47370 -14565
rect 47490 -14685 47535 -14565
rect 47655 -14685 47865 -14565
rect 47985 -14685 48040 -14565
rect 48160 -14685 48205 -14565
rect 48325 -14685 48370 -14565
rect 48490 -14685 48535 -14565
rect 48655 -14685 48710 -14565
rect 48830 -14685 48875 -14565
rect 48995 -14685 49040 -14565
rect 49160 -14685 49205 -14565
rect 49325 -14685 49380 -14565
rect 49500 -14685 49545 -14565
rect 49665 -14685 49710 -14565
rect 49830 -14685 49875 -14565
rect 49995 -14685 50050 -14565
rect 50170 -14685 50215 -14565
rect 50335 -14685 50380 -14565
rect 50500 -14685 50545 -14565
rect 50665 -14685 50720 -14565
rect 50840 -14685 50885 -14565
rect 51005 -14685 51050 -14565
rect 51170 -14685 51215 -14565
rect 51335 -14685 51390 -14565
rect 51510 -14685 51555 -14565
rect 51675 -14685 51720 -14565
rect 51840 -14685 51885 -14565
rect 52005 -14685 52060 -14565
rect 52180 -14685 52225 -14565
rect 52345 -14685 52390 -14565
rect 52510 -14685 52555 -14565
rect 52675 -14685 52730 -14565
rect 52850 -14685 52895 -14565
rect 53015 -14685 53060 -14565
rect 53180 -14685 53225 -14565
rect 53345 -14685 53370 -14565
rect 30770 -14740 53370 -14685
rect 30770 -14860 30795 -14740
rect 30915 -14860 30970 -14740
rect 31090 -14860 31135 -14740
rect 31255 -14860 31300 -14740
rect 31420 -14860 31465 -14740
rect 31585 -14860 31640 -14740
rect 31760 -14860 31805 -14740
rect 31925 -14860 31970 -14740
rect 32090 -14860 32135 -14740
rect 32255 -14860 32310 -14740
rect 32430 -14860 32475 -14740
rect 32595 -14860 32640 -14740
rect 32760 -14860 32805 -14740
rect 32925 -14860 32980 -14740
rect 33100 -14860 33145 -14740
rect 33265 -14860 33310 -14740
rect 33430 -14860 33475 -14740
rect 33595 -14860 33650 -14740
rect 33770 -14860 33815 -14740
rect 33935 -14860 33980 -14740
rect 34100 -14860 34145 -14740
rect 34265 -14860 34320 -14740
rect 34440 -14860 34485 -14740
rect 34605 -14860 34650 -14740
rect 34770 -14860 34815 -14740
rect 34935 -14860 34990 -14740
rect 35110 -14860 35155 -14740
rect 35275 -14860 35320 -14740
rect 35440 -14860 35485 -14740
rect 35605 -14860 35660 -14740
rect 35780 -14860 35825 -14740
rect 35945 -14860 35990 -14740
rect 36110 -14860 36155 -14740
rect 36275 -14860 36485 -14740
rect 36605 -14860 36660 -14740
rect 36780 -14860 36825 -14740
rect 36945 -14860 36990 -14740
rect 37110 -14860 37155 -14740
rect 37275 -14860 37330 -14740
rect 37450 -14860 37495 -14740
rect 37615 -14860 37660 -14740
rect 37780 -14860 37825 -14740
rect 37945 -14860 38000 -14740
rect 38120 -14860 38165 -14740
rect 38285 -14860 38330 -14740
rect 38450 -14860 38495 -14740
rect 38615 -14860 38670 -14740
rect 38790 -14860 38835 -14740
rect 38955 -14860 39000 -14740
rect 39120 -14860 39165 -14740
rect 39285 -14860 39340 -14740
rect 39460 -14860 39505 -14740
rect 39625 -14860 39670 -14740
rect 39790 -14860 39835 -14740
rect 39955 -14860 40010 -14740
rect 40130 -14860 40175 -14740
rect 40295 -14860 40340 -14740
rect 40460 -14860 40505 -14740
rect 40625 -14860 40680 -14740
rect 40800 -14860 40845 -14740
rect 40965 -14860 41010 -14740
rect 41130 -14860 41175 -14740
rect 41295 -14860 41350 -14740
rect 41470 -14860 41515 -14740
rect 41635 -14860 41680 -14740
rect 41800 -14860 41845 -14740
rect 41965 -14860 42175 -14740
rect 42295 -14860 42350 -14740
rect 42470 -14860 42515 -14740
rect 42635 -14860 42680 -14740
rect 42800 -14860 42845 -14740
rect 42965 -14860 43020 -14740
rect 43140 -14860 43185 -14740
rect 43305 -14860 43350 -14740
rect 43470 -14860 43515 -14740
rect 43635 -14860 43690 -14740
rect 43810 -14860 43855 -14740
rect 43975 -14860 44020 -14740
rect 44140 -14860 44185 -14740
rect 44305 -14860 44360 -14740
rect 44480 -14860 44525 -14740
rect 44645 -14860 44690 -14740
rect 44810 -14860 44855 -14740
rect 44975 -14860 45030 -14740
rect 45150 -14860 45195 -14740
rect 45315 -14860 45360 -14740
rect 45480 -14860 45525 -14740
rect 45645 -14860 45700 -14740
rect 45820 -14860 45865 -14740
rect 45985 -14860 46030 -14740
rect 46150 -14860 46195 -14740
rect 46315 -14860 46370 -14740
rect 46490 -14860 46535 -14740
rect 46655 -14860 46700 -14740
rect 46820 -14860 46865 -14740
rect 46985 -14860 47040 -14740
rect 47160 -14860 47205 -14740
rect 47325 -14860 47370 -14740
rect 47490 -14860 47535 -14740
rect 47655 -14860 47865 -14740
rect 47985 -14860 48040 -14740
rect 48160 -14860 48205 -14740
rect 48325 -14860 48370 -14740
rect 48490 -14860 48535 -14740
rect 48655 -14860 48710 -14740
rect 48830 -14860 48875 -14740
rect 48995 -14860 49040 -14740
rect 49160 -14860 49205 -14740
rect 49325 -14860 49380 -14740
rect 49500 -14860 49545 -14740
rect 49665 -14860 49710 -14740
rect 49830 -14860 49875 -14740
rect 49995 -14860 50050 -14740
rect 50170 -14860 50215 -14740
rect 50335 -14860 50380 -14740
rect 50500 -14860 50545 -14740
rect 50665 -14860 50720 -14740
rect 50840 -14860 50885 -14740
rect 51005 -14860 51050 -14740
rect 51170 -14860 51215 -14740
rect 51335 -14860 51390 -14740
rect 51510 -14860 51555 -14740
rect 51675 -14860 51720 -14740
rect 51840 -14860 51885 -14740
rect 52005 -14860 52060 -14740
rect 52180 -14860 52225 -14740
rect 52345 -14860 52390 -14740
rect 52510 -14860 52555 -14740
rect 52675 -14860 52730 -14740
rect 52850 -14860 52895 -14740
rect 53015 -14860 53060 -14740
rect 53180 -14860 53225 -14740
rect 53345 -14860 53370 -14740
rect 30770 -14905 53370 -14860
rect 30770 -15025 30795 -14905
rect 30915 -15025 30970 -14905
rect 31090 -15025 31135 -14905
rect 31255 -15025 31300 -14905
rect 31420 -15025 31465 -14905
rect 31585 -15025 31640 -14905
rect 31760 -15025 31805 -14905
rect 31925 -15025 31970 -14905
rect 32090 -15025 32135 -14905
rect 32255 -15025 32310 -14905
rect 32430 -15025 32475 -14905
rect 32595 -15025 32640 -14905
rect 32760 -15025 32805 -14905
rect 32925 -15025 32980 -14905
rect 33100 -15025 33145 -14905
rect 33265 -15025 33310 -14905
rect 33430 -15025 33475 -14905
rect 33595 -15025 33650 -14905
rect 33770 -15025 33815 -14905
rect 33935 -15025 33980 -14905
rect 34100 -15025 34145 -14905
rect 34265 -15025 34320 -14905
rect 34440 -15025 34485 -14905
rect 34605 -15025 34650 -14905
rect 34770 -15025 34815 -14905
rect 34935 -15025 34990 -14905
rect 35110 -15025 35155 -14905
rect 35275 -15025 35320 -14905
rect 35440 -15025 35485 -14905
rect 35605 -15025 35660 -14905
rect 35780 -15025 35825 -14905
rect 35945 -15025 35990 -14905
rect 36110 -15025 36155 -14905
rect 36275 -15025 36485 -14905
rect 36605 -15025 36660 -14905
rect 36780 -15025 36825 -14905
rect 36945 -15025 36990 -14905
rect 37110 -15025 37155 -14905
rect 37275 -15025 37330 -14905
rect 37450 -15025 37495 -14905
rect 37615 -15025 37660 -14905
rect 37780 -15025 37825 -14905
rect 37945 -15025 38000 -14905
rect 38120 -15025 38165 -14905
rect 38285 -15025 38330 -14905
rect 38450 -15025 38495 -14905
rect 38615 -15025 38670 -14905
rect 38790 -15025 38835 -14905
rect 38955 -15025 39000 -14905
rect 39120 -15025 39165 -14905
rect 39285 -15025 39340 -14905
rect 39460 -15025 39505 -14905
rect 39625 -15025 39670 -14905
rect 39790 -15025 39835 -14905
rect 39955 -15025 40010 -14905
rect 40130 -15025 40175 -14905
rect 40295 -15025 40340 -14905
rect 40460 -15025 40505 -14905
rect 40625 -15025 40680 -14905
rect 40800 -15025 40845 -14905
rect 40965 -15025 41010 -14905
rect 41130 -15025 41175 -14905
rect 41295 -15025 41350 -14905
rect 41470 -15025 41515 -14905
rect 41635 -15025 41680 -14905
rect 41800 -15025 41845 -14905
rect 41965 -15025 42175 -14905
rect 42295 -15025 42350 -14905
rect 42470 -15025 42515 -14905
rect 42635 -15025 42680 -14905
rect 42800 -15025 42845 -14905
rect 42965 -15025 43020 -14905
rect 43140 -15025 43185 -14905
rect 43305 -15025 43350 -14905
rect 43470 -15025 43515 -14905
rect 43635 -15025 43690 -14905
rect 43810 -15025 43855 -14905
rect 43975 -15025 44020 -14905
rect 44140 -15025 44185 -14905
rect 44305 -15025 44360 -14905
rect 44480 -15025 44525 -14905
rect 44645 -15025 44690 -14905
rect 44810 -15025 44855 -14905
rect 44975 -15025 45030 -14905
rect 45150 -15025 45195 -14905
rect 45315 -15025 45360 -14905
rect 45480 -15025 45525 -14905
rect 45645 -15025 45700 -14905
rect 45820 -15025 45865 -14905
rect 45985 -15025 46030 -14905
rect 46150 -15025 46195 -14905
rect 46315 -15025 46370 -14905
rect 46490 -15025 46535 -14905
rect 46655 -15025 46700 -14905
rect 46820 -15025 46865 -14905
rect 46985 -15025 47040 -14905
rect 47160 -15025 47205 -14905
rect 47325 -15025 47370 -14905
rect 47490 -15025 47535 -14905
rect 47655 -15025 47865 -14905
rect 47985 -15025 48040 -14905
rect 48160 -15025 48205 -14905
rect 48325 -15025 48370 -14905
rect 48490 -15025 48535 -14905
rect 48655 -15025 48710 -14905
rect 48830 -15025 48875 -14905
rect 48995 -15025 49040 -14905
rect 49160 -15025 49205 -14905
rect 49325 -15025 49380 -14905
rect 49500 -15025 49545 -14905
rect 49665 -15025 49710 -14905
rect 49830 -15025 49875 -14905
rect 49995 -15025 50050 -14905
rect 50170 -15025 50215 -14905
rect 50335 -15025 50380 -14905
rect 50500 -15025 50545 -14905
rect 50665 -15025 50720 -14905
rect 50840 -15025 50885 -14905
rect 51005 -15025 51050 -14905
rect 51170 -15025 51215 -14905
rect 51335 -15025 51390 -14905
rect 51510 -15025 51555 -14905
rect 51675 -15025 51720 -14905
rect 51840 -15025 51885 -14905
rect 52005 -15025 52060 -14905
rect 52180 -15025 52225 -14905
rect 52345 -15025 52390 -14905
rect 52510 -15025 52555 -14905
rect 52675 -15025 52730 -14905
rect 52850 -15025 52895 -14905
rect 53015 -15025 53060 -14905
rect 53180 -15025 53225 -14905
rect 53345 -15025 53370 -14905
rect 30770 -15070 53370 -15025
rect 30770 -15190 30795 -15070
rect 30915 -15190 30970 -15070
rect 31090 -15190 31135 -15070
rect 31255 -15190 31300 -15070
rect 31420 -15190 31465 -15070
rect 31585 -15190 31640 -15070
rect 31760 -15190 31805 -15070
rect 31925 -15190 31970 -15070
rect 32090 -15190 32135 -15070
rect 32255 -15190 32310 -15070
rect 32430 -15190 32475 -15070
rect 32595 -15190 32640 -15070
rect 32760 -15190 32805 -15070
rect 32925 -15190 32980 -15070
rect 33100 -15190 33145 -15070
rect 33265 -15190 33310 -15070
rect 33430 -15190 33475 -15070
rect 33595 -15190 33650 -15070
rect 33770 -15190 33815 -15070
rect 33935 -15190 33980 -15070
rect 34100 -15190 34145 -15070
rect 34265 -15190 34320 -15070
rect 34440 -15190 34485 -15070
rect 34605 -15190 34650 -15070
rect 34770 -15190 34815 -15070
rect 34935 -15190 34990 -15070
rect 35110 -15190 35155 -15070
rect 35275 -15190 35320 -15070
rect 35440 -15190 35485 -15070
rect 35605 -15190 35660 -15070
rect 35780 -15190 35825 -15070
rect 35945 -15190 35990 -15070
rect 36110 -15190 36155 -15070
rect 36275 -15190 36485 -15070
rect 36605 -15190 36660 -15070
rect 36780 -15190 36825 -15070
rect 36945 -15190 36990 -15070
rect 37110 -15190 37155 -15070
rect 37275 -15190 37330 -15070
rect 37450 -15190 37495 -15070
rect 37615 -15190 37660 -15070
rect 37780 -15190 37825 -15070
rect 37945 -15190 38000 -15070
rect 38120 -15190 38165 -15070
rect 38285 -15190 38330 -15070
rect 38450 -15190 38495 -15070
rect 38615 -15190 38670 -15070
rect 38790 -15190 38835 -15070
rect 38955 -15190 39000 -15070
rect 39120 -15190 39165 -15070
rect 39285 -15190 39340 -15070
rect 39460 -15190 39505 -15070
rect 39625 -15190 39670 -15070
rect 39790 -15190 39835 -15070
rect 39955 -15190 40010 -15070
rect 40130 -15190 40175 -15070
rect 40295 -15190 40340 -15070
rect 40460 -15190 40505 -15070
rect 40625 -15190 40680 -15070
rect 40800 -15190 40845 -15070
rect 40965 -15190 41010 -15070
rect 41130 -15190 41175 -15070
rect 41295 -15190 41350 -15070
rect 41470 -15190 41515 -15070
rect 41635 -15190 41680 -15070
rect 41800 -15190 41845 -15070
rect 41965 -15190 42175 -15070
rect 42295 -15190 42350 -15070
rect 42470 -15190 42515 -15070
rect 42635 -15190 42680 -15070
rect 42800 -15190 42845 -15070
rect 42965 -15190 43020 -15070
rect 43140 -15190 43185 -15070
rect 43305 -15190 43350 -15070
rect 43470 -15190 43515 -15070
rect 43635 -15190 43690 -15070
rect 43810 -15190 43855 -15070
rect 43975 -15190 44020 -15070
rect 44140 -15190 44185 -15070
rect 44305 -15190 44360 -15070
rect 44480 -15190 44525 -15070
rect 44645 -15190 44690 -15070
rect 44810 -15190 44855 -15070
rect 44975 -15190 45030 -15070
rect 45150 -15190 45195 -15070
rect 45315 -15190 45360 -15070
rect 45480 -15190 45525 -15070
rect 45645 -15190 45700 -15070
rect 45820 -15190 45865 -15070
rect 45985 -15190 46030 -15070
rect 46150 -15190 46195 -15070
rect 46315 -15190 46370 -15070
rect 46490 -15190 46535 -15070
rect 46655 -15190 46700 -15070
rect 46820 -15190 46865 -15070
rect 46985 -15190 47040 -15070
rect 47160 -15190 47205 -15070
rect 47325 -15190 47370 -15070
rect 47490 -15190 47535 -15070
rect 47655 -15190 47865 -15070
rect 47985 -15190 48040 -15070
rect 48160 -15190 48205 -15070
rect 48325 -15190 48370 -15070
rect 48490 -15190 48535 -15070
rect 48655 -15190 48710 -15070
rect 48830 -15190 48875 -15070
rect 48995 -15190 49040 -15070
rect 49160 -15190 49205 -15070
rect 49325 -15190 49380 -15070
rect 49500 -15190 49545 -15070
rect 49665 -15190 49710 -15070
rect 49830 -15190 49875 -15070
rect 49995 -15190 50050 -15070
rect 50170 -15190 50215 -15070
rect 50335 -15190 50380 -15070
rect 50500 -15190 50545 -15070
rect 50665 -15190 50720 -15070
rect 50840 -15190 50885 -15070
rect 51005 -15190 51050 -15070
rect 51170 -15190 51215 -15070
rect 51335 -15190 51390 -15070
rect 51510 -15190 51555 -15070
rect 51675 -15190 51720 -15070
rect 51840 -15190 51885 -15070
rect 52005 -15190 52060 -15070
rect 52180 -15190 52225 -15070
rect 52345 -15190 52390 -15070
rect 52510 -15190 52555 -15070
rect 52675 -15190 52730 -15070
rect 52850 -15190 52895 -15070
rect 53015 -15190 53060 -15070
rect 53180 -15190 53225 -15070
rect 53345 -15190 53370 -15070
rect 30770 -15235 53370 -15190
rect 30770 -15355 30795 -15235
rect 30915 -15355 30970 -15235
rect 31090 -15355 31135 -15235
rect 31255 -15355 31300 -15235
rect 31420 -15355 31465 -15235
rect 31585 -15355 31640 -15235
rect 31760 -15355 31805 -15235
rect 31925 -15355 31970 -15235
rect 32090 -15355 32135 -15235
rect 32255 -15355 32310 -15235
rect 32430 -15355 32475 -15235
rect 32595 -15355 32640 -15235
rect 32760 -15355 32805 -15235
rect 32925 -15355 32980 -15235
rect 33100 -15355 33145 -15235
rect 33265 -15355 33310 -15235
rect 33430 -15355 33475 -15235
rect 33595 -15355 33650 -15235
rect 33770 -15355 33815 -15235
rect 33935 -15355 33980 -15235
rect 34100 -15355 34145 -15235
rect 34265 -15355 34320 -15235
rect 34440 -15355 34485 -15235
rect 34605 -15355 34650 -15235
rect 34770 -15355 34815 -15235
rect 34935 -15355 34990 -15235
rect 35110 -15355 35155 -15235
rect 35275 -15355 35320 -15235
rect 35440 -15355 35485 -15235
rect 35605 -15355 35660 -15235
rect 35780 -15355 35825 -15235
rect 35945 -15355 35990 -15235
rect 36110 -15355 36155 -15235
rect 36275 -15355 36485 -15235
rect 36605 -15355 36660 -15235
rect 36780 -15355 36825 -15235
rect 36945 -15355 36990 -15235
rect 37110 -15355 37155 -15235
rect 37275 -15355 37330 -15235
rect 37450 -15355 37495 -15235
rect 37615 -15355 37660 -15235
rect 37780 -15355 37825 -15235
rect 37945 -15355 38000 -15235
rect 38120 -15355 38165 -15235
rect 38285 -15355 38330 -15235
rect 38450 -15355 38495 -15235
rect 38615 -15355 38670 -15235
rect 38790 -15355 38835 -15235
rect 38955 -15355 39000 -15235
rect 39120 -15355 39165 -15235
rect 39285 -15355 39340 -15235
rect 39460 -15355 39505 -15235
rect 39625 -15355 39670 -15235
rect 39790 -15355 39835 -15235
rect 39955 -15355 40010 -15235
rect 40130 -15355 40175 -15235
rect 40295 -15355 40340 -15235
rect 40460 -15355 40505 -15235
rect 40625 -15355 40680 -15235
rect 40800 -15355 40845 -15235
rect 40965 -15355 41010 -15235
rect 41130 -15355 41175 -15235
rect 41295 -15355 41350 -15235
rect 41470 -15355 41515 -15235
rect 41635 -15355 41680 -15235
rect 41800 -15355 41845 -15235
rect 41965 -15355 42175 -15235
rect 42295 -15355 42350 -15235
rect 42470 -15355 42515 -15235
rect 42635 -15355 42680 -15235
rect 42800 -15355 42845 -15235
rect 42965 -15355 43020 -15235
rect 43140 -15355 43185 -15235
rect 43305 -15355 43350 -15235
rect 43470 -15355 43515 -15235
rect 43635 -15355 43690 -15235
rect 43810 -15355 43855 -15235
rect 43975 -15355 44020 -15235
rect 44140 -15355 44185 -15235
rect 44305 -15355 44360 -15235
rect 44480 -15355 44525 -15235
rect 44645 -15355 44690 -15235
rect 44810 -15355 44855 -15235
rect 44975 -15355 45030 -15235
rect 45150 -15355 45195 -15235
rect 45315 -15355 45360 -15235
rect 45480 -15355 45525 -15235
rect 45645 -15355 45700 -15235
rect 45820 -15355 45865 -15235
rect 45985 -15355 46030 -15235
rect 46150 -15355 46195 -15235
rect 46315 -15355 46370 -15235
rect 46490 -15355 46535 -15235
rect 46655 -15355 46700 -15235
rect 46820 -15355 46865 -15235
rect 46985 -15355 47040 -15235
rect 47160 -15355 47205 -15235
rect 47325 -15355 47370 -15235
rect 47490 -15355 47535 -15235
rect 47655 -15355 47865 -15235
rect 47985 -15355 48040 -15235
rect 48160 -15355 48205 -15235
rect 48325 -15355 48370 -15235
rect 48490 -15355 48535 -15235
rect 48655 -15355 48710 -15235
rect 48830 -15355 48875 -15235
rect 48995 -15355 49040 -15235
rect 49160 -15355 49205 -15235
rect 49325 -15355 49380 -15235
rect 49500 -15355 49545 -15235
rect 49665 -15355 49710 -15235
rect 49830 -15355 49875 -15235
rect 49995 -15355 50050 -15235
rect 50170 -15355 50215 -15235
rect 50335 -15355 50380 -15235
rect 50500 -15355 50545 -15235
rect 50665 -15355 50720 -15235
rect 50840 -15355 50885 -15235
rect 51005 -15355 51050 -15235
rect 51170 -15355 51215 -15235
rect 51335 -15355 51390 -15235
rect 51510 -15355 51555 -15235
rect 51675 -15355 51720 -15235
rect 51840 -15355 51885 -15235
rect 52005 -15355 52060 -15235
rect 52180 -15355 52225 -15235
rect 52345 -15355 52390 -15235
rect 52510 -15355 52555 -15235
rect 52675 -15355 52730 -15235
rect 52850 -15355 52895 -15235
rect 53015 -15355 53060 -15235
rect 53180 -15355 53225 -15235
rect 53345 -15355 53370 -15235
rect 30770 -15410 53370 -15355
rect 30770 -15530 30795 -15410
rect 30915 -15530 30970 -15410
rect 31090 -15530 31135 -15410
rect 31255 -15530 31300 -15410
rect 31420 -15530 31465 -15410
rect 31585 -15530 31640 -15410
rect 31760 -15530 31805 -15410
rect 31925 -15530 31970 -15410
rect 32090 -15530 32135 -15410
rect 32255 -15530 32310 -15410
rect 32430 -15530 32475 -15410
rect 32595 -15530 32640 -15410
rect 32760 -15530 32805 -15410
rect 32925 -15530 32980 -15410
rect 33100 -15530 33145 -15410
rect 33265 -15530 33310 -15410
rect 33430 -15530 33475 -15410
rect 33595 -15530 33650 -15410
rect 33770 -15530 33815 -15410
rect 33935 -15530 33980 -15410
rect 34100 -15530 34145 -15410
rect 34265 -15530 34320 -15410
rect 34440 -15530 34485 -15410
rect 34605 -15530 34650 -15410
rect 34770 -15530 34815 -15410
rect 34935 -15530 34990 -15410
rect 35110 -15530 35155 -15410
rect 35275 -15530 35320 -15410
rect 35440 -15530 35485 -15410
rect 35605 -15530 35660 -15410
rect 35780 -15530 35825 -15410
rect 35945 -15530 35990 -15410
rect 36110 -15530 36155 -15410
rect 36275 -15530 36485 -15410
rect 36605 -15530 36660 -15410
rect 36780 -15530 36825 -15410
rect 36945 -15530 36990 -15410
rect 37110 -15530 37155 -15410
rect 37275 -15530 37330 -15410
rect 37450 -15530 37495 -15410
rect 37615 -15530 37660 -15410
rect 37780 -15530 37825 -15410
rect 37945 -15530 38000 -15410
rect 38120 -15530 38165 -15410
rect 38285 -15530 38330 -15410
rect 38450 -15530 38495 -15410
rect 38615 -15530 38670 -15410
rect 38790 -15530 38835 -15410
rect 38955 -15530 39000 -15410
rect 39120 -15530 39165 -15410
rect 39285 -15530 39340 -15410
rect 39460 -15530 39505 -15410
rect 39625 -15530 39670 -15410
rect 39790 -15530 39835 -15410
rect 39955 -15530 40010 -15410
rect 40130 -15530 40175 -15410
rect 40295 -15530 40340 -15410
rect 40460 -15530 40505 -15410
rect 40625 -15530 40680 -15410
rect 40800 -15530 40845 -15410
rect 40965 -15530 41010 -15410
rect 41130 -15530 41175 -15410
rect 41295 -15530 41350 -15410
rect 41470 -15530 41515 -15410
rect 41635 -15530 41680 -15410
rect 41800 -15530 41845 -15410
rect 41965 -15530 42175 -15410
rect 42295 -15530 42350 -15410
rect 42470 -15530 42515 -15410
rect 42635 -15530 42680 -15410
rect 42800 -15530 42845 -15410
rect 42965 -15530 43020 -15410
rect 43140 -15530 43185 -15410
rect 43305 -15530 43350 -15410
rect 43470 -15530 43515 -15410
rect 43635 -15530 43690 -15410
rect 43810 -15530 43855 -15410
rect 43975 -15530 44020 -15410
rect 44140 -15530 44185 -15410
rect 44305 -15530 44360 -15410
rect 44480 -15530 44525 -15410
rect 44645 -15530 44690 -15410
rect 44810 -15530 44855 -15410
rect 44975 -15530 45030 -15410
rect 45150 -15530 45195 -15410
rect 45315 -15530 45360 -15410
rect 45480 -15530 45525 -15410
rect 45645 -15530 45700 -15410
rect 45820 -15530 45865 -15410
rect 45985 -15530 46030 -15410
rect 46150 -15530 46195 -15410
rect 46315 -15530 46370 -15410
rect 46490 -15530 46535 -15410
rect 46655 -15530 46700 -15410
rect 46820 -15530 46865 -15410
rect 46985 -15530 47040 -15410
rect 47160 -15530 47205 -15410
rect 47325 -15530 47370 -15410
rect 47490 -15530 47535 -15410
rect 47655 -15530 47865 -15410
rect 47985 -15530 48040 -15410
rect 48160 -15530 48205 -15410
rect 48325 -15530 48370 -15410
rect 48490 -15530 48535 -15410
rect 48655 -15530 48710 -15410
rect 48830 -15530 48875 -15410
rect 48995 -15530 49040 -15410
rect 49160 -15530 49205 -15410
rect 49325 -15530 49380 -15410
rect 49500 -15530 49545 -15410
rect 49665 -15530 49710 -15410
rect 49830 -15530 49875 -15410
rect 49995 -15530 50050 -15410
rect 50170 -15530 50215 -15410
rect 50335 -15530 50380 -15410
rect 50500 -15530 50545 -15410
rect 50665 -15530 50720 -15410
rect 50840 -15530 50885 -15410
rect 51005 -15530 51050 -15410
rect 51170 -15530 51215 -15410
rect 51335 -15530 51390 -15410
rect 51510 -15530 51555 -15410
rect 51675 -15530 51720 -15410
rect 51840 -15530 51885 -15410
rect 52005 -15530 52060 -15410
rect 52180 -15530 52225 -15410
rect 52345 -15530 52390 -15410
rect 52510 -15530 52555 -15410
rect 52675 -15530 52730 -15410
rect 52850 -15530 52895 -15410
rect 53015 -15530 53060 -15410
rect 53180 -15530 53225 -15410
rect 53345 -15530 53370 -15410
rect 30770 -15555 53370 -15530
<< labels >>
rlabel metal4 30640 4460 30640 4460 1 VDD
port 1 n
rlabel metal4 30695 -2170 30695 -2170 1 VDD
rlabel metal4 30640 -14264 30640 -14264 1 VDD
rlabel metal5 30500 -10679 30500 -10679 1 GND
port 2 n
<< end >>
