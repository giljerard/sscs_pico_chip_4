magic
tech sky130A
timestamp 1636437882
<< metal3 >>
rect 7105 1610 12635 7185
rect 12795 1610 18325 7185
rect 18485 1610 24015 7185
rect 24175 1610 29705 7185
rect 7105 1590 29705 1610
rect 7105 1470 7170 1590
rect 7290 1470 7335 1590
rect 7455 1470 7500 1590
rect 7620 1470 7665 1590
rect 7785 1470 7830 1590
rect 7950 1470 7995 1590
rect 8115 1470 8160 1590
rect 8280 1470 8325 1590
rect 8445 1470 8490 1590
rect 8610 1470 8655 1590
rect 8775 1470 8820 1590
rect 8940 1470 8985 1590
rect 9105 1470 9150 1590
rect 9270 1470 9315 1590
rect 9435 1470 9480 1590
rect 9600 1470 9645 1590
rect 9765 1470 9810 1590
rect 9930 1470 9975 1590
rect 10095 1470 10140 1590
rect 10260 1470 10305 1590
rect 10425 1470 10470 1590
rect 10590 1470 10635 1590
rect 10755 1470 10800 1590
rect 10920 1470 10965 1590
rect 11085 1470 11130 1590
rect 11250 1470 11295 1590
rect 11415 1470 11460 1590
rect 11580 1470 11625 1590
rect 11745 1470 11790 1590
rect 11910 1470 11955 1590
rect 12075 1470 12120 1590
rect 12240 1470 12285 1590
rect 12405 1470 12450 1590
rect 12570 1470 12860 1590
rect 12980 1470 13025 1590
rect 13145 1470 13190 1590
rect 13310 1470 13355 1590
rect 13475 1470 13520 1590
rect 13640 1470 13685 1590
rect 13805 1470 13850 1590
rect 13970 1470 14015 1590
rect 14135 1470 14180 1590
rect 14300 1470 14345 1590
rect 14465 1470 14510 1590
rect 14630 1470 14675 1590
rect 14795 1470 14840 1590
rect 14960 1470 15005 1590
rect 15125 1470 15170 1590
rect 15290 1470 15335 1590
rect 15455 1470 15500 1590
rect 15620 1470 15665 1590
rect 15785 1470 15830 1590
rect 15950 1470 15995 1590
rect 16115 1470 16160 1590
rect 16280 1470 16325 1590
rect 16445 1470 16490 1590
rect 16610 1470 16655 1590
rect 16775 1470 16820 1590
rect 16940 1470 16985 1590
rect 17105 1470 17150 1590
rect 17270 1470 17315 1590
rect 17435 1470 17480 1590
rect 17600 1470 17645 1590
rect 17765 1470 17810 1590
rect 17930 1470 17975 1590
rect 18095 1470 18140 1590
rect 18260 1470 18550 1590
rect 18670 1470 18715 1590
rect 18835 1470 18880 1590
rect 19000 1470 19045 1590
rect 19165 1470 19210 1590
rect 19330 1470 19375 1590
rect 19495 1470 19540 1590
rect 19660 1470 19705 1590
rect 19825 1470 19870 1590
rect 19990 1470 20035 1590
rect 20155 1470 20200 1590
rect 20320 1470 20365 1590
rect 20485 1470 20530 1590
rect 20650 1470 20695 1590
rect 20815 1470 20860 1590
rect 20980 1470 21025 1590
rect 21145 1470 21190 1590
rect 21310 1470 21355 1590
rect 21475 1470 21520 1590
rect 21640 1470 21685 1590
rect 21805 1470 21850 1590
rect 21970 1470 22015 1590
rect 22135 1470 22180 1590
rect 22300 1470 22345 1590
rect 22465 1470 22510 1590
rect 22630 1470 22675 1590
rect 22795 1470 22840 1590
rect 22960 1470 23005 1590
rect 23125 1470 23170 1590
rect 23290 1470 23335 1590
rect 23455 1470 23500 1590
rect 23620 1470 23665 1590
rect 23785 1470 23830 1590
rect 23950 1470 24240 1590
rect 24360 1470 24405 1590
rect 24525 1470 24570 1590
rect 24690 1470 24735 1590
rect 24855 1470 24900 1590
rect 25020 1470 25065 1590
rect 25185 1470 25230 1590
rect 25350 1470 25395 1590
rect 25515 1470 25560 1590
rect 25680 1470 25725 1590
rect 25845 1470 25890 1590
rect 26010 1470 26055 1590
rect 26175 1470 26220 1590
rect 26340 1470 26385 1590
rect 26505 1470 26550 1590
rect 26670 1470 26715 1590
rect 26835 1470 26880 1590
rect 27000 1470 27045 1590
rect 27165 1470 27210 1590
rect 27330 1470 27375 1590
rect 27495 1470 27540 1590
rect 27660 1470 27705 1590
rect 27825 1470 27870 1590
rect 27990 1470 28035 1590
rect 28155 1470 28200 1590
rect 28320 1470 28365 1590
rect 28485 1470 28530 1590
rect 28650 1470 28695 1590
rect 28815 1470 28860 1590
rect 28980 1470 29025 1590
rect 29145 1470 29190 1590
rect 29310 1470 29355 1590
rect 29475 1470 29520 1590
rect 29640 1470 29705 1590
rect 7105 1450 29705 1470
rect 7105 -4125 12635 1450
rect 12795 -4125 18325 1450
rect 18485 -4125 24015 1450
rect 24175 -4125 29705 1450
rect 7105 -9860 12635 -4285
rect 12795 -9860 18325 -4285
rect 18485 -9860 24015 -4285
rect 24175 -9860 29705 -4285
rect 7105 -9880 29705 -9860
rect 7105 -10000 7170 -9880
rect 7290 -10000 7335 -9880
rect 7455 -10000 7500 -9880
rect 7620 -10000 7665 -9880
rect 7785 -10000 7830 -9880
rect 7950 -10000 7995 -9880
rect 8115 -10000 8160 -9880
rect 8280 -10000 8325 -9880
rect 8445 -10000 8490 -9880
rect 8610 -10000 8655 -9880
rect 8775 -10000 8820 -9880
rect 8940 -10000 8985 -9880
rect 9105 -10000 9150 -9880
rect 9270 -10000 9315 -9880
rect 9435 -10000 9480 -9880
rect 9600 -10000 9645 -9880
rect 9765 -10000 9810 -9880
rect 9930 -10000 9975 -9880
rect 10095 -10000 10140 -9880
rect 10260 -10000 10305 -9880
rect 10425 -10000 10470 -9880
rect 10590 -10000 10635 -9880
rect 10755 -10000 10800 -9880
rect 10920 -10000 10965 -9880
rect 11085 -10000 11130 -9880
rect 11250 -10000 11295 -9880
rect 11415 -10000 11460 -9880
rect 11580 -10000 11625 -9880
rect 11745 -10000 11790 -9880
rect 11910 -10000 11955 -9880
rect 12075 -10000 12120 -9880
rect 12240 -10000 12285 -9880
rect 12405 -10000 12450 -9880
rect 12570 -10000 12860 -9880
rect 12980 -10000 13025 -9880
rect 13145 -10000 13190 -9880
rect 13310 -10000 13355 -9880
rect 13475 -10000 13520 -9880
rect 13640 -10000 13685 -9880
rect 13805 -10000 13850 -9880
rect 13970 -10000 14015 -9880
rect 14135 -10000 14180 -9880
rect 14300 -10000 14345 -9880
rect 14465 -10000 14510 -9880
rect 14630 -10000 14675 -9880
rect 14795 -10000 14840 -9880
rect 14960 -10000 15005 -9880
rect 15125 -10000 15170 -9880
rect 15290 -10000 15335 -9880
rect 15455 -10000 15500 -9880
rect 15620 -10000 15665 -9880
rect 15785 -10000 15830 -9880
rect 15950 -10000 15995 -9880
rect 16115 -10000 16160 -9880
rect 16280 -10000 16325 -9880
rect 16445 -10000 16490 -9880
rect 16610 -10000 16655 -9880
rect 16775 -10000 16820 -9880
rect 16940 -10000 16985 -9880
rect 17105 -10000 17150 -9880
rect 17270 -10000 17315 -9880
rect 17435 -10000 17480 -9880
rect 17600 -10000 17645 -9880
rect 17765 -10000 17810 -9880
rect 17930 -10000 17975 -9880
rect 18095 -10000 18140 -9880
rect 18260 -10000 18550 -9880
rect 18670 -10000 18715 -9880
rect 18835 -10000 18880 -9880
rect 19000 -10000 19045 -9880
rect 19165 -10000 19210 -9880
rect 19330 -10000 19375 -9880
rect 19495 -10000 19540 -9880
rect 19660 -10000 19705 -9880
rect 19825 -10000 19870 -9880
rect 19990 -10000 20035 -9880
rect 20155 -10000 20200 -9880
rect 20320 -10000 20365 -9880
rect 20485 -10000 20530 -9880
rect 20650 -10000 20695 -9880
rect 20815 -10000 20860 -9880
rect 20980 -10000 21025 -9880
rect 21145 -10000 21190 -9880
rect 21310 -10000 21355 -9880
rect 21475 -10000 21520 -9880
rect 21640 -10000 21685 -9880
rect 21805 -10000 21850 -9880
rect 21970 -10000 22015 -9880
rect 22135 -10000 22180 -9880
rect 22300 -10000 22345 -9880
rect 22465 -10000 22510 -9880
rect 22630 -10000 22675 -9880
rect 22795 -10000 22840 -9880
rect 22960 -10000 23005 -9880
rect 23125 -10000 23170 -9880
rect 23290 -10000 23335 -9880
rect 23455 -10000 23500 -9880
rect 23620 -10000 23665 -9880
rect 23785 -10000 23830 -9880
rect 23950 -10000 24240 -9880
rect 24360 -10000 24405 -9880
rect 24525 -10000 24570 -9880
rect 24690 -10000 24735 -9880
rect 24855 -10000 24900 -9880
rect 25020 -10000 25065 -9880
rect 25185 -10000 25230 -9880
rect 25350 -10000 25395 -9880
rect 25515 -10000 25560 -9880
rect 25680 -10000 25725 -9880
rect 25845 -10000 25890 -9880
rect 26010 -10000 26055 -9880
rect 26175 -10000 26220 -9880
rect 26340 -10000 26385 -9880
rect 26505 -10000 26550 -9880
rect 26670 -10000 26715 -9880
rect 26835 -10000 26880 -9880
rect 27000 -10000 27045 -9880
rect 27165 -10000 27210 -9880
rect 27330 -10000 27375 -9880
rect 27495 -10000 27540 -9880
rect 27660 -10000 27705 -9880
rect 27825 -10000 27870 -9880
rect 27990 -10000 28035 -9880
rect 28155 -10000 28200 -9880
rect 28320 -10000 28365 -9880
rect 28485 -10000 28530 -9880
rect 28650 -10000 28695 -9880
rect 28815 -10000 28860 -9880
rect 28980 -10000 29025 -9880
rect 29145 -10000 29190 -9880
rect 29310 -10000 29355 -9880
rect 29475 -10000 29520 -9880
rect 29640 -10000 29705 -9880
rect 7105 -10020 29705 -10000
rect 7105 -15595 12635 -10020
rect 12795 -15595 18325 -10020
rect 18485 -15595 24015 -10020
rect 24175 -15595 29705 -10020
<< via3 >>
rect 7170 1470 7290 1590
rect 7335 1470 7455 1590
rect 7500 1470 7620 1590
rect 7665 1470 7785 1590
rect 7830 1470 7950 1590
rect 7995 1470 8115 1590
rect 8160 1470 8280 1590
rect 8325 1470 8445 1590
rect 8490 1470 8610 1590
rect 8655 1470 8775 1590
rect 8820 1470 8940 1590
rect 8985 1470 9105 1590
rect 9150 1470 9270 1590
rect 9315 1470 9435 1590
rect 9480 1470 9600 1590
rect 9645 1470 9765 1590
rect 9810 1470 9930 1590
rect 9975 1470 10095 1590
rect 10140 1470 10260 1590
rect 10305 1470 10425 1590
rect 10470 1470 10590 1590
rect 10635 1470 10755 1590
rect 10800 1470 10920 1590
rect 10965 1470 11085 1590
rect 11130 1470 11250 1590
rect 11295 1470 11415 1590
rect 11460 1470 11580 1590
rect 11625 1470 11745 1590
rect 11790 1470 11910 1590
rect 11955 1470 12075 1590
rect 12120 1470 12240 1590
rect 12285 1470 12405 1590
rect 12450 1470 12570 1590
rect 12860 1470 12980 1590
rect 13025 1470 13145 1590
rect 13190 1470 13310 1590
rect 13355 1470 13475 1590
rect 13520 1470 13640 1590
rect 13685 1470 13805 1590
rect 13850 1470 13970 1590
rect 14015 1470 14135 1590
rect 14180 1470 14300 1590
rect 14345 1470 14465 1590
rect 14510 1470 14630 1590
rect 14675 1470 14795 1590
rect 14840 1470 14960 1590
rect 15005 1470 15125 1590
rect 15170 1470 15290 1590
rect 15335 1470 15455 1590
rect 15500 1470 15620 1590
rect 15665 1470 15785 1590
rect 15830 1470 15950 1590
rect 15995 1470 16115 1590
rect 16160 1470 16280 1590
rect 16325 1470 16445 1590
rect 16490 1470 16610 1590
rect 16655 1470 16775 1590
rect 16820 1470 16940 1590
rect 16985 1470 17105 1590
rect 17150 1470 17270 1590
rect 17315 1470 17435 1590
rect 17480 1470 17600 1590
rect 17645 1470 17765 1590
rect 17810 1470 17930 1590
rect 17975 1470 18095 1590
rect 18140 1470 18260 1590
rect 18550 1470 18670 1590
rect 18715 1470 18835 1590
rect 18880 1470 19000 1590
rect 19045 1470 19165 1590
rect 19210 1470 19330 1590
rect 19375 1470 19495 1590
rect 19540 1470 19660 1590
rect 19705 1470 19825 1590
rect 19870 1470 19990 1590
rect 20035 1470 20155 1590
rect 20200 1470 20320 1590
rect 20365 1470 20485 1590
rect 20530 1470 20650 1590
rect 20695 1470 20815 1590
rect 20860 1470 20980 1590
rect 21025 1470 21145 1590
rect 21190 1470 21310 1590
rect 21355 1470 21475 1590
rect 21520 1470 21640 1590
rect 21685 1470 21805 1590
rect 21850 1470 21970 1590
rect 22015 1470 22135 1590
rect 22180 1470 22300 1590
rect 22345 1470 22465 1590
rect 22510 1470 22630 1590
rect 22675 1470 22795 1590
rect 22840 1470 22960 1590
rect 23005 1470 23125 1590
rect 23170 1470 23290 1590
rect 23335 1470 23455 1590
rect 23500 1470 23620 1590
rect 23665 1470 23785 1590
rect 23830 1470 23950 1590
rect 24240 1470 24360 1590
rect 24405 1470 24525 1590
rect 24570 1470 24690 1590
rect 24735 1470 24855 1590
rect 24900 1470 25020 1590
rect 25065 1470 25185 1590
rect 25230 1470 25350 1590
rect 25395 1470 25515 1590
rect 25560 1470 25680 1590
rect 25725 1470 25845 1590
rect 25890 1470 26010 1590
rect 26055 1470 26175 1590
rect 26220 1470 26340 1590
rect 26385 1470 26505 1590
rect 26550 1470 26670 1590
rect 26715 1470 26835 1590
rect 26880 1470 27000 1590
rect 27045 1470 27165 1590
rect 27210 1470 27330 1590
rect 27375 1470 27495 1590
rect 27540 1470 27660 1590
rect 27705 1470 27825 1590
rect 27870 1470 27990 1590
rect 28035 1470 28155 1590
rect 28200 1470 28320 1590
rect 28365 1470 28485 1590
rect 28530 1470 28650 1590
rect 28695 1470 28815 1590
rect 28860 1470 28980 1590
rect 29025 1470 29145 1590
rect 29190 1470 29310 1590
rect 29355 1470 29475 1590
rect 29520 1470 29640 1590
rect 7170 -10000 7290 -9880
rect 7335 -10000 7455 -9880
rect 7500 -10000 7620 -9880
rect 7665 -10000 7785 -9880
rect 7830 -10000 7950 -9880
rect 7995 -10000 8115 -9880
rect 8160 -10000 8280 -9880
rect 8325 -10000 8445 -9880
rect 8490 -10000 8610 -9880
rect 8655 -10000 8775 -9880
rect 8820 -10000 8940 -9880
rect 8985 -10000 9105 -9880
rect 9150 -10000 9270 -9880
rect 9315 -10000 9435 -9880
rect 9480 -10000 9600 -9880
rect 9645 -10000 9765 -9880
rect 9810 -10000 9930 -9880
rect 9975 -10000 10095 -9880
rect 10140 -10000 10260 -9880
rect 10305 -10000 10425 -9880
rect 10470 -10000 10590 -9880
rect 10635 -10000 10755 -9880
rect 10800 -10000 10920 -9880
rect 10965 -10000 11085 -9880
rect 11130 -10000 11250 -9880
rect 11295 -10000 11415 -9880
rect 11460 -10000 11580 -9880
rect 11625 -10000 11745 -9880
rect 11790 -10000 11910 -9880
rect 11955 -10000 12075 -9880
rect 12120 -10000 12240 -9880
rect 12285 -10000 12405 -9880
rect 12450 -10000 12570 -9880
rect 12860 -10000 12980 -9880
rect 13025 -10000 13145 -9880
rect 13190 -10000 13310 -9880
rect 13355 -10000 13475 -9880
rect 13520 -10000 13640 -9880
rect 13685 -10000 13805 -9880
rect 13850 -10000 13970 -9880
rect 14015 -10000 14135 -9880
rect 14180 -10000 14300 -9880
rect 14345 -10000 14465 -9880
rect 14510 -10000 14630 -9880
rect 14675 -10000 14795 -9880
rect 14840 -10000 14960 -9880
rect 15005 -10000 15125 -9880
rect 15170 -10000 15290 -9880
rect 15335 -10000 15455 -9880
rect 15500 -10000 15620 -9880
rect 15665 -10000 15785 -9880
rect 15830 -10000 15950 -9880
rect 15995 -10000 16115 -9880
rect 16160 -10000 16280 -9880
rect 16325 -10000 16445 -9880
rect 16490 -10000 16610 -9880
rect 16655 -10000 16775 -9880
rect 16820 -10000 16940 -9880
rect 16985 -10000 17105 -9880
rect 17150 -10000 17270 -9880
rect 17315 -10000 17435 -9880
rect 17480 -10000 17600 -9880
rect 17645 -10000 17765 -9880
rect 17810 -10000 17930 -9880
rect 17975 -10000 18095 -9880
rect 18140 -10000 18260 -9880
rect 18550 -10000 18670 -9880
rect 18715 -10000 18835 -9880
rect 18880 -10000 19000 -9880
rect 19045 -10000 19165 -9880
rect 19210 -10000 19330 -9880
rect 19375 -10000 19495 -9880
rect 19540 -10000 19660 -9880
rect 19705 -10000 19825 -9880
rect 19870 -10000 19990 -9880
rect 20035 -10000 20155 -9880
rect 20200 -10000 20320 -9880
rect 20365 -10000 20485 -9880
rect 20530 -10000 20650 -9880
rect 20695 -10000 20815 -9880
rect 20860 -10000 20980 -9880
rect 21025 -10000 21145 -9880
rect 21190 -10000 21310 -9880
rect 21355 -10000 21475 -9880
rect 21520 -10000 21640 -9880
rect 21685 -10000 21805 -9880
rect 21850 -10000 21970 -9880
rect 22015 -10000 22135 -9880
rect 22180 -10000 22300 -9880
rect 22345 -10000 22465 -9880
rect 22510 -10000 22630 -9880
rect 22675 -10000 22795 -9880
rect 22840 -10000 22960 -9880
rect 23005 -10000 23125 -9880
rect 23170 -10000 23290 -9880
rect 23335 -10000 23455 -9880
rect 23500 -10000 23620 -9880
rect 23665 -10000 23785 -9880
rect 23830 -10000 23950 -9880
rect 24240 -10000 24360 -9880
rect 24405 -10000 24525 -9880
rect 24570 -10000 24690 -9880
rect 24735 -10000 24855 -9880
rect 24900 -10000 25020 -9880
rect 25065 -10000 25185 -9880
rect 25230 -10000 25350 -9880
rect 25395 -10000 25515 -9880
rect 25560 -10000 25680 -9880
rect 25725 -10000 25845 -9880
rect 25890 -10000 26010 -9880
rect 26055 -10000 26175 -9880
rect 26220 -10000 26340 -9880
rect 26385 -10000 26505 -9880
rect 26550 -10000 26670 -9880
rect 26715 -10000 26835 -9880
rect 26880 -10000 27000 -9880
rect 27045 -10000 27165 -9880
rect 27210 -10000 27330 -9880
rect 27375 -10000 27495 -9880
rect 27540 -10000 27660 -9880
rect 27705 -10000 27825 -9880
rect 27870 -10000 27990 -9880
rect 28035 -10000 28155 -9880
rect 28200 -10000 28320 -9880
rect 28365 -10000 28485 -9880
rect 28530 -10000 28650 -9880
rect 28695 -10000 28815 -9880
rect 28860 -10000 28980 -9880
rect 29025 -10000 29145 -9880
rect 29190 -10000 29310 -9880
rect 29355 -10000 29475 -9880
rect 29520 -10000 29640 -9880
<< mimcap >>
rect 7120 7160 12620 7170
rect 7120 7040 7130 7160
rect 7250 7040 7295 7160
rect 7415 7040 7460 7160
rect 7580 7040 7625 7160
rect 7745 7040 7800 7160
rect 7920 7040 7965 7160
rect 8085 7040 8130 7160
rect 8250 7040 8295 7160
rect 8415 7040 8470 7160
rect 8590 7040 8635 7160
rect 8755 7040 8800 7160
rect 8920 7040 8965 7160
rect 9085 7040 9140 7160
rect 9260 7040 9305 7160
rect 9425 7040 9470 7160
rect 9590 7040 9635 7160
rect 9755 7040 9810 7160
rect 9930 7040 9975 7160
rect 10095 7040 10140 7160
rect 10260 7040 10305 7160
rect 10425 7040 10480 7160
rect 10600 7040 10645 7160
rect 10765 7040 10810 7160
rect 10930 7040 10975 7160
rect 11095 7040 11150 7160
rect 11270 7040 11315 7160
rect 11435 7040 11480 7160
rect 11600 7040 11645 7160
rect 11765 7040 11820 7160
rect 11940 7040 11985 7160
rect 12105 7040 12150 7160
rect 12270 7040 12315 7160
rect 12435 7040 12490 7160
rect 12610 7040 12620 7160
rect 7120 6985 12620 7040
rect 7120 6865 7130 6985
rect 7250 6865 7295 6985
rect 7415 6865 7460 6985
rect 7580 6865 7625 6985
rect 7745 6865 7800 6985
rect 7920 6865 7965 6985
rect 8085 6865 8130 6985
rect 8250 6865 8295 6985
rect 8415 6865 8470 6985
rect 8590 6865 8635 6985
rect 8755 6865 8800 6985
rect 8920 6865 8965 6985
rect 9085 6865 9140 6985
rect 9260 6865 9305 6985
rect 9425 6865 9470 6985
rect 9590 6865 9635 6985
rect 9755 6865 9810 6985
rect 9930 6865 9975 6985
rect 10095 6865 10140 6985
rect 10260 6865 10305 6985
rect 10425 6865 10480 6985
rect 10600 6865 10645 6985
rect 10765 6865 10810 6985
rect 10930 6865 10975 6985
rect 11095 6865 11150 6985
rect 11270 6865 11315 6985
rect 11435 6865 11480 6985
rect 11600 6865 11645 6985
rect 11765 6865 11820 6985
rect 11940 6865 11985 6985
rect 12105 6865 12150 6985
rect 12270 6865 12315 6985
rect 12435 6865 12490 6985
rect 12610 6865 12620 6985
rect 7120 6820 12620 6865
rect 7120 6700 7130 6820
rect 7250 6700 7295 6820
rect 7415 6700 7460 6820
rect 7580 6700 7625 6820
rect 7745 6700 7800 6820
rect 7920 6700 7965 6820
rect 8085 6700 8130 6820
rect 8250 6700 8295 6820
rect 8415 6700 8470 6820
rect 8590 6700 8635 6820
rect 8755 6700 8800 6820
rect 8920 6700 8965 6820
rect 9085 6700 9140 6820
rect 9260 6700 9305 6820
rect 9425 6700 9470 6820
rect 9590 6700 9635 6820
rect 9755 6700 9810 6820
rect 9930 6700 9975 6820
rect 10095 6700 10140 6820
rect 10260 6700 10305 6820
rect 10425 6700 10480 6820
rect 10600 6700 10645 6820
rect 10765 6700 10810 6820
rect 10930 6700 10975 6820
rect 11095 6700 11150 6820
rect 11270 6700 11315 6820
rect 11435 6700 11480 6820
rect 11600 6700 11645 6820
rect 11765 6700 11820 6820
rect 11940 6700 11985 6820
rect 12105 6700 12150 6820
rect 12270 6700 12315 6820
rect 12435 6700 12490 6820
rect 12610 6700 12620 6820
rect 7120 6655 12620 6700
rect 7120 6535 7130 6655
rect 7250 6535 7295 6655
rect 7415 6535 7460 6655
rect 7580 6535 7625 6655
rect 7745 6535 7800 6655
rect 7920 6535 7965 6655
rect 8085 6535 8130 6655
rect 8250 6535 8295 6655
rect 8415 6535 8470 6655
rect 8590 6535 8635 6655
rect 8755 6535 8800 6655
rect 8920 6535 8965 6655
rect 9085 6535 9140 6655
rect 9260 6535 9305 6655
rect 9425 6535 9470 6655
rect 9590 6535 9635 6655
rect 9755 6535 9810 6655
rect 9930 6535 9975 6655
rect 10095 6535 10140 6655
rect 10260 6535 10305 6655
rect 10425 6535 10480 6655
rect 10600 6535 10645 6655
rect 10765 6535 10810 6655
rect 10930 6535 10975 6655
rect 11095 6535 11150 6655
rect 11270 6535 11315 6655
rect 11435 6535 11480 6655
rect 11600 6535 11645 6655
rect 11765 6535 11820 6655
rect 11940 6535 11985 6655
rect 12105 6535 12150 6655
rect 12270 6535 12315 6655
rect 12435 6535 12490 6655
rect 12610 6535 12620 6655
rect 7120 6490 12620 6535
rect 7120 6370 7130 6490
rect 7250 6370 7295 6490
rect 7415 6370 7460 6490
rect 7580 6370 7625 6490
rect 7745 6370 7800 6490
rect 7920 6370 7965 6490
rect 8085 6370 8130 6490
rect 8250 6370 8295 6490
rect 8415 6370 8470 6490
rect 8590 6370 8635 6490
rect 8755 6370 8800 6490
rect 8920 6370 8965 6490
rect 9085 6370 9140 6490
rect 9260 6370 9305 6490
rect 9425 6370 9470 6490
rect 9590 6370 9635 6490
rect 9755 6370 9810 6490
rect 9930 6370 9975 6490
rect 10095 6370 10140 6490
rect 10260 6370 10305 6490
rect 10425 6370 10480 6490
rect 10600 6370 10645 6490
rect 10765 6370 10810 6490
rect 10930 6370 10975 6490
rect 11095 6370 11150 6490
rect 11270 6370 11315 6490
rect 11435 6370 11480 6490
rect 11600 6370 11645 6490
rect 11765 6370 11820 6490
rect 11940 6370 11985 6490
rect 12105 6370 12150 6490
rect 12270 6370 12315 6490
rect 12435 6370 12490 6490
rect 12610 6370 12620 6490
rect 7120 6315 12620 6370
rect 7120 6195 7130 6315
rect 7250 6195 7295 6315
rect 7415 6195 7460 6315
rect 7580 6195 7625 6315
rect 7745 6195 7800 6315
rect 7920 6195 7965 6315
rect 8085 6195 8130 6315
rect 8250 6195 8295 6315
rect 8415 6195 8470 6315
rect 8590 6195 8635 6315
rect 8755 6195 8800 6315
rect 8920 6195 8965 6315
rect 9085 6195 9140 6315
rect 9260 6195 9305 6315
rect 9425 6195 9470 6315
rect 9590 6195 9635 6315
rect 9755 6195 9810 6315
rect 9930 6195 9975 6315
rect 10095 6195 10140 6315
rect 10260 6195 10305 6315
rect 10425 6195 10480 6315
rect 10600 6195 10645 6315
rect 10765 6195 10810 6315
rect 10930 6195 10975 6315
rect 11095 6195 11150 6315
rect 11270 6195 11315 6315
rect 11435 6195 11480 6315
rect 11600 6195 11645 6315
rect 11765 6195 11820 6315
rect 11940 6195 11985 6315
rect 12105 6195 12150 6315
rect 12270 6195 12315 6315
rect 12435 6195 12490 6315
rect 12610 6195 12620 6315
rect 7120 6150 12620 6195
rect 7120 6030 7130 6150
rect 7250 6030 7295 6150
rect 7415 6030 7460 6150
rect 7580 6030 7625 6150
rect 7745 6030 7800 6150
rect 7920 6030 7965 6150
rect 8085 6030 8130 6150
rect 8250 6030 8295 6150
rect 8415 6030 8470 6150
rect 8590 6030 8635 6150
rect 8755 6030 8800 6150
rect 8920 6030 8965 6150
rect 9085 6030 9140 6150
rect 9260 6030 9305 6150
rect 9425 6030 9470 6150
rect 9590 6030 9635 6150
rect 9755 6030 9810 6150
rect 9930 6030 9975 6150
rect 10095 6030 10140 6150
rect 10260 6030 10305 6150
rect 10425 6030 10480 6150
rect 10600 6030 10645 6150
rect 10765 6030 10810 6150
rect 10930 6030 10975 6150
rect 11095 6030 11150 6150
rect 11270 6030 11315 6150
rect 11435 6030 11480 6150
rect 11600 6030 11645 6150
rect 11765 6030 11820 6150
rect 11940 6030 11985 6150
rect 12105 6030 12150 6150
rect 12270 6030 12315 6150
rect 12435 6030 12490 6150
rect 12610 6030 12620 6150
rect 7120 5985 12620 6030
rect 7120 5865 7130 5985
rect 7250 5865 7295 5985
rect 7415 5865 7460 5985
rect 7580 5865 7625 5985
rect 7745 5865 7800 5985
rect 7920 5865 7965 5985
rect 8085 5865 8130 5985
rect 8250 5865 8295 5985
rect 8415 5865 8470 5985
rect 8590 5865 8635 5985
rect 8755 5865 8800 5985
rect 8920 5865 8965 5985
rect 9085 5865 9140 5985
rect 9260 5865 9305 5985
rect 9425 5865 9470 5985
rect 9590 5865 9635 5985
rect 9755 5865 9810 5985
rect 9930 5865 9975 5985
rect 10095 5865 10140 5985
rect 10260 5865 10305 5985
rect 10425 5865 10480 5985
rect 10600 5865 10645 5985
rect 10765 5865 10810 5985
rect 10930 5865 10975 5985
rect 11095 5865 11150 5985
rect 11270 5865 11315 5985
rect 11435 5865 11480 5985
rect 11600 5865 11645 5985
rect 11765 5865 11820 5985
rect 11940 5865 11985 5985
rect 12105 5865 12150 5985
rect 12270 5865 12315 5985
rect 12435 5865 12490 5985
rect 12610 5865 12620 5985
rect 7120 5820 12620 5865
rect 7120 5700 7130 5820
rect 7250 5700 7295 5820
rect 7415 5700 7460 5820
rect 7580 5700 7625 5820
rect 7745 5700 7800 5820
rect 7920 5700 7965 5820
rect 8085 5700 8130 5820
rect 8250 5700 8295 5820
rect 8415 5700 8470 5820
rect 8590 5700 8635 5820
rect 8755 5700 8800 5820
rect 8920 5700 8965 5820
rect 9085 5700 9140 5820
rect 9260 5700 9305 5820
rect 9425 5700 9470 5820
rect 9590 5700 9635 5820
rect 9755 5700 9810 5820
rect 9930 5700 9975 5820
rect 10095 5700 10140 5820
rect 10260 5700 10305 5820
rect 10425 5700 10480 5820
rect 10600 5700 10645 5820
rect 10765 5700 10810 5820
rect 10930 5700 10975 5820
rect 11095 5700 11150 5820
rect 11270 5700 11315 5820
rect 11435 5700 11480 5820
rect 11600 5700 11645 5820
rect 11765 5700 11820 5820
rect 11940 5700 11985 5820
rect 12105 5700 12150 5820
rect 12270 5700 12315 5820
rect 12435 5700 12490 5820
rect 12610 5700 12620 5820
rect 7120 5645 12620 5700
rect 7120 5525 7130 5645
rect 7250 5525 7295 5645
rect 7415 5525 7460 5645
rect 7580 5525 7625 5645
rect 7745 5525 7800 5645
rect 7920 5525 7965 5645
rect 8085 5525 8130 5645
rect 8250 5525 8295 5645
rect 8415 5525 8470 5645
rect 8590 5525 8635 5645
rect 8755 5525 8800 5645
rect 8920 5525 8965 5645
rect 9085 5525 9140 5645
rect 9260 5525 9305 5645
rect 9425 5525 9470 5645
rect 9590 5525 9635 5645
rect 9755 5525 9810 5645
rect 9930 5525 9975 5645
rect 10095 5525 10140 5645
rect 10260 5525 10305 5645
rect 10425 5525 10480 5645
rect 10600 5525 10645 5645
rect 10765 5525 10810 5645
rect 10930 5525 10975 5645
rect 11095 5525 11150 5645
rect 11270 5525 11315 5645
rect 11435 5525 11480 5645
rect 11600 5525 11645 5645
rect 11765 5525 11820 5645
rect 11940 5525 11985 5645
rect 12105 5525 12150 5645
rect 12270 5525 12315 5645
rect 12435 5525 12490 5645
rect 12610 5525 12620 5645
rect 7120 5480 12620 5525
rect 7120 5360 7130 5480
rect 7250 5360 7295 5480
rect 7415 5360 7460 5480
rect 7580 5360 7625 5480
rect 7745 5360 7800 5480
rect 7920 5360 7965 5480
rect 8085 5360 8130 5480
rect 8250 5360 8295 5480
rect 8415 5360 8470 5480
rect 8590 5360 8635 5480
rect 8755 5360 8800 5480
rect 8920 5360 8965 5480
rect 9085 5360 9140 5480
rect 9260 5360 9305 5480
rect 9425 5360 9470 5480
rect 9590 5360 9635 5480
rect 9755 5360 9810 5480
rect 9930 5360 9975 5480
rect 10095 5360 10140 5480
rect 10260 5360 10305 5480
rect 10425 5360 10480 5480
rect 10600 5360 10645 5480
rect 10765 5360 10810 5480
rect 10930 5360 10975 5480
rect 11095 5360 11150 5480
rect 11270 5360 11315 5480
rect 11435 5360 11480 5480
rect 11600 5360 11645 5480
rect 11765 5360 11820 5480
rect 11940 5360 11985 5480
rect 12105 5360 12150 5480
rect 12270 5360 12315 5480
rect 12435 5360 12490 5480
rect 12610 5360 12620 5480
rect 7120 5315 12620 5360
rect 7120 5195 7130 5315
rect 7250 5195 7295 5315
rect 7415 5195 7460 5315
rect 7580 5195 7625 5315
rect 7745 5195 7800 5315
rect 7920 5195 7965 5315
rect 8085 5195 8130 5315
rect 8250 5195 8295 5315
rect 8415 5195 8470 5315
rect 8590 5195 8635 5315
rect 8755 5195 8800 5315
rect 8920 5195 8965 5315
rect 9085 5195 9140 5315
rect 9260 5195 9305 5315
rect 9425 5195 9470 5315
rect 9590 5195 9635 5315
rect 9755 5195 9810 5315
rect 9930 5195 9975 5315
rect 10095 5195 10140 5315
rect 10260 5195 10305 5315
rect 10425 5195 10480 5315
rect 10600 5195 10645 5315
rect 10765 5195 10810 5315
rect 10930 5195 10975 5315
rect 11095 5195 11150 5315
rect 11270 5195 11315 5315
rect 11435 5195 11480 5315
rect 11600 5195 11645 5315
rect 11765 5195 11820 5315
rect 11940 5195 11985 5315
rect 12105 5195 12150 5315
rect 12270 5195 12315 5315
rect 12435 5195 12490 5315
rect 12610 5195 12620 5315
rect 7120 5150 12620 5195
rect 7120 5030 7130 5150
rect 7250 5030 7295 5150
rect 7415 5030 7460 5150
rect 7580 5030 7625 5150
rect 7745 5030 7800 5150
rect 7920 5030 7965 5150
rect 8085 5030 8130 5150
rect 8250 5030 8295 5150
rect 8415 5030 8470 5150
rect 8590 5030 8635 5150
rect 8755 5030 8800 5150
rect 8920 5030 8965 5150
rect 9085 5030 9140 5150
rect 9260 5030 9305 5150
rect 9425 5030 9470 5150
rect 9590 5030 9635 5150
rect 9755 5030 9810 5150
rect 9930 5030 9975 5150
rect 10095 5030 10140 5150
rect 10260 5030 10305 5150
rect 10425 5030 10480 5150
rect 10600 5030 10645 5150
rect 10765 5030 10810 5150
rect 10930 5030 10975 5150
rect 11095 5030 11150 5150
rect 11270 5030 11315 5150
rect 11435 5030 11480 5150
rect 11600 5030 11645 5150
rect 11765 5030 11820 5150
rect 11940 5030 11985 5150
rect 12105 5030 12150 5150
rect 12270 5030 12315 5150
rect 12435 5030 12490 5150
rect 12610 5030 12620 5150
rect 7120 4975 12620 5030
rect 7120 4855 7130 4975
rect 7250 4855 7295 4975
rect 7415 4855 7460 4975
rect 7580 4855 7625 4975
rect 7745 4855 7800 4975
rect 7920 4855 7965 4975
rect 8085 4855 8130 4975
rect 8250 4855 8295 4975
rect 8415 4855 8470 4975
rect 8590 4855 8635 4975
rect 8755 4855 8800 4975
rect 8920 4855 8965 4975
rect 9085 4855 9140 4975
rect 9260 4855 9305 4975
rect 9425 4855 9470 4975
rect 9590 4855 9635 4975
rect 9755 4855 9810 4975
rect 9930 4855 9975 4975
rect 10095 4855 10140 4975
rect 10260 4855 10305 4975
rect 10425 4855 10480 4975
rect 10600 4855 10645 4975
rect 10765 4855 10810 4975
rect 10930 4855 10975 4975
rect 11095 4855 11150 4975
rect 11270 4855 11315 4975
rect 11435 4855 11480 4975
rect 11600 4855 11645 4975
rect 11765 4855 11820 4975
rect 11940 4855 11985 4975
rect 12105 4855 12150 4975
rect 12270 4855 12315 4975
rect 12435 4855 12490 4975
rect 12610 4855 12620 4975
rect 7120 4810 12620 4855
rect 7120 4690 7130 4810
rect 7250 4690 7295 4810
rect 7415 4690 7460 4810
rect 7580 4690 7625 4810
rect 7745 4690 7800 4810
rect 7920 4690 7965 4810
rect 8085 4690 8130 4810
rect 8250 4690 8295 4810
rect 8415 4690 8470 4810
rect 8590 4690 8635 4810
rect 8755 4690 8800 4810
rect 8920 4690 8965 4810
rect 9085 4690 9140 4810
rect 9260 4690 9305 4810
rect 9425 4690 9470 4810
rect 9590 4690 9635 4810
rect 9755 4690 9810 4810
rect 9930 4690 9975 4810
rect 10095 4690 10140 4810
rect 10260 4690 10305 4810
rect 10425 4690 10480 4810
rect 10600 4690 10645 4810
rect 10765 4690 10810 4810
rect 10930 4690 10975 4810
rect 11095 4690 11150 4810
rect 11270 4690 11315 4810
rect 11435 4690 11480 4810
rect 11600 4690 11645 4810
rect 11765 4690 11820 4810
rect 11940 4690 11985 4810
rect 12105 4690 12150 4810
rect 12270 4690 12315 4810
rect 12435 4690 12490 4810
rect 12610 4690 12620 4810
rect 7120 4645 12620 4690
rect 7120 4525 7130 4645
rect 7250 4525 7295 4645
rect 7415 4525 7460 4645
rect 7580 4525 7625 4645
rect 7745 4525 7800 4645
rect 7920 4525 7965 4645
rect 8085 4525 8130 4645
rect 8250 4525 8295 4645
rect 8415 4525 8470 4645
rect 8590 4525 8635 4645
rect 8755 4525 8800 4645
rect 8920 4525 8965 4645
rect 9085 4525 9140 4645
rect 9260 4525 9305 4645
rect 9425 4525 9470 4645
rect 9590 4525 9635 4645
rect 9755 4525 9810 4645
rect 9930 4525 9975 4645
rect 10095 4525 10140 4645
rect 10260 4525 10305 4645
rect 10425 4525 10480 4645
rect 10600 4525 10645 4645
rect 10765 4525 10810 4645
rect 10930 4525 10975 4645
rect 11095 4525 11150 4645
rect 11270 4525 11315 4645
rect 11435 4525 11480 4645
rect 11600 4525 11645 4645
rect 11765 4525 11820 4645
rect 11940 4525 11985 4645
rect 12105 4525 12150 4645
rect 12270 4525 12315 4645
rect 12435 4525 12490 4645
rect 12610 4525 12620 4645
rect 7120 4480 12620 4525
rect 7120 4360 7130 4480
rect 7250 4360 7295 4480
rect 7415 4360 7460 4480
rect 7580 4360 7625 4480
rect 7745 4360 7800 4480
rect 7920 4360 7965 4480
rect 8085 4360 8130 4480
rect 8250 4360 8295 4480
rect 8415 4360 8470 4480
rect 8590 4360 8635 4480
rect 8755 4360 8800 4480
rect 8920 4360 8965 4480
rect 9085 4360 9140 4480
rect 9260 4360 9305 4480
rect 9425 4360 9470 4480
rect 9590 4360 9635 4480
rect 9755 4360 9810 4480
rect 9930 4360 9975 4480
rect 10095 4360 10140 4480
rect 10260 4360 10305 4480
rect 10425 4360 10480 4480
rect 10600 4360 10645 4480
rect 10765 4360 10810 4480
rect 10930 4360 10975 4480
rect 11095 4360 11150 4480
rect 11270 4360 11315 4480
rect 11435 4360 11480 4480
rect 11600 4360 11645 4480
rect 11765 4360 11820 4480
rect 11940 4360 11985 4480
rect 12105 4360 12150 4480
rect 12270 4360 12315 4480
rect 12435 4360 12490 4480
rect 12610 4360 12620 4480
rect 7120 4305 12620 4360
rect 7120 4185 7130 4305
rect 7250 4185 7295 4305
rect 7415 4185 7460 4305
rect 7580 4185 7625 4305
rect 7745 4185 7800 4305
rect 7920 4185 7965 4305
rect 8085 4185 8130 4305
rect 8250 4185 8295 4305
rect 8415 4185 8470 4305
rect 8590 4185 8635 4305
rect 8755 4185 8800 4305
rect 8920 4185 8965 4305
rect 9085 4185 9140 4305
rect 9260 4185 9305 4305
rect 9425 4185 9470 4305
rect 9590 4185 9635 4305
rect 9755 4185 9810 4305
rect 9930 4185 9975 4305
rect 10095 4185 10140 4305
rect 10260 4185 10305 4305
rect 10425 4185 10480 4305
rect 10600 4185 10645 4305
rect 10765 4185 10810 4305
rect 10930 4185 10975 4305
rect 11095 4185 11150 4305
rect 11270 4185 11315 4305
rect 11435 4185 11480 4305
rect 11600 4185 11645 4305
rect 11765 4185 11820 4305
rect 11940 4185 11985 4305
rect 12105 4185 12150 4305
rect 12270 4185 12315 4305
rect 12435 4185 12490 4305
rect 12610 4185 12620 4305
rect 7120 4140 12620 4185
rect 7120 4020 7130 4140
rect 7250 4020 7295 4140
rect 7415 4020 7460 4140
rect 7580 4020 7625 4140
rect 7745 4020 7800 4140
rect 7920 4020 7965 4140
rect 8085 4020 8130 4140
rect 8250 4020 8295 4140
rect 8415 4020 8470 4140
rect 8590 4020 8635 4140
rect 8755 4020 8800 4140
rect 8920 4020 8965 4140
rect 9085 4020 9140 4140
rect 9260 4020 9305 4140
rect 9425 4020 9470 4140
rect 9590 4020 9635 4140
rect 9755 4020 9810 4140
rect 9930 4020 9975 4140
rect 10095 4020 10140 4140
rect 10260 4020 10305 4140
rect 10425 4020 10480 4140
rect 10600 4020 10645 4140
rect 10765 4020 10810 4140
rect 10930 4020 10975 4140
rect 11095 4020 11150 4140
rect 11270 4020 11315 4140
rect 11435 4020 11480 4140
rect 11600 4020 11645 4140
rect 11765 4020 11820 4140
rect 11940 4020 11985 4140
rect 12105 4020 12150 4140
rect 12270 4020 12315 4140
rect 12435 4020 12490 4140
rect 12610 4020 12620 4140
rect 7120 3975 12620 4020
rect 7120 3855 7130 3975
rect 7250 3855 7295 3975
rect 7415 3855 7460 3975
rect 7580 3855 7625 3975
rect 7745 3855 7800 3975
rect 7920 3855 7965 3975
rect 8085 3855 8130 3975
rect 8250 3855 8295 3975
rect 8415 3855 8470 3975
rect 8590 3855 8635 3975
rect 8755 3855 8800 3975
rect 8920 3855 8965 3975
rect 9085 3855 9140 3975
rect 9260 3855 9305 3975
rect 9425 3855 9470 3975
rect 9590 3855 9635 3975
rect 9755 3855 9810 3975
rect 9930 3855 9975 3975
rect 10095 3855 10140 3975
rect 10260 3855 10305 3975
rect 10425 3855 10480 3975
rect 10600 3855 10645 3975
rect 10765 3855 10810 3975
rect 10930 3855 10975 3975
rect 11095 3855 11150 3975
rect 11270 3855 11315 3975
rect 11435 3855 11480 3975
rect 11600 3855 11645 3975
rect 11765 3855 11820 3975
rect 11940 3855 11985 3975
rect 12105 3855 12150 3975
rect 12270 3855 12315 3975
rect 12435 3855 12490 3975
rect 12610 3855 12620 3975
rect 7120 3810 12620 3855
rect 7120 3690 7130 3810
rect 7250 3690 7295 3810
rect 7415 3690 7460 3810
rect 7580 3690 7625 3810
rect 7745 3690 7800 3810
rect 7920 3690 7965 3810
rect 8085 3690 8130 3810
rect 8250 3690 8295 3810
rect 8415 3690 8470 3810
rect 8590 3690 8635 3810
rect 8755 3690 8800 3810
rect 8920 3690 8965 3810
rect 9085 3690 9140 3810
rect 9260 3690 9305 3810
rect 9425 3690 9470 3810
rect 9590 3690 9635 3810
rect 9755 3690 9810 3810
rect 9930 3690 9975 3810
rect 10095 3690 10140 3810
rect 10260 3690 10305 3810
rect 10425 3690 10480 3810
rect 10600 3690 10645 3810
rect 10765 3690 10810 3810
rect 10930 3690 10975 3810
rect 11095 3690 11150 3810
rect 11270 3690 11315 3810
rect 11435 3690 11480 3810
rect 11600 3690 11645 3810
rect 11765 3690 11820 3810
rect 11940 3690 11985 3810
rect 12105 3690 12150 3810
rect 12270 3690 12315 3810
rect 12435 3690 12490 3810
rect 12610 3690 12620 3810
rect 7120 3635 12620 3690
rect 7120 3515 7130 3635
rect 7250 3515 7295 3635
rect 7415 3515 7460 3635
rect 7580 3515 7625 3635
rect 7745 3515 7800 3635
rect 7920 3515 7965 3635
rect 8085 3515 8130 3635
rect 8250 3515 8295 3635
rect 8415 3515 8470 3635
rect 8590 3515 8635 3635
rect 8755 3515 8800 3635
rect 8920 3515 8965 3635
rect 9085 3515 9140 3635
rect 9260 3515 9305 3635
rect 9425 3515 9470 3635
rect 9590 3515 9635 3635
rect 9755 3515 9810 3635
rect 9930 3515 9975 3635
rect 10095 3515 10140 3635
rect 10260 3515 10305 3635
rect 10425 3515 10480 3635
rect 10600 3515 10645 3635
rect 10765 3515 10810 3635
rect 10930 3515 10975 3635
rect 11095 3515 11150 3635
rect 11270 3515 11315 3635
rect 11435 3515 11480 3635
rect 11600 3515 11645 3635
rect 11765 3515 11820 3635
rect 11940 3515 11985 3635
rect 12105 3515 12150 3635
rect 12270 3515 12315 3635
rect 12435 3515 12490 3635
rect 12610 3515 12620 3635
rect 7120 3470 12620 3515
rect 7120 3350 7130 3470
rect 7250 3350 7295 3470
rect 7415 3350 7460 3470
rect 7580 3350 7625 3470
rect 7745 3350 7800 3470
rect 7920 3350 7965 3470
rect 8085 3350 8130 3470
rect 8250 3350 8295 3470
rect 8415 3350 8470 3470
rect 8590 3350 8635 3470
rect 8755 3350 8800 3470
rect 8920 3350 8965 3470
rect 9085 3350 9140 3470
rect 9260 3350 9305 3470
rect 9425 3350 9470 3470
rect 9590 3350 9635 3470
rect 9755 3350 9810 3470
rect 9930 3350 9975 3470
rect 10095 3350 10140 3470
rect 10260 3350 10305 3470
rect 10425 3350 10480 3470
rect 10600 3350 10645 3470
rect 10765 3350 10810 3470
rect 10930 3350 10975 3470
rect 11095 3350 11150 3470
rect 11270 3350 11315 3470
rect 11435 3350 11480 3470
rect 11600 3350 11645 3470
rect 11765 3350 11820 3470
rect 11940 3350 11985 3470
rect 12105 3350 12150 3470
rect 12270 3350 12315 3470
rect 12435 3350 12490 3470
rect 12610 3350 12620 3470
rect 7120 3305 12620 3350
rect 7120 3185 7130 3305
rect 7250 3185 7295 3305
rect 7415 3185 7460 3305
rect 7580 3185 7625 3305
rect 7745 3185 7800 3305
rect 7920 3185 7965 3305
rect 8085 3185 8130 3305
rect 8250 3185 8295 3305
rect 8415 3185 8470 3305
rect 8590 3185 8635 3305
rect 8755 3185 8800 3305
rect 8920 3185 8965 3305
rect 9085 3185 9140 3305
rect 9260 3185 9305 3305
rect 9425 3185 9470 3305
rect 9590 3185 9635 3305
rect 9755 3185 9810 3305
rect 9930 3185 9975 3305
rect 10095 3185 10140 3305
rect 10260 3185 10305 3305
rect 10425 3185 10480 3305
rect 10600 3185 10645 3305
rect 10765 3185 10810 3305
rect 10930 3185 10975 3305
rect 11095 3185 11150 3305
rect 11270 3185 11315 3305
rect 11435 3185 11480 3305
rect 11600 3185 11645 3305
rect 11765 3185 11820 3305
rect 11940 3185 11985 3305
rect 12105 3185 12150 3305
rect 12270 3185 12315 3305
rect 12435 3185 12490 3305
rect 12610 3185 12620 3305
rect 7120 3140 12620 3185
rect 7120 3020 7130 3140
rect 7250 3020 7295 3140
rect 7415 3020 7460 3140
rect 7580 3020 7625 3140
rect 7745 3020 7800 3140
rect 7920 3020 7965 3140
rect 8085 3020 8130 3140
rect 8250 3020 8295 3140
rect 8415 3020 8470 3140
rect 8590 3020 8635 3140
rect 8755 3020 8800 3140
rect 8920 3020 8965 3140
rect 9085 3020 9140 3140
rect 9260 3020 9305 3140
rect 9425 3020 9470 3140
rect 9590 3020 9635 3140
rect 9755 3020 9810 3140
rect 9930 3020 9975 3140
rect 10095 3020 10140 3140
rect 10260 3020 10305 3140
rect 10425 3020 10480 3140
rect 10600 3020 10645 3140
rect 10765 3020 10810 3140
rect 10930 3020 10975 3140
rect 11095 3020 11150 3140
rect 11270 3020 11315 3140
rect 11435 3020 11480 3140
rect 11600 3020 11645 3140
rect 11765 3020 11820 3140
rect 11940 3020 11985 3140
rect 12105 3020 12150 3140
rect 12270 3020 12315 3140
rect 12435 3020 12490 3140
rect 12610 3020 12620 3140
rect 7120 2965 12620 3020
rect 7120 2845 7130 2965
rect 7250 2845 7295 2965
rect 7415 2845 7460 2965
rect 7580 2845 7625 2965
rect 7745 2845 7800 2965
rect 7920 2845 7965 2965
rect 8085 2845 8130 2965
rect 8250 2845 8295 2965
rect 8415 2845 8470 2965
rect 8590 2845 8635 2965
rect 8755 2845 8800 2965
rect 8920 2845 8965 2965
rect 9085 2845 9140 2965
rect 9260 2845 9305 2965
rect 9425 2845 9470 2965
rect 9590 2845 9635 2965
rect 9755 2845 9810 2965
rect 9930 2845 9975 2965
rect 10095 2845 10140 2965
rect 10260 2845 10305 2965
rect 10425 2845 10480 2965
rect 10600 2845 10645 2965
rect 10765 2845 10810 2965
rect 10930 2845 10975 2965
rect 11095 2845 11150 2965
rect 11270 2845 11315 2965
rect 11435 2845 11480 2965
rect 11600 2845 11645 2965
rect 11765 2845 11820 2965
rect 11940 2845 11985 2965
rect 12105 2845 12150 2965
rect 12270 2845 12315 2965
rect 12435 2845 12490 2965
rect 12610 2845 12620 2965
rect 7120 2800 12620 2845
rect 7120 2680 7130 2800
rect 7250 2680 7295 2800
rect 7415 2680 7460 2800
rect 7580 2680 7625 2800
rect 7745 2680 7800 2800
rect 7920 2680 7965 2800
rect 8085 2680 8130 2800
rect 8250 2680 8295 2800
rect 8415 2680 8470 2800
rect 8590 2680 8635 2800
rect 8755 2680 8800 2800
rect 8920 2680 8965 2800
rect 9085 2680 9140 2800
rect 9260 2680 9305 2800
rect 9425 2680 9470 2800
rect 9590 2680 9635 2800
rect 9755 2680 9810 2800
rect 9930 2680 9975 2800
rect 10095 2680 10140 2800
rect 10260 2680 10305 2800
rect 10425 2680 10480 2800
rect 10600 2680 10645 2800
rect 10765 2680 10810 2800
rect 10930 2680 10975 2800
rect 11095 2680 11150 2800
rect 11270 2680 11315 2800
rect 11435 2680 11480 2800
rect 11600 2680 11645 2800
rect 11765 2680 11820 2800
rect 11940 2680 11985 2800
rect 12105 2680 12150 2800
rect 12270 2680 12315 2800
rect 12435 2680 12490 2800
rect 12610 2680 12620 2800
rect 7120 2635 12620 2680
rect 7120 2515 7130 2635
rect 7250 2515 7295 2635
rect 7415 2515 7460 2635
rect 7580 2515 7625 2635
rect 7745 2515 7800 2635
rect 7920 2515 7965 2635
rect 8085 2515 8130 2635
rect 8250 2515 8295 2635
rect 8415 2515 8470 2635
rect 8590 2515 8635 2635
rect 8755 2515 8800 2635
rect 8920 2515 8965 2635
rect 9085 2515 9140 2635
rect 9260 2515 9305 2635
rect 9425 2515 9470 2635
rect 9590 2515 9635 2635
rect 9755 2515 9810 2635
rect 9930 2515 9975 2635
rect 10095 2515 10140 2635
rect 10260 2515 10305 2635
rect 10425 2515 10480 2635
rect 10600 2515 10645 2635
rect 10765 2515 10810 2635
rect 10930 2515 10975 2635
rect 11095 2515 11150 2635
rect 11270 2515 11315 2635
rect 11435 2515 11480 2635
rect 11600 2515 11645 2635
rect 11765 2515 11820 2635
rect 11940 2515 11985 2635
rect 12105 2515 12150 2635
rect 12270 2515 12315 2635
rect 12435 2515 12490 2635
rect 12610 2515 12620 2635
rect 7120 2470 12620 2515
rect 7120 2350 7130 2470
rect 7250 2350 7295 2470
rect 7415 2350 7460 2470
rect 7580 2350 7625 2470
rect 7745 2350 7800 2470
rect 7920 2350 7965 2470
rect 8085 2350 8130 2470
rect 8250 2350 8295 2470
rect 8415 2350 8470 2470
rect 8590 2350 8635 2470
rect 8755 2350 8800 2470
rect 8920 2350 8965 2470
rect 9085 2350 9140 2470
rect 9260 2350 9305 2470
rect 9425 2350 9470 2470
rect 9590 2350 9635 2470
rect 9755 2350 9810 2470
rect 9930 2350 9975 2470
rect 10095 2350 10140 2470
rect 10260 2350 10305 2470
rect 10425 2350 10480 2470
rect 10600 2350 10645 2470
rect 10765 2350 10810 2470
rect 10930 2350 10975 2470
rect 11095 2350 11150 2470
rect 11270 2350 11315 2470
rect 11435 2350 11480 2470
rect 11600 2350 11645 2470
rect 11765 2350 11820 2470
rect 11940 2350 11985 2470
rect 12105 2350 12150 2470
rect 12270 2350 12315 2470
rect 12435 2350 12490 2470
rect 12610 2350 12620 2470
rect 7120 2295 12620 2350
rect 7120 2175 7130 2295
rect 7250 2175 7295 2295
rect 7415 2175 7460 2295
rect 7580 2175 7625 2295
rect 7745 2175 7800 2295
rect 7920 2175 7965 2295
rect 8085 2175 8130 2295
rect 8250 2175 8295 2295
rect 8415 2175 8470 2295
rect 8590 2175 8635 2295
rect 8755 2175 8800 2295
rect 8920 2175 8965 2295
rect 9085 2175 9140 2295
rect 9260 2175 9305 2295
rect 9425 2175 9470 2295
rect 9590 2175 9635 2295
rect 9755 2175 9810 2295
rect 9930 2175 9975 2295
rect 10095 2175 10140 2295
rect 10260 2175 10305 2295
rect 10425 2175 10480 2295
rect 10600 2175 10645 2295
rect 10765 2175 10810 2295
rect 10930 2175 10975 2295
rect 11095 2175 11150 2295
rect 11270 2175 11315 2295
rect 11435 2175 11480 2295
rect 11600 2175 11645 2295
rect 11765 2175 11820 2295
rect 11940 2175 11985 2295
rect 12105 2175 12150 2295
rect 12270 2175 12315 2295
rect 12435 2175 12490 2295
rect 12610 2175 12620 2295
rect 7120 2130 12620 2175
rect 7120 2010 7130 2130
rect 7250 2010 7295 2130
rect 7415 2010 7460 2130
rect 7580 2010 7625 2130
rect 7745 2010 7800 2130
rect 7920 2010 7965 2130
rect 8085 2010 8130 2130
rect 8250 2010 8295 2130
rect 8415 2010 8470 2130
rect 8590 2010 8635 2130
rect 8755 2010 8800 2130
rect 8920 2010 8965 2130
rect 9085 2010 9140 2130
rect 9260 2010 9305 2130
rect 9425 2010 9470 2130
rect 9590 2010 9635 2130
rect 9755 2010 9810 2130
rect 9930 2010 9975 2130
rect 10095 2010 10140 2130
rect 10260 2010 10305 2130
rect 10425 2010 10480 2130
rect 10600 2010 10645 2130
rect 10765 2010 10810 2130
rect 10930 2010 10975 2130
rect 11095 2010 11150 2130
rect 11270 2010 11315 2130
rect 11435 2010 11480 2130
rect 11600 2010 11645 2130
rect 11765 2010 11820 2130
rect 11940 2010 11985 2130
rect 12105 2010 12150 2130
rect 12270 2010 12315 2130
rect 12435 2010 12490 2130
rect 12610 2010 12620 2130
rect 7120 1965 12620 2010
rect 7120 1845 7130 1965
rect 7250 1845 7295 1965
rect 7415 1845 7460 1965
rect 7580 1845 7625 1965
rect 7745 1845 7800 1965
rect 7920 1845 7965 1965
rect 8085 1845 8130 1965
rect 8250 1845 8295 1965
rect 8415 1845 8470 1965
rect 8590 1845 8635 1965
rect 8755 1845 8800 1965
rect 8920 1845 8965 1965
rect 9085 1845 9140 1965
rect 9260 1845 9305 1965
rect 9425 1845 9470 1965
rect 9590 1845 9635 1965
rect 9755 1845 9810 1965
rect 9930 1845 9975 1965
rect 10095 1845 10140 1965
rect 10260 1845 10305 1965
rect 10425 1845 10480 1965
rect 10600 1845 10645 1965
rect 10765 1845 10810 1965
rect 10930 1845 10975 1965
rect 11095 1845 11150 1965
rect 11270 1845 11315 1965
rect 11435 1845 11480 1965
rect 11600 1845 11645 1965
rect 11765 1845 11820 1965
rect 11940 1845 11985 1965
rect 12105 1845 12150 1965
rect 12270 1845 12315 1965
rect 12435 1845 12490 1965
rect 12610 1845 12620 1965
rect 7120 1800 12620 1845
rect 7120 1680 7130 1800
rect 7250 1680 7295 1800
rect 7415 1680 7460 1800
rect 7580 1680 7625 1800
rect 7745 1680 7800 1800
rect 7920 1680 7965 1800
rect 8085 1680 8130 1800
rect 8250 1680 8295 1800
rect 8415 1680 8470 1800
rect 8590 1680 8635 1800
rect 8755 1680 8800 1800
rect 8920 1680 8965 1800
rect 9085 1680 9140 1800
rect 9260 1680 9305 1800
rect 9425 1680 9470 1800
rect 9590 1680 9635 1800
rect 9755 1680 9810 1800
rect 9930 1680 9975 1800
rect 10095 1680 10140 1800
rect 10260 1680 10305 1800
rect 10425 1680 10480 1800
rect 10600 1680 10645 1800
rect 10765 1680 10810 1800
rect 10930 1680 10975 1800
rect 11095 1680 11150 1800
rect 11270 1680 11315 1800
rect 11435 1680 11480 1800
rect 11600 1680 11645 1800
rect 11765 1680 11820 1800
rect 11940 1680 11985 1800
rect 12105 1680 12150 1800
rect 12270 1680 12315 1800
rect 12435 1680 12490 1800
rect 12610 1680 12620 1800
rect 7120 1670 12620 1680
rect 12810 7160 18310 7170
rect 12810 7040 12820 7160
rect 12940 7040 12985 7160
rect 13105 7040 13150 7160
rect 13270 7040 13315 7160
rect 13435 7040 13490 7160
rect 13610 7040 13655 7160
rect 13775 7040 13820 7160
rect 13940 7040 13985 7160
rect 14105 7040 14160 7160
rect 14280 7040 14325 7160
rect 14445 7040 14490 7160
rect 14610 7040 14655 7160
rect 14775 7040 14830 7160
rect 14950 7040 14995 7160
rect 15115 7040 15160 7160
rect 15280 7040 15325 7160
rect 15445 7040 15500 7160
rect 15620 7040 15665 7160
rect 15785 7040 15830 7160
rect 15950 7040 15995 7160
rect 16115 7040 16170 7160
rect 16290 7040 16335 7160
rect 16455 7040 16500 7160
rect 16620 7040 16665 7160
rect 16785 7040 16840 7160
rect 16960 7040 17005 7160
rect 17125 7040 17170 7160
rect 17290 7040 17335 7160
rect 17455 7040 17510 7160
rect 17630 7040 17675 7160
rect 17795 7040 17840 7160
rect 17960 7040 18005 7160
rect 18125 7040 18180 7160
rect 18300 7040 18310 7160
rect 12810 6985 18310 7040
rect 12810 6865 12820 6985
rect 12940 6865 12985 6985
rect 13105 6865 13150 6985
rect 13270 6865 13315 6985
rect 13435 6865 13490 6985
rect 13610 6865 13655 6985
rect 13775 6865 13820 6985
rect 13940 6865 13985 6985
rect 14105 6865 14160 6985
rect 14280 6865 14325 6985
rect 14445 6865 14490 6985
rect 14610 6865 14655 6985
rect 14775 6865 14830 6985
rect 14950 6865 14995 6985
rect 15115 6865 15160 6985
rect 15280 6865 15325 6985
rect 15445 6865 15500 6985
rect 15620 6865 15665 6985
rect 15785 6865 15830 6985
rect 15950 6865 15995 6985
rect 16115 6865 16170 6985
rect 16290 6865 16335 6985
rect 16455 6865 16500 6985
rect 16620 6865 16665 6985
rect 16785 6865 16840 6985
rect 16960 6865 17005 6985
rect 17125 6865 17170 6985
rect 17290 6865 17335 6985
rect 17455 6865 17510 6985
rect 17630 6865 17675 6985
rect 17795 6865 17840 6985
rect 17960 6865 18005 6985
rect 18125 6865 18180 6985
rect 18300 6865 18310 6985
rect 12810 6820 18310 6865
rect 12810 6700 12820 6820
rect 12940 6700 12985 6820
rect 13105 6700 13150 6820
rect 13270 6700 13315 6820
rect 13435 6700 13490 6820
rect 13610 6700 13655 6820
rect 13775 6700 13820 6820
rect 13940 6700 13985 6820
rect 14105 6700 14160 6820
rect 14280 6700 14325 6820
rect 14445 6700 14490 6820
rect 14610 6700 14655 6820
rect 14775 6700 14830 6820
rect 14950 6700 14995 6820
rect 15115 6700 15160 6820
rect 15280 6700 15325 6820
rect 15445 6700 15500 6820
rect 15620 6700 15665 6820
rect 15785 6700 15830 6820
rect 15950 6700 15995 6820
rect 16115 6700 16170 6820
rect 16290 6700 16335 6820
rect 16455 6700 16500 6820
rect 16620 6700 16665 6820
rect 16785 6700 16840 6820
rect 16960 6700 17005 6820
rect 17125 6700 17170 6820
rect 17290 6700 17335 6820
rect 17455 6700 17510 6820
rect 17630 6700 17675 6820
rect 17795 6700 17840 6820
rect 17960 6700 18005 6820
rect 18125 6700 18180 6820
rect 18300 6700 18310 6820
rect 12810 6655 18310 6700
rect 12810 6535 12820 6655
rect 12940 6535 12985 6655
rect 13105 6535 13150 6655
rect 13270 6535 13315 6655
rect 13435 6535 13490 6655
rect 13610 6535 13655 6655
rect 13775 6535 13820 6655
rect 13940 6535 13985 6655
rect 14105 6535 14160 6655
rect 14280 6535 14325 6655
rect 14445 6535 14490 6655
rect 14610 6535 14655 6655
rect 14775 6535 14830 6655
rect 14950 6535 14995 6655
rect 15115 6535 15160 6655
rect 15280 6535 15325 6655
rect 15445 6535 15500 6655
rect 15620 6535 15665 6655
rect 15785 6535 15830 6655
rect 15950 6535 15995 6655
rect 16115 6535 16170 6655
rect 16290 6535 16335 6655
rect 16455 6535 16500 6655
rect 16620 6535 16665 6655
rect 16785 6535 16840 6655
rect 16960 6535 17005 6655
rect 17125 6535 17170 6655
rect 17290 6535 17335 6655
rect 17455 6535 17510 6655
rect 17630 6535 17675 6655
rect 17795 6535 17840 6655
rect 17960 6535 18005 6655
rect 18125 6535 18180 6655
rect 18300 6535 18310 6655
rect 12810 6490 18310 6535
rect 12810 6370 12820 6490
rect 12940 6370 12985 6490
rect 13105 6370 13150 6490
rect 13270 6370 13315 6490
rect 13435 6370 13490 6490
rect 13610 6370 13655 6490
rect 13775 6370 13820 6490
rect 13940 6370 13985 6490
rect 14105 6370 14160 6490
rect 14280 6370 14325 6490
rect 14445 6370 14490 6490
rect 14610 6370 14655 6490
rect 14775 6370 14830 6490
rect 14950 6370 14995 6490
rect 15115 6370 15160 6490
rect 15280 6370 15325 6490
rect 15445 6370 15500 6490
rect 15620 6370 15665 6490
rect 15785 6370 15830 6490
rect 15950 6370 15995 6490
rect 16115 6370 16170 6490
rect 16290 6370 16335 6490
rect 16455 6370 16500 6490
rect 16620 6370 16665 6490
rect 16785 6370 16840 6490
rect 16960 6370 17005 6490
rect 17125 6370 17170 6490
rect 17290 6370 17335 6490
rect 17455 6370 17510 6490
rect 17630 6370 17675 6490
rect 17795 6370 17840 6490
rect 17960 6370 18005 6490
rect 18125 6370 18180 6490
rect 18300 6370 18310 6490
rect 12810 6315 18310 6370
rect 12810 6195 12820 6315
rect 12940 6195 12985 6315
rect 13105 6195 13150 6315
rect 13270 6195 13315 6315
rect 13435 6195 13490 6315
rect 13610 6195 13655 6315
rect 13775 6195 13820 6315
rect 13940 6195 13985 6315
rect 14105 6195 14160 6315
rect 14280 6195 14325 6315
rect 14445 6195 14490 6315
rect 14610 6195 14655 6315
rect 14775 6195 14830 6315
rect 14950 6195 14995 6315
rect 15115 6195 15160 6315
rect 15280 6195 15325 6315
rect 15445 6195 15500 6315
rect 15620 6195 15665 6315
rect 15785 6195 15830 6315
rect 15950 6195 15995 6315
rect 16115 6195 16170 6315
rect 16290 6195 16335 6315
rect 16455 6195 16500 6315
rect 16620 6195 16665 6315
rect 16785 6195 16840 6315
rect 16960 6195 17005 6315
rect 17125 6195 17170 6315
rect 17290 6195 17335 6315
rect 17455 6195 17510 6315
rect 17630 6195 17675 6315
rect 17795 6195 17840 6315
rect 17960 6195 18005 6315
rect 18125 6195 18180 6315
rect 18300 6195 18310 6315
rect 12810 6150 18310 6195
rect 12810 6030 12820 6150
rect 12940 6030 12985 6150
rect 13105 6030 13150 6150
rect 13270 6030 13315 6150
rect 13435 6030 13490 6150
rect 13610 6030 13655 6150
rect 13775 6030 13820 6150
rect 13940 6030 13985 6150
rect 14105 6030 14160 6150
rect 14280 6030 14325 6150
rect 14445 6030 14490 6150
rect 14610 6030 14655 6150
rect 14775 6030 14830 6150
rect 14950 6030 14995 6150
rect 15115 6030 15160 6150
rect 15280 6030 15325 6150
rect 15445 6030 15500 6150
rect 15620 6030 15665 6150
rect 15785 6030 15830 6150
rect 15950 6030 15995 6150
rect 16115 6030 16170 6150
rect 16290 6030 16335 6150
rect 16455 6030 16500 6150
rect 16620 6030 16665 6150
rect 16785 6030 16840 6150
rect 16960 6030 17005 6150
rect 17125 6030 17170 6150
rect 17290 6030 17335 6150
rect 17455 6030 17510 6150
rect 17630 6030 17675 6150
rect 17795 6030 17840 6150
rect 17960 6030 18005 6150
rect 18125 6030 18180 6150
rect 18300 6030 18310 6150
rect 12810 5985 18310 6030
rect 12810 5865 12820 5985
rect 12940 5865 12985 5985
rect 13105 5865 13150 5985
rect 13270 5865 13315 5985
rect 13435 5865 13490 5985
rect 13610 5865 13655 5985
rect 13775 5865 13820 5985
rect 13940 5865 13985 5985
rect 14105 5865 14160 5985
rect 14280 5865 14325 5985
rect 14445 5865 14490 5985
rect 14610 5865 14655 5985
rect 14775 5865 14830 5985
rect 14950 5865 14995 5985
rect 15115 5865 15160 5985
rect 15280 5865 15325 5985
rect 15445 5865 15500 5985
rect 15620 5865 15665 5985
rect 15785 5865 15830 5985
rect 15950 5865 15995 5985
rect 16115 5865 16170 5985
rect 16290 5865 16335 5985
rect 16455 5865 16500 5985
rect 16620 5865 16665 5985
rect 16785 5865 16840 5985
rect 16960 5865 17005 5985
rect 17125 5865 17170 5985
rect 17290 5865 17335 5985
rect 17455 5865 17510 5985
rect 17630 5865 17675 5985
rect 17795 5865 17840 5985
rect 17960 5865 18005 5985
rect 18125 5865 18180 5985
rect 18300 5865 18310 5985
rect 12810 5820 18310 5865
rect 12810 5700 12820 5820
rect 12940 5700 12985 5820
rect 13105 5700 13150 5820
rect 13270 5700 13315 5820
rect 13435 5700 13490 5820
rect 13610 5700 13655 5820
rect 13775 5700 13820 5820
rect 13940 5700 13985 5820
rect 14105 5700 14160 5820
rect 14280 5700 14325 5820
rect 14445 5700 14490 5820
rect 14610 5700 14655 5820
rect 14775 5700 14830 5820
rect 14950 5700 14995 5820
rect 15115 5700 15160 5820
rect 15280 5700 15325 5820
rect 15445 5700 15500 5820
rect 15620 5700 15665 5820
rect 15785 5700 15830 5820
rect 15950 5700 15995 5820
rect 16115 5700 16170 5820
rect 16290 5700 16335 5820
rect 16455 5700 16500 5820
rect 16620 5700 16665 5820
rect 16785 5700 16840 5820
rect 16960 5700 17005 5820
rect 17125 5700 17170 5820
rect 17290 5700 17335 5820
rect 17455 5700 17510 5820
rect 17630 5700 17675 5820
rect 17795 5700 17840 5820
rect 17960 5700 18005 5820
rect 18125 5700 18180 5820
rect 18300 5700 18310 5820
rect 12810 5645 18310 5700
rect 12810 5525 12820 5645
rect 12940 5525 12985 5645
rect 13105 5525 13150 5645
rect 13270 5525 13315 5645
rect 13435 5525 13490 5645
rect 13610 5525 13655 5645
rect 13775 5525 13820 5645
rect 13940 5525 13985 5645
rect 14105 5525 14160 5645
rect 14280 5525 14325 5645
rect 14445 5525 14490 5645
rect 14610 5525 14655 5645
rect 14775 5525 14830 5645
rect 14950 5525 14995 5645
rect 15115 5525 15160 5645
rect 15280 5525 15325 5645
rect 15445 5525 15500 5645
rect 15620 5525 15665 5645
rect 15785 5525 15830 5645
rect 15950 5525 15995 5645
rect 16115 5525 16170 5645
rect 16290 5525 16335 5645
rect 16455 5525 16500 5645
rect 16620 5525 16665 5645
rect 16785 5525 16840 5645
rect 16960 5525 17005 5645
rect 17125 5525 17170 5645
rect 17290 5525 17335 5645
rect 17455 5525 17510 5645
rect 17630 5525 17675 5645
rect 17795 5525 17840 5645
rect 17960 5525 18005 5645
rect 18125 5525 18180 5645
rect 18300 5525 18310 5645
rect 12810 5480 18310 5525
rect 12810 5360 12820 5480
rect 12940 5360 12985 5480
rect 13105 5360 13150 5480
rect 13270 5360 13315 5480
rect 13435 5360 13490 5480
rect 13610 5360 13655 5480
rect 13775 5360 13820 5480
rect 13940 5360 13985 5480
rect 14105 5360 14160 5480
rect 14280 5360 14325 5480
rect 14445 5360 14490 5480
rect 14610 5360 14655 5480
rect 14775 5360 14830 5480
rect 14950 5360 14995 5480
rect 15115 5360 15160 5480
rect 15280 5360 15325 5480
rect 15445 5360 15500 5480
rect 15620 5360 15665 5480
rect 15785 5360 15830 5480
rect 15950 5360 15995 5480
rect 16115 5360 16170 5480
rect 16290 5360 16335 5480
rect 16455 5360 16500 5480
rect 16620 5360 16665 5480
rect 16785 5360 16840 5480
rect 16960 5360 17005 5480
rect 17125 5360 17170 5480
rect 17290 5360 17335 5480
rect 17455 5360 17510 5480
rect 17630 5360 17675 5480
rect 17795 5360 17840 5480
rect 17960 5360 18005 5480
rect 18125 5360 18180 5480
rect 18300 5360 18310 5480
rect 12810 5315 18310 5360
rect 12810 5195 12820 5315
rect 12940 5195 12985 5315
rect 13105 5195 13150 5315
rect 13270 5195 13315 5315
rect 13435 5195 13490 5315
rect 13610 5195 13655 5315
rect 13775 5195 13820 5315
rect 13940 5195 13985 5315
rect 14105 5195 14160 5315
rect 14280 5195 14325 5315
rect 14445 5195 14490 5315
rect 14610 5195 14655 5315
rect 14775 5195 14830 5315
rect 14950 5195 14995 5315
rect 15115 5195 15160 5315
rect 15280 5195 15325 5315
rect 15445 5195 15500 5315
rect 15620 5195 15665 5315
rect 15785 5195 15830 5315
rect 15950 5195 15995 5315
rect 16115 5195 16170 5315
rect 16290 5195 16335 5315
rect 16455 5195 16500 5315
rect 16620 5195 16665 5315
rect 16785 5195 16840 5315
rect 16960 5195 17005 5315
rect 17125 5195 17170 5315
rect 17290 5195 17335 5315
rect 17455 5195 17510 5315
rect 17630 5195 17675 5315
rect 17795 5195 17840 5315
rect 17960 5195 18005 5315
rect 18125 5195 18180 5315
rect 18300 5195 18310 5315
rect 12810 5150 18310 5195
rect 12810 5030 12820 5150
rect 12940 5030 12985 5150
rect 13105 5030 13150 5150
rect 13270 5030 13315 5150
rect 13435 5030 13490 5150
rect 13610 5030 13655 5150
rect 13775 5030 13820 5150
rect 13940 5030 13985 5150
rect 14105 5030 14160 5150
rect 14280 5030 14325 5150
rect 14445 5030 14490 5150
rect 14610 5030 14655 5150
rect 14775 5030 14830 5150
rect 14950 5030 14995 5150
rect 15115 5030 15160 5150
rect 15280 5030 15325 5150
rect 15445 5030 15500 5150
rect 15620 5030 15665 5150
rect 15785 5030 15830 5150
rect 15950 5030 15995 5150
rect 16115 5030 16170 5150
rect 16290 5030 16335 5150
rect 16455 5030 16500 5150
rect 16620 5030 16665 5150
rect 16785 5030 16840 5150
rect 16960 5030 17005 5150
rect 17125 5030 17170 5150
rect 17290 5030 17335 5150
rect 17455 5030 17510 5150
rect 17630 5030 17675 5150
rect 17795 5030 17840 5150
rect 17960 5030 18005 5150
rect 18125 5030 18180 5150
rect 18300 5030 18310 5150
rect 12810 4975 18310 5030
rect 12810 4855 12820 4975
rect 12940 4855 12985 4975
rect 13105 4855 13150 4975
rect 13270 4855 13315 4975
rect 13435 4855 13490 4975
rect 13610 4855 13655 4975
rect 13775 4855 13820 4975
rect 13940 4855 13985 4975
rect 14105 4855 14160 4975
rect 14280 4855 14325 4975
rect 14445 4855 14490 4975
rect 14610 4855 14655 4975
rect 14775 4855 14830 4975
rect 14950 4855 14995 4975
rect 15115 4855 15160 4975
rect 15280 4855 15325 4975
rect 15445 4855 15500 4975
rect 15620 4855 15665 4975
rect 15785 4855 15830 4975
rect 15950 4855 15995 4975
rect 16115 4855 16170 4975
rect 16290 4855 16335 4975
rect 16455 4855 16500 4975
rect 16620 4855 16665 4975
rect 16785 4855 16840 4975
rect 16960 4855 17005 4975
rect 17125 4855 17170 4975
rect 17290 4855 17335 4975
rect 17455 4855 17510 4975
rect 17630 4855 17675 4975
rect 17795 4855 17840 4975
rect 17960 4855 18005 4975
rect 18125 4855 18180 4975
rect 18300 4855 18310 4975
rect 12810 4810 18310 4855
rect 12810 4690 12820 4810
rect 12940 4690 12985 4810
rect 13105 4690 13150 4810
rect 13270 4690 13315 4810
rect 13435 4690 13490 4810
rect 13610 4690 13655 4810
rect 13775 4690 13820 4810
rect 13940 4690 13985 4810
rect 14105 4690 14160 4810
rect 14280 4690 14325 4810
rect 14445 4690 14490 4810
rect 14610 4690 14655 4810
rect 14775 4690 14830 4810
rect 14950 4690 14995 4810
rect 15115 4690 15160 4810
rect 15280 4690 15325 4810
rect 15445 4690 15500 4810
rect 15620 4690 15665 4810
rect 15785 4690 15830 4810
rect 15950 4690 15995 4810
rect 16115 4690 16170 4810
rect 16290 4690 16335 4810
rect 16455 4690 16500 4810
rect 16620 4690 16665 4810
rect 16785 4690 16840 4810
rect 16960 4690 17005 4810
rect 17125 4690 17170 4810
rect 17290 4690 17335 4810
rect 17455 4690 17510 4810
rect 17630 4690 17675 4810
rect 17795 4690 17840 4810
rect 17960 4690 18005 4810
rect 18125 4690 18180 4810
rect 18300 4690 18310 4810
rect 12810 4645 18310 4690
rect 12810 4525 12820 4645
rect 12940 4525 12985 4645
rect 13105 4525 13150 4645
rect 13270 4525 13315 4645
rect 13435 4525 13490 4645
rect 13610 4525 13655 4645
rect 13775 4525 13820 4645
rect 13940 4525 13985 4645
rect 14105 4525 14160 4645
rect 14280 4525 14325 4645
rect 14445 4525 14490 4645
rect 14610 4525 14655 4645
rect 14775 4525 14830 4645
rect 14950 4525 14995 4645
rect 15115 4525 15160 4645
rect 15280 4525 15325 4645
rect 15445 4525 15500 4645
rect 15620 4525 15665 4645
rect 15785 4525 15830 4645
rect 15950 4525 15995 4645
rect 16115 4525 16170 4645
rect 16290 4525 16335 4645
rect 16455 4525 16500 4645
rect 16620 4525 16665 4645
rect 16785 4525 16840 4645
rect 16960 4525 17005 4645
rect 17125 4525 17170 4645
rect 17290 4525 17335 4645
rect 17455 4525 17510 4645
rect 17630 4525 17675 4645
rect 17795 4525 17840 4645
rect 17960 4525 18005 4645
rect 18125 4525 18180 4645
rect 18300 4525 18310 4645
rect 12810 4480 18310 4525
rect 12810 4360 12820 4480
rect 12940 4360 12985 4480
rect 13105 4360 13150 4480
rect 13270 4360 13315 4480
rect 13435 4360 13490 4480
rect 13610 4360 13655 4480
rect 13775 4360 13820 4480
rect 13940 4360 13985 4480
rect 14105 4360 14160 4480
rect 14280 4360 14325 4480
rect 14445 4360 14490 4480
rect 14610 4360 14655 4480
rect 14775 4360 14830 4480
rect 14950 4360 14995 4480
rect 15115 4360 15160 4480
rect 15280 4360 15325 4480
rect 15445 4360 15500 4480
rect 15620 4360 15665 4480
rect 15785 4360 15830 4480
rect 15950 4360 15995 4480
rect 16115 4360 16170 4480
rect 16290 4360 16335 4480
rect 16455 4360 16500 4480
rect 16620 4360 16665 4480
rect 16785 4360 16840 4480
rect 16960 4360 17005 4480
rect 17125 4360 17170 4480
rect 17290 4360 17335 4480
rect 17455 4360 17510 4480
rect 17630 4360 17675 4480
rect 17795 4360 17840 4480
rect 17960 4360 18005 4480
rect 18125 4360 18180 4480
rect 18300 4360 18310 4480
rect 12810 4305 18310 4360
rect 12810 4185 12820 4305
rect 12940 4185 12985 4305
rect 13105 4185 13150 4305
rect 13270 4185 13315 4305
rect 13435 4185 13490 4305
rect 13610 4185 13655 4305
rect 13775 4185 13820 4305
rect 13940 4185 13985 4305
rect 14105 4185 14160 4305
rect 14280 4185 14325 4305
rect 14445 4185 14490 4305
rect 14610 4185 14655 4305
rect 14775 4185 14830 4305
rect 14950 4185 14995 4305
rect 15115 4185 15160 4305
rect 15280 4185 15325 4305
rect 15445 4185 15500 4305
rect 15620 4185 15665 4305
rect 15785 4185 15830 4305
rect 15950 4185 15995 4305
rect 16115 4185 16170 4305
rect 16290 4185 16335 4305
rect 16455 4185 16500 4305
rect 16620 4185 16665 4305
rect 16785 4185 16840 4305
rect 16960 4185 17005 4305
rect 17125 4185 17170 4305
rect 17290 4185 17335 4305
rect 17455 4185 17510 4305
rect 17630 4185 17675 4305
rect 17795 4185 17840 4305
rect 17960 4185 18005 4305
rect 18125 4185 18180 4305
rect 18300 4185 18310 4305
rect 12810 4140 18310 4185
rect 12810 4020 12820 4140
rect 12940 4020 12985 4140
rect 13105 4020 13150 4140
rect 13270 4020 13315 4140
rect 13435 4020 13490 4140
rect 13610 4020 13655 4140
rect 13775 4020 13820 4140
rect 13940 4020 13985 4140
rect 14105 4020 14160 4140
rect 14280 4020 14325 4140
rect 14445 4020 14490 4140
rect 14610 4020 14655 4140
rect 14775 4020 14830 4140
rect 14950 4020 14995 4140
rect 15115 4020 15160 4140
rect 15280 4020 15325 4140
rect 15445 4020 15500 4140
rect 15620 4020 15665 4140
rect 15785 4020 15830 4140
rect 15950 4020 15995 4140
rect 16115 4020 16170 4140
rect 16290 4020 16335 4140
rect 16455 4020 16500 4140
rect 16620 4020 16665 4140
rect 16785 4020 16840 4140
rect 16960 4020 17005 4140
rect 17125 4020 17170 4140
rect 17290 4020 17335 4140
rect 17455 4020 17510 4140
rect 17630 4020 17675 4140
rect 17795 4020 17840 4140
rect 17960 4020 18005 4140
rect 18125 4020 18180 4140
rect 18300 4020 18310 4140
rect 12810 3975 18310 4020
rect 12810 3855 12820 3975
rect 12940 3855 12985 3975
rect 13105 3855 13150 3975
rect 13270 3855 13315 3975
rect 13435 3855 13490 3975
rect 13610 3855 13655 3975
rect 13775 3855 13820 3975
rect 13940 3855 13985 3975
rect 14105 3855 14160 3975
rect 14280 3855 14325 3975
rect 14445 3855 14490 3975
rect 14610 3855 14655 3975
rect 14775 3855 14830 3975
rect 14950 3855 14995 3975
rect 15115 3855 15160 3975
rect 15280 3855 15325 3975
rect 15445 3855 15500 3975
rect 15620 3855 15665 3975
rect 15785 3855 15830 3975
rect 15950 3855 15995 3975
rect 16115 3855 16170 3975
rect 16290 3855 16335 3975
rect 16455 3855 16500 3975
rect 16620 3855 16665 3975
rect 16785 3855 16840 3975
rect 16960 3855 17005 3975
rect 17125 3855 17170 3975
rect 17290 3855 17335 3975
rect 17455 3855 17510 3975
rect 17630 3855 17675 3975
rect 17795 3855 17840 3975
rect 17960 3855 18005 3975
rect 18125 3855 18180 3975
rect 18300 3855 18310 3975
rect 12810 3810 18310 3855
rect 12810 3690 12820 3810
rect 12940 3690 12985 3810
rect 13105 3690 13150 3810
rect 13270 3690 13315 3810
rect 13435 3690 13490 3810
rect 13610 3690 13655 3810
rect 13775 3690 13820 3810
rect 13940 3690 13985 3810
rect 14105 3690 14160 3810
rect 14280 3690 14325 3810
rect 14445 3690 14490 3810
rect 14610 3690 14655 3810
rect 14775 3690 14830 3810
rect 14950 3690 14995 3810
rect 15115 3690 15160 3810
rect 15280 3690 15325 3810
rect 15445 3690 15500 3810
rect 15620 3690 15665 3810
rect 15785 3690 15830 3810
rect 15950 3690 15995 3810
rect 16115 3690 16170 3810
rect 16290 3690 16335 3810
rect 16455 3690 16500 3810
rect 16620 3690 16665 3810
rect 16785 3690 16840 3810
rect 16960 3690 17005 3810
rect 17125 3690 17170 3810
rect 17290 3690 17335 3810
rect 17455 3690 17510 3810
rect 17630 3690 17675 3810
rect 17795 3690 17840 3810
rect 17960 3690 18005 3810
rect 18125 3690 18180 3810
rect 18300 3690 18310 3810
rect 12810 3635 18310 3690
rect 12810 3515 12820 3635
rect 12940 3515 12985 3635
rect 13105 3515 13150 3635
rect 13270 3515 13315 3635
rect 13435 3515 13490 3635
rect 13610 3515 13655 3635
rect 13775 3515 13820 3635
rect 13940 3515 13985 3635
rect 14105 3515 14160 3635
rect 14280 3515 14325 3635
rect 14445 3515 14490 3635
rect 14610 3515 14655 3635
rect 14775 3515 14830 3635
rect 14950 3515 14995 3635
rect 15115 3515 15160 3635
rect 15280 3515 15325 3635
rect 15445 3515 15500 3635
rect 15620 3515 15665 3635
rect 15785 3515 15830 3635
rect 15950 3515 15995 3635
rect 16115 3515 16170 3635
rect 16290 3515 16335 3635
rect 16455 3515 16500 3635
rect 16620 3515 16665 3635
rect 16785 3515 16840 3635
rect 16960 3515 17005 3635
rect 17125 3515 17170 3635
rect 17290 3515 17335 3635
rect 17455 3515 17510 3635
rect 17630 3515 17675 3635
rect 17795 3515 17840 3635
rect 17960 3515 18005 3635
rect 18125 3515 18180 3635
rect 18300 3515 18310 3635
rect 12810 3470 18310 3515
rect 12810 3350 12820 3470
rect 12940 3350 12985 3470
rect 13105 3350 13150 3470
rect 13270 3350 13315 3470
rect 13435 3350 13490 3470
rect 13610 3350 13655 3470
rect 13775 3350 13820 3470
rect 13940 3350 13985 3470
rect 14105 3350 14160 3470
rect 14280 3350 14325 3470
rect 14445 3350 14490 3470
rect 14610 3350 14655 3470
rect 14775 3350 14830 3470
rect 14950 3350 14995 3470
rect 15115 3350 15160 3470
rect 15280 3350 15325 3470
rect 15445 3350 15500 3470
rect 15620 3350 15665 3470
rect 15785 3350 15830 3470
rect 15950 3350 15995 3470
rect 16115 3350 16170 3470
rect 16290 3350 16335 3470
rect 16455 3350 16500 3470
rect 16620 3350 16665 3470
rect 16785 3350 16840 3470
rect 16960 3350 17005 3470
rect 17125 3350 17170 3470
rect 17290 3350 17335 3470
rect 17455 3350 17510 3470
rect 17630 3350 17675 3470
rect 17795 3350 17840 3470
rect 17960 3350 18005 3470
rect 18125 3350 18180 3470
rect 18300 3350 18310 3470
rect 12810 3305 18310 3350
rect 12810 3185 12820 3305
rect 12940 3185 12985 3305
rect 13105 3185 13150 3305
rect 13270 3185 13315 3305
rect 13435 3185 13490 3305
rect 13610 3185 13655 3305
rect 13775 3185 13820 3305
rect 13940 3185 13985 3305
rect 14105 3185 14160 3305
rect 14280 3185 14325 3305
rect 14445 3185 14490 3305
rect 14610 3185 14655 3305
rect 14775 3185 14830 3305
rect 14950 3185 14995 3305
rect 15115 3185 15160 3305
rect 15280 3185 15325 3305
rect 15445 3185 15500 3305
rect 15620 3185 15665 3305
rect 15785 3185 15830 3305
rect 15950 3185 15995 3305
rect 16115 3185 16170 3305
rect 16290 3185 16335 3305
rect 16455 3185 16500 3305
rect 16620 3185 16665 3305
rect 16785 3185 16840 3305
rect 16960 3185 17005 3305
rect 17125 3185 17170 3305
rect 17290 3185 17335 3305
rect 17455 3185 17510 3305
rect 17630 3185 17675 3305
rect 17795 3185 17840 3305
rect 17960 3185 18005 3305
rect 18125 3185 18180 3305
rect 18300 3185 18310 3305
rect 12810 3140 18310 3185
rect 12810 3020 12820 3140
rect 12940 3020 12985 3140
rect 13105 3020 13150 3140
rect 13270 3020 13315 3140
rect 13435 3020 13490 3140
rect 13610 3020 13655 3140
rect 13775 3020 13820 3140
rect 13940 3020 13985 3140
rect 14105 3020 14160 3140
rect 14280 3020 14325 3140
rect 14445 3020 14490 3140
rect 14610 3020 14655 3140
rect 14775 3020 14830 3140
rect 14950 3020 14995 3140
rect 15115 3020 15160 3140
rect 15280 3020 15325 3140
rect 15445 3020 15500 3140
rect 15620 3020 15665 3140
rect 15785 3020 15830 3140
rect 15950 3020 15995 3140
rect 16115 3020 16170 3140
rect 16290 3020 16335 3140
rect 16455 3020 16500 3140
rect 16620 3020 16665 3140
rect 16785 3020 16840 3140
rect 16960 3020 17005 3140
rect 17125 3020 17170 3140
rect 17290 3020 17335 3140
rect 17455 3020 17510 3140
rect 17630 3020 17675 3140
rect 17795 3020 17840 3140
rect 17960 3020 18005 3140
rect 18125 3020 18180 3140
rect 18300 3020 18310 3140
rect 12810 2965 18310 3020
rect 12810 2845 12820 2965
rect 12940 2845 12985 2965
rect 13105 2845 13150 2965
rect 13270 2845 13315 2965
rect 13435 2845 13490 2965
rect 13610 2845 13655 2965
rect 13775 2845 13820 2965
rect 13940 2845 13985 2965
rect 14105 2845 14160 2965
rect 14280 2845 14325 2965
rect 14445 2845 14490 2965
rect 14610 2845 14655 2965
rect 14775 2845 14830 2965
rect 14950 2845 14995 2965
rect 15115 2845 15160 2965
rect 15280 2845 15325 2965
rect 15445 2845 15500 2965
rect 15620 2845 15665 2965
rect 15785 2845 15830 2965
rect 15950 2845 15995 2965
rect 16115 2845 16170 2965
rect 16290 2845 16335 2965
rect 16455 2845 16500 2965
rect 16620 2845 16665 2965
rect 16785 2845 16840 2965
rect 16960 2845 17005 2965
rect 17125 2845 17170 2965
rect 17290 2845 17335 2965
rect 17455 2845 17510 2965
rect 17630 2845 17675 2965
rect 17795 2845 17840 2965
rect 17960 2845 18005 2965
rect 18125 2845 18180 2965
rect 18300 2845 18310 2965
rect 12810 2800 18310 2845
rect 12810 2680 12820 2800
rect 12940 2680 12985 2800
rect 13105 2680 13150 2800
rect 13270 2680 13315 2800
rect 13435 2680 13490 2800
rect 13610 2680 13655 2800
rect 13775 2680 13820 2800
rect 13940 2680 13985 2800
rect 14105 2680 14160 2800
rect 14280 2680 14325 2800
rect 14445 2680 14490 2800
rect 14610 2680 14655 2800
rect 14775 2680 14830 2800
rect 14950 2680 14995 2800
rect 15115 2680 15160 2800
rect 15280 2680 15325 2800
rect 15445 2680 15500 2800
rect 15620 2680 15665 2800
rect 15785 2680 15830 2800
rect 15950 2680 15995 2800
rect 16115 2680 16170 2800
rect 16290 2680 16335 2800
rect 16455 2680 16500 2800
rect 16620 2680 16665 2800
rect 16785 2680 16840 2800
rect 16960 2680 17005 2800
rect 17125 2680 17170 2800
rect 17290 2680 17335 2800
rect 17455 2680 17510 2800
rect 17630 2680 17675 2800
rect 17795 2680 17840 2800
rect 17960 2680 18005 2800
rect 18125 2680 18180 2800
rect 18300 2680 18310 2800
rect 12810 2635 18310 2680
rect 12810 2515 12820 2635
rect 12940 2515 12985 2635
rect 13105 2515 13150 2635
rect 13270 2515 13315 2635
rect 13435 2515 13490 2635
rect 13610 2515 13655 2635
rect 13775 2515 13820 2635
rect 13940 2515 13985 2635
rect 14105 2515 14160 2635
rect 14280 2515 14325 2635
rect 14445 2515 14490 2635
rect 14610 2515 14655 2635
rect 14775 2515 14830 2635
rect 14950 2515 14995 2635
rect 15115 2515 15160 2635
rect 15280 2515 15325 2635
rect 15445 2515 15500 2635
rect 15620 2515 15665 2635
rect 15785 2515 15830 2635
rect 15950 2515 15995 2635
rect 16115 2515 16170 2635
rect 16290 2515 16335 2635
rect 16455 2515 16500 2635
rect 16620 2515 16665 2635
rect 16785 2515 16840 2635
rect 16960 2515 17005 2635
rect 17125 2515 17170 2635
rect 17290 2515 17335 2635
rect 17455 2515 17510 2635
rect 17630 2515 17675 2635
rect 17795 2515 17840 2635
rect 17960 2515 18005 2635
rect 18125 2515 18180 2635
rect 18300 2515 18310 2635
rect 12810 2470 18310 2515
rect 12810 2350 12820 2470
rect 12940 2350 12985 2470
rect 13105 2350 13150 2470
rect 13270 2350 13315 2470
rect 13435 2350 13490 2470
rect 13610 2350 13655 2470
rect 13775 2350 13820 2470
rect 13940 2350 13985 2470
rect 14105 2350 14160 2470
rect 14280 2350 14325 2470
rect 14445 2350 14490 2470
rect 14610 2350 14655 2470
rect 14775 2350 14830 2470
rect 14950 2350 14995 2470
rect 15115 2350 15160 2470
rect 15280 2350 15325 2470
rect 15445 2350 15500 2470
rect 15620 2350 15665 2470
rect 15785 2350 15830 2470
rect 15950 2350 15995 2470
rect 16115 2350 16170 2470
rect 16290 2350 16335 2470
rect 16455 2350 16500 2470
rect 16620 2350 16665 2470
rect 16785 2350 16840 2470
rect 16960 2350 17005 2470
rect 17125 2350 17170 2470
rect 17290 2350 17335 2470
rect 17455 2350 17510 2470
rect 17630 2350 17675 2470
rect 17795 2350 17840 2470
rect 17960 2350 18005 2470
rect 18125 2350 18180 2470
rect 18300 2350 18310 2470
rect 12810 2295 18310 2350
rect 12810 2175 12820 2295
rect 12940 2175 12985 2295
rect 13105 2175 13150 2295
rect 13270 2175 13315 2295
rect 13435 2175 13490 2295
rect 13610 2175 13655 2295
rect 13775 2175 13820 2295
rect 13940 2175 13985 2295
rect 14105 2175 14160 2295
rect 14280 2175 14325 2295
rect 14445 2175 14490 2295
rect 14610 2175 14655 2295
rect 14775 2175 14830 2295
rect 14950 2175 14995 2295
rect 15115 2175 15160 2295
rect 15280 2175 15325 2295
rect 15445 2175 15500 2295
rect 15620 2175 15665 2295
rect 15785 2175 15830 2295
rect 15950 2175 15995 2295
rect 16115 2175 16170 2295
rect 16290 2175 16335 2295
rect 16455 2175 16500 2295
rect 16620 2175 16665 2295
rect 16785 2175 16840 2295
rect 16960 2175 17005 2295
rect 17125 2175 17170 2295
rect 17290 2175 17335 2295
rect 17455 2175 17510 2295
rect 17630 2175 17675 2295
rect 17795 2175 17840 2295
rect 17960 2175 18005 2295
rect 18125 2175 18180 2295
rect 18300 2175 18310 2295
rect 12810 2130 18310 2175
rect 12810 2010 12820 2130
rect 12940 2010 12985 2130
rect 13105 2010 13150 2130
rect 13270 2010 13315 2130
rect 13435 2010 13490 2130
rect 13610 2010 13655 2130
rect 13775 2010 13820 2130
rect 13940 2010 13985 2130
rect 14105 2010 14160 2130
rect 14280 2010 14325 2130
rect 14445 2010 14490 2130
rect 14610 2010 14655 2130
rect 14775 2010 14830 2130
rect 14950 2010 14995 2130
rect 15115 2010 15160 2130
rect 15280 2010 15325 2130
rect 15445 2010 15500 2130
rect 15620 2010 15665 2130
rect 15785 2010 15830 2130
rect 15950 2010 15995 2130
rect 16115 2010 16170 2130
rect 16290 2010 16335 2130
rect 16455 2010 16500 2130
rect 16620 2010 16665 2130
rect 16785 2010 16840 2130
rect 16960 2010 17005 2130
rect 17125 2010 17170 2130
rect 17290 2010 17335 2130
rect 17455 2010 17510 2130
rect 17630 2010 17675 2130
rect 17795 2010 17840 2130
rect 17960 2010 18005 2130
rect 18125 2010 18180 2130
rect 18300 2010 18310 2130
rect 12810 1965 18310 2010
rect 12810 1845 12820 1965
rect 12940 1845 12985 1965
rect 13105 1845 13150 1965
rect 13270 1845 13315 1965
rect 13435 1845 13490 1965
rect 13610 1845 13655 1965
rect 13775 1845 13820 1965
rect 13940 1845 13985 1965
rect 14105 1845 14160 1965
rect 14280 1845 14325 1965
rect 14445 1845 14490 1965
rect 14610 1845 14655 1965
rect 14775 1845 14830 1965
rect 14950 1845 14995 1965
rect 15115 1845 15160 1965
rect 15280 1845 15325 1965
rect 15445 1845 15500 1965
rect 15620 1845 15665 1965
rect 15785 1845 15830 1965
rect 15950 1845 15995 1965
rect 16115 1845 16170 1965
rect 16290 1845 16335 1965
rect 16455 1845 16500 1965
rect 16620 1845 16665 1965
rect 16785 1845 16840 1965
rect 16960 1845 17005 1965
rect 17125 1845 17170 1965
rect 17290 1845 17335 1965
rect 17455 1845 17510 1965
rect 17630 1845 17675 1965
rect 17795 1845 17840 1965
rect 17960 1845 18005 1965
rect 18125 1845 18180 1965
rect 18300 1845 18310 1965
rect 12810 1800 18310 1845
rect 12810 1680 12820 1800
rect 12940 1680 12985 1800
rect 13105 1680 13150 1800
rect 13270 1680 13315 1800
rect 13435 1680 13490 1800
rect 13610 1680 13655 1800
rect 13775 1680 13820 1800
rect 13940 1680 13985 1800
rect 14105 1680 14160 1800
rect 14280 1680 14325 1800
rect 14445 1680 14490 1800
rect 14610 1680 14655 1800
rect 14775 1680 14830 1800
rect 14950 1680 14995 1800
rect 15115 1680 15160 1800
rect 15280 1680 15325 1800
rect 15445 1680 15500 1800
rect 15620 1680 15665 1800
rect 15785 1680 15830 1800
rect 15950 1680 15995 1800
rect 16115 1680 16170 1800
rect 16290 1680 16335 1800
rect 16455 1680 16500 1800
rect 16620 1680 16665 1800
rect 16785 1680 16840 1800
rect 16960 1680 17005 1800
rect 17125 1680 17170 1800
rect 17290 1680 17335 1800
rect 17455 1680 17510 1800
rect 17630 1680 17675 1800
rect 17795 1680 17840 1800
rect 17960 1680 18005 1800
rect 18125 1680 18180 1800
rect 18300 1680 18310 1800
rect 12810 1670 18310 1680
rect 18500 7160 24000 7170
rect 18500 7040 18510 7160
rect 18630 7040 18675 7160
rect 18795 7040 18840 7160
rect 18960 7040 19005 7160
rect 19125 7040 19180 7160
rect 19300 7040 19345 7160
rect 19465 7040 19510 7160
rect 19630 7040 19675 7160
rect 19795 7040 19850 7160
rect 19970 7040 20015 7160
rect 20135 7040 20180 7160
rect 20300 7040 20345 7160
rect 20465 7040 20520 7160
rect 20640 7040 20685 7160
rect 20805 7040 20850 7160
rect 20970 7040 21015 7160
rect 21135 7040 21190 7160
rect 21310 7040 21355 7160
rect 21475 7040 21520 7160
rect 21640 7040 21685 7160
rect 21805 7040 21860 7160
rect 21980 7040 22025 7160
rect 22145 7040 22190 7160
rect 22310 7040 22355 7160
rect 22475 7040 22530 7160
rect 22650 7040 22695 7160
rect 22815 7040 22860 7160
rect 22980 7040 23025 7160
rect 23145 7040 23200 7160
rect 23320 7040 23365 7160
rect 23485 7040 23530 7160
rect 23650 7040 23695 7160
rect 23815 7040 23870 7160
rect 23990 7040 24000 7160
rect 18500 6985 24000 7040
rect 18500 6865 18510 6985
rect 18630 6865 18675 6985
rect 18795 6865 18840 6985
rect 18960 6865 19005 6985
rect 19125 6865 19180 6985
rect 19300 6865 19345 6985
rect 19465 6865 19510 6985
rect 19630 6865 19675 6985
rect 19795 6865 19850 6985
rect 19970 6865 20015 6985
rect 20135 6865 20180 6985
rect 20300 6865 20345 6985
rect 20465 6865 20520 6985
rect 20640 6865 20685 6985
rect 20805 6865 20850 6985
rect 20970 6865 21015 6985
rect 21135 6865 21190 6985
rect 21310 6865 21355 6985
rect 21475 6865 21520 6985
rect 21640 6865 21685 6985
rect 21805 6865 21860 6985
rect 21980 6865 22025 6985
rect 22145 6865 22190 6985
rect 22310 6865 22355 6985
rect 22475 6865 22530 6985
rect 22650 6865 22695 6985
rect 22815 6865 22860 6985
rect 22980 6865 23025 6985
rect 23145 6865 23200 6985
rect 23320 6865 23365 6985
rect 23485 6865 23530 6985
rect 23650 6865 23695 6985
rect 23815 6865 23870 6985
rect 23990 6865 24000 6985
rect 18500 6820 24000 6865
rect 18500 6700 18510 6820
rect 18630 6700 18675 6820
rect 18795 6700 18840 6820
rect 18960 6700 19005 6820
rect 19125 6700 19180 6820
rect 19300 6700 19345 6820
rect 19465 6700 19510 6820
rect 19630 6700 19675 6820
rect 19795 6700 19850 6820
rect 19970 6700 20015 6820
rect 20135 6700 20180 6820
rect 20300 6700 20345 6820
rect 20465 6700 20520 6820
rect 20640 6700 20685 6820
rect 20805 6700 20850 6820
rect 20970 6700 21015 6820
rect 21135 6700 21190 6820
rect 21310 6700 21355 6820
rect 21475 6700 21520 6820
rect 21640 6700 21685 6820
rect 21805 6700 21860 6820
rect 21980 6700 22025 6820
rect 22145 6700 22190 6820
rect 22310 6700 22355 6820
rect 22475 6700 22530 6820
rect 22650 6700 22695 6820
rect 22815 6700 22860 6820
rect 22980 6700 23025 6820
rect 23145 6700 23200 6820
rect 23320 6700 23365 6820
rect 23485 6700 23530 6820
rect 23650 6700 23695 6820
rect 23815 6700 23870 6820
rect 23990 6700 24000 6820
rect 18500 6655 24000 6700
rect 18500 6535 18510 6655
rect 18630 6535 18675 6655
rect 18795 6535 18840 6655
rect 18960 6535 19005 6655
rect 19125 6535 19180 6655
rect 19300 6535 19345 6655
rect 19465 6535 19510 6655
rect 19630 6535 19675 6655
rect 19795 6535 19850 6655
rect 19970 6535 20015 6655
rect 20135 6535 20180 6655
rect 20300 6535 20345 6655
rect 20465 6535 20520 6655
rect 20640 6535 20685 6655
rect 20805 6535 20850 6655
rect 20970 6535 21015 6655
rect 21135 6535 21190 6655
rect 21310 6535 21355 6655
rect 21475 6535 21520 6655
rect 21640 6535 21685 6655
rect 21805 6535 21860 6655
rect 21980 6535 22025 6655
rect 22145 6535 22190 6655
rect 22310 6535 22355 6655
rect 22475 6535 22530 6655
rect 22650 6535 22695 6655
rect 22815 6535 22860 6655
rect 22980 6535 23025 6655
rect 23145 6535 23200 6655
rect 23320 6535 23365 6655
rect 23485 6535 23530 6655
rect 23650 6535 23695 6655
rect 23815 6535 23870 6655
rect 23990 6535 24000 6655
rect 18500 6490 24000 6535
rect 18500 6370 18510 6490
rect 18630 6370 18675 6490
rect 18795 6370 18840 6490
rect 18960 6370 19005 6490
rect 19125 6370 19180 6490
rect 19300 6370 19345 6490
rect 19465 6370 19510 6490
rect 19630 6370 19675 6490
rect 19795 6370 19850 6490
rect 19970 6370 20015 6490
rect 20135 6370 20180 6490
rect 20300 6370 20345 6490
rect 20465 6370 20520 6490
rect 20640 6370 20685 6490
rect 20805 6370 20850 6490
rect 20970 6370 21015 6490
rect 21135 6370 21190 6490
rect 21310 6370 21355 6490
rect 21475 6370 21520 6490
rect 21640 6370 21685 6490
rect 21805 6370 21860 6490
rect 21980 6370 22025 6490
rect 22145 6370 22190 6490
rect 22310 6370 22355 6490
rect 22475 6370 22530 6490
rect 22650 6370 22695 6490
rect 22815 6370 22860 6490
rect 22980 6370 23025 6490
rect 23145 6370 23200 6490
rect 23320 6370 23365 6490
rect 23485 6370 23530 6490
rect 23650 6370 23695 6490
rect 23815 6370 23870 6490
rect 23990 6370 24000 6490
rect 18500 6315 24000 6370
rect 18500 6195 18510 6315
rect 18630 6195 18675 6315
rect 18795 6195 18840 6315
rect 18960 6195 19005 6315
rect 19125 6195 19180 6315
rect 19300 6195 19345 6315
rect 19465 6195 19510 6315
rect 19630 6195 19675 6315
rect 19795 6195 19850 6315
rect 19970 6195 20015 6315
rect 20135 6195 20180 6315
rect 20300 6195 20345 6315
rect 20465 6195 20520 6315
rect 20640 6195 20685 6315
rect 20805 6195 20850 6315
rect 20970 6195 21015 6315
rect 21135 6195 21190 6315
rect 21310 6195 21355 6315
rect 21475 6195 21520 6315
rect 21640 6195 21685 6315
rect 21805 6195 21860 6315
rect 21980 6195 22025 6315
rect 22145 6195 22190 6315
rect 22310 6195 22355 6315
rect 22475 6195 22530 6315
rect 22650 6195 22695 6315
rect 22815 6195 22860 6315
rect 22980 6195 23025 6315
rect 23145 6195 23200 6315
rect 23320 6195 23365 6315
rect 23485 6195 23530 6315
rect 23650 6195 23695 6315
rect 23815 6195 23870 6315
rect 23990 6195 24000 6315
rect 18500 6150 24000 6195
rect 18500 6030 18510 6150
rect 18630 6030 18675 6150
rect 18795 6030 18840 6150
rect 18960 6030 19005 6150
rect 19125 6030 19180 6150
rect 19300 6030 19345 6150
rect 19465 6030 19510 6150
rect 19630 6030 19675 6150
rect 19795 6030 19850 6150
rect 19970 6030 20015 6150
rect 20135 6030 20180 6150
rect 20300 6030 20345 6150
rect 20465 6030 20520 6150
rect 20640 6030 20685 6150
rect 20805 6030 20850 6150
rect 20970 6030 21015 6150
rect 21135 6030 21190 6150
rect 21310 6030 21355 6150
rect 21475 6030 21520 6150
rect 21640 6030 21685 6150
rect 21805 6030 21860 6150
rect 21980 6030 22025 6150
rect 22145 6030 22190 6150
rect 22310 6030 22355 6150
rect 22475 6030 22530 6150
rect 22650 6030 22695 6150
rect 22815 6030 22860 6150
rect 22980 6030 23025 6150
rect 23145 6030 23200 6150
rect 23320 6030 23365 6150
rect 23485 6030 23530 6150
rect 23650 6030 23695 6150
rect 23815 6030 23870 6150
rect 23990 6030 24000 6150
rect 18500 5985 24000 6030
rect 18500 5865 18510 5985
rect 18630 5865 18675 5985
rect 18795 5865 18840 5985
rect 18960 5865 19005 5985
rect 19125 5865 19180 5985
rect 19300 5865 19345 5985
rect 19465 5865 19510 5985
rect 19630 5865 19675 5985
rect 19795 5865 19850 5985
rect 19970 5865 20015 5985
rect 20135 5865 20180 5985
rect 20300 5865 20345 5985
rect 20465 5865 20520 5985
rect 20640 5865 20685 5985
rect 20805 5865 20850 5985
rect 20970 5865 21015 5985
rect 21135 5865 21190 5985
rect 21310 5865 21355 5985
rect 21475 5865 21520 5985
rect 21640 5865 21685 5985
rect 21805 5865 21860 5985
rect 21980 5865 22025 5985
rect 22145 5865 22190 5985
rect 22310 5865 22355 5985
rect 22475 5865 22530 5985
rect 22650 5865 22695 5985
rect 22815 5865 22860 5985
rect 22980 5865 23025 5985
rect 23145 5865 23200 5985
rect 23320 5865 23365 5985
rect 23485 5865 23530 5985
rect 23650 5865 23695 5985
rect 23815 5865 23870 5985
rect 23990 5865 24000 5985
rect 18500 5820 24000 5865
rect 18500 5700 18510 5820
rect 18630 5700 18675 5820
rect 18795 5700 18840 5820
rect 18960 5700 19005 5820
rect 19125 5700 19180 5820
rect 19300 5700 19345 5820
rect 19465 5700 19510 5820
rect 19630 5700 19675 5820
rect 19795 5700 19850 5820
rect 19970 5700 20015 5820
rect 20135 5700 20180 5820
rect 20300 5700 20345 5820
rect 20465 5700 20520 5820
rect 20640 5700 20685 5820
rect 20805 5700 20850 5820
rect 20970 5700 21015 5820
rect 21135 5700 21190 5820
rect 21310 5700 21355 5820
rect 21475 5700 21520 5820
rect 21640 5700 21685 5820
rect 21805 5700 21860 5820
rect 21980 5700 22025 5820
rect 22145 5700 22190 5820
rect 22310 5700 22355 5820
rect 22475 5700 22530 5820
rect 22650 5700 22695 5820
rect 22815 5700 22860 5820
rect 22980 5700 23025 5820
rect 23145 5700 23200 5820
rect 23320 5700 23365 5820
rect 23485 5700 23530 5820
rect 23650 5700 23695 5820
rect 23815 5700 23870 5820
rect 23990 5700 24000 5820
rect 18500 5645 24000 5700
rect 18500 5525 18510 5645
rect 18630 5525 18675 5645
rect 18795 5525 18840 5645
rect 18960 5525 19005 5645
rect 19125 5525 19180 5645
rect 19300 5525 19345 5645
rect 19465 5525 19510 5645
rect 19630 5525 19675 5645
rect 19795 5525 19850 5645
rect 19970 5525 20015 5645
rect 20135 5525 20180 5645
rect 20300 5525 20345 5645
rect 20465 5525 20520 5645
rect 20640 5525 20685 5645
rect 20805 5525 20850 5645
rect 20970 5525 21015 5645
rect 21135 5525 21190 5645
rect 21310 5525 21355 5645
rect 21475 5525 21520 5645
rect 21640 5525 21685 5645
rect 21805 5525 21860 5645
rect 21980 5525 22025 5645
rect 22145 5525 22190 5645
rect 22310 5525 22355 5645
rect 22475 5525 22530 5645
rect 22650 5525 22695 5645
rect 22815 5525 22860 5645
rect 22980 5525 23025 5645
rect 23145 5525 23200 5645
rect 23320 5525 23365 5645
rect 23485 5525 23530 5645
rect 23650 5525 23695 5645
rect 23815 5525 23870 5645
rect 23990 5525 24000 5645
rect 18500 5480 24000 5525
rect 18500 5360 18510 5480
rect 18630 5360 18675 5480
rect 18795 5360 18840 5480
rect 18960 5360 19005 5480
rect 19125 5360 19180 5480
rect 19300 5360 19345 5480
rect 19465 5360 19510 5480
rect 19630 5360 19675 5480
rect 19795 5360 19850 5480
rect 19970 5360 20015 5480
rect 20135 5360 20180 5480
rect 20300 5360 20345 5480
rect 20465 5360 20520 5480
rect 20640 5360 20685 5480
rect 20805 5360 20850 5480
rect 20970 5360 21015 5480
rect 21135 5360 21190 5480
rect 21310 5360 21355 5480
rect 21475 5360 21520 5480
rect 21640 5360 21685 5480
rect 21805 5360 21860 5480
rect 21980 5360 22025 5480
rect 22145 5360 22190 5480
rect 22310 5360 22355 5480
rect 22475 5360 22530 5480
rect 22650 5360 22695 5480
rect 22815 5360 22860 5480
rect 22980 5360 23025 5480
rect 23145 5360 23200 5480
rect 23320 5360 23365 5480
rect 23485 5360 23530 5480
rect 23650 5360 23695 5480
rect 23815 5360 23870 5480
rect 23990 5360 24000 5480
rect 18500 5315 24000 5360
rect 18500 5195 18510 5315
rect 18630 5195 18675 5315
rect 18795 5195 18840 5315
rect 18960 5195 19005 5315
rect 19125 5195 19180 5315
rect 19300 5195 19345 5315
rect 19465 5195 19510 5315
rect 19630 5195 19675 5315
rect 19795 5195 19850 5315
rect 19970 5195 20015 5315
rect 20135 5195 20180 5315
rect 20300 5195 20345 5315
rect 20465 5195 20520 5315
rect 20640 5195 20685 5315
rect 20805 5195 20850 5315
rect 20970 5195 21015 5315
rect 21135 5195 21190 5315
rect 21310 5195 21355 5315
rect 21475 5195 21520 5315
rect 21640 5195 21685 5315
rect 21805 5195 21860 5315
rect 21980 5195 22025 5315
rect 22145 5195 22190 5315
rect 22310 5195 22355 5315
rect 22475 5195 22530 5315
rect 22650 5195 22695 5315
rect 22815 5195 22860 5315
rect 22980 5195 23025 5315
rect 23145 5195 23200 5315
rect 23320 5195 23365 5315
rect 23485 5195 23530 5315
rect 23650 5195 23695 5315
rect 23815 5195 23870 5315
rect 23990 5195 24000 5315
rect 18500 5150 24000 5195
rect 18500 5030 18510 5150
rect 18630 5030 18675 5150
rect 18795 5030 18840 5150
rect 18960 5030 19005 5150
rect 19125 5030 19180 5150
rect 19300 5030 19345 5150
rect 19465 5030 19510 5150
rect 19630 5030 19675 5150
rect 19795 5030 19850 5150
rect 19970 5030 20015 5150
rect 20135 5030 20180 5150
rect 20300 5030 20345 5150
rect 20465 5030 20520 5150
rect 20640 5030 20685 5150
rect 20805 5030 20850 5150
rect 20970 5030 21015 5150
rect 21135 5030 21190 5150
rect 21310 5030 21355 5150
rect 21475 5030 21520 5150
rect 21640 5030 21685 5150
rect 21805 5030 21860 5150
rect 21980 5030 22025 5150
rect 22145 5030 22190 5150
rect 22310 5030 22355 5150
rect 22475 5030 22530 5150
rect 22650 5030 22695 5150
rect 22815 5030 22860 5150
rect 22980 5030 23025 5150
rect 23145 5030 23200 5150
rect 23320 5030 23365 5150
rect 23485 5030 23530 5150
rect 23650 5030 23695 5150
rect 23815 5030 23870 5150
rect 23990 5030 24000 5150
rect 18500 4975 24000 5030
rect 18500 4855 18510 4975
rect 18630 4855 18675 4975
rect 18795 4855 18840 4975
rect 18960 4855 19005 4975
rect 19125 4855 19180 4975
rect 19300 4855 19345 4975
rect 19465 4855 19510 4975
rect 19630 4855 19675 4975
rect 19795 4855 19850 4975
rect 19970 4855 20015 4975
rect 20135 4855 20180 4975
rect 20300 4855 20345 4975
rect 20465 4855 20520 4975
rect 20640 4855 20685 4975
rect 20805 4855 20850 4975
rect 20970 4855 21015 4975
rect 21135 4855 21190 4975
rect 21310 4855 21355 4975
rect 21475 4855 21520 4975
rect 21640 4855 21685 4975
rect 21805 4855 21860 4975
rect 21980 4855 22025 4975
rect 22145 4855 22190 4975
rect 22310 4855 22355 4975
rect 22475 4855 22530 4975
rect 22650 4855 22695 4975
rect 22815 4855 22860 4975
rect 22980 4855 23025 4975
rect 23145 4855 23200 4975
rect 23320 4855 23365 4975
rect 23485 4855 23530 4975
rect 23650 4855 23695 4975
rect 23815 4855 23870 4975
rect 23990 4855 24000 4975
rect 18500 4810 24000 4855
rect 18500 4690 18510 4810
rect 18630 4690 18675 4810
rect 18795 4690 18840 4810
rect 18960 4690 19005 4810
rect 19125 4690 19180 4810
rect 19300 4690 19345 4810
rect 19465 4690 19510 4810
rect 19630 4690 19675 4810
rect 19795 4690 19850 4810
rect 19970 4690 20015 4810
rect 20135 4690 20180 4810
rect 20300 4690 20345 4810
rect 20465 4690 20520 4810
rect 20640 4690 20685 4810
rect 20805 4690 20850 4810
rect 20970 4690 21015 4810
rect 21135 4690 21190 4810
rect 21310 4690 21355 4810
rect 21475 4690 21520 4810
rect 21640 4690 21685 4810
rect 21805 4690 21860 4810
rect 21980 4690 22025 4810
rect 22145 4690 22190 4810
rect 22310 4690 22355 4810
rect 22475 4690 22530 4810
rect 22650 4690 22695 4810
rect 22815 4690 22860 4810
rect 22980 4690 23025 4810
rect 23145 4690 23200 4810
rect 23320 4690 23365 4810
rect 23485 4690 23530 4810
rect 23650 4690 23695 4810
rect 23815 4690 23870 4810
rect 23990 4690 24000 4810
rect 18500 4645 24000 4690
rect 18500 4525 18510 4645
rect 18630 4525 18675 4645
rect 18795 4525 18840 4645
rect 18960 4525 19005 4645
rect 19125 4525 19180 4645
rect 19300 4525 19345 4645
rect 19465 4525 19510 4645
rect 19630 4525 19675 4645
rect 19795 4525 19850 4645
rect 19970 4525 20015 4645
rect 20135 4525 20180 4645
rect 20300 4525 20345 4645
rect 20465 4525 20520 4645
rect 20640 4525 20685 4645
rect 20805 4525 20850 4645
rect 20970 4525 21015 4645
rect 21135 4525 21190 4645
rect 21310 4525 21355 4645
rect 21475 4525 21520 4645
rect 21640 4525 21685 4645
rect 21805 4525 21860 4645
rect 21980 4525 22025 4645
rect 22145 4525 22190 4645
rect 22310 4525 22355 4645
rect 22475 4525 22530 4645
rect 22650 4525 22695 4645
rect 22815 4525 22860 4645
rect 22980 4525 23025 4645
rect 23145 4525 23200 4645
rect 23320 4525 23365 4645
rect 23485 4525 23530 4645
rect 23650 4525 23695 4645
rect 23815 4525 23870 4645
rect 23990 4525 24000 4645
rect 18500 4480 24000 4525
rect 18500 4360 18510 4480
rect 18630 4360 18675 4480
rect 18795 4360 18840 4480
rect 18960 4360 19005 4480
rect 19125 4360 19180 4480
rect 19300 4360 19345 4480
rect 19465 4360 19510 4480
rect 19630 4360 19675 4480
rect 19795 4360 19850 4480
rect 19970 4360 20015 4480
rect 20135 4360 20180 4480
rect 20300 4360 20345 4480
rect 20465 4360 20520 4480
rect 20640 4360 20685 4480
rect 20805 4360 20850 4480
rect 20970 4360 21015 4480
rect 21135 4360 21190 4480
rect 21310 4360 21355 4480
rect 21475 4360 21520 4480
rect 21640 4360 21685 4480
rect 21805 4360 21860 4480
rect 21980 4360 22025 4480
rect 22145 4360 22190 4480
rect 22310 4360 22355 4480
rect 22475 4360 22530 4480
rect 22650 4360 22695 4480
rect 22815 4360 22860 4480
rect 22980 4360 23025 4480
rect 23145 4360 23200 4480
rect 23320 4360 23365 4480
rect 23485 4360 23530 4480
rect 23650 4360 23695 4480
rect 23815 4360 23870 4480
rect 23990 4360 24000 4480
rect 18500 4305 24000 4360
rect 18500 4185 18510 4305
rect 18630 4185 18675 4305
rect 18795 4185 18840 4305
rect 18960 4185 19005 4305
rect 19125 4185 19180 4305
rect 19300 4185 19345 4305
rect 19465 4185 19510 4305
rect 19630 4185 19675 4305
rect 19795 4185 19850 4305
rect 19970 4185 20015 4305
rect 20135 4185 20180 4305
rect 20300 4185 20345 4305
rect 20465 4185 20520 4305
rect 20640 4185 20685 4305
rect 20805 4185 20850 4305
rect 20970 4185 21015 4305
rect 21135 4185 21190 4305
rect 21310 4185 21355 4305
rect 21475 4185 21520 4305
rect 21640 4185 21685 4305
rect 21805 4185 21860 4305
rect 21980 4185 22025 4305
rect 22145 4185 22190 4305
rect 22310 4185 22355 4305
rect 22475 4185 22530 4305
rect 22650 4185 22695 4305
rect 22815 4185 22860 4305
rect 22980 4185 23025 4305
rect 23145 4185 23200 4305
rect 23320 4185 23365 4305
rect 23485 4185 23530 4305
rect 23650 4185 23695 4305
rect 23815 4185 23870 4305
rect 23990 4185 24000 4305
rect 18500 4140 24000 4185
rect 18500 4020 18510 4140
rect 18630 4020 18675 4140
rect 18795 4020 18840 4140
rect 18960 4020 19005 4140
rect 19125 4020 19180 4140
rect 19300 4020 19345 4140
rect 19465 4020 19510 4140
rect 19630 4020 19675 4140
rect 19795 4020 19850 4140
rect 19970 4020 20015 4140
rect 20135 4020 20180 4140
rect 20300 4020 20345 4140
rect 20465 4020 20520 4140
rect 20640 4020 20685 4140
rect 20805 4020 20850 4140
rect 20970 4020 21015 4140
rect 21135 4020 21190 4140
rect 21310 4020 21355 4140
rect 21475 4020 21520 4140
rect 21640 4020 21685 4140
rect 21805 4020 21860 4140
rect 21980 4020 22025 4140
rect 22145 4020 22190 4140
rect 22310 4020 22355 4140
rect 22475 4020 22530 4140
rect 22650 4020 22695 4140
rect 22815 4020 22860 4140
rect 22980 4020 23025 4140
rect 23145 4020 23200 4140
rect 23320 4020 23365 4140
rect 23485 4020 23530 4140
rect 23650 4020 23695 4140
rect 23815 4020 23870 4140
rect 23990 4020 24000 4140
rect 18500 3975 24000 4020
rect 18500 3855 18510 3975
rect 18630 3855 18675 3975
rect 18795 3855 18840 3975
rect 18960 3855 19005 3975
rect 19125 3855 19180 3975
rect 19300 3855 19345 3975
rect 19465 3855 19510 3975
rect 19630 3855 19675 3975
rect 19795 3855 19850 3975
rect 19970 3855 20015 3975
rect 20135 3855 20180 3975
rect 20300 3855 20345 3975
rect 20465 3855 20520 3975
rect 20640 3855 20685 3975
rect 20805 3855 20850 3975
rect 20970 3855 21015 3975
rect 21135 3855 21190 3975
rect 21310 3855 21355 3975
rect 21475 3855 21520 3975
rect 21640 3855 21685 3975
rect 21805 3855 21860 3975
rect 21980 3855 22025 3975
rect 22145 3855 22190 3975
rect 22310 3855 22355 3975
rect 22475 3855 22530 3975
rect 22650 3855 22695 3975
rect 22815 3855 22860 3975
rect 22980 3855 23025 3975
rect 23145 3855 23200 3975
rect 23320 3855 23365 3975
rect 23485 3855 23530 3975
rect 23650 3855 23695 3975
rect 23815 3855 23870 3975
rect 23990 3855 24000 3975
rect 18500 3810 24000 3855
rect 18500 3690 18510 3810
rect 18630 3690 18675 3810
rect 18795 3690 18840 3810
rect 18960 3690 19005 3810
rect 19125 3690 19180 3810
rect 19300 3690 19345 3810
rect 19465 3690 19510 3810
rect 19630 3690 19675 3810
rect 19795 3690 19850 3810
rect 19970 3690 20015 3810
rect 20135 3690 20180 3810
rect 20300 3690 20345 3810
rect 20465 3690 20520 3810
rect 20640 3690 20685 3810
rect 20805 3690 20850 3810
rect 20970 3690 21015 3810
rect 21135 3690 21190 3810
rect 21310 3690 21355 3810
rect 21475 3690 21520 3810
rect 21640 3690 21685 3810
rect 21805 3690 21860 3810
rect 21980 3690 22025 3810
rect 22145 3690 22190 3810
rect 22310 3690 22355 3810
rect 22475 3690 22530 3810
rect 22650 3690 22695 3810
rect 22815 3690 22860 3810
rect 22980 3690 23025 3810
rect 23145 3690 23200 3810
rect 23320 3690 23365 3810
rect 23485 3690 23530 3810
rect 23650 3690 23695 3810
rect 23815 3690 23870 3810
rect 23990 3690 24000 3810
rect 18500 3635 24000 3690
rect 18500 3515 18510 3635
rect 18630 3515 18675 3635
rect 18795 3515 18840 3635
rect 18960 3515 19005 3635
rect 19125 3515 19180 3635
rect 19300 3515 19345 3635
rect 19465 3515 19510 3635
rect 19630 3515 19675 3635
rect 19795 3515 19850 3635
rect 19970 3515 20015 3635
rect 20135 3515 20180 3635
rect 20300 3515 20345 3635
rect 20465 3515 20520 3635
rect 20640 3515 20685 3635
rect 20805 3515 20850 3635
rect 20970 3515 21015 3635
rect 21135 3515 21190 3635
rect 21310 3515 21355 3635
rect 21475 3515 21520 3635
rect 21640 3515 21685 3635
rect 21805 3515 21860 3635
rect 21980 3515 22025 3635
rect 22145 3515 22190 3635
rect 22310 3515 22355 3635
rect 22475 3515 22530 3635
rect 22650 3515 22695 3635
rect 22815 3515 22860 3635
rect 22980 3515 23025 3635
rect 23145 3515 23200 3635
rect 23320 3515 23365 3635
rect 23485 3515 23530 3635
rect 23650 3515 23695 3635
rect 23815 3515 23870 3635
rect 23990 3515 24000 3635
rect 18500 3470 24000 3515
rect 18500 3350 18510 3470
rect 18630 3350 18675 3470
rect 18795 3350 18840 3470
rect 18960 3350 19005 3470
rect 19125 3350 19180 3470
rect 19300 3350 19345 3470
rect 19465 3350 19510 3470
rect 19630 3350 19675 3470
rect 19795 3350 19850 3470
rect 19970 3350 20015 3470
rect 20135 3350 20180 3470
rect 20300 3350 20345 3470
rect 20465 3350 20520 3470
rect 20640 3350 20685 3470
rect 20805 3350 20850 3470
rect 20970 3350 21015 3470
rect 21135 3350 21190 3470
rect 21310 3350 21355 3470
rect 21475 3350 21520 3470
rect 21640 3350 21685 3470
rect 21805 3350 21860 3470
rect 21980 3350 22025 3470
rect 22145 3350 22190 3470
rect 22310 3350 22355 3470
rect 22475 3350 22530 3470
rect 22650 3350 22695 3470
rect 22815 3350 22860 3470
rect 22980 3350 23025 3470
rect 23145 3350 23200 3470
rect 23320 3350 23365 3470
rect 23485 3350 23530 3470
rect 23650 3350 23695 3470
rect 23815 3350 23870 3470
rect 23990 3350 24000 3470
rect 18500 3305 24000 3350
rect 18500 3185 18510 3305
rect 18630 3185 18675 3305
rect 18795 3185 18840 3305
rect 18960 3185 19005 3305
rect 19125 3185 19180 3305
rect 19300 3185 19345 3305
rect 19465 3185 19510 3305
rect 19630 3185 19675 3305
rect 19795 3185 19850 3305
rect 19970 3185 20015 3305
rect 20135 3185 20180 3305
rect 20300 3185 20345 3305
rect 20465 3185 20520 3305
rect 20640 3185 20685 3305
rect 20805 3185 20850 3305
rect 20970 3185 21015 3305
rect 21135 3185 21190 3305
rect 21310 3185 21355 3305
rect 21475 3185 21520 3305
rect 21640 3185 21685 3305
rect 21805 3185 21860 3305
rect 21980 3185 22025 3305
rect 22145 3185 22190 3305
rect 22310 3185 22355 3305
rect 22475 3185 22530 3305
rect 22650 3185 22695 3305
rect 22815 3185 22860 3305
rect 22980 3185 23025 3305
rect 23145 3185 23200 3305
rect 23320 3185 23365 3305
rect 23485 3185 23530 3305
rect 23650 3185 23695 3305
rect 23815 3185 23870 3305
rect 23990 3185 24000 3305
rect 18500 3140 24000 3185
rect 18500 3020 18510 3140
rect 18630 3020 18675 3140
rect 18795 3020 18840 3140
rect 18960 3020 19005 3140
rect 19125 3020 19180 3140
rect 19300 3020 19345 3140
rect 19465 3020 19510 3140
rect 19630 3020 19675 3140
rect 19795 3020 19850 3140
rect 19970 3020 20015 3140
rect 20135 3020 20180 3140
rect 20300 3020 20345 3140
rect 20465 3020 20520 3140
rect 20640 3020 20685 3140
rect 20805 3020 20850 3140
rect 20970 3020 21015 3140
rect 21135 3020 21190 3140
rect 21310 3020 21355 3140
rect 21475 3020 21520 3140
rect 21640 3020 21685 3140
rect 21805 3020 21860 3140
rect 21980 3020 22025 3140
rect 22145 3020 22190 3140
rect 22310 3020 22355 3140
rect 22475 3020 22530 3140
rect 22650 3020 22695 3140
rect 22815 3020 22860 3140
rect 22980 3020 23025 3140
rect 23145 3020 23200 3140
rect 23320 3020 23365 3140
rect 23485 3020 23530 3140
rect 23650 3020 23695 3140
rect 23815 3020 23870 3140
rect 23990 3020 24000 3140
rect 18500 2965 24000 3020
rect 18500 2845 18510 2965
rect 18630 2845 18675 2965
rect 18795 2845 18840 2965
rect 18960 2845 19005 2965
rect 19125 2845 19180 2965
rect 19300 2845 19345 2965
rect 19465 2845 19510 2965
rect 19630 2845 19675 2965
rect 19795 2845 19850 2965
rect 19970 2845 20015 2965
rect 20135 2845 20180 2965
rect 20300 2845 20345 2965
rect 20465 2845 20520 2965
rect 20640 2845 20685 2965
rect 20805 2845 20850 2965
rect 20970 2845 21015 2965
rect 21135 2845 21190 2965
rect 21310 2845 21355 2965
rect 21475 2845 21520 2965
rect 21640 2845 21685 2965
rect 21805 2845 21860 2965
rect 21980 2845 22025 2965
rect 22145 2845 22190 2965
rect 22310 2845 22355 2965
rect 22475 2845 22530 2965
rect 22650 2845 22695 2965
rect 22815 2845 22860 2965
rect 22980 2845 23025 2965
rect 23145 2845 23200 2965
rect 23320 2845 23365 2965
rect 23485 2845 23530 2965
rect 23650 2845 23695 2965
rect 23815 2845 23870 2965
rect 23990 2845 24000 2965
rect 18500 2800 24000 2845
rect 18500 2680 18510 2800
rect 18630 2680 18675 2800
rect 18795 2680 18840 2800
rect 18960 2680 19005 2800
rect 19125 2680 19180 2800
rect 19300 2680 19345 2800
rect 19465 2680 19510 2800
rect 19630 2680 19675 2800
rect 19795 2680 19850 2800
rect 19970 2680 20015 2800
rect 20135 2680 20180 2800
rect 20300 2680 20345 2800
rect 20465 2680 20520 2800
rect 20640 2680 20685 2800
rect 20805 2680 20850 2800
rect 20970 2680 21015 2800
rect 21135 2680 21190 2800
rect 21310 2680 21355 2800
rect 21475 2680 21520 2800
rect 21640 2680 21685 2800
rect 21805 2680 21860 2800
rect 21980 2680 22025 2800
rect 22145 2680 22190 2800
rect 22310 2680 22355 2800
rect 22475 2680 22530 2800
rect 22650 2680 22695 2800
rect 22815 2680 22860 2800
rect 22980 2680 23025 2800
rect 23145 2680 23200 2800
rect 23320 2680 23365 2800
rect 23485 2680 23530 2800
rect 23650 2680 23695 2800
rect 23815 2680 23870 2800
rect 23990 2680 24000 2800
rect 18500 2635 24000 2680
rect 18500 2515 18510 2635
rect 18630 2515 18675 2635
rect 18795 2515 18840 2635
rect 18960 2515 19005 2635
rect 19125 2515 19180 2635
rect 19300 2515 19345 2635
rect 19465 2515 19510 2635
rect 19630 2515 19675 2635
rect 19795 2515 19850 2635
rect 19970 2515 20015 2635
rect 20135 2515 20180 2635
rect 20300 2515 20345 2635
rect 20465 2515 20520 2635
rect 20640 2515 20685 2635
rect 20805 2515 20850 2635
rect 20970 2515 21015 2635
rect 21135 2515 21190 2635
rect 21310 2515 21355 2635
rect 21475 2515 21520 2635
rect 21640 2515 21685 2635
rect 21805 2515 21860 2635
rect 21980 2515 22025 2635
rect 22145 2515 22190 2635
rect 22310 2515 22355 2635
rect 22475 2515 22530 2635
rect 22650 2515 22695 2635
rect 22815 2515 22860 2635
rect 22980 2515 23025 2635
rect 23145 2515 23200 2635
rect 23320 2515 23365 2635
rect 23485 2515 23530 2635
rect 23650 2515 23695 2635
rect 23815 2515 23870 2635
rect 23990 2515 24000 2635
rect 18500 2470 24000 2515
rect 18500 2350 18510 2470
rect 18630 2350 18675 2470
rect 18795 2350 18840 2470
rect 18960 2350 19005 2470
rect 19125 2350 19180 2470
rect 19300 2350 19345 2470
rect 19465 2350 19510 2470
rect 19630 2350 19675 2470
rect 19795 2350 19850 2470
rect 19970 2350 20015 2470
rect 20135 2350 20180 2470
rect 20300 2350 20345 2470
rect 20465 2350 20520 2470
rect 20640 2350 20685 2470
rect 20805 2350 20850 2470
rect 20970 2350 21015 2470
rect 21135 2350 21190 2470
rect 21310 2350 21355 2470
rect 21475 2350 21520 2470
rect 21640 2350 21685 2470
rect 21805 2350 21860 2470
rect 21980 2350 22025 2470
rect 22145 2350 22190 2470
rect 22310 2350 22355 2470
rect 22475 2350 22530 2470
rect 22650 2350 22695 2470
rect 22815 2350 22860 2470
rect 22980 2350 23025 2470
rect 23145 2350 23200 2470
rect 23320 2350 23365 2470
rect 23485 2350 23530 2470
rect 23650 2350 23695 2470
rect 23815 2350 23870 2470
rect 23990 2350 24000 2470
rect 18500 2295 24000 2350
rect 18500 2175 18510 2295
rect 18630 2175 18675 2295
rect 18795 2175 18840 2295
rect 18960 2175 19005 2295
rect 19125 2175 19180 2295
rect 19300 2175 19345 2295
rect 19465 2175 19510 2295
rect 19630 2175 19675 2295
rect 19795 2175 19850 2295
rect 19970 2175 20015 2295
rect 20135 2175 20180 2295
rect 20300 2175 20345 2295
rect 20465 2175 20520 2295
rect 20640 2175 20685 2295
rect 20805 2175 20850 2295
rect 20970 2175 21015 2295
rect 21135 2175 21190 2295
rect 21310 2175 21355 2295
rect 21475 2175 21520 2295
rect 21640 2175 21685 2295
rect 21805 2175 21860 2295
rect 21980 2175 22025 2295
rect 22145 2175 22190 2295
rect 22310 2175 22355 2295
rect 22475 2175 22530 2295
rect 22650 2175 22695 2295
rect 22815 2175 22860 2295
rect 22980 2175 23025 2295
rect 23145 2175 23200 2295
rect 23320 2175 23365 2295
rect 23485 2175 23530 2295
rect 23650 2175 23695 2295
rect 23815 2175 23870 2295
rect 23990 2175 24000 2295
rect 18500 2130 24000 2175
rect 18500 2010 18510 2130
rect 18630 2010 18675 2130
rect 18795 2010 18840 2130
rect 18960 2010 19005 2130
rect 19125 2010 19180 2130
rect 19300 2010 19345 2130
rect 19465 2010 19510 2130
rect 19630 2010 19675 2130
rect 19795 2010 19850 2130
rect 19970 2010 20015 2130
rect 20135 2010 20180 2130
rect 20300 2010 20345 2130
rect 20465 2010 20520 2130
rect 20640 2010 20685 2130
rect 20805 2010 20850 2130
rect 20970 2010 21015 2130
rect 21135 2010 21190 2130
rect 21310 2010 21355 2130
rect 21475 2010 21520 2130
rect 21640 2010 21685 2130
rect 21805 2010 21860 2130
rect 21980 2010 22025 2130
rect 22145 2010 22190 2130
rect 22310 2010 22355 2130
rect 22475 2010 22530 2130
rect 22650 2010 22695 2130
rect 22815 2010 22860 2130
rect 22980 2010 23025 2130
rect 23145 2010 23200 2130
rect 23320 2010 23365 2130
rect 23485 2010 23530 2130
rect 23650 2010 23695 2130
rect 23815 2010 23870 2130
rect 23990 2010 24000 2130
rect 18500 1965 24000 2010
rect 18500 1845 18510 1965
rect 18630 1845 18675 1965
rect 18795 1845 18840 1965
rect 18960 1845 19005 1965
rect 19125 1845 19180 1965
rect 19300 1845 19345 1965
rect 19465 1845 19510 1965
rect 19630 1845 19675 1965
rect 19795 1845 19850 1965
rect 19970 1845 20015 1965
rect 20135 1845 20180 1965
rect 20300 1845 20345 1965
rect 20465 1845 20520 1965
rect 20640 1845 20685 1965
rect 20805 1845 20850 1965
rect 20970 1845 21015 1965
rect 21135 1845 21190 1965
rect 21310 1845 21355 1965
rect 21475 1845 21520 1965
rect 21640 1845 21685 1965
rect 21805 1845 21860 1965
rect 21980 1845 22025 1965
rect 22145 1845 22190 1965
rect 22310 1845 22355 1965
rect 22475 1845 22530 1965
rect 22650 1845 22695 1965
rect 22815 1845 22860 1965
rect 22980 1845 23025 1965
rect 23145 1845 23200 1965
rect 23320 1845 23365 1965
rect 23485 1845 23530 1965
rect 23650 1845 23695 1965
rect 23815 1845 23870 1965
rect 23990 1845 24000 1965
rect 18500 1800 24000 1845
rect 18500 1680 18510 1800
rect 18630 1680 18675 1800
rect 18795 1680 18840 1800
rect 18960 1680 19005 1800
rect 19125 1680 19180 1800
rect 19300 1680 19345 1800
rect 19465 1680 19510 1800
rect 19630 1680 19675 1800
rect 19795 1680 19850 1800
rect 19970 1680 20015 1800
rect 20135 1680 20180 1800
rect 20300 1680 20345 1800
rect 20465 1680 20520 1800
rect 20640 1680 20685 1800
rect 20805 1680 20850 1800
rect 20970 1680 21015 1800
rect 21135 1680 21190 1800
rect 21310 1680 21355 1800
rect 21475 1680 21520 1800
rect 21640 1680 21685 1800
rect 21805 1680 21860 1800
rect 21980 1680 22025 1800
rect 22145 1680 22190 1800
rect 22310 1680 22355 1800
rect 22475 1680 22530 1800
rect 22650 1680 22695 1800
rect 22815 1680 22860 1800
rect 22980 1680 23025 1800
rect 23145 1680 23200 1800
rect 23320 1680 23365 1800
rect 23485 1680 23530 1800
rect 23650 1680 23695 1800
rect 23815 1680 23870 1800
rect 23990 1680 24000 1800
rect 18500 1670 24000 1680
rect 24190 7160 29690 7170
rect 24190 7040 24200 7160
rect 24320 7040 24365 7160
rect 24485 7040 24530 7160
rect 24650 7040 24695 7160
rect 24815 7040 24870 7160
rect 24990 7040 25035 7160
rect 25155 7040 25200 7160
rect 25320 7040 25365 7160
rect 25485 7040 25540 7160
rect 25660 7040 25705 7160
rect 25825 7040 25870 7160
rect 25990 7040 26035 7160
rect 26155 7040 26210 7160
rect 26330 7040 26375 7160
rect 26495 7040 26540 7160
rect 26660 7040 26705 7160
rect 26825 7040 26880 7160
rect 27000 7040 27045 7160
rect 27165 7040 27210 7160
rect 27330 7040 27375 7160
rect 27495 7040 27550 7160
rect 27670 7040 27715 7160
rect 27835 7040 27880 7160
rect 28000 7040 28045 7160
rect 28165 7040 28220 7160
rect 28340 7040 28385 7160
rect 28505 7040 28550 7160
rect 28670 7040 28715 7160
rect 28835 7040 28890 7160
rect 29010 7040 29055 7160
rect 29175 7040 29220 7160
rect 29340 7040 29385 7160
rect 29505 7040 29560 7160
rect 29680 7040 29690 7160
rect 24190 6985 29690 7040
rect 24190 6865 24200 6985
rect 24320 6865 24365 6985
rect 24485 6865 24530 6985
rect 24650 6865 24695 6985
rect 24815 6865 24870 6985
rect 24990 6865 25035 6985
rect 25155 6865 25200 6985
rect 25320 6865 25365 6985
rect 25485 6865 25540 6985
rect 25660 6865 25705 6985
rect 25825 6865 25870 6985
rect 25990 6865 26035 6985
rect 26155 6865 26210 6985
rect 26330 6865 26375 6985
rect 26495 6865 26540 6985
rect 26660 6865 26705 6985
rect 26825 6865 26880 6985
rect 27000 6865 27045 6985
rect 27165 6865 27210 6985
rect 27330 6865 27375 6985
rect 27495 6865 27550 6985
rect 27670 6865 27715 6985
rect 27835 6865 27880 6985
rect 28000 6865 28045 6985
rect 28165 6865 28220 6985
rect 28340 6865 28385 6985
rect 28505 6865 28550 6985
rect 28670 6865 28715 6985
rect 28835 6865 28890 6985
rect 29010 6865 29055 6985
rect 29175 6865 29220 6985
rect 29340 6865 29385 6985
rect 29505 6865 29560 6985
rect 29680 6865 29690 6985
rect 24190 6820 29690 6865
rect 24190 6700 24200 6820
rect 24320 6700 24365 6820
rect 24485 6700 24530 6820
rect 24650 6700 24695 6820
rect 24815 6700 24870 6820
rect 24990 6700 25035 6820
rect 25155 6700 25200 6820
rect 25320 6700 25365 6820
rect 25485 6700 25540 6820
rect 25660 6700 25705 6820
rect 25825 6700 25870 6820
rect 25990 6700 26035 6820
rect 26155 6700 26210 6820
rect 26330 6700 26375 6820
rect 26495 6700 26540 6820
rect 26660 6700 26705 6820
rect 26825 6700 26880 6820
rect 27000 6700 27045 6820
rect 27165 6700 27210 6820
rect 27330 6700 27375 6820
rect 27495 6700 27550 6820
rect 27670 6700 27715 6820
rect 27835 6700 27880 6820
rect 28000 6700 28045 6820
rect 28165 6700 28220 6820
rect 28340 6700 28385 6820
rect 28505 6700 28550 6820
rect 28670 6700 28715 6820
rect 28835 6700 28890 6820
rect 29010 6700 29055 6820
rect 29175 6700 29220 6820
rect 29340 6700 29385 6820
rect 29505 6700 29560 6820
rect 29680 6700 29690 6820
rect 24190 6655 29690 6700
rect 24190 6535 24200 6655
rect 24320 6535 24365 6655
rect 24485 6535 24530 6655
rect 24650 6535 24695 6655
rect 24815 6535 24870 6655
rect 24990 6535 25035 6655
rect 25155 6535 25200 6655
rect 25320 6535 25365 6655
rect 25485 6535 25540 6655
rect 25660 6535 25705 6655
rect 25825 6535 25870 6655
rect 25990 6535 26035 6655
rect 26155 6535 26210 6655
rect 26330 6535 26375 6655
rect 26495 6535 26540 6655
rect 26660 6535 26705 6655
rect 26825 6535 26880 6655
rect 27000 6535 27045 6655
rect 27165 6535 27210 6655
rect 27330 6535 27375 6655
rect 27495 6535 27550 6655
rect 27670 6535 27715 6655
rect 27835 6535 27880 6655
rect 28000 6535 28045 6655
rect 28165 6535 28220 6655
rect 28340 6535 28385 6655
rect 28505 6535 28550 6655
rect 28670 6535 28715 6655
rect 28835 6535 28890 6655
rect 29010 6535 29055 6655
rect 29175 6535 29220 6655
rect 29340 6535 29385 6655
rect 29505 6535 29560 6655
rect 29680 6535 29690 6655
rect 24190 6490 29690 6535
rect 24190 6370 24200 6490
rect 24320 6370 24365 6490
rect 24485 6370 24530 6490
rect 24650 6370 24695 6490
rect 24815 6370 24870 6490
rect 24990 6370 25035 6490
rect 25155 6370 25200 6490
rect 25320 6370 25365 6490
rect 25485 6370 25540 6490
rect 25660 6370 25705 6490
rect 25825 6370 25870 6490
rect 25990 6370 26035 6490
rect 26155 6370 26210 6490
rect 26330 6370 26375 6490
rect 26495 6370 26540 6490
rect 26660 6370 26705 6490
rect 26825 6370 26880 6490
rect 27000 6370 27045 6490
rect 27165 6370 27210 6490
rect 27330 6370 27375 6490
rect 27495 6370 27550 6490
rect 27670 6370 27715 6490
rect 27835 6370 27880 6490
rect 28000 6370 28045 6490
rect 28165 6370 28220 6490
rect 28340 6370 28385 6490
rect 28505 6370 28550 6490
rect 28670 6370 28715 6490
rect 28835 6370 28890 6490
rect 29010 6370 29055 6490
rect 29175 6370 29220 6490
rect 29340 6370 29385 6490
rect 29505 6370 29560 6490
rect 29680 6370 29690 6490
rect 24190 6315 29690 6370
rect 24190 6195 24200 6315
rect 24320 6195 24365 6315
rect 24485 6195 24530 6315
rect 24650 6195 24695 6315
rect 24815 6195 24870 6315
rect 24990 6195 25035 6315
rect 25155 6195 25200 6315
rect 25320 6195 25365 6315
rect 25485 6195 25540 6315
rect 25660 6195 25705 6315
rect 25825 6195 25870 6315
rect 25990 6195 26035 6315
rect 26155 6195 26210 6315
rect 26330 6195 26375 6315
rect 26495 6195 26540 6315
rect 26660 6195 26705 6315
rect 26825 6195 26880 6315
rect 27000 6195 27045 6315
rect 27165 6195 27210 6315
rect 27330 6195 27375 6315
rect 27495 6195 27550 6315
rect 27670 6195 27715 6315
rect 27835 6195 27880 6315
rect 28000 6195 28045 6315
rect 28165 6195 28220 6315
rect 28340 6195 28385 6315
rect 28505 6195 28550 6315
rect 28670 6195 28715 6315
rect 28835 6195 28890 6315
rect 29010 6195 29055 6315
rect 29175 6195 29220 6315
rect 29340 6195 29385 6315
rect 29505 6195 29560 6315
rect 29680 6195 29690 6315
rect 24190 6150 29690 6195
rect 24190 6030 24200 6150
rect 24320 6030 24365 6150
rect 24485 6030 24530 6150
rect 24650 6030 24695 6150
rect 24815 6030 24870 6150
rect 24990 6030 25035 6150
rect 25155 6030 25200 6150
rect 25320 6030 25365 6150
rect 25485 6030 25540 6150
rect 25660 6030 25705 6150
rect 25825 6030 25870 6150
rect 25990 6030 26035 6150
rect 26155 6030 26210 6150
rect 26330 6030 26375 6150
rect 26495 6030 26540 6150
rect 26660 6030 26705 6150
rect 26825 6030 26880 6150
rect 27000 6030 27045 6150
rect 27165 6030 27210 6150
rect 27330 6030 27375 6150
rect 27495 6030 27550 6150
rect 27670 6030 27715 6150
rect 27835 6030 27880 6150
rect 28000 6030 28045 6150
rect 28165 6030 28220 6150
rect 28340 6030 28385 6150
rect 28505 6030 28550 6150
rect 28670 6030 28715 6150
rect 28835 6030 28890 6150
rect 29010 6030 29055 6150
rect 29175 6030 29220 6150
rect 29340 6030 29385 6150
rect 29505 6030 29560 6150
rect 29680 6030 29690 6150
rect 24190 5985 29690 6030
rect 24190 5865 24200 5985
rect 24320 5865 24365 5985
rect 24485 5865 24530 5985
rect 24650 5865 24695 5985
rect 24815 5865 24870 5985
rect 24990 5865 25035 5985
rect 25155 5865 25200 5985
rect 25320 5865 25365 5985
rect 25485 5865 25540 5985
rect 25660 5865 25705 5985
rect 25825 5865 25870 5985
rect 25990 5865 26035 5985
rect 26155 5865 26210 5985
rect 26330 5865 26375 5985
rect 26495 5865 26540 5985
rect 26660 5865 26705 5985
rect 26825 5865 26880 5985
rect 27000 5865 27045 5985
rect 27165 5865 27210 5985
rect 27330 5865 27375 5985
rect 27495 5865 27550 5985
rect 27670 5865 27715 5985
rect 27835 5865 27880 5985
rect 28000 5865 28045 5985
rect 28165 5865 28220 5985
rect 28340 5865 28385 5985
rect 28505 5865 28550 5985
rect 28670 5865 28715 5985
rect 28835 5865 28890 5985
rect 29010 5865 29055 5985
rect 29175 5865 29220 5985
rect 29340 5865 29385 5985
rect 29505 5865 29560 5985
rect 29680 5865 29690 5985
rect 24190 5820 29690 5865
rect 24190 5700 24200 5820
rect 24320 5700 24365 5820
rect 24485 5700 24530 5820
rect 24650 5700 24695 5820
rect 24815 5700 24870 5820
rect 24990 5700 25035 5820
rect 25155 5700 25200 5820
rect 25320 5700 25365 5820
rect 25485 5700 25540 5820
rect 25660 5700 25705 5820
rect 25825 5700 25870 5820
rect 25990 5700 26035 5820
rect 26155 5700 26210 5820
rect 26330 5700 26375 5820
rect 26495 5700 26540 5820
rect 26660 5700 26705 5820
rect 26825 5700 26880 5820
rect 27000 5700 27045 5820
rect 27165 5700 27210 5820
rect 27330 5700 27375 5820
rect 27495 5700 27550 5820
rect 27670 5700 27715 5820
rect 27835 5700 27880 5820
rect 28000 5700 28045 5820
rect 28165 5700 28220 5820
rect 28340 5700 28385 5820
rect 28505 5700 28550 5820
rect 28670 5700 28715 5820
rect 28835 5700 28890 5820
rect 29010 5700 29055 5820
rect 29175 5700 29220 5820
rect 29340 5700 29385 5820
rect 29505 5700 29560 5820
rect 29680 5700 29690 5820
rect 24190 5645 29690 5700
rect 24190 5525 24200 5645
rect 24320 5525 24365 5645
rect 24485 5525 24530 5645
rect 24650 5525 24695 5645
rect 24815 5525 24870 5645
rect 24990 5525 25035 5645
rect 25155 5525 25200 5645
rect 25320 5525 25365 5645
rect 25485 5525 25540 5645
rect 25660 5525 25705 5645
rect 25825 5525 25870 5645
rect 25990 5525 26035 5645
rect 26155 5525 26210 5645
rect 26330 5525 26375 5645
rect 26495 5525 26540 5645
rect 26660 5525 26705 5645
rect 26825 5525 26880 5645
rect 27000 5525 27045 5645
rect 27165 5525 27210 5645
rect 27330 5525 27375 5645
rect 27495 5525 27550 5645
rect 27670 5525 27715 5645
rect 27835 5525 27880 5645
rect 28000 5525 28045 5645
rect 28165 5525 28220 5645
rect 28340 5525 28385 5645
rect 28505 5525 28550 5645
rect 28670 5525 28715 5645
rect 28835 5525 28890 5645
rect 29010 5525 29055 5645
rect 29175 5525 29220 5645
rect 29340 5525 29385 5645
rect 29505 5525 29560 5645
rect 29680 5525 29690 5645
rect 24190 5480 29690 5525
rect 24190 5360 24200 5480
rect 24320 5360 24365 5480
rect 24485 5360 24530 5480
rect 24650 5360 24695 5480
rect 24815 5360 24870 5480
rect 24990 5360 25035 5480
rect 25155 5360 25200 5480
rect 25320 5360 25365 5480
rect 25485 5360 25540 5480
rect 25660 5360 25705 5480
rect 25825 5360 25870 5480
rect 25990 5360 26035 5480
rect 26155 5360 26210 5480
rect 26330 5360 26375 5480
rect 26495 5360 26540 5480
rect 26660 5360 26705 5480
rect 26825 5360 26880 5480
rect 27000 5360 27045 5480
rect 27165 5360 27210 5480
rect 27330 5360 27375 5480
rect 27495 5360 27550 5480
rect 27670 5360 27715 5480
rect 27835 5360 27880 5480
rect 28000 5360 28045 5480
rect 28165 5360 28220 5480
rect 28340 5360 28385 5480
rect 28505 5360 28550 5480
rect 28670 5360 28715 5480
rect 28835 5360 28890 5480
rect 29010 5360 29055 5480
rect 29175 5360 29220 5480
rect 29340 5360 29385 5480
rect 29505 5360 29560 5480
rect 29680 5360 29690 5480
rect 24190 5315 29690 5360
rect 24190 5195 24200 5315
rect 24320 5195 24365 5315
rect 24485 5195 24530 5315
rect 24650 5195 24695 5315
rect 24815 5195 24870 5315
rect 24990 5195 25035 5315
rect 25155 5195 25200 5315
rect 25320 5195 25365 5315
rect 25485 5195 25540 5315
rect 25660 5195 25705 5315
rect 25825 5195 25870 5315
rect 25990 5195 26035 5315
rect 26155 5195 26210 5315
rect 26330 5195 26375 5315
rect 26495 5195 26540 5315
rect 26660 5195 26705 5315
rect 26825 5195 26880 5315
rect 27000 5195 27045 5315
rect 27165 5195 27210 5315
rect 27330 5195 27375 5315
rect 27495 5195 27550 5315
rect 27670 5195 27715 5315
rect 27835 5195 27880 5315
rect 28000 5195 28045 5315
rect 28165 5195 28220 5315
rect 28340 5195 28385 5315
rect 28505 5195 28550 5315
rect 28670 5195 28715 5315
rect 28835 5195 28890 5315
rect 29010 5195 29055 5315
rect 29175 5195 29220 5315
rect 29340 5195 29385 5315
rect 29505 5195 29560 5315
rect 29680 5195 29690 5315
rect 24190 5150 29690 5195
rect 24190 5030 24200 5150
rect 24320 5030 24365 5150
rect 24485 5030 24530 5150
rect 24650 5030 24695 5150
rect 24815 5030 24870 5150
rect 24990 5030 25035 5150
rect 25155 5030 25200 5150
rect 25320 5030 25365 5150
rect 25485 5030 25540 5150
rect 25660 5030 25705 5150
rect 25825 5030 25870 5150
rect 25990 5030 26035 5150
rect 26155 5030 26210 5150
rect 26330 5030 26375 5150
rect 26495 5030 26540 5150
rect 26660 5030 26705 5150
rect 26825 5030 26880 5150
rect 27000 5030 27045 5150
rect 27165 5030 27210 5150
rect 27330 5030 27375 5150
rect 27495 5030 27550 5150
rect 27670 5030 27715 5150
rect 27835 5030 27880 5150
rect 28000 5030 28045 5150
rect 28165 5030 28220 5150
rect 28340 5030 28385 5150
rect 28505 5030 28550 5150
rect 28670 5030 28715 5150
rect 28835 5030 28890 5150
rect 29010 5030 29055 5150
rect 29175 5030 29220 5150
rect 29340 5030 29385 5150
rect 29505 5030 29560 5150
rect 29680 5030 29690 5150
rect 24190 4975 29690 5030
rect 24190 4855 24200 4975
rect 24320 4855 24365 4975
rect 24485 4855 24530 4975
rect 24650 4855 24695 4975
rect 24815 4855 24870 4975
rect 24990 4855 25035 4975
rect 25155 4855 25200 4975
rect 25320 4855 25365 4975
rect 25485 4855 25540 4975
rect 25660 4855 25705 4975
rect 25825 4855 25870 4975
rect 25990 4855 26035 4975
rect 26155 4855 26210 4975
rect 26330 4855 26375 4975
rect 26495 4855 26540 4975
rect 26660 4855 26705 4975
rect 26825 4855 26880 4975
rect 27000 4855 27045 4975
rect 27165 4855 27210 4975
rect 27330 4855 27375 4975
rect 27495 4855 27550 4975
rect 27670 4855 27715 4975
rect 27835 4855 27880 4975
rect 28000 4855 28045 4975
rect 28165 4855 28220 4975
rect 28340 4855 28385 4975
rect 28505 4855 28550 4975
rect 28670 4855 28715 4975
rect 28835 4855 28890 4975
rect 29010 4855 29055 4975
rect 29175 4855 29220 4975
rect 29340 4855 29385 4975
rect 29505 4855 29560 4975
rect 29680 4855 29690 4975
rect 24190 4810 29690 4855
rect 24190 4690 24200 4810
rect 24320 4690 24365 4810
rect 24485 4690 24530 4810
rect 24650 4690 24695 4810
rect 24815 4690 24870 4810
rect 24990 4690 25035 4810
rect 25155 4690 25200 4810
rect 25320 4690 25365 4810
rect 25485 4690 25540 4810
rect 25660 4690 25705 4810
rect 25825 4690 25870 4810
rect 25990 4690 26035 4810
rect 26155 4690 26210 4810
rect 26330 4690 26375 4810
rect 26495 4690 26540 4810
rect 26660 4690 26705 4810
rect 26825 4690 26880 4810
rect 27000 4690 27045 4810
rect 27165 4690 27210 4810
rect 27330 4690 27375 4810
rect 27495 4690 27550 4810
rect 27670 4690 27715 4810
rect 27835 4690 27880 4810
rect 28000 4690 28045 4810
rect 28165 4690 28220 4810
rect 28340 4690 28385 4810
rect 28505 4690 28550 4810
rect 28670 4690 28715 4810
rect 28835 4690 28890 4810
rect 29010 4690 29055 4810
rect 29175 4690 29220 4810
rect 29340 4690 29385 4810
rect 29505 4690 29560 4810
rect 29680 4690 29690 4810
rect 24190 4645 29690 4690
rect 24190 4525 24200 4645
rect 24320 4525 24365 4645
rect 24485 4525 24530 4645
rect 24650 4525 24695 4645
rect 24815 4525 24870 4645
rect 24990 4525 25035 4645
rect 25155 4525 25200 4645
rect 25320 4525 25365 4645
rect 25485 4525 25540 4645
rect 25660 4525 25705 4645
rect 25825 4525 25870 4645
rect 25990 4525 26035 4645
rect 26155 4525 26210 4645
rect 26330 4525 26375 4645
rect 26495 4525 26540 4645
rect 26660 4525 26705 4645
rect 26825 4525 26880 4645
rect 27000 4525 27045 4645
rect 27165 4525 27210 4645
rect 27330 4525 27375 4645
rect 27495 4525 27550 4645
rect 27670 4525 27715 4645
rect 27835 4525 27880 4645
rect 28000 4525 28045 4645
rect 28165 4525 28220 4645
rect 28340 4525 28385 4645
rect 28505 4525 28550 4645
rect 28670 4525 28715 4645
rect 28835 4525 28890 4645
rect 29010 4525 29055 4645
rect 29175 4525 29220 4645
rect 29340 4525 29385 4645
rect 29505 4525 29560 4645
rect 29680 4525 29690 4645
rect 24190 4480 29690 4525
rect 24190 4360 24200 4480
rect 24320 4360 24365 4480
rect 24485 4360 24530 4480
rect 24650 4360 24695 4480
rect 24815 4360 24870 4480
rect 24990 4360 25035 4480
rect 25155 4360 25200 4480
rect 25320 4360 25365 4480
rect 25485 4360 25540 4480
rect 25660 4360 25705 4480
rect 25825 4360 25870 4480
rect 25990 4360 26035 4480
rect 26155 4360 26210 4480
rect 26330 4360 26375 4480
rect 26495 4360 26540 4480
rect 26660 4360 26705 4480
rect 26825 4360 26880 4480
rect 27000 4360 27045 4480
rect 27165 4360 27210 4480
rect 27330 4360 27375 4480
rect 27495 4360 27550 4480
rect 27670 4360 27715 4480
rect 27835 4360 27880 4480
rect 28000 4360 28045 4480
rect 28165 4360 28220 4480
rect 28340 4360 28385 4480
rect 28505 4360 28550 4480
rect 28670 4360 28715 4480
rect 28835 4360 28890 4480
rect 29010 4360 29055 4480
rect 29175 4360 29220 4480
rect 29340 4360 29385 4480
rect 29505 4360 29560 4480
rect 29680 4360 29690 4480
rect 24190 4305 29690 4360
rect 24190 4185 24200 4305
rect 24320 4185 24365 4305
rect 24485 4185 24530 4305
rect 24650 4185 24695 4305
rect 24815 4185 24870 4305
rect 24990 4185 25035 4305
rect 25155 4185 25200 4305
rect 25320 4185 25365 4305
rect 25485 4185 25540 4305
rect 25660 4185 25705 4305
rect 25825 4185 25870 4305
rect 25990 4185 26035 4305
rect 26155 4185 26210 4305
rect 26330 4185 26375 4305
rect 26495 4185 26540 4305
rect 26660 4185 26705 4305
rect 26825 4185 26880 4305
rect 27000 4185 27045 4305
rect 27165 4185 27210 4305
rect 27330 4185 27375 4305
rect 27495 4185 27550 4305
rect 27670 4185 27715 4305
rect 27835 4185 27880 4305
rect 28000 4185 28045 4305
rect 28165 4185 28220 4305
rect 28340 4185 28385 4305
rect 28505 4185 28550 4305
rect 28670 4185 28715 4305
rect 28835 4185 28890 4305
rect 29010 4185 29055 4305
rect 29175 4185 29220 4305
rect 29340 4185 29385 4305
rect 29505 4185 29560 4305
rect 29680 4185 29690 4305
rect 24190 4140 29690 4185
rect 24190 4020 24200 4140
rect 24320 4020 24365 4140
rect 24485 4020 24530 4140
rect 24650 4020 24695 4140
rect 24815 4020 24870 4140
rect 24990 4020 25035 4140
rect 25155 4020 25200 4140
rect 25320 4020 25365 4140
rect 25485 4020 25540 4140
rect 25660 4020 25705 4140
rect 25825 4020 25870 4140
rect 25990 4020 26035 4140
rect 26155 4020 26210 4140
rect 26330 4020 26375 4140
rect 26495 4020 26540 4140
rect 26660 4020 26705 4140
rect 26825 4020 26880 4140
rect 27000 4020 27045 4140
rect 27165 4020 27210 4140
rect 27330 4020 27375 4140
rect 27495 4020 27550 4140
rect 27670 4020 27715 4140
rect 27835 4020 27880 4140
rect 28000 4020 28045 4140
rect 28165 4020 28220 4140
rect 28340 4020 28385 4140
rect 28505 4020 28550 4140
rect 28670 4020 28715 4140
rect 28835 4020 28890 4140
rect 29010 4020 29055 4140
rect 29175 4020 29220 4140
rect 29340 4020 29385 4140
rect 29505 4020 29560 4140
rect 29680 4020 29690 4140
rect 24190 3975 29690 4020
rect 24190 3855 24200 3975
rect 24320 3855 24365 3975
rect 24485 3855 24530 3975
rect 24650 3855 24695 3975
rect 24815 3855 24870 3975
rect 24990 3855 25035 3975
rect 25155 3855 25200 3975
rect 25320 3855 25365 3975
rect 25485 3855 25540 3975
rect 25660 3855 25705 3975
rect 25825 3855 25870 3975
rect 25990 3855 26035 3975
rect 26155 3855 26210 3975
rect 26330 3855 26375 3975
rect 26495 3855 26540 3975
rect 26660 3855 26705 3975
rect 26825 3855 26880 3975
rect 27000 3855 27045 3975
rect 27165 3855 27210 3975
rect 27330 3855 27375 3975
rect 27495 3855 27550 3975
rect 27670 3855 27715 3975
rect 27835 3855 27880 3975
rect 28000 3855 28045 3975
rect 28165 3855 28220 3975
rect 28340 3855 28385 3975
rect 28505 3855 28550 3975
rect 28670 3855 28715 3975
rect 28835 3855 28890 3975
rect 29010 3855 29055 3975
rect 29175 3855 29220 3975
rect 29340 3855 29385 3975
rect 29505 3855 29560 3975
rect 29680 3855 29690 3975
rect 24190 3810 29690 3855
rect 24190 3690 24200 3810
rect 24320 3690 24365 3810
rect 24485 3690 24530 3810
rect 24650 3690 24695 3810
rect 24815 3690 24870 3810
rect 24990 3690 25035 3810
rect 25155 3690 25200 3810
rect 25320 3690 25365 3810
rect 25485 3690 25540 3810
rect 25660 3690 25705 3810
rect 25825 3690 25870 3810
rect 25990 3690 26035 3810
rect 26155 3690 26210 3810
rect 26330 3690 26375 3810
rect 26495 3690 26540 3810
rect 26660 3690 26705 3810
rect 26825 3690 26880 3810
rect 27000 3690 27045 3810
rect 27165 3690 27210 3810
rect 27330 3690 27375 3810
rect 27495 3690 27550 3810
rect 27670 3690 27715 3810
rect 27835 3690 27880 3810
rect 28000 3690 28045 3810
rect 28165 3690 28220 3810
rect 28340 3690 28385 3810
rect 28505 3690 28550 3810
rect 28670 3690 28715 3810
rect 28835 3690 28890 3810
rect 29010 3690 29055 3810
rect 29175 3690 29220 3810
rect 29340 3690 29385 3810
rect 29505 3690 29560 3810
rect 29680 3690 29690 3810
rect 24190 3635 29690 3690
rect 24190 3515 24200 3635
rect 24320 3515 24365 3635
rect 24485 3515 24530 3635
rect 24650 3515 24695 3635
rect 24815 3515 24870 3635
rect 24990 3515 25035 3635
rect 25155 3515 25200 3635
rect 25320 3515 25365 3635
rect 25485 3515 25540 3635
rect 25660 3515 25705 3635
rect 25825 3515 25870 3635
rect 25990 3515 26035 3635
rect 26155 3515 26210 3635
rect 26330 3515 26375 3635
rect 26495 3515 26540 3635
rect 26660 3515 26705 3635
rect 26825 3515 26880 3635
rect 27000 3515 27045 3635
rect 27165 3515 27210 3635
rect 27330 3515 27375 3635
rect 27495 3515 27550 3635
rect 27670 3515 27715 3635
rect 27835 3515 27880 3635
rect 28000 3515 28045 3635
rect 28165 3515 28220 3635
rect 28340 3515 28385 3635
rect 28505 3515 28550 3635
rect 28670 3515 28715 3635
rect 28835 3515 28890 3635
rect 29010 3515 29055 3635
rect 29175 3515 29220 3635
rect 29340 3515 29385 3635
rect 29505 3515 29560 3635
rect 29680 3515 29690 3635
rect 24190 3470 29690 3515
rect 24190 3350 24200 3470
rect 24320 3350 24365 3470
rect 24485 3350 24530 3470
rect 24650 3350 24695 3470
rect 24815 3350 24870 3470
rect 24990 3350 25035 3470
rect 25155 3350 25200 3470
rect 25320 3350 25365 3470
rect 25485 3350 25540 3470
rect 25660 3350 25705 3470
rect 25825 3350 25870 3470
rect 25990 3350 26035 3470
rect 26155 3350 26210 3470
rect 26330 3350 26375 3470
rect 26495 3350 26540 3470
rect 26660 3350 26705 3470
rect 26825 3350 26880 3470
rect 27000 3350 27045 3470
rect 27165 3350 27210 3470
rect 27330 3350 27375 3470
rect 27495 3350 27550 3470
rect 27670 3350 27715 3470
rect 27835 3350 27880 3470
rect 28000 3350 28045 3470
rect 28165 3350 28220 3470
rect 28340 3350 28385 3470
rect 28505 3350 28550 3470
rect 28670 3350 28715 3470
rect 28835 3350 28890 3470
rect 29010 3350 29055 3470
rect 29175 3350 29220 3470
rect 29340 3350 29385 3470
rect 29505 3350 29560 3470
rect 29680 3350 29690 3470
rect 24190 3305 29690 3350
rect 24190 3185 24200 3305
rect 24320 3185 24365 3305
rect 24485 3185 24530 3305
rect 24650 3185 24695 3305
rect 24815 3185 24870 3305
rect 24990 3185 25035 3305
rect 25155 3185 25200 3305
rect 25320 3185 25365 3305
rect 25485 3185 25540 3305
rect 25660 3185 25705 3305
rect 25825 3185 25870 3305
rect 25990 3185 26035 3305
rect 26155 3185 26210 3305
rect 26330 3185 26375 3305
rect 26495 3185 26540 3305
rect 26660 3185 26705 3305
rect 26825 3185 26880 3305
rect 27000 3185 27045 3305
rect 27165 3185 27210 3305
rect 27330 3185 27375 3305
rect 27495 3185 27550 3305
rect 27670 3185 27715 3305
rect 27835 3185 27880 3305
rect 28000 3185 28045 3305
rect 28165 3185 28220 3305
rect 28340 3185 28385 3305
rect 28505 3185 28550 3305
rect 28670 3185 28715 3305
rect 28835 3185 28890 3305
rect 29010 3185 29055 3305
rect 29175 3185 29220 3305
rect 29340 3185 29385 3305
rect 29505 3185 29560 3305
rect 29680 3185 29690 3305
rect 24190 3140 29690 3185
rect 24190 3020 24200 3140
rect 24320 3020 24365 3140
rect 24485 3020 24530 3140
rect 24650 3020 24695 3140
rect 24815 3020 24870 3140
rect 24990 3020 25035 3140
rect 25155 3020 25200 3140
rect 25320 3020 25365 3140
rect 25485 3020 25540 3140
rect 25660 3020 25705 3140
rect 25825 3020 25870 3140
rect 25990 3020 26035 3140
rect 26155 3020 26210 3140
rect 26330 3020 26375 3140
rect 26495 3020 26540 3140
rect 26660 3020 26705 3140
rect 26825 3020 26880 3140
rect 27000 3020 27045 3140
rect 27165 3020 27210 3140
rect 27330 3020 27375 3140
rect 27495 3020 27550 3140
rect 27670 3020 27715 3140
rect 27835 3020 27880 3140
rect 28000 3020 28045 3140
rect 28165 3020 28220 3140
rect 28340 3020 28385 3140
rect 28505 3020 28550 3140
rect 28670 3020 28715 3140
rect 28835 3020 28890 3140
rect 29010 3020 29055 3140
rect 29175 3020 29220 3140
rect 29340 3020 29385 3140
rect 29505 3020 29560 3140
rect 29680 3020 29690 3140
rect 24190 2965 29690 3020
rect 24190 2845 24200 2965
rect 24320 2845 24365 2965
rect 24485 2845 24530 2965
rect 24650 2845 24695 2965
rect 24815 2845 24870 2965
rect 24990 2845 25035 2965
rect 25155 2845 25200 2965
rect 25320 2845 25365 2965
rect 25485 2845 25540 2965
rect 25660 2845 25705 2965
rect 25825 2845 25870 2965
rect 25990 2845 26035 2965
rect 26155 2845 26210 2965
rect 26330 2845 26375 2965
rect 26495 2845 26540 2965
rect 26660 2845 26705 2965
rect 26825 2845 26880 2965
rect 27000 2845 27045 2965
rect 27165 2845 27210 2965
rect 27330 2845 27375 2965
rect 27495 2845 27550 2965
rect 27670 2845 27715 2965
rect 27835 2845 27880 2965
rect 28000 2845 28045 2965
rect 28165 2845 28220 2965
rect 28340 2845 28385 2965
rect 28505 2845 28550 2965
rect 28670 2845 28715 2965
rect 28835 2845 28890 2965
rect 29010 2845 29055 2965
rect 29175 2845 29220 2965
rect 29340 2845 29385 2965
rect 29505 2845 29560 2965
rect 29680 2845 29690 2965
rect 24190 2800 29690 2845
rect 24190 2680 24200 2800
rect 24320 2680 24365 2800
rect 24485 2680 24530 2800
rect 24650 2680 24695 2800
rect 24815 2680 24870 2800
rect 24990 2680 25035 2800
rect 25155 2680 25200 2800
rect 25320 2680 25365 2800
rect 25485 2680 25540 2800
rect 25660 2680 25705 2800
rect 25825 2680 25870 2800
rect 25990 2680 26035 2800
rect 26155 2680 26210 2800
rect 26330 2680 26375 2800
rect 26495 2680 26540 2800
rect 26660 2680 26705 2800
rect 26825 2680 26880 2800
rect 27000 2680 27045 2800
rect 27165 2680 27210 2800
rect 27330 2680 27375 2800
rect 27495 2680 27550 2800
rect 27670 2680 27715 2800
rect 27835 2680 27880 2800
rect 28000 2680 28045 2800
rect 28165 2680 28220 2800
rect 28340 2680 28385 2800
rect 28505 2680 28550 2800
rect 28670 2680 28715 2800
rect 28835 2680 28890 2800
rect 29010 2680 29055 2800
rect 29175 2680 29220 2800
rect 29340 2680 29385 2800
rect 29505 2680 29560 2800
rect 29680 2680 29690 2800
rect 24190 2635 29690 2680
rect 24190 2515 24200 2635
rect 24320 2515 24365 2635
rect 24485 2515 24530 2635
rect 24650 2515 24695 2635
rect 24815 2515 24870 2635
rect 24990 2515 25035 2635
rect 25155 2515 25200 2635
rect 25320 2515 25365 2635
rect 25485 2515 25540 2635
rect 25660 2515 25705 2635
rect 25825 2515 25870 2635
rect 25990 2515 26035 2635
rect 26155 2515 26210 2635
rect 26330 2515 26375 2635
rect 26495 2515 26540 2635
rect 26660 2515 26705 2635
rect 26825 2515 26880 2635
rect 27000 2515 27045 2635
rect 27165 2515 27210 2635
rect 27330 2515 27375 2635
rect 27495 2515 27550 2635
rect 27670 2515 27715 2635
rect 27835 2515 27880 2635
rect 28000 2515 28045 2635
rect 28165 2515 28220 2635
rect 28340 2515 28385 2635
rect 28505 2515 28550 2635
rect 28670 2515 28715 2635
rect 28835 2515 28890 2635
rect 29010 2515 29055 2635
rect 29175 2515 29220 2635
rect 29340 2515 29385 2635
rect 29505 2515 29560 2635
rect 29680 2515 29690 2635
rect 24190 2470 29690 2515
rect 24190 2350 24200 2470
rect 24320 2350 24365 2470
rect 24485 2350 24530 2470
rect 24650 2350 24695 2470
rect 24815 2350 24870 2470
rect 24990 2350 25035 2470
rect 25155 2350 25200 2470
rect 25320 2350 25365 2470
rect 25485 2350 25540 2470
rect 25660 2350 25705 2470
rect 25825 2350 25870 2470
rect 25990 2350 26035 2470
rect 26155 2350 26210 2470
rect 26330 2350 26375 2470
rect 26495 2350 26540 2470
rect 26660 2350 26705 2470
rect 26825 2350 26880 2470
rect 27000 2350 27045 2470
rect 27165 2350 27210 2470
rect 27330 2350 27375 2470
rect 27495 2350 27550 2470
rect 27670 2350 27715 2470
rect 27835 2350 27880 2470
rect 28000 2350 28045 2470
rect 28165 2350 28220 2470
rect 28340 2350 28385 2470
rect 28505 2350 28550 2470
rect 28670 2350 28715 2470
rect 28835 2350 28890 2470
rect 29010 2350 29055 2470
rect 29175 2350 29220 2470
rect 29340 2350 29385 2470
rect 29505 2350 29560 2470
rect 29680 2350 29690 2470
rect 24190 2295 29690 2350
rect 24190 2175 24200 2295
rect 24320 2175 24365 2295
rect 24485 2175 24530 2295
rect 24650 2175 24695 2295
rect 24815 2175 24870 2295
rect 24990 2175 25035 2295
rect 25155 2175 25200 2295
rect 25320 2175 25365 2295
rect 25485 2175 25540 2295
rect 25660 2175 25705 2295
rect 25825 2175 25870 2295
rect 25990 2175 26035 2295
rect 26155 2175 26210 2295
rect 26330 2175 26375 2295
rect 26495 2175 26540 2295
rect 26660 2175 26705 2295
rect 26825 2175 26880 2295
rect 27000 2175 27045 2295
rect 27165 2175 27210 2295
rect 27330 2175 27375 2295
rect 27495 2175 27550 2295
rect 27670 2175 27715 2295
rect 27835 2175 27880 2295
rect 28000 2175 28045 2295
rect 28165 2175 28220 2295
rect 28340 2175 28385 2295
rect 28505 2175 28550 2295
rect 28670 2175 28715 2295
rect 28835 2175 28890 2295
rect 29010 2175 29055 2295
rect 29175 2175 29220 2295
rect 29340 2175 29385 2295
rect 29505 2175 29560 2295
rect 29680 2175 29690 2295
rect 24190 2130 29690 2175
rect 24190 2010 24200 2130
rect 24320 2010 24365 2130
rect 24485 2010 24530 2130
rect 24650 2010 24695 2130
rect 24815 2010 24870 2130
rect 24990 2010 25035 2130
rect 25155 2010 25200 2130
rect 25320 2010 25365 2130
rect 25485 2010 25540 2130
rect 25660 2010 25705 2130
rect 25825 2010 25870 2130
rect 25990 2010 26035 2130
rect 26155 2010 26210 2130
rect 26330 2010 26375 2130
rect 26495 2010 26540 2130
rect 26660 2010 26705 2130
rect 26825 2010 26880 2130
rect 27000 2010 27045 2130
rect 27165 2010 27210 2130
rect 27330 2010 27375 2130
rect 27495 2010 27550 2130
rect 27670 2010 27715 2130
rect 27835 2010 27880 2130
rect 28000 2010 28045 2130
rect 28165 2010 28220 2130
rect 28340 2010 28385 2130
rect 28505 2010 28550 2130
rect 28670 2010 28715 2130
rect 28835 2010 28890 2130
rect 29010 2010 29055 2130
rect 29175 2010 29220 2130
rect 29340 2010 29385 2130
rect 29505 2010 29560 2130
rect 29680 2010 29690 2130
rect 24190 1965 29690 2010
rect 24190 1845 24200 1965
rect 24320 1845 24365 1965
rect 24485 1845 24530 1965
rect 24650 1845 24695 1965
rect 24815 1845 24870 1965
rect 24990 1845 25035 1965
rect 25155 1845 25200 1965
rect 25320 1845 25365 1965
rect 25485 1845 25540 1965
rect 25660 1845 25705 1965
rect 25825 1845 25870 1965
rect 25990 1845 26035 1965
rect 26155 1845 26210 1965
rect 26330 1845 26375 1965
rect 26495 1845 26540 1965
rect 26660 1845 26705 1965
rect 26825 1845 26880 1965
rect 27000 1845 27045 1965
rect 27165 1845 27210 1965
rect 27330 1845 27375 1965
rect 27495 1845 27550 1965
rect 27670 1845 27715 1965
rect 27835 1845 27880 1965
rect 28000 1845 28045 1965
rect 28165 1845 28220 1965
rect 28340 1845 28385 1965
rect 28505 1845 28550 1965
rect 28670 1845 28715 1965
rect 28835 1845 28890 1965
rect 29010 1845 29055 1965
rect 29175 1845 29220 1965
rect 29340 1845 29385 1965
rect 29505 1845 29560 1965
rect 29680 1845 29690 1965
rect 24190 1800 29690 1845
rect 24190 1680 24200 1800
rect 24320 1680 24365 1800
rect 24485 1680 24530 1800
rect 24650 1680 24695 1800
rect 24815 1680 24870 1800
rect 24990 1680 25035 1800
rect 25155 1680 25200 1800
rect 25320 1680 25365 1800
rect 25485 1680 25540 1800
rect 25660 1680 25705 1800
rect 25825 1680 25870 1800
rect 25990 1680 26035 1800
rect 26155 1680 26210 1800
rect 26330 1680 26375 1800
rect 26495 1680 26540 1800
rect 26660 1680 26705 1800
rect 26825 1680 26880 1800
rect 27000 1680 27045 1800
rect 27165 1680 27210 1800
rect 27330 1680 27375 1800
rect 27495 1680 27550 1800
rect 27670 1680 27715 1800
rect 27835 1680 27880 1800
rect 28000 1680 28045 1800
rect 28165 1680 28220 1800
rect 28340 1680 28385 1800
rect 28505 1680 28550 1800
rect 28670 1680 28715 1800
rect 28835 1680 28890 1800
rect 29010 1680 29055 1800
rect 29175 1680 29220 1800
rect 29340 1680 29385 1800
rect 29505 1680 29560 1800
rect 29680 1680 29690 1800
rect 24190 1670 29690 1680
rect 7120 1380 12620 1390
rect 7120 1260 7130 1380
rect 7250 1260 7305 1380
rect 7425 1260 7470 1380
rect 7590 1260 7635 1380
rect 7755 1260 7800 1380
rect 7920 1260 7975 1380
rect 8095 1260 8140 1380
rect 8260 1260 8305 1380
rect 8425 1260 8470 1380
rect 8590 1260 8645 1380
rect 8765 1260 8810 1380
rect 8930 1260 8975 1380
rect 9095 1260 9140 1380
rect 9260 1260 9315 1380
rect 9435 1260 9480 1380
rect 9600 1260 9645 1380
rect 9765 1260 9810 1380
rect 9930 1260 9985 1380
rect 10105 1260 10150 1380
rect 10270 1260 10315 1380
rect 10435 1260 10480 1380
rect 10600 1260 10655 1380
rect 10775 1260 10820 1380
rect 10940 1260 10985 1380
rect 11105 1260 11150 1380
rect 11270 1260 11325 1380
rect 11445 1260 11490 1380
rect 11610 1260 11655 1380
rect 11775 1260 11820 1380
rect 11940 1260 11995 1380
rect 12115 1260 12160 1380
rect 12280 1260 12325 1380
rect 12445 1260 12490 1380
rect 12610 1260 12620 1380
rect 7120 1215 12620 1260
rect 7120 1095 7130 1215
rect 7250 1095 7305 1215
rect 7425 1095 7470 1215
rect 7590 1095 7635 1215
rect 7755 1095 7800 1215
rect 7920 1095 7975 1215
rect 8095 1095 8140 1215
rect 8260 1095 8305 1215
rect 8425 1095 8470 1215
rect 8590 1095 8645 1215
rect 8765 1095 8810 1215
rect 8930 1095 8975 1215
rect 9095 1095 9140 1215
rect 9260 1095 9315 1215
rect 9435 1095 9480 1215
rect 9600 1095 9645 1215
rect 9765 1095 9810 1215
rect 9930 1095 9985 1215
rect 10105 1095 10150 1215
rect 10270 1095 10315 1215
rect 10435 1095 10480 1215
rect 10600 1095 10655 1215
rect 10775 1095 10820 1215
rect 10940 1095 10985 1215
rect 11105 1095 11150 1215
rect 11270 1095 11325 1215
rect 11445 1095 11490 1215
rect 11610 1095 11655 1215
rect 11775 1095 11820 1215
rect 11940 1095 11995 1215
rect 12115 1095 12160 1215
rect 12280 1095 12325 1215
rect 12445 1095 12490 1215
rect 12610 1095 12620 1215
rect 7120 1050 12620 1095
rect 7120 930 7130 1050
rect 7250 930 7305 1050
rect 7425 930 7470 1050
rect 7590 930 7635 1050
rect 7755 930 7800 1050
rect 7920 930 7975 1050
rect 8095 930 8140 1050
rect 8260 930 8305 1050
rect 8425 930 8470 1050
rect 8590 930 8645 1050
rect 8765 930 8810 1050
rect 8930 930 8975 1050
rect 9095 930 9140 1050
rect 9260 930 9315 1050
rect 9435 930 9480 1050
rect 9600 930 9645 1050
rect 9765 930 9810 1050
rect 9930 930 9985 1050
rect 10105 930 10150 1050
rect 10270 930 10315 1050
rect 10435 930 10480 1050
rect 10600 930 10655 1050
rect 10775 930 10820 1050
rect 10940 930 10985 1050
rect 11105 930 11150 1050
rect 11270 930 11325 1050
rect 11445 930 11490 1050
rect 11610 930 11655 1050
rect 11775 930 11820 1050
rect 11940 930 11995 1050
rect 12115 930 12160 1050
rect 12280 930 12325 1050
rect 12445 930 12490 1050
rect 12610 930 12620 1050
rect 7120 885 12620 930
rect 7120 765 7130 885
rect 7250 765 7305 885
rect 7425 765 7470 885
rect 7590 765 7635 885
rect 7755 765 7800 885
rect 7920 765 7975 885
rect 8095 765 8140 885
rect 8260 765 8305 885
rect 8425 765 8470 885
rect 8590 765 8645 885
rect 8765 765 8810 885
rect 8930 765 8975 885
rect 9095 765 9140 885
rect 9260 765 9315 885
rect 9435 765 9480 885
rect 9600 765 9645 885
rect 9765 765 9810 885
rect 9930 765 9985 885
rect 10105 765 10150 885
rect 10270 765 10315 885
rect 10435 765 10480 885
rect 10600 765 10655 885
rect 10775 765 10820 885
rect 10940 765 10985 885
rect 11105 765 11150 885
rect 11270 765 11325 885
rect 11445 765 11490 885
rect 11610 765 11655 885
rect 11775 765 11820 885
rect 11940 765 11995 885
rect 12115 765 12160 885
rect 12280 765 12325 885
rect 12445 765 12490 885
rect 12610 765 12620 885
rect 7120 710 12620 765
rect 7120 590 7130 710
rect 7250 590 7305 710
rect 7425 590 7470 710
rect 7590 590 7635 710
rect 7755 590 7800 710
rect 7920 590 7975 710
rect 8095 590 8140 710
rect 8260 590 8305 710
rect 8425 590 8470 710
rect 8590 590 8645 710
rect 8765 590 8810 710
rect 8930 590 8975 710
rect 9095 590 9140 710
rect 9260 590 9315 710
rect 9435 590 9480 710
rect 9600 590 9645 710
rect 9765 590 9810 710
rect 9930 590 9985 710
rect 10105 590 10150 710
rect 10270 590 10315 710
rect 10435 590 10480 710
rect 10600 590 10655 710
rect 10775 590 10820 710
rect 10940 590 10985 710
rect 11105 590 11150 710
rect 11270 590 11325 710
rect 11445 590 11490 710
rect 11610 590 11655 710
rect 11775 590 11820 710
rect 11940 590 11995 710
rect 12115 590 12160 710
rect 12280 590 12325 710
rect 12445 590 12490 710
rect 12610 590 12620 710
rect 7120 545 12620 590
rect 7120 425 7130 545
rect 7250 425 7305 545
rect 7425 425 7470 545
rect 7590 425 7635 545
rect 7755 425 7800 545
rect 7920 425 7975 545
rect 8095 425 8140 545
rect 8260 425 8305 545
rect 8425 425 8470 545
rect 8590 425 8645 545
rect 8765 425 8810 545
rect 8930 425 8975 545
rect 9095 425 9140 545
rect 9260 425 9315 545
rect 9435 425 9480 545
rect 9600 425 9645 545
rect 9765 425 9810 545
rect 9930 425 9985 545
rect 10105 425 10150 545
rect 10270 425 10315 545
rect 10435 425 10480 545
rect 10600 425 10655 545
rect 10775 425 10820 545
rect 10940 425 10985 545
rect 11105 425 11150 545
rect 11270 425 11325 545
rect 11445 425 11490 545
rect 11610 425 11655 545
rect 11775 425 11820 545
rect 11940 425 11995 545
rect 12115 425 12160 545
rect 12280 425 12325 545
rect 12445 425 12490 545
rect 12610 425 12620 545
rect 7120 380 12620 425
rect 7120 260 7130 380
rect 7250 260 7305 380
rect 7425 260 7470 380
rect 7590 260 7635 380
rect 7755 260 7800 380
rect 7920 260 7975 380
rect 8095 260 8140 380
rect 8260 260 8305 380
rect 8425 260 8470 380
rect 8590 260 8645 380
rect 8765 260 8810 380
rect 8930 260 8975 380
rect 9095 260 9140 380
rect 9260 260 9315 380
rect 9435 260 9480 380
rect 9600 260 9645 380
rect 9765 260 9810 380
rect 9930 260 9985 380
rect 10105 260 10150 380
rect 10270 260 10315 380
rect 10435 260 10480 380
rect 10600 260 10655 380
rect 10775 260 10820 380
rect 10940 260 10985 380
rect 11105 260 11150 380
rect 11270 260 11325 380
rect 11445 260 11490 380
rect 11610 260 11655 380
rect 11775 260 11820 380
rect 11940 260 11995 380
rect 12115 260 12160 380
rect 12280 260 12325 380
rect 12445 260 12490 380
rect 12610 260 12620 380
rect 7120 215 12620 260
rect 7120 95 7130 215
rect 7250 95 7305 215
rect 7425 95 7470 215
rect 7590 95 7635 215
rect 7755 95 7800 215
rect 7920 95 7975 215
rect 8095 95 8140 215
rect 8260 95 8305 215
rect 8425 95 8470 215
rect 8590 95 8645 215
rect 8765 95 8810 215
rect 8930 95 8975 215
rect 9095 95 9140 215
rect 9260 95 9315 215
rect 9435 95 9480 215
rect 9600 95 9645 215
rect 9765 95 9810 215
rect 9930 95 9985 215
rect 10105 95 10150 215
rect 10270 95 10315 215
rect 10435 95 10480 215
rect 10600 95 10655 215
rect 10775 95 10820 215
rect 10940 95 10985 215
rect 11105 95 11150 215
rect 11270 95 11325 215
rect 11445 95 11490 215
rect 11610 95 11655 215
rect 11775 95 11820 215
rect 11940 95 11995 215
rect 12115 95 12160 215
rect 12280 95 12325 215
rect 12445 95 12490 215
rect 12610 95 12620 215
rect 7120 40 12620 95
rect 7120 -80 7130 40
rect 7250 -80 7305 40
rect 7425 -80 7470 40
rect 7590 -80 7635 40
rect 7755 -80 7800 40
rect 7920 -80 7975 40
rect 8095 -80 8140 40
rect 8260 -80 8305 40
rect 8425 -80 8470 40
rect 8590 -80 8645 40
rect 8765 -80 8810 40
rect 8930 -80 8975 40
rect 9095 -80 9140 40
rect 9260 -80 9315 40
rect 9435 -80 9480 40
rect 9600 -80 9645 40
rect 9765 -80 9810 40
rect 9930 -80 9985 40
rect 10105 -80 10150 40
rect 10270 -80 10315 40
rect 10435 -80 10480 40
rect 10600 -80 10655 40
rect 10775 -80 10820 40
rect 10940 -80 10985 40
rect 11105 -80 11150 40
rect 11270 -80 11325 40
rect 11445 -80 11490 40
rect 11610 -80 11655 40
rect 11775 -80 11820 40
rect 11940 -80 11995 40
rect 12115 -80 12160 40
rect 12280 -80 12325 40
rect 12445 -80 12490 40
rect 12610 -80 12620 40
rect 7120 -125 12620 -80
rect 7120 -245 7130 -125
rect 7250 -245 7305 -125
rect 7425 -245 7470 -125
rect 7590 -245 7635 -125
rect 7755 -245 7800 -125
rect 7920 -245 7975 -125
rect 8095 -245 8140 -125
rect 8260 -245 8305 -125
rect 8425 -245 8470 -125
rect 8590 -245 8645 -125
rect 8765 -245 8810 -125
rect 8930 -245 8975 -125
rect 9095 -245 9140 -125
rect 9260 -245 9315 -125
rect 9435 -245 9480 -125
rect 9600 -245 9645 -125
rect 9765 -245 9810 -125
rect 9930 -245 9985 -125
rect 10105 -245 10150 -125
rect 10270 -245 10315 -125
rect 10435 -245 10480 -125
rect 10600 -245 10655 -125
rect 10775 -245 10820 -125
rect 10940 -245 10985 -125
rect 11105 -245 11150 -125
rect 11270 -245 11325 -125
rect 11445 -245 11490 -125
rect 11610 -245 11655 -125
rect 11775 -245 11820 -125
rect 11940 -245 11995 -125
rect 12115 -245 12160 -125
rect 12280 -245 12325 -125
rect 12445 -245 12490 -125
rect 12610 -245 12620 -125
rect 7120 -290 12620 -245
rect 7120 -410 7130 -290
rect 7250 -410 7305 -290
rect 7425 -410 7470 -290
rect 7590 -410 7635 -290
rect 7755 -410 7800 -290
rect 7920 -410 7975 -290
rect 8095 -410 8140 -290
rect 8260 -410 8305 -290
rect 8425 -410 8470 -290
rect 8590 -410 8645 -290
rect 8765 -410 8810 -290
rect 8930 -410 8975 -290
rect 9095 -410 9140 -290
rect 9260 -410 9315 -290
rect 9435 -410 9480 -290
rect 9600 -410 9645 -290
rect 9765 -410 9810 -290
rect 9930 -410 9985 -290
rect 10105 -410 10150 -290
rect 10270 -410 10315 -290
rect 10435 -410 10480 -290
rect 10600 -410 10655 -290
rect 10775 -410 10820 -290
rect 10940 -410 10985 -290
rect 11105 -410 11150 -290
rect 11270 -410 11325 -290
rect 11445 -410 11490 -290
rect 11610 -410 11655 -290
rect 11775 -410 11820 -290
rect 11940 -410 11995 -290
rect 12115 -410 12160 -290
rect 12280 -410 12325 -290
rect 12445 -410 12490 -290
rect 12610 -410 12620 -290
rect 7120 -455 12620 -410
rect 7120 -575 7130 -455
rect 7250 -575 7305 -455
rect 7425 -575 7470 -455
rect 7590 -575 7635 -455
rect 7755 -575 7800 -455
rect 7920 -575 7975 -455
rect 8095 -575 8140 -455
rect 8260 -575 8305 -455
rect 8425 -575 8470 -455
rect 8590 -575 8645 -455
rect 8765 -575 8810 -455
rect 8930 -575 8975 -455
rect 9095 -575 9140 -455
rect 9260 -575 9315 -455
rect 9435 -575 9480 -455
rect 9600 -575 9645 -455
rect 9765 -575 9810 -455
rect 9930 -575 9985 -455
rect 10105 -575 10150 -455
rect 10270 -575 10315 -455
rect 10435 -575 10480 -455
rect 10600 -575 10655 -455
rect 10775 -575 10820 -455
rect 10940 -575 10985 -455
rect 11105 -575 11150 -455
rect 11270 -575 11325 -455
rect 11445 -575 11490 -455
rect 11610 -575 11655 -455
rect 11775 -575 11820 -455
rect 11940 -575 11995 -455
rect 12115 -575 12160 -455
rect 12280 -575 12325 -455
rect 12445 -575 12490 -455
rect 12610 -575 12620 -455
rect 7120 -630 12620 -575
rect 7120 -750 7130 -630
rect 7250 -750 7305 -630
rect 7425 -750 7470 -630
rect 7590 -750 7635 -630
rect 7755 -750 7800 -630
rect 7920 -750 7975 -630
rect 8095 -750 8140 -630
rect 8260 -750 8305 -630
rect 8425 -750 8470 -630
rect 8590 -750 8645 -630
rect 8765 -750 8810 -630
rect 8930 -750 8975 -630
rect 9095 -750 9140 -630
rect 9260 -750 9315 -630
rect 9435 -750 9480 -630
rect 9600 -750 9645 -630
rect 9765 -750 9810 -630
rect 9930 -750 9985 -630
rect 10105 -750 10150 -630
rect 10270 -750 10315 -630
rect 10435 -750 10480 -630
rect 10600 -750 10655 -630
rect 10775 -750 10820 -630
rect 10940 -750 10985 -630
rect 11105 -750 11150 -630
rect 11270 -750 11325 -630
rect 11445 -750 11490 -630
rect 11610 -750 11655 -630
rect 11775 -750 11820 -630
rect 11940 -750 11995 -630
rect 12115 -750 12160 -630
rect 12280 -750 12325 -630
rect 12445 -750 12490 -630
rect 12610 -750 12620 -630
rect 7120 -795 12620 -750
rect 7120 -915 7130 -795
rect 7250 -915 7305 -795
rect 7425 -915 7470 -795
rect 7590 -915 7635 -795
rect 7755 -915 7800 -795
rect 7920 -915 7975 -795
rect 8095 -915 8140 -795
rect 8260 -915 8305 -795
rect 8425 -915 8470 -795
rect 8590 -915 8645 -795
rect 8765 -915 8810 -795
rect 8930 -915 8975 -795
rect 9095 -915 9140 -795
rect 9260 -915 9315 -795
rect 9435 -915 9480 -795
rect 9600 -915 9645 -795
rect 9765 -915 9810 -795
rect 9930 -915 9985 -795
rect 10105 -915 10150 -795
rect 10270 -915 10315 -795
rect 10435 -915 10480 -795
rect 10600 -915 10655 -795
rect 10775 -915 10820 -795
rect 10940 -915 10985 -795
rect 11105 -915 11150 -795
rect 11270 -915 11325 -795
rect 11445 -915 11490 -795
rect 11610 -915 11655 -795
rect 11775 -915 11820 -795
rect 11940 -915 11995 -795
rect 12115 -915 12160 -795
rect 12280 -915 12325 -795
rect 12445 -915 12490 -795
rect 12610 -915 12620 -795
rect 7120 -960 12620 -915
rect 7120 -1080 7130 -960
rect 7250 -1080 7305 -960
rect 7425 -1080 7470 -960
rect 7590 -1080 7635 -960
rect 7755 -1080 7800 -960
rect 7920 -1080 7975 -960
rect 8095 -1080 8140 -960
rect 8260 -1080 8305 -960
rect 8425 -1080 8470 -960
rect 8590 -1080 8645 -960
rect 8765 -1080 8810 -960
rect 8930 -1080 8975 -960
rect 9095 -1080 9140 -960
rect 9260 -1080 9315 -960
rect 9435 -1080 9480 -960
rect 9600 -1080 9645 -960
rect 9765 -1080 9810 -960
rect 9930 -1080 9985 -960
rect 10105 -1080 10150 -960
rect 10270 -1080 10315 -960
rect 10435 -1080 10480 -960
rect 10600 -1080 10655 -960
rect 10775 -1080 10820 -960
rect 10940 -1080 10985 -960
rect 11105 -1080 11150 -960
rect 11270 -1080 11325 -960
rect 11445 -1080 11490 -960
rect 11610 -1080 11655 -960
rect 11775 -1080 11820 -960
rect 11940 -1080 11995 -960
rect 12115 -1080 12160 -960
rect 12280 -1080 12325 -960
rect 12445 -1080 12490 -960
rect 12610 -1080 12620 -960
rect 7120 -1125 12620 -1080
rect 7120 -1245 7130 -1125
rect 7250 -1245 7305 -1125
rect 7425 -1245 7470 -1125
rect 7590 -1245 7635 -1125
rect 7755 -1245 7800 -1125
rect 7920 -1245 7975 -1125
rect 8095 -1245 8140 -1125
rect 8260 -1245 8305 -1125
rect 8425 -1245 8470 -1125
rect 8590 -1245 8645 -1125
rect 8765 -1245 8810 -1125
rect 8930 -1245 8975 -1125
rect 9095 -1245 9140 -1125
rect 9260 -1245 9315 -1125
rect 9435 -1245 9480 -1125
rect 9600 -1245 9645 -1125
rect 9765 -1245 9810 -1125
rect 9930 -1245 9985 -1125
rect 10105 -1245 10150 -1125
rect 10270 -1245 10315 -1125
rect 10435 -1245 10480 -1125
rect 10600 -1245 10655 -1125
rect 10775 -1245 10820 -1125
rect 10940 -1245 10985 -1125
rect 11105 -1245 11150 -1125
rect 11270 -1245 11325 -1125
rect 11445 -1245 11490 -1125
rect 11610 -1245 11655 -1125
rect 11775 -1245 11820 -1125
rect 11940 -1245 11995 -1125
rect 12115 -1245 12160 -1125
rect 12280 -1245 12325 -1125
rect 12445 -1245 12490 -1125
rect 12610 -1245 12620 -1125
rect 7120 -1300 12620 -1245
rect 7120 -1420 7130 -1300
rect 7250 -1420 7305 -1300
rect 7425 -1420 7470 -1300
rect 7590 -1420 7635 -1300
rect 7755 -1420 7800 -1300
rect 7920 -1420 7975 -1300
rect 8095 -1420 8140 -1300
rect 8260 -1420 8305 -1300
rect 8425 -1420 8470 -1300
rect 8590 -1420 8645 -1300
rect 8765 -1420 8810 -1300
rect 8930 -1420 8975 -1300
rect 9095 -1420 9140 -1300
rect 9260 -1420 9315 -1300
rect 9435 -1420 9480 -1300
rect 9600 -1420 9645 -1300
rect 9765 -1420 9810 -1300
rect 9930 -1420 9985 -1300
rect 10105 -1420 10150 -1300
rect 10270 -1420 10315 -1300
rect 10435 -1420 10480 -1300
rect 10600 -1420 10655 -1300
rect 10775 -1420 10820 -1300
rect 10940 -1420 10985 -1300
rect 11105 -1420 11150 -1300
rect 11270 -1420 11325 -1300
rect 11445 -1420 11490 -1300
rect 11610 -1420 11655 -1300
rect 11775 -1420 11820 -1300
rect 11940 -1420 11995 -1300
rect 12115 -1420 12160 -1300
rect 12280 -1420 12325 -1300
rect 12445 -1420 12490 -1300
rect 12610 -1420 12620 -1300
rect 7120 -1465 12620 -1420
rect 7120 -1585 7130 -1465
rect 7250 -1585 7305 -1465
rect 7425 -1585 7470 -1465
rect 7590 -1585 7635 -1465
rect 7755 -1585 7800 -1465
rect 7920 -1585 7975 -1465
rect 8095 -1585 8140 -1465
rect 8260 -1585 8305 -1465
rect 8425 -1585 8470 -1465
rect 8590 -1585 8645 -1465
rect 8765 -1585 8810 -1465
rect 8930 -1585 8975 -1465
rect 9095 -1585 9140 -1465
rect 9260 -1585 9315 -1465
rect 9435 -1585 9480 -1465
rect 9600 -1585 9645 -1465
rect 9765 -1585 9810 -1465
rect 9930 -1585 9985 -1465
rect 10105 -1585 10150 -1465
rect 10270 -1585 10315 -1465
rect 10435 -1585 10480 -1465
rect 10600 -1585 10655 -1465
rect 10775 -1585 10820 -1465
rect 10940 -1585 10985 -1465
rect 11105 -1585 11150 -1465
rect 11270 -1585 11325 -1465
rect 11445 -1585 11490 -1465
rect 11610 -1585 11655 -1465
rect 11775 -1585 11820 -1465
rect 11940 -1585 11995 -1465
rect 12115 -1585 12160 -1465
rect 12280 -1585 12325 -1465
rect 12445 -1585 12490 -1465
rect 12610 -1585 12620 -1465
rect 7120 -1630 12620 -1585
rect 7120 -1750 7130 -1630
rect 7250 -1750 7305 -1630
rect 7425 -1750 7470 -1630
rect 7590 -1750 7635 -1630
rect 7755 -1750 7800 -1630
rect 7920 -1750 7975 -1630
rect 8095 -1750 8140 -1630
rect 8260 -1750 8305 -1630
rect 8425 -1750 8470 -1630
rect 8590 -1750 8645 -1630
rect 8765 -1750 8810 -1630
rect 8930 -1750 8975 -1630
rect 9095 -1750 9140 -1630
rect 9260 -1750 9315 -1630
rect 9435 -1750 9480 -1630
rect 9600 -1750 9645 -1630
rect 9765 -1750 9810 -1630
rect 9930 -1750 9985 -1630
rect 10105 -1750 10150 -1630
rect 10270 -1750 10315 -1630
rect 10435 -1750 10480 -1630
rect 10600 -1750 10655 -1630
rect 10775 -1750 10820 -1630
rect 10940 -1750 10985 -1630
rect 11105 -1750 11150 -1630
rect 11270 -1750 11325 -1630
rect 11445 -1750 11490 -1630
rect 11610 -1750 11655 -1630
rect 11775 -1750 11820 -1630
rect 11940 -1750 11995 -1630
rect 12115 -1750 12160 -1630
rect 12280 -1750 12325 -1630
rect 12445 -1750 12490 -1630
rect 12610 -1750 12620 -1630
rect 7120 -1795 12620 -1750
rect 7120 -1915 7130 -1795
rect 7250 -1915 7305 -1795
rect 7425 -1915 7470 -1795
rect 7590 -1915 7635 -1795
rect 7755 -1915 7800 -1795
rect 7920 -1915 7975 -1795
rect 8095 -1915 8140 -1795
rect 8260 -1915 8305 -1795
rect 8425 -1915 8470 -1795
rect 8590 -1915 8645 -1795
rect 8765 -1915 8810 -1795
rect 8930 -1915 8975 -1795
rect 9095 -1915 9140 -1795
rect 9260 -1915 9315 -1795
rect 9435 -1915 9480 -1795
rect 9600 -1915 9645 -1795
rect 9765 -1915 9810 -1795
rect 9930 -1915 9985 -1795
rect 10105 -1915 10150 -1795
rect 10270 -1915 10315 -1795
rect 10435 -1915 10480 -1795
rect 10600 -1915 10655 -1795
rect 10775 -1915 10820 -1795
rect 10940 -1915 10985 -1795
rect 11105 -1915 11150 -1795
rect 11270 -1915 11325 -1795
rect 11445 -1915 11490 -1795
rect 11610 -1915 11655 -1795
rect 11775 -1915 11820 -1795
rect 11940 -1915 11995 -1795
rect 12115 -1915 12160 -1795
rect 12280 -1915 12325 -1795
rect 12445 -1915 12490 -1795
rect 12610 -1915 12620 -1795
rect 7120 -1970 12620 -1915
rect 7120 -2090 7130 -1970
rect 7250 -2090 7305 -1970
rect 7425 -2090 7470 -1970
rect 7590 -2090 7635 -1970
rect 7755 -2090 7800 -1970
rect 7920 -2090 7975 -1970
rect 8095 -2090 8140 -1970
rect 8260 -2090 8305 -1970
rect 8425 -2090 8470 -1970
rect 8590 -2090 8645 -1970
rect 8765 -2090 8810 -1970
rect 8930 -2090 8975 -1970
rect 9095 -2090 9140 -1970
rect 9260 -2090 9315 -1970
rect 9435 -2090 9480 -1970
rect 9600 -2090 9645 -1970
rect 9765 -2090 9810 -1970
rect 9930 -2090 9985 -1970
rect 10105 -2090 10150 -1970
rect 10270 -2090 10315 -1970
rect 10435 -2090 10480 -1970
rect 10600 -2090 10655 -1970
rect 10775 -2090 10820 -1970
rect 10940 -2090 10985 -1970
rect 11105 -2090 11150 -1970
rect 11270 -2090 11325 -1970
rect 11445 -2090 11490 -1970
rect 11610 -2090 11655 -1970
rect 11775 -2090 11820 -1970
rect 11940 -2090 11995 -1970
rect 12115 -2090 12160 -1970
rect 12280 -2090 12325 -1970
rect 12445 -2090 12490 -1970
rect 12610 -2090 12620 -1970
rect 7120 -2135 12620 -2090
rect 7120 -2255 7130 -2135
rect 7250 -2255 7305 -2135
rect 7425 -2255 7470 -2135
rect 7590 -2255 7635 -2135
rect 7755 -2255 7800 -2135
rect 7920 -2255 7975 -2135
rect 8095 -2255 8140 -2135
rect 8260 -2255 8305 -2135
rect 8425 -2255 8470 -2135
rect 8590 -2255 8645 -2135
rect 8765 -2255 8810 -2135
rect 8930 -2255 8975 -2135
rect 9095 -2255 9140 -2135
rect 9260 -2255 9315 -2135
rect 9435 -2255 9480 -2135
rect 9600 -2255 9645 -2135
rect 9765 -2255 9810 -2135
rect 9930 -2255 9985 -2135
rect 10105 -2255 10150 -2135
rect 10270 -2255 10315 -2135
rect 10435 -2255 10480 -2135
rect 10600 -2255 10655 -2135
rect 10775 -2255 10820 -2135
rect 10940 -2255 10985 -2135
rect 11105 -2255 11150 -2135
rect 11270 -2255 11325 -2135
rect 11445 -2255 11490 -2135
rect 11610 -2255 11655 -2135
rect 11775 -2255 11820 -2135
rect 11940 -2255 11995 -2135
rect 12115 -2255 12160 -2135
rect 12280 -2255 12325 -2135
rect 12445 -2255 12490 -2135
rect 12610 -2255 12620 -2135
rect 7120 -2300 12620 -2255
rect 7120 -2420 7130 -2300
rect 7250 -2420 7305 -2300
rect 7425 -2420 7470 -2300
rect 7590 -2420 7635 -2300
rect 7755 -2420 7800 -2300
rect 7920 -2420 7975 -2300
rect 8095 -2420 8140 -2300
rect 8260 -2420 8305 -2300
rect 8425 -2420 8470 -2300
rect 8590 -2420 8645 -2300
rect 8765 -2420 8810 -2300
rect 8930 -2420 8975 -2300
rect 9095 -2420 9140 -2300
rect 9260 -2420 9315 -2300
rect 9435 -2420 9480 -2300
rect 9600 -2420 9645 -2300
rect 9765 -2420 9810 -2300
rect 9930 -2420 9985 -2300
rect 10105 -2420 10150 -2300
rect 10270 -2420 10315 -2300
rect 10435 -2420 10480 -2300
rect 10600 -2420 10655 -2300
rect 10775 -2420 10820 -2300
rect 10940 -2420 10985 -2300
rect 11105 -2420 11150 -2300
rect 11270 -2420 11325 -2300
rect 11445 -2420 11490 -2300
rect 11610 -2420 11655 -2300
rect 11775 -2420 11820 -2300
rect 11940 -2420 11995 -2300
rect 12115 -2420 12160 -2300
rect 12280 -2420 12325 -2300
rect 12445 -2420 12490 -2300
rect 12610 -2420 12620 -2300
rect 7120 -2465 12620 -2420
rect 7120 -2585 7130 -2465
rect 7250 -2585 7305 -2465
rect 7425 -2585 7470 -2465
rect 7590 -2585 7635 -2465
rect 7755 -2585 7800 -2465
rect 7920 -2585 7975 -2465
rect 8095 -2585 8140 -2465
rect 8260 -2585 8305 -2465
rect 8425 -2585 8470 -2465
rect 8590 -2585 8645 -2465
rect 8765 -2585 8810 -2465
rect 8930 -2585 8975 -2465
rect 9095 -2585 9140 -2465
rect 9260 -2585 9315 -2465
rect 9435 -2585 9480 -2465
rect 9600 -2585 9645 -2465
rect 9765 -2585 9810 -2465
rect 9930 -2585 9985 -2465
rect 10105 -2585 10150 -2465
rect 10270 -2585 10315 -2465
rect 10435 -2585 10480 -2465
rect 10600 -2585 10655 -2465
rect 10775 -2585 10820 -2465
rect 10940 -2585 10985 -2465
rect 11105 -2585 11150 -2465
rect 11270 -2585 11325 -2465
rect 11445 -2585 11490 -2465
rect 11610 -2585 11655 -2465
rect 11775 -2585 11820 -2465
rect 11940 -2585 11995 -2465
rect 12115 -2585 12160 -2465
rect 12280 -2585 12325 -2465
rect 12445 -2585 12490 -2465
rect 12610 -2585 12620 -2465
rect 7120 -2640 12620 -2585
rect 7120 -2760 7130 -2640
rect 7250 -2760 7305 -2640
rect 7425 -2760 7470 -2640
rect 7590 -2760 7635 -2640
rect 7755 -2760 7800 -2640
rect 7920 -2760 7975 -2640
rect 8095 -2760 8140 -2640
rect 8260 -2760 8305 -2640
rect 8425 -2760 8470 -2640
rect 8590 -2760 8645 -2640
rect 8765 -2760 8810 -2640
rect 8930 -2760 8975 -2640
rect 9095 -2760 9140 -2640
rect 9260 -2760 9315 -2640
rect 9435 -2760 9480 -2640
rect 9600 -2760 9645 -2640
rect 9765 -2760 9810 -2640
rect 9930 -2760 9985 -2640
rect 10105 -2760 10150 -2640
rect 10270 -2760 10315 -2640
rect 10435 -2760 10480 -2640
rect 10600 -2760 10655 -2640
rect 10775 -2760 10820 -2640
rect 10940 -2760 10985 -2640
rect 11105 -2760 11150 -2640
rect 11270 -2760 11325 -2640
rect 11445 -2760 11490 -2640
rect 11610 -2760 11655 -2640
rect 11775 -2760 11820 -2640
rect 11940 -2760 11995 -2640
rect 12115 -2760 12160 -2640
rect 12280 -2760 12325 -2640
rect 12445 -2760 12490 -2640
rect 12610 -2760 12620 -2640
rect 7120 -2805 12620 -2760
rect 7120 -2925 7130 -2805
rect 7250 -2925 7305 -2805
rect 7425 -2925 7470 -2805
rect 7590 -2925 7635 -2805
rect 7755 -2925 7800 -2805
rect 7920 -2925 7975 -2805
rect 8095 -2925 8140 -2805
rect 8260 -2925 8305 -2805
rect 8425 -2925 8470 -2805
rect 8590 -2925 8645 -2805
rect 8765 -2925 8810 -2805
rect 8930 -2925 8975 -2805
rect 9095 -2925 9140 -2805
rect 9260 -2925 9315 -2805
rect 9435 -2925 9480 -2805
rect 9600 -2925 9645 -2805
rect 9765 -2925 9810 -2805
rect 9930 -2925 9985 -2805
rect 10105 -2925 10150 -2805
rect 10270 -2925 10315 -2805
rect 10435 -2925 10480 -2805
rect 10600 -2925 10655 -2805
rect 10775 -2925 10820 -2805
rect 10940 -2925 10985 -2805
rect 11105 -2925 11150 -2805
rect 11270 -2925 11325 -2805
rect 11445 -2925 11490 -2805
rect 11610 -2925 11655 -2805
rect 11775 -2925 11820 -2805
rect 11940 -2925 11995 -2805
rect 12115 -2925 12160 -2805
rect 12280 -2925 12325 -2805
rect 12445 -2925 12490 -2805
rect 12610 -2925 12620 -2805
rect 7120 -2970 12620 -2925
rect 7120 -3090 7130 -2970
rect 7250 -3090 7305 -2970
rect 7425 -3090 7470 -2970
rect 7590 -3090 7635 -2970
rect 7755 -3090 7800 -2970
rect 7920 -3090 7975 -2970
rect 8095 -3090 8140 -2970
rect 8260 -3090 8305 -2970
rect 8425 -3090 8470 -2970
rect 8590 -3090 8645 -2970
rect 8765 -3090 8810 -2970
rect 8930 -3090 8975 -2970
rect 9095 -3090 9140 -2970
rect 9260 -3090 9315 -2970
rect 9435 -3090 9480 -2970
rect 9600 -3090 9645 -2970
rect 9765 -3090 9810 -2970
rect 9930 -3090 9985 -2970
rect 10105 -3090 10150 -2970
rect 10270 -3090 10315 -2970
rect 10435 -3090 10480 -2970
rect 10600 -3090 10655 -2970
rect 10775 -3090 10820 -2970
rect 10940 -3090 10985 -2970
rect 11105 -3090 11150 -2970
rect 11270 -3090 11325 -2970
rect 11445 -3090 11490 -2970
rect 11610 -3090 11655 -2970
rect 11775 -3090 11820 -2970
rect 11940 -3090 11995 -2970
rect 12115 -3090 12160 -2970
rect 12280 -3090 12325 -2970
rect 12445 -3090 12490 -2970
rect 12610 -3090 12620 -2970
rect 7120 -3135 12620 -3090
rect 7120 -3255 7130 -3135
rect 7250 -3255 7305 -3135
rect 7425 -3255 7470 -3135
rect 7590 -3255 7635 -3135
rect 7755 -3255 7800 -3135
rect 7920 -3255 7975 -3135
rect 8095 -3255 8140 -3135
rect 8260 -3255 8305 -3135
rect 8425 -3255 8470 -3135
rect 8590 -3255 8645 -3135
rect 8765 -3255 8810 -3135
rect 8930 -3255 8975 -3135
rect 9095 -3255 9140 -3135
rect 9260 -3255 9315 -3135
rect 9435 -3255 9480 -3135
rect 9600 -3255 9645 -3135
rect 9765 -3255 9810 -3135
rect 9930 -3255 9985 -3135
rect 10105 -3255 10150 -3135
rect 10270 -3255 10315 -3135
rect 10435 -3255 10480 -3135
rect 10600 -3255 10655 -3135
rect 10775 -3255 10820 -3135
rect 10940 -3255 10985 -3135
rect 11105 -3255 11150 -3135
rect 11270 -3255 11325 -3135
rect 11445 -3255 11490 -3135
rect 11610 -3255 11655 -3135
rect 11775 -3255 11820 -3135
rect 11940 -3255 11995 -3135
rect 12115 -3255 12160 -3135
rect 12280 -3255 12325 -3135
rect 12445 -3255 12490 -3135
rect 12610 -3255 12620 -3135
rect 7120 -3310 12620 -3255
rect 7120 -3430 7130 -3310
rect 7250 -3430 7305 -3310
rect 7425 -3430 7470 -3310
rect 7590 -3430 7635 -3310
rect 7755 -3430 7800 -3310
rect 7920 -3430 7975 -3310
rect 8095 -3430 8140 -3310
rect 8260 -3430 8305 -3310
rect 8425 -3430 8470 -3310
rect 8590 -3430 8645 -3310
rect 8765 -3430 8810 -3310
rect 8930 -3430 8975 -3310
rect 9095 -3430 9140 -3310
rect 9260 -3430 9315 -3310
rect 9435 -3430 9480 -3310
rect 9600 -3430 9645 -3310
rect 9765 -3430 9810 -3310
rect 9930 -3430 9985 -3310
rect 10105 -3430 10150 -3310
rect 10270 -3430 10315 -3310
rect 10435 -3430 10480 -3310
rect 10600 -3430 10655 -3310
rect 10775 -3430 10820 -3310
rect 10940 -3430 10985 -3310
rect 11105 -3430 11150 -3310
rect 11270 -3430 11325 -3310
rect 11445 -3430 11490 -3310
rect 11610 -3430 11655 -3310
rect 11775 -3430 11820 -3310
rect 11940 -3430 11995 -3310
rect 12115 -3430 12160 -3310
rect 12280 -3430 12325 -3310
rect 12445 -3430 12490 -3310
rect 12610 -3430 12620 -3310
rect 7120 -3475 12620 -3430
rect 7120 -3595 7130 -3475
rect 7250 -3595 7305 -3475
rect 7425 -3595 7470 -3475
rect 7590 -3595 7635 -3475
rect 7755 -3595 7800 -3475
rect 7920 -3595 7975 -3475
rect 8095 -3595 8140 -3475
rect 8260 -3595 8305 -3475
rect 8425 -3595 8470 -3475
rect 8590 -3595 8645 -3475
rect 8765 -3595 8810 -3475
rect 8930 -3595 8975 -3475
rect 9095 -3595 9140 -3475
rect 9260 -3595 9315 -3475
rect 9435 -3595 9480 -3475
rect 9600 -3595 9645 -3475
rect 9765 -3595 9810 -3475
rect 9930 -3595 9985 -3475
rect 10105 -3595 10150 -3475
rect 10270 -3595 10315 -3475
rect 10435 -3595 10480 -3475
rect 10600 -3595 10655 -3475
rect 10775 -3595 10820 -3475
rect 10940 -3595 10985 -3475
rect 11105 -3595 11150 -3475
rect 11270 -3595 11325 -3475
rect 11445 -3595 11490 -3475
rect 11610 -3595 11655 -3475
rect 11775 -3595 11820 -3475
rect 11940 -3595 11995 -3475
rect 12115 -3595 12160 -3475
rect 12280 -3595 12325 -3475
rect 12445 -3595 12490 -3475
rect 12610 -3595 12620 -3475
rect 7120 -3640 12620 -3595
rect 7120 -3760 7130 -3640
rect 7250 -3760 7305 -3640
rect 7425 -3760 7470 -3640
rect 7590 -3760 7635 -3640
rect 7755 -3760 7800 -3640
rect 7920 -3760 7975 -3640
rect 8095 -3760 8140 -3640
rect 8260 -3760 8305 -3640
rect 8425 -3760 8470 -3640
rect 8590 -3760 8645 -3640
rect 8765 -3760 8810 -3640
rect 8930 -3760 8975 -3640
rect 9095 -3760 9140 -3640
rect 9260 -3760 9315 -3640
rect 9435 -3760 9480 -3640
rect 9600 -3760 9645 -3640
rect 9765 -3760 9810 -3640
rect 9930 -3760 9985 -3640
rect 10105 -3760 10150 -3640
rect 10270 -3760 10315 -3640
rect 10435 -3760 10480 -3640
rect 10600 -3760 10655 -3640
rect 10775 -3760 10820 -3640
rect 10940 -3760 10985 -3640
rect 11105 -3760 11150 -3640
rect 11270 -3760 11325 -3640
rect 11445 -3760 11490 -3640
rect 11610 -3760 11655 -3640
rect 11775 -3760 11820 -3640
rect 11940 -3760 11995 -3640
rect 12115 -3760 12160 -3640
rect 12280 -3760 12325 -3640
rect 12445 -3760 12490 -3640
rect 12610 -3760 12620 -3640
rect 7120 -3805 12620 -3760
rect 7120 -3925 7130 -3805
rect 7250 -3925 7305 -3805
rect 7425 -3925 7470 -3805
rect 7590 -3925 7635 -3805
rect 7755 -3925 7800 -3805
rect 7920 -3925 7975 -3805
rect 8095 -3925 8140 -3805
rect 8260 -3925 8305 -3805
rect 8425 -3925 8470 -3805
rect 8590 -3925 8645 -3805
rect 8765 -3925 8810 -3805
rect 8930 -3925 8975 -3805
rect 9095 -3925 9140 -3805
rect 9260 -3925 9315 -3805
rect 9435 -3925 9480 -3805
rect 9600 -3925 9645 -3805
rect 9765 -3925 9810 -3805
rect 9930 -3925 9985 -3805
rect 10105 -3925 10150 -3805
rect 10270 -3925 10315 -3805
rect 10435 -3925 10480 -3805
rect 10600 -3925 10655 -3805
rect 10775 -3925 10820 -3805
rect 10940 -3925 10985 -3805
rect 11105 -3925 11150 -3805
rect 11270 -3925 11325 -3805
rect 11445 -3925 11490 -3805
rect 11610 -3925 11655 -3805
rect 11775 -3925 11820 -3805
rect 11940 -3925 11995 -3805
rect 12115 -3925 12160 -3805
rect 12280 -3925 12325 -3805
rect 12445 -3925 12490 -3805
rect 12610 -3925 12620 -3805
rect 7120 -3980 12620 -3925
rect 7120 -4100 7130 -3980
rect 7250 -4100 7305 -3980
rect 7425 -4100 7470 -3980
rect 7590 -4100 7635 -3980
rect 7755 -4100 7800 -3980
rect 7920 -4100 7975 -3980
rect 8095 -4100 8140 -3980
rect 8260 -4100 8305 -3980
rect 8425 -4100 8470 -3980
rect 8590 -4100 8645 -3980
rect 8765 -4100 8810 -3980
rect 8930 -4100 8975 -3980
rect 9095 -4100 9140 -3980
rect 9260 -4100 9315 -3980
rect 9435 -4100 9480 -3980
rect 9600 -4100 9645 -3980
rect 9765 -4100 9810 -3980
rect 9930 -4100 9985 -3980
rect 10105 -4100 10150 -3980
rect 10270 -4100 10315 -3980
rect 10435 -4100 10480 -3980
rect 10600 -4100 10655 -3980
rect 10775 -4100 10820 -3980
rect 10940 -4100 10985 -3980
rect 11105 -4100 11150 -3980
rect 11270 -4100 11325 -3980
rect 11445 -4100 11490 -3980
rect 11610 -4100 11655 -3980
rect 11775 -4100 11820 -3980
rect 11940 -4100 11995 -3980
rect 12115 -4100 12160 -3980
rect 12280 -4100 12325 -3980
rect 12445 -4100 12490 -3980
rect 12610 -4100 12620 -3980
rect 7120 -4110 12620 -4100
rect 12810 1380 18310 1390
rect 12810 1260 12820 1380
rect 12940 1260 12995 1380
rect 13115 1260 13160 1380
rect 13280 1260 13325 1380
rect 13445 1260 13490 1380
rect 13610 1260 13665 1380
rect 13785 1260 13830 1380
rect 13950 1260 13995 1380
rect 14115 1260 14160 1380
rect 14280 1260 14335 1380
rect 14455 1260 14500 1380
rect 14620 1260 14665 1380
rect 14785 1260 14830 1380
rect 14950 1260 15005 1380
rect 15125 1260 15170 1380
rect 15290 1260 15335 1380
rect 15455 1260 15500 1380
rect 15620 1260 15675 1380
rect 15795 1260 15840 1380
rect 15960 1260 16005 1380
rect 16125 1260 16170 1380
rect 16290 1260 16345 1380
rect 16465 1260 16510 1380
rect 16630 1260 16675 1380
rect 16795 1260 16840 1380
rect 16960 1260 17015 1380
rect 17135 1260 17180 1380
rect 17300 1260 17345 1380
rect 17465 1260 17510 1380
rect 17630 1260 17685 1380
rect 17805 1260 17850 1380
rect 17970 1260 18015 1380
rect 18135 1260 18180 1380
rect 18300 1260 18310 1380
rect 12810 1215 18310 1260
rect 12810 1095 12820 1215
rect 12940 1095 12995 1215
rect 13115 1095 13160 1215
rect 13280 1095 13325 1215
rect 13445 1095 13490 1215
rect 13610 1095 13665 1215
rect 13785 1095 13830 1215
rect 13950 1095 13995 1215
rect 14115 1095 14160 1215
rect 14280 1095 14335 1215
rect 14455 1095 14500 1215
rect 14620 1095 14665 1215
rect 14785 1095 14830 1215
rect 14950 1095 15005 1215
rect 15125 1095 15170 1215
rect 15290 1095 15335 1215
rect 15455 1095 15500 1215
rect 15620 1095 15675 1215
rect 15795 1095 15840 1215
rect 15960 1095 16005 1215
rect 16125 1095 16170 1215
rect 16290 1095 16345 1215
rect 16465 1095 16510 1215
rect 16630 1095 16675 1215
rect 16795 1095 16840 1215
rect 16960 1095 17015 1215
rect 17135 1095 17180 1215
rect 17300 1095 17345 1215
rect 17465 1095 17510 1215
rect 17630 1095 17685 1215
rect 17805 1095 17850 1215
rect 17970 1095 18015 1215
rect 18135 1095 18180 1215
rect 18300 1095 18310 1215
rect 12810 1050 18310 1095
rect 12810 930 12820 1050
rect 12940 930 12995 1050
rect 13115 930 13160 1050
rect 13280 930 13325 1050
rect 13445 930 13490 1050
rect 13610 930 13665 1050
rect 13785 930 13830 1050
rect 13950 930 13995 1050
rect 14115 930 14160 1050
rect 14280 930 14335 1050
rect 14455 930 14500 1050
rect 14620 930 14665 1050
rect 14785 930 14830 1050
rect 14950 930 15005 1050
rect 15125 930 15170 1050
rect 15290 930 15335 1050
rect 15455 930 15500 1050
rect 15620 930 15675 1050
rect 15795 930 15840 1050
rect 15960 930 16005 1050
rect 16125 930 16170 1050
rect 16290 930 16345 1050
rect 16465 930 16510 1050
rect 16630 930 16675 1050
rect 16795 930 16840 1050
rect 16960 930 17015 1050
rect 17135 930 17180 1050
rect 17300 930 17345 1050
rect 17465 930 17510 1050
rect 17630 930 17685 1050
rect 17805 930 17850 1050
rect 17970 930 18015 1050
rect 18135 930 18180 1050
rect 18300 930 18310 1050
rect 12810 885 18310 930
rect 12810 765 12820 885
rect 12940 765 12995 885
rect 13115 765 13160 885
rect 13280 765 13325 885
rect 13445 765 13490 885
rect 13610 765 13665 885
rect 13785 765 13830 885
rect 13950 765 13995 885
rect 14115 765 14160 885
rect 14280 765 14335 885
rect 14455 765 14500 885
rect 14620 765 14665 885
rect 14785 765 14830 885
rect 14950 765 15005 885
rect 15125 765 15170 885
rect 15290 765 15335 885
rect 15455 765 15500 885
rect 15620 765 15675 885
rect 15795 765 15840 885
rect 15960 765 16005 885
rect 16125 765 16170 885
rect 16290 765 16345 885
rect 16465 765 16510 885
rect 16630 765 16675 885
rect 16795 765 16840 885
rect 16960 765 17015 885
rect 17135 765 17180 885
rect 17300 765 17345 885
rect 17465 765 17510 885
rect 17630 765 17685 885
rect 17805 765 17850 885
rect 17970 765 18015 885
rect 18135 765 18180 885
rect 18300 765 18310 885
rect 12810 710 18310 765
rect 12810 590 12820 710
rect 12940 590 12995 710
rect 13115 590 13160 710
rect 13280 590 13325 710
rect 13445 590 13490 710
rect 13610 590 13665 710
rect 13785 590 13830 710
rect 13950 590 13995 710
rect 14115 590 14160 710
rect 14280 590 14335 710
rect 14455 590 14500 710
rect 14620 590 14665 710
rect 14785 590 14830 710
rect 14950 590 15005 710
rect 15125 590 15170 710
rect 15290 590 15335 710
rect 15455 590 15500 710
rect 15620 590 15675 710
rect 15795 590 15840 710
rect 15960 590 16005 710
rect 16125 590 16170 710
rect 16290 590 16345 710
rect 16465 590 16510 710
rect 16630 590 16675 710
rect 16795 590 16840 710
rect 16960 590 17015 710
rect 17135 590 17180 710
rect 17300 590 17345 710
rect 17465 590 17510 710
rect 17630 590 17685 710
rect 17805 590 17850 710
rect 17970 590 18015 710
rect 18135 590 18180 710
rect 18300 590 18310 710
rect 12810 545 18310 590
rect 12810 425 12820 545
rect 12940 425 12995 545
rect 13115 425 13160 545
rect 13280 425 13325 545
rect 13445 425 13490 545
rect 13610 425 13665 545
rect 13785 425 13830 545
rect 13950 425 13995 545
rect 14115 425 14160 545
rect 14280 425 14335 545
rect 14455 425 14500 545
rect 14620 425 14665 545
rect 14785 425 14830 545
rect 14950 425 15005 545
rect 15125 425 15170 545
rect 15290 425 15335 545
rect 15455 425 15500 545
rect 15620 425 15675 545
rect 15795 425 15840 545
rect 15960 425 16005 545
rect 16125 425 16170 545
rect 16290 425 16345 545
rect 16465 425 16510 545
rect 16630 425 16675 545
rect 16795 425 16840 545
rect 16960 425 17015 545
rect 17135 425 17180 545
rect 17300 425 17345 545
rect 17465 425 17510 545
rect 17630 425 17685 545
rect 17805 425 17850 545
rect 17970 425 18015 545
rect 18135 425 18180 545
rect 18300 425 18310 545
rect 12810 380 18310 425
rect 12810 260 12820 380
rect 12940 260 12995 380
rect 13115 260 13160 380
rect 13280 260 13325 380
rect 13445 260 13490 380
rect 13610 260 13665 380
rect 13785 260 13830 380
rect 13950 260 13995 380
rect 14115 260 14160 380
rect 14280 260 14335 380
rect 14455 260 14500 380
rect 14620 260 14665 380
rect 14785 260 14830 380
rect 14950 260 15005 380
rect 15125 260 15170 380
rect 15290 260 15335 380
rect 15455 260 15500 380
rect 15620 260 15675 380
rect 15795 260 15840 380
rect 15960 260 16005 380
rect 16125 260 16170 380
rect 16290 260 16345 380
rect 16465 260 16510 380
rect 16630 260 16675 380
rect 16795 260 16840 380
rect 16960 260 17015 380
rect 17135 260 17180 380
rect 17300 260 17345 380
rect 17465 260 17510 380
rect 17630 260 17685 380
rect 17805 260 17850 380
rect 17970 260 18015 380
rect 18135 260 18180 380
rect 18300 260 18310 380
rect 12810 215 18310 260
rect 12810 95 12820 215
rect 12940 95 12995 215
rect 13115 95 13160 215
rect 13280 95 13325 215
rect 13445 95 13490 215
rect 13610 95 13665 215
rect 13785 95 13830 215
rect 13950 95 13995 215
rect 14115 95 14160 215
rect 14280 95 14335 215
rect 14455 95 14500 215
rect 14620 95 14665 215
rect 14785 95 14830 215
rect 14950 95 15005 215
rect 15125 95 15170 215
rect 15290 95 15335 215
rect 15455 95 15500 215
rect 15620 95 15675 215
rect 15795 95 15840 215
rect 15960 95 16005 215
rect 16125 95 16170 215
rect 16290 95 16345 215
rect 16465 95 16510 215
rect 16630 95 16675 215
rect 16795 95 16840 215
rect 16960 95 17015 215
rect 17135 95 17180 215
rect 17300 95 17345 215
rect 17465 95 17510 215
rect 17630 95 17685 215
rect 17805 95 17850 215
rect 17970 95 18015 215
rect 18135 95 18180 215
rect 18300 95 18310 215
rect 12810 40 18310 95
rect 12810 -80 12820 40
rect 12940 -80 12995 40
rect 13115 -80 13160 40
rect 13280 -80 13325 40
rect 13445 -80 13490 40
rect 13610 -80 13665 40
rect 13785 -80 13830 40
rect 13950 -80 13995 40
rect 14115 -80 14160 40
rect 14280 -80 14335 40
rect 14455 -80 14500 40
rect 14620 -80 14665 40
rect 14785 -80 14830 40
rect 14950 -80 15005 40
rect 15125 -80 15170 40
rect 15290 -80 15335 40
rect 15455 -80 15500 40
rect 15620 -80 15675 40
rect 15795 -80 15840 40
rect 15960 -80 16005 40
rect 16125 -80 16170 40
rect 16290 -80 16345 40
rect 16465 -80 16510 40
rect 16630 -80 16675 40
rect 16795 -80 16840 40
rect 16960 -80 17015 40
rect 17135 -80 17180 40
rect 17300 -80 17345 40
rect 17465 -80 17510 40
rect 17630 -80 17685 40
rect 17805 -80 17850 40
rect 17970 -80 18015 40
rect 18135 -80 18180 40
rect 18300 -80 18310 40
rect 12810 -125 18310 -80
rect 12810 -245 12820 -125
rect 12940 -245 12995 -125
rect 13115 -245 13160 -125
rect 13280 -245 13325 -125
rect 13445 -245 13490 -125
rect 13610 -245 13665 -125
rect 13785 -245 13830 -125
rect 13950 -245 13995 -125
rect 14115 -245 14160 -125
rect 14280 -245 14335 -125
rect 14455 -245 14500 -125
rect 14620 -245 14665 -125
rect 14785 -245 14830 -125
rect 14950 -245 15005 -125
rect 15125 -245 15170 -125
rect 15290 -245 15335 -125
rect 15455 -245 15500 -125
rect 15620 -245 15675 -125
rect 15795 -245 15840 -125
rect 15960 -245 16005 -125
rect 16125 -245 16170 -125
rect 16290 -245 16345 -125
rect 16465 -245 16510 -125
rect 16630 -245 16675 -125
rect 16795 -245 16840 -125
rect 16960 -245 17015 -125
rect 17135 -245 17180 -125
rect 17300 -245 17345 -125
rect 17465 -245 17510 -125
rect 17630 -245 17685 -125
rect 17805 -245 17850 -125
rect 17970 -245 18015 -125
rect 18135 -245 18180 -125
rect 18300 -245 18310 -125
rect 12810 -290 18310 -245
rect 12810 -410 12820 -290
rect 12940 -410 12995 -290
rect 13115 -410 13160 -290
rect 13280 -410 13325 -290
rect 13445 -410 13490 -290
rect 13610 -410 13665 -290
rect 13785 -410 13830 -290
rect 13950 -410 13995 -290
rect 14115 -410 14160 -290
rect 14280 -410 14335 -290
rect 14455 -410 14500 -290
rect 14620 -410 14665 -290
rect 14785 -410 14830 -290
rect 14950 -410 15005 -290
rect 15125 -410 15170 -290
rect 15290 -410 15335 -290
rect 15455 -410 15500 -290
rect 15620 -410 15675 -290
rect 15795 -410 15840 -290
rect 15960 -410 16005 -290
rect 16125 -410 16170 -290
rect 16290 -410 16345 -290
rect 16465 -410 16510 -290
rect 16630 -410 16675 -290
rect 16795 -410 16840 -290
rect 16960 -410 17015 -290
rect 17135 -410 17180 -290
rect 17300 -410 17345 -290
rect 17465 -410 17510 -290
rect 17630 -410 17685 -290
rect 17805 -410 17850 -290
rect 17970 -410 18015 -290
rect 18135 -410 18180 -290
rect 18300 -410 18310 -290
rect 12810 -455 18310 -410
rect 12810 -575 12820 -455
rect 12940 -575 12995 -455
rect 13115 -575 13160 -455
rect 13280 -575 13325 -455
rect 13445 -575 13490 -455
rect 13610 -575 13665 -455
rect 13785 -575 13830 -455
rect 13950 -575 13995 -455
rect 14115 -575 14160 -455
rect 14280 -575 14335 -455
rect 14455 -575 14500 -455
rect 14620 -575 14665 -455
rect 14785 -575 14830 -455
rect 14950 -575 15005 -455
rect 15125 -575 15170 -455
rect 15290 -575 15335 -455
rect 15455 -575 15500 -455
rect 15620 -575 15675 -455
rect 15795 -575 15840 -455
rect 15960 -575 16005 -455
rect 16125 -575 16170 -455
rect 16290 -575 16345 -455
rect 16465 -575 16510 -455
rect 16630 -575 16675 -455
rect 16795 -575 16840 -455
rect 16960 -575 17015 -455
rect 17135 -575 17180 -455
rect 17300 -575 17345 -455
rect 17465 -575 17510 -455
rect 17630 -575 17685 -455
rect 17805 -575 17850 -455
rect 17970 -575 18015 -455
rect 18135 -575 18180 -455
rect 18300 -575 18310 -455
rect 12810 -630 18310 -575
rect 12810 -750 12820 -630
rect 12940 -750 12995 -630
rect 13115 -750 13160 -630
rect 13280 -750 13325 -630
rect 13445 -750 13490 -630
rect 13610 -750 13665 -630
rect 13785 -750 13830 -630
rect 13950 -750 13995 -630
rect 14115 -750 14160 -630
rect 14280 -750 14335 -630
rect 14455 -750 14500 -630
rect 14620 -750 14665 -630
rect 14785 -750 14830 -630
rect 14950 -750 15005 -630
rect 15125 -750 15170 -630
rect 15290 -750 15335 -630
rect 15455 -750 15500 -630
rect 15620 -750 15675 -630
rect 15795 -750 15840 -630
rect 15960 -750 16005 -630
rect 16125 -750 16170 -630
rect 16290 -750 16345 -630
rect 16465 -750 16510 -630
rect 16630 -750 16675 -630
rect 16795 -750 16840 -630
rect 16960 -750 17015 -630
rect 17135 -750 17180 -630
rect 17300 -750 17345 -630
rect 17465 -750 17510 -630
rect 17630 -750 17685 -630
rect 17805 -750 17850 -630
rect 17970 -750 18015 -630
rect 18135 -750 18180 -630
rect 18300 -750 18310 -630
rect 12810 -795 18310 -750
rect 12810 -915 12820 -795
rect 12940 -915 12995 -795
rect 13115 -915 13160 -795
rect 13280 -915 13325 -795
rect 13445 -915 13490 -795
rect 13610 -915 13665 -795
rect 13785 -915 13830 -795
rect 13950 -915 13995 -795
rect 14115 -915 14160 -795
rect 14280 -915 14335 -795
rect 14455 -915 14500 -795
rect 14620 -915 14665 -795
rect 14785 -915 14830 -795
rect 14950 -915 15005 -795
rect 15125 -915 15170 -795
rect 15290 -915 15335 -795
rect 15455 -915 15500 -795
rect 15620 -915 15675 -795
rect 15795 -915 15840 -795
rect 15960 -915 16005 -795
rect 16125 -915 16170 -795
rect 16290 -915 16345 -795
rect 16465 -915 16510 -795
rect 16630 -915 16675 -795
rect 16795 -915 16840 -795
rect 16960 -915 17015 -795
rect 17135 -915 17180 -795
rect 17300 -915 17345 -795
rect 17465 -915 17510 -795
rect 17630 -915 17685 -795
rect 17805 -915 17850 -795
rect 17970 -915 18015 -795
rect 18135 -915 18180 -795
rect 18300 -915 18310 -795
rect 12810 -960 18310 -915
rect 12810 -1080 12820 -960
rect 12940 -1080 12995 -960
rect 13115 -1080 13160 -960
rect 13280 -1080 13325 -960
rect 13445 -1080 13490 -960
rect 13610 -1080 13665 -960
rect 13785 -1080 13830 -960
rect 13950 -1080 13995 -960
rect 14115 -1080 14160 -960
rect 14280 -1080 14335 -960
rect 14455 -1080 14500 -960
rect 14620 -1080 14665 -960
rect 14785 -1080 14830 -960
rect 14950 -1080 15005 -960
rect 15125 -1080 15170 -960
rect 15290 -1080 15335 -960
rect 15455 -1080 15500 -960
rect 15620 -1080 15675 -960
rect 15795 -1080 15840 -960
rect 15960 -1080 16005 -960
rect 16125 -1080 16170 -960
rect 16290 -1080 16345 -960
rect 16465 -1080 16510 -960
rect 16630 -1080 16675 -960
rect 16795 -1080 16840 -960
rect 16960 -1080 17015 -960
rect 17135 -1080 17180 -960
rect 17300 -1080 17345 -960
rect 17465 -1080 17510 -960
rect 17630 -1080 17685 -960
rect 17805 -1080 17850 -960
rect 17970 -1080 18015 -960
rect 18135 -1080 18180 -960
rect 18300 -1080 18310 -960
rect 12810 -1125 18310 -1080
rect 12810 -1245 12820 -1125
rect 12940 -1245 12995 -1125
rect 13115 -1245 13160 -1125
rect 13280 -1245 13325 -1125
rect 13445 -1245 13490 -1125
rect 13610 -1245 13665 -1125
rect 13785 -1245 13830 -1125
rect 13950 -1245 13995 -1125
rect 14115 -1245 14160 -1125
rect 14280 -1245 14335 -1125
rect 14455 -1245 14500 -1125
rect 14620 -1245 14665 -1125
rect 14785 -1245 14830 -1125
rect 14950 -1245 15005 -1125
rect 15125 -1245 15170 -1125
rect 15290 -1245 15335 -1125
rect 15455 -1245 15500 -1125
rect 15620 -1245 15675 -1125
rect 15795 -1245 15840 -1125
rect 15960 -1245 16005 -1125
rect 16125 -1245 16170 -1125
rect 16290 -1245 16345 -1125
rect 16465 -1245 16510 -1125
rect 16630 -1245 16675 -1125
rect 16795 -1245 16840 -1125
rect 16960 -1245 17015 -1125
rect 17135 -1245 17180 -1125
rect 17300 -1245 17345 -1125
rect 17465 -1245 17510 -1125
rect 17630 -1245 17685 -1125
rect 17805 -1245 17850 -1125
rect 17970 -1245 18015 -1125
rect 18135 -1245 18180 -1125
rect 18300 -1245 18310 -1125
rect 12810 -1300 18310 -1245
rect 12810 -1420 12820 -1300
rect 12940 -1420 12995 -1300
rect 13115 -1420 13160 -1300
rect 13280 -1420 13325 -1300
rect 13445 -1420 13490 -1300
rect 13610 -1420 13665 -1300
rect 13785 -1420 13830 -1300
rect 13950 -1420 13995 -1300
rect 14115 -1420 14160 -1300
rect 14280 -1420 14335 -1300
rect 14455 -1420 14500 -1300
rect 14620 -1420 14665 -1300
rect 14785 -1420 14830 -1300
rect 14950 -1420 15005 -1300
rect 15125 -1420 15170 -1300
rect 15290 -1420 15335 -1300
rect 15455 -1420 15500 -1300
rect 15620 -1420 15675 -1300
rect 15795 -1420 15840 -1300
rect 15960 -1420 16005 -1300
rect 16125 -1420 16170 -1300
rect 16290 -1420 16345 -1300
rect 16465 -1420 16510 -1300
rect 16630 -1420 16675 -1300
rect 16795 -1420 16840 -1300
rect 16960 -1420 17015 -1300
rect 17135 -1420 17180 -1300
rect 17300 -1420 17345 -1300
rect 17465 -1420 17510 -1300
rect 17630 -1420 17685 -1300
rect 17805 -1420 17850 -1300
rect 17970 -1420 18015 -1300
rect 18135 -1420 18180 -1300
rect 18300 -1420 18310 -1300
rect 12810 -1465 18310 -1420
rect 12810 -1585 12820 -1465
rect 12940 -1585 12995 -1465
rect 13115 -1585 13160 -1465
rect 13280 -1585 13325 -1465
rect 13445 -1585 13490 -1465
rect 13610 -1585 13665 -1465
rect 13785 -1585 13830 -1465
rect 13950 -1585 13995 -1465
rect 14115 -1585 14160 -1465
rect 14280 -1585 14335 -1465
rect 14455 -1585 14500 -1465
rect 14620 -1585 14665 -1465
rect 14785 -1585 14830 -1465
rect 14950 -1585 15005 -1465
rect 15125 -1585 15170 -1465
rect 15290 -1585 15335 -1465
rect 15455 -1585 15500 -1465
rect 15620 -1585 15675 -1465
rect 15795 -1585 15840 -1465
rect 15960 -1585 16005 -1465
rect 16125 -1585 16170 -1465
rect 16290 -1585 16345 -1465
rect 16465 -1585 16510 -1465
rect 16630 -1585 16675 -1465
rect 16795 -1585 16840 -1465
rect 16960 -1585 17015 -1465
rect 17135 -1585 17180 -1465
rect 17300 -1585 17345 -1465
rect 17465 -1585 17510 -1465
rect 17630 -1585 17685 -1465
rect 17805 -1585 17850 -1465
rect 17970 -1585 18015 -1465
rect 18135 -1585 18180 -1465
rect 18300 -1585 18310 -1465
rect 12810 -1630 18310 -1585
rect 12810 -1750 12820 -1630
rect 12940 -1750 12995 -1630
rect 13115 -1750 13160 -1630
rect 13280 -1750 13325 -1630
rect 13445 -1750 13490 -1630
rect 13610 -1750 13665 -1630
rect 13785 -1750 13830 -1630
rect 13950 -1750 13995 -1630
rect 14115 -1750 14160 -1630
rect 14280 -1750 14335 -1630
rect 14455 -1750 14500 -1630
rect 14620 -1750 14665 -1630
rect 14785 -1750 14830 -1630
rect 14950 -1750 15005 -1630
rect 15125 -1750 15170 -1630
rect 15290 -1750 15335 -1630
rect 15455 -1750 15500 -1630
rect 15620 -1750 15675 -1630
rect 15795 -1750 15840 -1630
rect 15960 -1750 16005 -1630
rect 16125 -1750 16170 -1630
rect 16290 -1750 16345 -1630
rect 16465 -1750 16510 -1630
rect 16630 -1750 16675 -1630
rect 16795 -1750 16840 -1630
rect 16960 -1750 17015 -1630
rect 17135 -1750 17180 -1630
rect 17300 -1750 17345 -1630
rect 17465 -1750 17510 -1630
rect 17630 -1750 17685 -1630
rect 17805 -1750 17850 -1630
rect 17970 -1750 18015 -1630
rect 18135 -1750 18180 -1630
rect 18300 -1750 18310 -1630
rect 12810 -1795 18310 -1750
rect 12810 -1915 12820 -1795
rect 12940 -1915 12995 -1795
rect 13115 -1915 13160 -1795
rect 13280 -1915 13325 -1795
rect 13445 -1915 13490 -1795
rect 13610 -1915 13665 -1795
rect 13785 -1915 13830 -1795
rect 13950 -1915 13995 -1795
rect 14115 -1915 14160 -1795
rect 14280 -1915 14335 -1795
rect 14455 -1915 14500 -1795
rect 14620 -1915 14665 -1795
rect 14785 -1915 14830 -1795
rect 14950 -1915 15005 -1795
rect 15125 -1915 15170 -1795
rect 15290 -1915 15335 -1795
rect 15455 -1915 15500 -1795
rect 15620 -1915 15675 -1795
rect 15795 -1915 15840 -1795
rect 15960 -1915 16005 -1795
rect 16125 -1915 16170 -1795
rect 16290 -1915 16345 -1795
rect 16465 -1915 16510 -1795
rect 16630 -1915 16675 -1795
rect 16795 -1915 16840 -1795
rect 16960 -1915 17015 -1795
rect 17135 -1915 17180 -1795
rect 17300 -1915 17345 -1795
rect 17465 -1915 17510 -1795
rect 17630 -1915 17685 -1795
rect 17805 -1915 17850 -1795
rect 17970 -1915 18015 -1795
rect 18135 -1915 18180 -1795
rect 18300 -1915 18310 -1795
rect 12810 -1970 18310 -1915
rect 12810 -2090 12820 -1970
rect 12940 -2090 12995 -1970
rect 13115 -2090 13160 -1970
rect 13280 -2090 13325 -1970
rect 13445 -2090 13490 -1970
rect 13610 -2090 13665 -1970
rect 13785 -2090 13830 -1970
rect 13950 -2090 13995 -1970
rect 14115 -2090 14160 -1970
rect 14280 -2090 14335 -1970
rect 14455 -2090 14500 -1970
rect 14620 -2090 14665 -1970
rect 14785 -2090 14830 -1970
rect 14950 -2090 15005 -1970
rect 15125 -2090 15170 -1970
rect 15290 -2090 15335 -1970
rect 15455 -2090 15500 -1970
rect 15620 -2090 15675 -1970
rect 15795 -2090 15840 -1970
rect 15960 -2090 16005 -1970
rect 16125 -2090 16170 -1970
rect 16290 -2090 16345 -1970
rect 16465 -2090 16510 -1970
rect 16630 -2090 16675 -1970
rect 16795 -2090 16840 -1970
rect 16960 -2090 17015 -1970
rect 17135 -2090 17180 -1970
rect 17300 -2090 17345 -1970
rect 17465 -2090 17510 -1970
rect 17630 -2090 17685 -1970
rect 17805 -2090 17850 -1970
rect 17970 -2090 18015 -1970
rect 18135 -2090 18180 -1970
rect 18300 -2090 18310 -1970
rect 12810 -2135 18310 -2090
rect 12810 -2255 12820 -2135
rect 12940 -2255 12995 -2135
rect 13115 -2255 13160 -2135
rect 13280 -2255 13325 -2135
rect 13445 -2255 13490 -2135
rect 13610 -2255 13665 -2135
rect 13785 -2255 13830 -2135
rect 13950 -2255 13995 -2135
rect 14115 -2255 14160 -2135
rect 14280 -2255 14335 -2135
rect 14455 -2255 14500 -2135
rect 14620 -2255 14665 -2135
rect 14785 -2255 14830 -2135
rect 14950 -2255 15005 -2135
rect 15125 -2255 15170 -2135
rect 15290 -2255 15335 -2135
rect 15455 -2255 15500 -2135
rect 15620 -2255 15675 -2135
rect 15795 -2255 15840 -2135
rect 15960 -2255 16005 -2135
rect 16125 -2255 16170 -2135
rect 16290 -2255 16345 -2135
rect 16465 -2255 16510 -2135
rect 16630 -2255 16675 -2135
rect 16795 -2255 16840 -2135
rect 16960 -2255 17015 -2135
rect 17135 -2255 17180 -2135
rect 17300 -2255 17345 -2135
rect 17465 -2255 17510 -2135
rect 17630 -2255 17685 -2135
rect 17805 -2255 17850 -2135
rect 17970 -2255 18015 -2135
rect 18135 -2255 18180 -2135
rect 18300 -2255 18310 -2135
rect 12810 -2300 18310 -2255
rect 12810 -2420 12820 -2300
rect 12940 -2420 12995 -2300
rect 13115 -2420 13160 -2300
rect 13280 -2420 13325 -2300
rect 13445 -2420 13490 -2300
rect 13610 -2420 13665 -2300
rect 13785 -2420 13830 -2300
rect 13950 -2420 13995 -2300
rect 14115 -2420 14160 -2300
rect 14280 -2420 14335 -2300
rect 14455 -2420 14500 -2300
rect 14620 -2420 14665 -2300
rect 14785 -2420 14830 -2300
rect 14950 -2420 15005 -2300
rect 15125 -2420 15170 -2300
rect 15290 -2420 15335 -2300
rect 15455 -2420 15500 -2300
rect 15620 -2420 15675 -2300
rect 15795 -2420 15840 -2300
rect 15960 -2420 16005 -2300
rect 16125 -2420 16170 -2300
rect 16290 -2420 16345 -2300
rect 16465 -2420 16510 -2300
rect 16630 -2420 16675 -2300
rect 16795 -2420 16840 -2300
rect 16960 -2420 17015 -2300
rect 17135 -2420 17180 -2300
rect 17300 -2420 17345 -2300
rect 17465 -2420 17510 -2300
rect 17630 -2420 17685 -2300
rect 17805 -2420 17850 -2300
rect 17970 -2420 18015 -2300
rect 18135 -2420 18180 -2300
rect 18300 -2420 18310 -2300
rect 12810 -2465 18310 -2420
rect 12810 -2585 12820 -2465
rect 12940 -2585 12995 -2465
rect 13115 -2585 13160 -2465
rect 13280 -2585 13325 -2465
rect 13445 -2585 13490 -2465
rect 13610 -2585 13665 -2465
rect 13785 -2585 13830 -2465
rect 13950 -2585 13995 -2465
rect 14115 -2585 14160 -2465
rect 14280 -2585 14335 -2465
rect 14455 -2585 14500 -2465
rect 14620 -2585 14665 -2465
rect 14785 -2585 14830 -2465
rect 14950 -2585 15005 -2465
rect 15125 -2585 15170 -2465
rect 15290 -2585 15335 -2465
rect 15455 -2585 15500 -2465
rect 15620 -2585 15675 -2465
rect 15795 -2585 15840 -2465
rect 15960 -2585 16005 -2465
rect 16125 -2585 16170 -2465
rect 16290 -2585 16345 -2465
rect 16465 -2585 16510 -2465
rect 16630 -2585 16675 -2465
rect 16795 -2585 16840 -2465
rect 16960 -2585 17015 -2465
rect 17135 -2585 17180 -2465
rect 17300 -2585 17345 -2465
rect 17465 -2585 17510 -2465
rect 17630 -2585 17685 -2465
rect 17805 -2585 17850 -2465
rect 17970 -2585 18015 -2465
rect 18135 -2585 18180 -2465
rect 18300 -2585 18310 -2465
rect 12810 -2640 18310 -2585
rect 12810 -2760 12820 -2640
rect 12940 -2760 12995 -2640
rect 13115 -2760 13160 -2640
rect 13280 -2760 13325 -2640
rect 13445 -2760 13490 -2640
rect 13610 -2760 13665 -2640
rect 13785 -2760 13830 -2640
rect 13950 -2760 13995 -2640
rect 14115 -2760 14160 -2640
rect 14280 -2760 14335 -2640
rect 14455 -2760 14500 -2640
rect 14620 -2760 14665 -2640
rect 14785 -2760 14830 -2640
rect 14950 -2760 15005 -2640
rect 15125 -2760 15170 -2640
rect 15290 -2760 15335 -2640
rect 15455 -2760 15500 -2640
rect 15620 -2760 15675 -2640
rect 15795 -2760 15840 -2640
rect 15960 -2760 16005 -2640
rect 16125 -2760 16170 -2640
rect 16290 -2760 16345 -2640
rect 16465 -2760 16510 -2640
rect 16630 -2760 16675 -2640
rect 16795 -2760 16840 -2640
rect 16960 -2760 17015 -2640
rect 17135 -2760 17180 -2640
rect 17300 -2760 17345 -2640
rect 17465 -2760 17510 -2640
rect 17630 -2760 17685 -2640
rect 17805 -2760 17850 -2640
rect 17970 -2760 18015 -2640
rect 18135 -2760 18180 -2640
rect 18300 -2760 18310 -2640
rect 12810 -2805 18310 -2760
rect 12810 -2925 12820 -2805
rect 12940 -2925 12995 -2805
rect 13115 -2925 13160 -2805
rect 13280 -2925 13325 -2805
rect 13445 -2925 13490 -2805
rect 13610 -2925 13665 -2805
rect 13785 -2925 13830 -2805
rect 13950 -2925 13995 -2805
rect 14115 -2925 14160 -2805
rect 14280 -2925 14335 -2805
rect 14455 -2925 14500 -2805
rect 14620 -2925 14665 -2805
rect 14785 -2925 14830 -2805
rect 14950 -2925 15005 -2805
rect 15125 -2925 15170 -2805
rect 15290 -2925 15335 -2805
rect 15455 -2925 15500 -2805
rect 15620 -2925 15675 -2805
rect 15795 -2925 15840 -2805
rect 15960 -2925 16005 -2805
rect 16125 -2925 16170 -2805
rect 16290 -2925 16345 -2805
rect 16465 -2925 16510 -2805
rect 16630 -2925 16675 -2805
rect 16795 -2925 16840 -2805
rect 16960 -2925 17015 -2805
rect 17135 -2925 17180 -2805
rect 17300 -2925 17345 -2805
rect 17465 -2925 17510 -2805
rect 17630 -2925 17685 -2805
rect 17805 -2925 17850 -2805
rect 17970 -2925 18015 -2805
rect 18135 -2925 18180 -2805
rect 18300 -2925 18310 -2805
rect 12810 -2970 18310 -2925
rect 12810 -3090 12820 -2970
rect 12940 -3090 12995 -2970
rect 13115 -3090 13160 -2970
rect 13280 -3090 13325 -2970
rect 13445 -3090 13490 -2970
rect 13610 -3090 13665 -2970
rect 13785 -3090 13830 -2970
rect 13950 -3090 13995 -2970
rect 14115 -3090 14160 -2970
rect 14280 -3090 14335 -2970
rect 14455 -3090 14500 -2970
rect 14620 -3090 14665 -2970
rect 14785 -3090 14830 -2970
rect 14950 -3090 15005 -2970
rect 15125 -3090 15170 -2970
rect 15290 -3090 15335 -2970
rect 15455 -3090 15500 -2970
rect 15620 -3090 15675 -2970
rect 15795 -3090 15840 -2970
rect 15960 -3090 16005 -2970
rect 16125 -3090 16170 -2970
rect 16290 -3090 16345 -2970
rect 16465 -3090 16510 -2970
rect 16630 -3090 16675 -2970
rect 16795 -3090 16840 -2970
rect 16960 -3090 17015 -2970
rect 17135 -3090 17180 -2970
rect 17300 -3090 17345 -2970
rect 17465 -3090 17510 -2970
rect 17630 -3090 17685 -2970
rect 17805 -3090 17850 -2970
rect 17970 -3090 18015 -2970
rect 18135 -3090 18180 -2970
rect 18300 -3090 18310 -2970
rect 12810 -3135 18310 -3090
rect 12810 -3255 12820 -3135
rect 12940 -3255 12995 -3135
rect 13115 -3255 13160 -3135
rect 13280 -3255 13325 -3135
rect 13445 -3255 13490 -3135
rect 13610 -3255 13665 -3135
rect 13785 -3255 13830 -3135
rect 13950 -3255 13995 -3135
rect 14115 -3255 14160 -3135
rect 14280 -3255 14335 -3135
rect 14455 -3255 14500 -3135
rect 14620 -3255 14665 -3135
rect 14785 -3255 14830 -3135
rect 14950 -3255 15005 -3135
rect 15125 -3255 15170 -3135
rect 15290 -3255 15335 -3135
rect 15455 -3255 15500 -3135
rect 15620 -3255 15675 -3135
rect 15795 -3255 15840 -3135
rect 15960 -3255 16005 -3135
rect 16125 -3255 16170 -3135
rect 16290 -3255 16345 -3135
rect 16465 -3255 16510 -3135
rect 16630 -3255 16675 -3135
rect 16795 -3255 16840 -3135
rect 16960 -3255 17015 -3135
rect 17135 -3255 17180 -3135
rect 17300 -3255 17345 -3135
rect 17465 -3255 17510 -3135
rect 17630 -3255 17685 -3135
rect 17805 -3255 17850 -3135
rect 17970 -3255 18015 -3135
rect 18135 -3255 18180 -3135
rect 18300 -3255 18310 -3135
rect 12810 -3310 18310 -3255
rect 12810 -3430 12820 -3310
rect 12940 -3430 12995 -3310
rect 13115 -3430 13160 -3310
rect 13280 -3430 13325 -3310
rect 13445 -3430 13490 -3310
rect 13610 -3430 13665 -3310
rect 13785 -3430 13830 -3310
rect 13950 -3430 13995 -3310
rect 14115 -3430 14160 -3310
rect 14280 -3430 14335 -3310
rect 14455 -3430 14500 -3310
rect 14620 -3430 14665 -3310
rect 14785 -3430 14830 -3310
rect 14950 -3430 15005 -3310
rect 15125 -3430 15170 -3310
rect 15290 -3430 15335 -3310
rect 15455 -3430 15500 -3310
rect 15620 -3430 15675 -3310
rect 15795 -3430 15840 -3310
rect 15960 -3430 16005 -3310
rect 16125 -3430 16170 -3310
rect 16290 -3430 16345 -3310
rect 16465 -3430 16510 -3310
rect 16630 -3430 16675 -3310
rect 16795 -3430 16840 -3310
rect 16960 -3430 17015 -3310
rect 17135 -3430 17180 -3310
rect 17300 -3430 17345 -3310
rect 17465 -3430 17510 -3310
rect 17630 -3430 17685 -3310
rect 17805 -3430 17850 -3310
rect 17970 -3430 18015 -3310
rect 18135 -3430 18180 -3310
rect 18300 -3430 18310 -3310
rect 12810 -3475 18310 -3430
rect 12810 -3595 12820 -3475
rect 12940 -3595 12995 -3475
rect 13115 -3595 13160 -3475
rect 13280 -3595 13325 -3475
rect 13445 -3595 13490 -3475
rect 13610 -3595 13665 -3475
rect 13785 -3595 13830 -3475
rect 13950 -3595 13995 -3475
rect 14115 -3595 14160 -3475
rect 14280 -3595 14335 -3475
rect 14455 -3595 14500 -3475
rect 14620 -3595 14665 -3475
rect 14785 -3595 14830 -3475
rect 14950 -3595 15005 -3475
rect 15125 -3595 15170 -3475
rect 15290 -3595 15335 -3475
rect 15455 -3595 15500 -3475
rect 15620 -3595 15675 -3475
rect 15795 -3595 15840 -3475
rect 15960 -3595 16005 -3475
rect 16125 -3595 16170 -3475
rect 16290 -3595 16345 -3475
rect 16465 -3595 16510 -3475
rect 16630 -3595 16675 -3475
rect 16795 -3595 16840 -3475
rect 16960 -3595 17015 -3475
rect 17135 -3595 17180 -3475
rect 17300 -3595 17345 -3475
rect 17465 -3595 17510 -3475
rect 17630 -3595 17685 -3475
rect 17805 -3595 17850 -3475
rect 17970 -3595 18015 -3475
rect 18135 -3595 18180 -3475
rect 18300 -3595 18310 -3475
rect 12810 -3640 18310 -3595
rect 12810 -3760 12820 -3640
rect 12940 -3760 12995 -3640
rect 13115 -3760 13160 -3640
rect 13280 -3760 13325 -3640
rect 13445 -3760 13490 -3640
rect 13610 -3760 13665 -3640
rect 13785 -3760 13830 -3640
rect 13950 -3760 13995 -3640
rect 14115 -3760 14160 -3640
rect 14280 -3760 14335 -3640
rect 14455 -3760 14500 -3640
rect 14620 -3760 14665 -3640
rect 14785 -3760 14830 -3640
rect 14950 -3760 15005 -3640
rect 15125 -3760 15170 -3640
rect 15290 -3760 15335 -3640
rect 15455 -3760 15500 -3640
rect 15620 -3760 15675 -3640
rect 15795 -3760 15840 -3640
rect 15960 -3760 16005 -3640
rect 16125 -3760 16170 -3640
rect 16290 -3760 16345 -3640
rect 16465 -3760 16510 -3640
rect 16630 -3760 16675 -3640
rect 16795 -3760 16840 -3640
rect 16960 -3760 17015 -3640
rect 17135 -3760 17180 -3640
rect 17300 -3760 17345 -3640
rect 17465 -3760 17510 -3640
rect 17630 -3760 17685 -3640
rect 17805 -3760 17850 -3640
rect 17970 -3760 18015 -3640
rect 18135 -3760 18180 -3640
rect 18300 -3760 18310 -3640
rect 12810 -3805 18310 -3760
rect 12810 -3925 12820 -3805
rect 12940 -3925 12995 -3805
rect 13115 -3925 13160 -3805
rect 13280 -3925 13325 -3805
rect 13445 -3925 13490 -3805
rect 13610 -3925 13665 -3805
rect 13785 -3925 13830 -3805
rect 13950 -3925 13995 -3805
rect 14115 -3925 14160 -3805
rect 14280 -3925 14335 -3805
rect 14455 -3925 14500 -3805
rect 14620 -3925 14665 -3805
rect 14785 -3925 14830 -3805
rect 14950 -3925 15005 -3805
rect 15125 -3925 15170 -3805
rect 15290 -3925 15335 -3805
rect 15455 -3925 15500 -3805
rect 15620 -3925 15675 -3805
rect 15795 -3925 15840 -3805
rect 15960 -3925 16005 -3805
rect 16125 -3925 16170 -3805
rect 16290 -3925 16345 -3805
rect 16465 -3925 16510 -3805
rect 16630 -3925 16675 -3805
rect 16795 -3925 16840 -3805
rect 16960 -3925 17015 -3805
rect 17135 -3925 17180 -3805
rect 17300 -3925 17345 -3805
rect 17465 -3925 17510 -3805
rect 17630 -3925 17685 -3805
rect 17805 -3925 17850 -3805
rect 17970 -3925 18015 -3805
rect 18135 -3925 18180 -3805
rect 18300 -3925 18310 -3805
rect 12810 -3980 18310 -3925
rect 12810 -4100 12820 -3980
rect 12940 -4100 12995 -3980
rect 13115 -4100 13160 -3980
rect 13280 -4100 13325 -3980
rect 13445 -4100 13490 -3980
rect 13610 -4100 13665 -3980
rect 13785 -4100 13830 -3980
rect 13950 -4100 13995 -3980
rect 14115 -4100 14160 -3980
rect 14280 -4100 14335 -3980
rect 14455 -4100 14500 -3980
rect 14620 -4100 14665 -3980
rect 14785 -4100 14830 -3980
rect 14950 -4100 15005 -3980
rect 15125 -4100 15170 -3980
rect 15290 -4100 15335 -3980
rect 15455 -4100 15500 -3980
rect 15620 -4100 15675 -3980
rect 15795 -4100 15840 -3980
rect 15960 -4100 16005 -3980
rect 16125 -4100 16170 -3980
rect 16290 -4100 16345 -3980
rect 16465 -4100 16510 -3980
rect 16630 -4100 16675 -3980
rect 16795 -4100 16840 -3980
rect 16960 -4100 17015 -3980
rect 17135 -4100 17180 -3980
rect 17300 -4100 17345 -3980
rect 17465 -4100 17510 -3980
rect 17630 -4100 17685 -3980
rect 17805 -4100 17850 -3980
rect 17970 -4100 18015 -3980
rect 18135 -4100 18180 -3980
rect 18300 -4100 18310 -3980
rect 12810 -4110 18310 -4100
rect 18500 1380 24000 1390
rect 18500 1260 18510 1380
rect 18630 1260 18685 1380
rect 18805 1260 18850 1380
rect 18970 1260 19015 1380
rect 19135 1260 19180 1380
rect 19300 1260 19355 1380
rect 19475 1260 19520 1380
rect 19640 1260 19685 1380
rect 19805 1260 19850 1380
rect 19970 1260 20025 1380
rect 20145 1260 20190 1380
rect 20310 1260 20355 1380
rect 20475 1260 20520 1380
rect 20640 1260 20695 1380
rect 20815 1260 20860 1380
rect 20980 1260 21025 1380
rect 21145 1260 21190 1380
rect 21310 1260 21365 1380
rect 21485 1260 21530 1380
rect 21650 1260 21695 1380
rect 21815 1260 21860 1380
rect 21980 1260 22035 1380
rect 22155 1260 22200 1380
rect 22320 1260 22365 1380
rect 22485 1260 22530 1380
rect 22650 1260 22705 1380
rect 22825 1260 22870 1380
rect 22990 1260 23035 1380
rect 23155 1260 23200 1380
rect 23320 1260 23375 1380
rect 23495 1260 23540 1380
rect 23660 1260 23705 1380
rect 23825 1260 23870 1380
rect 23990 1260 24000 1380
rect 18500 1215 24000 1260
rect 18500 1095 18510 1215
rect 18630 1095 18685 1215
rect 18805 1095 18850 1215
rect 18970 1095 19015 1215
rect 19135 1095 19180 1215
rect 19300 1095 19355 1215
rect 19475 1095 19520 1215
rect 19640 1095 19685 1215
rect 19805 1095 19850 1215
rect 19970 1095 20025 1215
rect 20145 1095 20190 1215
rect 20310 1095 20355 1215
rect 20475 1095 20520 1215
rect 20640 1095 20695 1215
rect 20815 1095 20860 1215
rect 20980 1095 21025 1215
rect 21145 1095 21190 1215
rect 21310 1095 21365 1215
rect 21485 1095 21530 1215
rect 21650 1095 21695 1215
rect 21815 1095 21860 1215
rect 21980 1095 22035 1215
rect 22155 1095 22200 1215
rect 22320 1095 22365 1215
rect 22485 1095 22530 1215
rect 22650 1095 22705 1215
rect 22825 1095 22870 1215
rect 22990 1095 23035 1215
rect 23155 1095 23200 1215
rect 23320 1095 23375 1215
rect 23495 1095 23540 1215
rect 23660 1095 23705 1215
rect 23825 1095 23870 1215
rect 23990 1095 24000 1215
rect 18500 1050 24000 1095
rect 18500 930 18510 1050
rect 18630 930 18685 1050
rect 18805 930 18850 1050
rect 18970 930 19015 1050
rect 19135 930 19180 1050
rect 19300 930 19355 1050
rect 19475 930 19520 1050
rect 19640 930 19685 1050
rect 19805 930 19850 1050
rect 19970 930 20025 1050
rect 20145 930 20190 1050
rect 20310 930 20355 1050
rect 20475 930 20520 1050
rect 20640 930 20695 1050
rect 20815 930 20860 1050
rect 20980 930 21025 1050
rect 21145 930 21190 1050
rect 21310 930 21365 1050
rect 21485 930 21530 1050
rect 21650 930 21695 1050
rect 21815 930 21860 1050
rect 21980 930 22035 1050
rect 22155 930 22200 1050
rect 22320 930 22365 1050
rect 22485 930 22530 1050
rect 22650 930 22705 1050
rect 22825 930 22870 1050
rect 22990 930 23035 1050
rect 23155 930 23200 1050
rect 23320 930 23375 1050
rect 23495 930 23540 1050
rect 23660 930 23705 1050
rect 23825 930 23870 1050
rect 23990 930 24000 1050
rect 18500 885 24000 930
rect 18500 765 18510 885
rect 18630 765 18685 885
rect 18805 765 18850 885
rect 18970 765 19015 885
rect 19135 765 19180 885
rect 19300 765 19355 885
rect 19475 765 19520 885
rect 19640 765 19685 885
rect 19805 765 19850 885
rect 19970 765 20025 885
rect 20145 765 20190 885
rect 20310 765 20355 885
rect 20475 765 20520 885
rect 20640 765 20695 885
rect 20815 765 20860 885
rect 20980 765 21025 885
rect 21145 765 21190 885
rect 21310 765 21365 885
rect 21485 765 21530 885
rect 21650 765 21695 885
rect 21815 765 21860 885
rect 21980 765 22035 885
rect 22155 765 22200 885
rect 22320 765 22365 885
rect 22485 765 22530 885
rect 22650 765 22705 885
rect 22825 765 22870 885
rect 22990 765 23035 885
rect 23155 765 23200 885
rect 23320 765 23375 885
rect 23495 765 23540 885
rect 23660 765 23705 885
rect 23825 765 23870 885
rect 23990 765 24000 885
rect 18500 710 24000 765
rect 18500 590 18510 710
rect 18630 590 18685 710
rect 18805 590 18850 710
rect 18970 590 19015 710
rect 19135 590 19180 710
rect 19300 590 19355 710
rect 19475 590 19520 710
rect 19640 590 19685 710
rect 19805 590 19850 710
rect 19970 590 20025 710
rect 20145 590 20190 710
rect 20310 590 20355 710
rect 20475 590 20520 710
rect 20640 590 20695 710
rect 20815 590 20860 710
rect 20980 590 21025 710
rect 21145 590 21190 710
rect 21310 590 21365 710
rect 21485 590 21530 710
rect 21650 590 21695 710
rect 21815 590 21860 710
rect 21980 590 22035 710
rect 22155 590 22200 710
rect 22320 590 22365 710
rect 22485 590 22530 710
rect 22650 590 22705 710
rect 22825 590 22870 710
rect 22990 590 23035 710
rect 23155 590 23200 710
rect 23320 590 23375 710
rect 23495 590 23540 710
rect 23660 590 23705 710
rect 23825 590 23870 710
rect 23990 590 24000 710
rect 18500 545 24000 590
rect 18500 425 18510 545
rect 18630 425 18685 545
rect 18805 425 18850 545
rect 18970 425 19015 545
rect 19135 425 19180 545
rect 19300 425 19355 545
rect 19475 425 19520 545
rect 19640 425 19685 545
rect 19805 425 19850 545
rect 19970 425 20025 545
rect 20145 425 20190 545
rect 20310 425 20355 545
rect 20475 425 20520 545
rect 20640 425 20695 545
rect 20815 425 20860 545
rect 20980 425 21025 545
rect 21145 425 21190 545
rect 21310 425 21365 545
rect 21485 425 21530 545
rect 21650 425 21695 545
rect 21815 425 21860 545
rect 21980 425 22035 545
rect 22155 425 22200 545
rect 22320 425 22365 545
rect 22485 425 22530 545
rect 22650 425 22705 545
rect 22825 425 22870 545
rect 22990 425 23035 545
rect 23155 425 23200 545
rect 23320 425 23375 545
rect 23495 425 23540 545
rect 23660 425 23705 545
rect 23825 425 23870 545
rect 23990 425 24000 545
rect 18500 380 24000 425
rect 18500 260 18510 380
rect 18630 260 18685 380
rect 18805 260 18850 380
rect 18970 260 19015 380
rect 19135 260 19180 380
rect 19300 260 19355 380
rect 19475 260 19520 380
rect 19640 260 19685 380
rect 19805 260 19850 380
rect 19970 260 20025 380
rect 20145 260 20190 380
rect 20310 260 20355 380
rect 20475 260 20520 380
rect 20640 260 20695 380
rect 20815 260 20860 380
rect 20980 260 21025 380
rect 21145 260 21190 380
rect 21310 260 21365 380
rect 21485 260 21530 380
rect 21650 260 21695 380
rect 21815 260 21860 380
rect 21980 260 22035 380
rect 22155 260 22200 380
rect 22320 260 22365 380
rect 22485 260 22530 380
rect 22650 260 22705 380
rect 22825 260 22870 380
rect 22990 260 23035 380
rect 23155 260 23200 380
rect 23320 260 23375 380
rect 23495 260 23540 380
rect 23660 260 23705 380
rect 23825 260 23870 380
rect 23990 260 24000 380
rect 18500 215 24000 260
rect 18500 95 18510 215
rect 18630 95 18685 215
rect 18805 95 18850 215
rect 18970 95 19015 215
rect 19135 95 19180 215
rect 19300 95 19355 215
rect 19475 95 19520 215
rect 19640 95 19685 215
rect 19805 95 19850 215
rect 19970 95 20025 215
rect 20145 95 20190 215
rect 20310 95 20355 215
rect 20475 95 20520 215
rect 20640 95 20695 215
rect 20815 95 20860 215
rect 20980 95 21025 215
rect 21145 95 21190 215
rect 21310 95 21365 215
rect 21485 95 21530 215
rect 21650 95 21695 215
rect 21815 95 21860 215
rect 21980 95 22035 215
rect 22155 95 22200 215
rect 22320 95 22365 215
rect 22485 95 22530 215
rect 22650 95 22705 215
rect 22825 95 22870 215
rect 22990 95 23035 215
rect 23155 95 23200 215
rect 23320 95 23375 215
rect 23495 95 23540 215
rect 23660 95 23705 215
rect 23825 95 23870 215
rect 23990 95 24000 215
rect 18500 40 24000 95
rect 18500 -80 18510 40
rect 18630 -80 18685 40
rect 18805 -80 18850 40
rect 18970 -80 19015 40
rect 19135 -80 19180 40
rect 19300 -80 19355 40
rect 19475 -80 19520 40
rect 19640 -80 19685 40
rect 19805 -80 19850 40
rect 19970 -80 20025 40
rect 20145 -80 20190 40
rect 20310 -80 20355 40
rect 20475 -80 20520 40
rect 20640 -80 20695 40
rect 20815 -80 20860 40
rect 20980 -80 21025 40
rect 21145 -80 21190 40
rect 21310 -80 21365 40
rect 21485 -80 21530 40
rect 21650 -80 21695 40
rect 21815 -80 21860 40
rect 21980 -80 22035 40
rect 22155 -80 22200 40
rect 22320 -80 22365 40
rect 22485 -80 22530 40
rect 22650 -80 22705 40
rect 22825 -80 22870 40
rect 22990 -80 23035 40
rect 23155 -80 23200 40
rect 23320 -80 23375 40
rect 23495 -80 23540 40
rect 23660 -80 23705 40
rect 23825 -80 23870 40
rect 23990 -80 24000 40
rect 18500 -125 24000 -80
rect 18500 -245 18510 -125
rect 18630 -245 18685 -125
rect 18805 -245 18850 -125
rect 18970 -245 19015 -125
rect 19135 -245 19180 -125
rect 19300 -245 19355 -125
rect 19475 -245 19520 -125
rect 19640 -245 19685 -125
rect 19805 -245 19850 -125
rect 19970 -245 20025 -125
rect 20145 -245 20190 -125
rect 20310 -245 20355 -125
rect 20475 -245 20520 -125
rect 20640 -245 20695 -125
rect 20815 -245 20860 -125
rect 20980 -245 21025 -125
rect 21145 -245 21190 -125
rect 21310 -245 21365 -125
rect 21485 -245 21530 -125
rect 21650 -245 21695 -125
rect 21815 -245 21860 -125
rect 21980 -245 22035 -125
rect 22155 -245 22200 -125
rect 22320 -245 22365 -125
rect 22485 -245 22530 -125
rect 22650 -245 22705 -125
rect 22825 -245 22870 -125
rect 22990 -245 23035 -125
rect 23155 -245 23200 -125
rect 23320 -245 23375 -125
rect 23495 -245 23540 -125
rect 23660 -245 23705 -125
rect 23825 -245 23870 -125
rect 23990 -245 24000 -125
rect 18500 -290 24000 -245
rect 18500 -410 18510 -290
rect 18630 -410 18685 -290
rect 18805 -410 18850 -290
rect 18970 -410 19015 -290
rect 19135 -410 19180 -290
rect 19300 -410 19355 -290
rect 19475 -410 19520 -290
rect 19640 -410 19685 -290
rect 19805 -410 19850 -290
rect 19970 -410 20025 -290
rect 20145 -410 20190 -290
rect 20310 -410 20355 -290
rect 20475 -410 20520 -290
rect 20640 -410 20695 -290
rect 20815 -410 20860 -290
rect 20980 -410 21025 -290
rect 21145 -410 21190 -290
rect 21310 -410 21365 -290
rect 21485 -410 21530 -290
rect 21650 -410 21695 -290
rect 21815 -410 21860 -290
rect 21980 -410 22035 -290
rect 22155 -410 22200 -290
rect 22320 -410 22365 -290
rect 22485 -410 22530 -290
rect 22650 -410 22705 -290
rect 22825 -410 22870 -290
rect 22990 -410 23035 -290
rect 23155 -410 23200 -290
rect 23320 -410 23375 -290
rect 23495 -410 23540 -290
rect 23660 -410 23705 -290
rect 23825 -410 23870 -290
rect 23990 -410 24000 -290
rect 18500 -455 24000 -410
rect 18500 -575 18510 -455
rect 18630 -575 18685 -455
rect 18805 -575 18850 -455
rect 18970 -575 19015 -455
rect 19135 -575 19180 -455
rect 19300 -575 19355 -455
rect 19475 -575 19520 -455
rect 19640 -575 19685 -455
rect 19805 -575 19850 -455
rect 19970 -575 20025 -455
rect 20145 -575 20190 -455
rect 20310 -575 20355 -455
rect 20475 -575 20520 -455
rect 20640 -575 20695 -455
rect 20815 -575 20860 -455
rect 20980 -575 21025 -455
rect 21145 -575 21190 -455
rect 21310 -575 21365 -455
rect 21485 -575 21530 -455
rect 21650 -575 21695 -455
rect 21815 -575 21860 -455
rect 21980 -575 22035 -455
rect 22155 -575 22200 -455
rect 22320 -575 22365 -455
rect 22485 -575 22530 -455
rect 22650 -575 22705 -455
rect 22825 -575 22870 -455
rect 22990 -575 23035 -455
rect 23155 -575 23200 -455
rect 23320 -575 23375 -455
rect 23495 -575 23540 -455
rect 23660 -575 23705 -455
rect 23825 -575 23870 -455
rect 23990 -575 24000 -455
rect 18500 -630 24000 -575
rect 18500 -750 18510 -630
rect 18630 -750 18685 -630
rect 18805 -750 18850 -630
rect 18970 -750 19015 -630
rect 19135 -750 19180 -630
rect 19300 -750 19355 -630
rect 19475 -750 19520 -630
rect 19640 -750 19685 -630
rect 19805 -750 19850 -630
rect 19970 -750 20025 -630
rect 20145 -750 20190 -630
rect 20310 -750 20355 -630
rect 20475 -750 20520 -630
rect 20640 -750 20695 -630
rect 20815 -750 20860 -630
rect 20980 -750 21025 -630
rect 21145 -750 21190 -630
rect 21310 -750 21365 -630
rect 21485 -750 21530 -630
rect 21650 -750 21695 -630
rect 21815 -750 21860 -630
rect 21980 -750 22035 -630
rect 22155 -750 22200 -630
rect 22320 -750 22365 -630
rect 22485 -750 22530 -630
rect 22650 -750 22705 -630
rect 22825 -750 22870 -630
rect 22990 -750 23035 -630
rect 23155 -750 23200 -630
rect 23320 -750 23375 -630
rect 23495 -750 23540 -630
rect 23660 -750 23705 -630
rect 23825 -750 23870 -630
rect 23990 -750 24000 -630
rect 18500 -795 24000 -750
rect 18500 -915 18510 -795
rect 18630 -915 18685 -795
rect 18805 -915 18850 -795
rect 18970 -915 19015 -795
rect 19135 -915 19180 -795
rect 19300 -915 19355 -795
rect 19475 -915 19520 -795
rect 19640 -915 19685 -795
rect 19805 -915 19850 -795
rect 19970 -915 20025 -795
rect 20145 -915 20190 -795
rect 20310 -915 20355 -795
rect 20475 -915 20520 -795
rect 20640 -915 20695 -795
rect 20815 -915 20860 -795
rect 20980 -915 21025 -795
rect 21145 -915 21190 -795
rect 21310 -915 21365 -795
rect 21485 -915 21530 -795
rect 21650 -915 21695 -795
rect 21815 -915 21860 -795
rect 21980 -915 22035 -795
rect 22155 -915 22200 -795
rect 22320 -915 22365 -795
rect 22485 -915 22530 -795
rect 22650 -915 22705 -795
rect 22825 -915 22870 -795
rect 22990 -915 23035 -795
rect 23155 -915 23200 -795
rect 23320 -915 23375 -795
rect 23495 -915 23540 -795
rect 23660 -915 23705 -795
rect 23825 -915 23870 -795
rect 23990 -915 24000 -795
rect 18500 -960 24000 -915
rect 18500 -1080 18510 -960
rect 18630 -1080 18685 -960
rect 18805 -1080 18850 -960
rect 18970 -1080 19015 -960
rect 19135 -1080 19180 -960
rect 19300 -1080 19355 -960
rect 19475 -1080 19520 -960
rect 19640 -1080 19685 -960
rect 19805 -1080 19850 -960
rect 19970 -1080 20025 -960
rect 20145 -1080 20190 -960
rect 20310 -1080 20355 -960
rect 20475 -1080 20520 -960
rect 20640 -1080 20695 -960
rect 20815 -1080 20860 -960
rect 20980 -1080 21025 -960
rect 21145 -1080 21190 -960
rect 21310 -1080 21365 -960
rect 21485 -1080 21530 -960
rect 21650 -1080 21695 -960
rect 21815 -1080 21860 -960
rect 21980 -1080 22035 -960
rect 22155 -1080 22200 -960
rect 22320 -1080 22365 -960
rect 22485 -1080 22530 -960
rect 22650 -1080 22705 -960
rect 22825 -1080 22870 -960
rect 22990 -1080 23035 -960
rect 23155 -1080 23200 -960
rect 23320 -1080 23375 -960
rect 23495 -1080 23540 -960
rect 23660 -1080 23705 -960
rect 23825 -1080 23870 -960
rect 23990 -1080 24000 -960
rect 18500 -1125 24000 -1080
rect 18500 -1245 18510 -1125
rect 18630 -1245 18685 -1125
rect 18805 -1245 18850 -1125
rect 18970 -1245 19015 -1125
rect 19135 -1245 19180 -1125
rect 19300 -1245 19355 -1125
rect 19475 -1245 19520 -1125
rect 19640 -1245 19685 -1125
rect 19805 -1245 19850 -1125
rect 19970 -1245 20025 -1125
rect 20145 -1245 20190 -1125
rect 20310 -1245 20355 -1125
rect 20475 -1245 20520 -1125
rect 20640 -1245 20695 -1125
rect 20815 -1245 20860 -1125
rect 20980 -1245 21025 -1125
rect 21145 -1245 21190 -1125
rect 21310 -1245 21365 -1125
rect 21485 -1245 21530 -1125
rect 21650 -1245 21695 -1125
rect 21815 -1245 21860 -1125
rect 21980 -1245 22035 -1125
rect 22155 -1245 22200 -1125
rect 22320 -1245 22365 -1125
rect 22485 -1245 22530 -1125
rect 22650 -1245 22705 -1125
rect 22825 -1245 22870 -1125
rect 22990 -1245 23035 -1125
rect 23155 -1245 23200 -1125
rect 23320 -1245 23375 -1125
rect 23495 -1245 23540 -1125
rect 23660 -1245 23705 -1125
rect 23825 -1245 23870 -1125
rect 23990 -1245 24000 -1125
rect 18500 -1300 24000 -1245
rect 18500 -1420 18510 -1300
rect 18630 -1420 18685 -1300
rect 18805 -1420 18850 -1300
rect 18970 -1420 19015 -1300
rect 19135 -1420 19180 -1300
rect 19300 -1420 19355 -1300
rect 19475 -1420 19520 -1300
rect 19640 -1420 19685 -1300
rect 19805 -1420 19850 -1300
rect 19970 -1420 20025 -1300
rect 20145 -1420 20190 -1300
rect 20310 -1420 20355 -1300
rect 20475 -1420 20520 -1300
rect 20640 -1420 20695 -1300
rect 20815 -1420 20860 -1300
rect 20980 -1420 21025 -1300
rect 21145 -1420 21190 -1300
rect 21310 -1420 21365 -1300
rect 21485 -1420 21530 -1300
rect 21650 -1420 21695 -1300
rect 21815 -1420 21860 -1300
rect 21980 -1420 22035 -1300
rect 22155 -1420 22200 -1300
rect 22320 -1420 22365 -1300
rect 22485 -1420 22530 -1300
rect 22650 -1420 22705 -1300
rect 22825 -1420 22870 -1300
rect 22990 -1420 23035 -1300
rect 23155 -1420 23200 -1300
rect 23320 -1420 23375 -1300
rect 23495 -1420 23540 -1300
rect 23660 -1420 23705 -1300
rect 23825 -1420 23870 -1300
rect 23990 -1420 24000 -1300
rect 18500 -1465 24000 -1420
rect 18500 -1585 18510 -1465
rect 18630 -1585 18685 -1465
rect 18805 -1585 18850 -1465
rect 18970 -1585 19015 -1465
rect 19135 -1585 19180 -1465
rect 19300 -1585 19355 -1465
rect 19475 -1585 19520 -1465
rect 19640 -1585 19685 -1465
rect 19805 -1585 19850 -1465
rect 19970 -1585 20025 -1465
rect 20145 -1585 20190 -1465
rect 20310 -1585 20355 -1465
rect 20475 -1585 20520 -1465
rect 20640 -1585 20695 -1465
rect 20815 -1585 20860 -1465
rect 20980 -1585 21025 -1465
rect 21145 -1585 21190 -1465
rect 21310 -1585 21365 -1465
rect 21485 -1585 21530 -1465
rect 21650 -1585 21695 -1465
rect 21815 -1585 21860 -1465
rect 21980 -1585 22035 -1465
rect 22155 -1585 22200 -1465
rect 22320 -1585 22365 -1465
rect 22485 -1585 22530 -1465
rect 22650 -1585 22705 -1465
rect 22825 -1585 22870 -1465
rect 22990 -1585 23035 -1465
rect 23155 -1585 23200 -1465
rect 23320 -1585 23375 -1465
rect 23495 -1585 23540 -1465
rect 23660 -1585 23705 -1465
rect 23825 -1585 23870 -1465
rect 23990 -1585 24000 -1465
rect 18500 -1630 24000 -1585
rect 18500 -1750 18510 -1630
rect 18630 -1750 18685 -1630
rect 18805 -1750 18850 -1630
rect 18970 -1750 19015 -1630
rect 19135 -1750 19180 -1630
rect 19300 -1750 19355 -1630
rect 19475 -1750 19520 -1630
rect 19640 -1750 19685 -1630
rect 19805 -1750 19850 -1630
rect 19970 -1750 20025 -1630
rect 20145 -1750 20190 -1630
rect 20310 -1750 20355 -1630
rect 20475 -1750 20520 -1630
rect 20640 -1750 20695 -1630
rect 20815 -1750 20860 -1630
rect 20980 -1750 21025 -1630
rect 21145 -1750 21190 -1630
rect 21310 -1750 21365 -1630
rect 21485 -1750 21530 -1630
rect 21650 -1750 21695 -1630
rect 21815 -1750 21860 -1630
rect 21980 -1750 22035 -1630
rect 22155 -1750 22200 -1630
rect 22320 -1750 22365 -1630
rect 22485 -1750 22530 -1630
rect 22650 -1750 22705 -1630
rect 22825 -1750 22870 -1630
rect 22990 -1750 23035 -1630
rect 23155 -1750 23200 -1630
rect 23320 -1750 23375 -1630
rect 23495 -1750 23540 -1630
rect 23660 -1750 23705 -1630
rect 23825 -1750 23870 -1630
rect 23990 -1750 24000 -1630
rect 18500 -1795 24000 -1750
rect 18500 -1915 18510 -1795
rect 18630 -1915 18685 -1795
rect 18805 -1915 18850 -1795
rect 18970 -1915 19015 -1795
rect 19135 -1915 19180 -1795
rect 19300 -1915 19355 -1795
rect 19475 -1915 19520 -1795
rect 19640 -1915 19685 -1795
rect 19805 -1915 19850 -1795
rect 19970 -1915 20025 -1795
rect 20145 -1915 20190 -1795
rect 20310 -1915 20355 -1795
rect 20475 -1915 20520 -1795
rect 20640 -1915 20695 -1795
rect 20815 -1915 20860 -1795
rect 20980 -1915 21025 -1795
rect 21145 -1915 21190 -1795
rect 21310 -1915 21365 -1795
rect 21485 -1915 21530 -1795
rect 21650 -1915 21695 -1795
rect 21815 -1915 21860 -1795
rect 21980 -1915 22035 -1795
rect 22155 -1915 22200 -1795
rect 22320 -1915 22365 -1795
rect 22485 -1915 22530 -1795
rect 22650 -1915 22705 -1795
rect 22825 -1915 22870 -1795
rect 22990 -1915 23035 -1795
rect 23155 -1915 23200 -1795
rect 23320 -1915 23375 -1795
rect 23495 -1915 23540 -1795
rect 23660 -1915 23705 -1795
rect 23825 -1915 23870 -1795
rect 23990 -1915 24000 -1795
rect 18500 -1970 24000 -1915
rect 18500 -2090 18510 -1970
rect 18630 -2090 18685 -1970
rect 18805 -2090 18850 -1970
rect 18970 -2090 19015 -1970
rect 19135 -2090 19180 -1970
rect 19300 -2090 19355 -1970
rect 19475 -2090 19520 -1970
rect 19640 -2090 19685 -1970
rect 19805 -2090 19850 -1970
rect 19970 -2090 20025 -1970
rect 20145 -2090 20190 -1970
rect 20310 -2090 20355 -1970
rect 20475 -2090 20520 -1970
rect 20640 -2090 20695 -1970
rect 20815 -2090 20860 -1970
rect 20980 -2090 21025 -1970
rect 21145 -2090 21190 -1970
rect 21310 -2090 21365 -1970
rect 21485 -2090 21530 -1970
rect 21650 -2090 21695 -1970
rect 21815 -2090 21860 -1970
rect 21980 -2090 22035 -1970
rect 22155 -2090 22200 -1970
rect 22320 -2090 22365 -1970
rect 22485 -2090 22530 -1970
rect 22650 -2090 22705 -1970
rect 22825 -2090 22870 -1970
rect 22990 -2090 23035 -1970
rect 23155 -2090 23200 -1970
rect 23320 -2090 23375 -1970
rect 23495 -2090 23540 -1970
rect 23660 -2090 23705 -1970
rect 23825 -2090 23870 -1970
rect 23990 -2090 24000 -1970
rect 18500 -2135 24000 -2090
rect 18500 -2255 18510 -2135
rect 18630 -2255 18685 -2135
rect 18805 -2255 18850 -2135
rect 18970 -2255 19015 -2135
rect 19135 -2255 19180 -2135
rect 19300 -2255 19355 -2135
rect 19475 -2255 19520 -2135
rect 19640 -2255 19685 -2135
rect 19805 -2255 19850 -2135
rect 19970 -2255 20025 -2135
rect 20145 -2255 20190 -2135
rect 20310 -2255 20355 -2135
rect 20475 -2255 20520 -2135
rect 20640 -2255 20695 -2135
rect 20815 -2255 20860 -2135
rect 20980 -2255 21025 -2135
rect 21145 -2255 21190 -2135
rect 21310 -2255 21365 -2135
rect 21485 -2255 21530 -2135
rect 21650 -2255 21695 -2135
rect 21815 -2255 21860 -2135
rect 21980 -2255 22035 -2135
rect 22155 -2255 22200 -2135
rect 22320 -2255 22365 -2135
rect 22485 -2255 22530 -2135
rect 22650 -2255 22705 -2135
rect 22825 -2255 22870 -2135
rect 22990 -2255 23035 -2135
rect 23155 -2255 23200 -2135
rect 23320 -2255 23375 -2135
rect 23495 -2255 23540 -2135
rect 23660 -2255 23705 -2135
rect 23825 -2255 23870 -2135
rect 23990 -2255 24000 -2135
rect 18500 -2300 24000 -2255
rect 18500 -2420 18510 -2300
rect 18630 -2420 18685 -2300
rect 18805 -2420 18850 -2300
rect 18970 -2420 19015 -2300
rect 19135 -2420 19180 -2300
rect 19300 -2420 19355 -2300
rect 19475 -2420 19520 -2300
rect 19640 -2420 19685 -2300
rect 19805 -2420 19850 -2300
rect 19970 -2420 20025 -2300
rect 20145 -2420 20190 -2300
rect 20310 -2420 20355 -2300
rect 20475 -2420 20520 -2300
rect 20640 -2420 20695 -2300
rect 20815 -2420 20860 -2300
rect 20980 -2420 21025 -2300
rect 21145 -2420 21190 -2300
rect 21310 -2420 21365 -2300
rect 21485 -2420 21530 -2300
rect 21650 -2420 21695 -2300
rect 21815 -2420 21860 -2300
rect 21980 -2420 22035 -2300
rect 22155 -2420 22200 -2300
rect 22320 -2420 22365 -2300
rect 22485 -2420 22530 -2300
rect 22650 -2420 22705 -2300
rect 22825 -2420 22870 -2300
rect 22990 -2420 23035 -2300
rect 23155 -2420 23200 -2300
rect 23320 -2420 23375 -2300
rect 23495 -2420 23540 -2300
rect 23660 -2420 23705 -2300
rect 23825 -2420 23870 -2300
rect 23990 -2420 24000 -2300
rect 18500 -2465 24000 -2420
rect 18500 -2585 18510 -2465
rect 18630 -2585 18685 -2465
rect 18805 -2585 18850 -2465
rect 18970 -2585 19015 -2465
rect 19135 -2585 19180 -2465
rect 19300 -2585 19355 -2465
rect 19475 -2585 19520 -2465
rect 19640 -2585 19685 -2465
rect 19805 -2585 19850 -2465
rect 19970 -2585 20025 -2465
rect 20145 -2585 20190 -2465
rect 20310 -2585 20355 -2465
rect 20475 -2585 20520 -2465
rect 20640 -2585 20695 -2465
rect 20815 -2585 20860 -2465
rect 20980 -2585 21025 -2465
rect 21145 -2585 21190 -2465
rect 21310 -2585 21365 -2465
rect 21485 -2585 21530 -2465
rect 21650 -2585 21695 -2465
rect 21815 -2585 21860 -2465
rect 21980 -2585 22035 -2465
rect 22155 -2585 22200 -2465
rect 22320 -2585 22365 -2465
rect 22485 -2585 22530 -2465
rect 22650 -2585 22705 -2465
rect 22825 -2585 22870 -2465
rect 22990 -2585 23035 -2465
rect 23155 -2585 23200 -2465
rect 23320 -2585 23375 -2465
rect 23495 -2585 23540 -2465
rect 23660 -2585 23705 -2465
rect 23825 -2585 23870 -2465
rect 23990 -2585 24000 -2465
rect 18500 -2640 24000 -2585
rect 18500 -2760 18510 -2640
rect 18630 -2760 18685 -2640
rect 18805 -2760 18850 -2640
rect 18970 -2760 19015 -2640
rect 19135 -2760 19180 -2640
rect 19300 -2760 19355 -2640
rect 19475 -2760 19520 -2640
rect 19640 -2760 19685 -2640
rect 19805 -2760 19850 -2640
rect 19970 -2760 20025 -2640
rect 20145 -2760 20190 -2640
rect 20310 -2760 20355 -2640
rect 20475 -2760 20520 -2640
rect 20640 -2760 20695 -2640
rect 20815 -2760 20860 -2640
rect 20980 -2760 21025 -2640
rect 21145 -2760 21190 -2640
rect 21310 -2760 21365 -2640
rect 21485 -2760 21530 -2640
rect 21650 -2760 21695 -2640
rect 21815 -2760 21860 -2640
rect 21980 -2760 22035 -2640
rect 22155 -2760 22200 -2640
rect 22320 -2760 22365 -2640
rect 22485 -2760 22530 -2640
rect 22650 -2760 22705 -2640
rect 22825 -2760 22870 -2640
rect 22990 -2760 23035 -2640
rect 23155 -2760 23200 -2640
rect 23320 -2760 23375 -2640
rect 23495 -2760 23540 -2640
rect 23660 -2760 23705 -2640
rect 23825 -2760 23870 -2640
rect 23990 -2760 24000 -2640
rect 18500 -2805 24000 -2760
rect 18500 -2925 18510 -2805
rect 18630 -2925 18685 -2805
rect 18805 -2925 18850 -2805
rect 18970 -2925 19015 -2805
rect 19135 -2925 19180 -2805
rect 19300 -2925 19355 -2805
rect 19475 -2925 19520 -2805
rect 19640 -2925 19685 -2805
rect 19805 -2925 19850 -2805
rect 19970 -2925 20025 -2805
rect 20145 -2925 20190 -2805
rect 20310 -2925 20355 -2805
rect 20475 -2925 20520 -2805
rect 20640 -2925 20695 -2805
rect 20815 -2925 20860 -2805
rect 20980 -2925 21025 -2805
rect 21145 -2925 21190 -2805
rect 21310 -2925 21365 -2805
rect 21485 -2925 21530 -2805
rect 21650 -2925 21695 -2805
rect 21815 -2925 21860 -2805
rect 21980 -2925 22035 -2805
rect 22155 -2925 22200 -2805
rect 22320 -2925 22365 -2805
rect 22485 -2925 22530 -2805
rect 22650 -2925 22705 -2805
rect 22825 -2925 22870 -2805
rect 22990 -2925 23035 -2805
rect 23155 -2925 23200 -2805
rect 23320 -2925 23375 -2805
rect 23495 -2925 23540 -2805
rect 23660 -2925 23705 -2805
rect 23825 -2925 23870 -2805
rect 23990 -2925 24000 -2805
rect 18500 -2970 24000 -2925
rect 18500 -3090 18510 -2970
rect 18630 -3090 18685 -2970
rect 18805 -3090 18850 -2970
rect 18970 -3090 19015 -2970
rect 19135 -3090 19180 -2970
rect 19300 -3090 19355 -2970
rect 19475 -3090 19520 -2970
rect 19640 -3090 19685 -2970
rect 19805 -3090 19850 -2970
rect 19970 -3090 20025 -2970
rect 20145 -3090 20190 -2970
rect 20310 -3090 20355 -2970
rect 20475 -3090 20520 -2970
rect 20640 -3090 20695 -2970
rect 20815 -3090 20860 -2970
rect 20980 -3090 21025 -2970
rect 21145 -3090 21190 -2970
rect 21310 -3090 21365 -2970
rect 21485 -3090 21530 -2970
rect 21650 -3090 21695 -2970
rect 21815 -3090 21860 -2970
rect 21980 -3090 22035 -2970
rect 22155 -3090 22200 -2970
rect 22320 -3090 22365 -2970
rect 22485 -3090 22530 -2970
rect 22650 -3090 22705 -2970
rect 22825 -3090 22870 -2970
rect 22990 -3090 23035 -2970
rect 23155 -3090 23200 -2970
rect 23320 -3090 23375 -2970
rect 23495 -3090 23540 -2970
rect 23660 -3090 23705 -2970
rect 23825 -3090 23870 -2970
rect 23990 -3090 24000 -2970
rect 18500 -3135 24000 -3090
rect 18500 -3255 18510 -3135
rect 18630 -3255 18685 -3135
rect 18805 -3255 18850 -3135
rect 18970 -3255 19015 -3135
rect 19135 -3255 19180 -3135
rect 19300 -3255 19355 -3135
rect 19475 -3255 19520 -3135
rect 19640 -3255 19685 -3135
rect 19805 -3255 19850 -3135
rect 19970 -3255 20025 -3135
rect 20145 -3255 20190 -3135
rect 20310 -3255 20355 -3135
rect 20475 -3255 20520 -3135
rect 20640 -3255 20695 -3135
rect 20815 -3255 20860 -3135
rect 20980 -3255 21025 -3135
rect 21145 -3255 21190 -3135
rect 21310 -3255 21365 -3135
rect 21485 -3255 21530 -3135
rect 21650 -3255 21695 -3135
rect 21815 -3255 21860 -3135
rect 21980 -3255 22035 -3135
rect 22155 -3255 22200 -3135
rect 22320 -3255 22365 -3135
rect 22485 -3255 22530 -3135
rect 22650 -3255 22705 -3135
rect 22825 -3255 22870 -3135
rect 22990 -3255 23035 -3135
rect 23155 -3255 23200 -3135
rect 23320 -3255 23375 -3135
rect 23495 -3255 23540 -3135
rect 23660 -3255 23705 -3135
rect 23825 -3255 23870 -3135
rect 23990 -3255 24000 -3135
rect 18500 -3310 24000 -3255
rect 18500 -3430 18510 -3310
rect 18630 -3430 18685 -3310
rect 18805 -3430 18850 -3310
rect 18970 -3430 19015 -3310
rect 19135 -3430 19180 -3310
rect 19300 -3430 19355 -3310
rect 19475 -3430 19520 -3310
rect 19640 -3430 19685 -3310
rect 19805 -3430 19850 -3310
rect 19970 -3430 20025 -3310
rect 20145 -3430 20190 -3310
rect 20310 -3430 20355 -3310
rect 20475 -3430 20520 -3310
rect 20640 -3430 20695 -3310
rect 20815 -3430 20860 -3310
rect 20980 -3430 21025 -3310
rect 21145 -3430 21190 -3310
rect 21310 -3430 21365 -3310
rect 21485 -3430 21530 -3310
rect 21650 -3430 21695 -3310
rect 21815 -3430 21860 -3310
rect 21980 -3430 22035 -3310
rect 22155 -3430 22200 -3310
rect 22320 -3430 22365 -3310
rect 22485 -3430 22530 -3310
rect 22650 -3430 22705 -3310
rect 22825 -3430 22870 -3310
rect 22990 -3430 23035 -3310
rect 23155 -3430 23200 -3310
rect 23320 -3430 23375 -3310
rect 23495 -3430 23540 -3310
rect 23660 -3430 23705 -3310
rect 23825 -3430 23870 -3310
rect 23990 -3430 24000 -3310
rect 18500 -3475 24000 -3430
rect 18500 -3595 18510 -3475
rect 18630 -3595 18685 -3475
rect 18805 -3595 18850 -3475
rect 18970 -3595 19015 -3475
rect 19135 -3595 19180 -3475
rect 19300 -3595 19355 -3475
rect 19475 -3595 19520 -3475
rect 19640 -3595 19685 -3475
rect 19805 -3595 19850 -3475
rect 19970 -3595 20025 -3475
rect 20145 -3595 20190 -3475
rect 20310 -3595 20355 -3475
rect 20475 -3595 20520 -3475
rect 20640 -3595 20695 -3475
rect 20815 -3595 20860 -3475
rect 20980 -3595 21025 -3475
rect 21145 -3595 21190 -3475
rect 21310 -3595 21365 -3475
rect 21485 -3595 21530 -3475
rect 21650 -3595 21695 -3475
rect 21815 -3595 21860 -3475
rect 21980 -3595 22035 -3475
rect 22155 -3595 22200 -3475
rect 22320 -3595 22365 -3475
rect 22485 -3595 22530 -3475
rect 22650 -3595 22705 -3475
rect 22825 -3595 22870 -3475
rect 22990 -3595 23035 -3475
rect 23155 -3595 23200 -3475
rect 23320 -3595 23375 -3475
rect 23495 -3595 23540 -3475
rect 23660 -3595 23705 -3475
rect 23825 -3595 23870 -3475
rect 23990 -3595 24000 -3475
rect 18500 -3640 24000 -3595
rect 18500 -3760 18510 -3640
rect 18630 -3760 18685 -3640
rect 18805 -3760 18850 -3640
rect 18970 -3760 19015 -3640
rect 19135 -3760 19180 -3640
rect 19300 -3760 19355 -3640
rect 19475 -3760 19520 -3640
rect 19640 -3760 19685 -3640
rect 19805 -3760 19850 -3640
rect 19970 -3760 20025 -3640
rect 20145 -3760 20190 -3640
rect 20310 -3760 20355 -3640
rect 20475 -3760 20520 -3640
rect 20640 -3760 20695 -3640
rect 20815 -3760 20860 -3640
rect 20980 -3760 21025 -3640
rect 21145 -3760 21190 -3640
rect 21310 -3760 21365 -3640
rect 21485 -3760 21530 -3640
rect 21650 -3760 21695 -3640
rect 21815 -3760 21860 -3640
rect 21980 -3760 22035 -3640
rect 22155 -3760 22200 -3640
rect 22320 -3760 22365 -3640
rect 22485 -3760 22530 -3640
rect 22650 -3760 22705 -3640
rect 22825 -3760 22870 -3640
rect 22990 -3760 23035 -3640
rect 23155 -3760 23200 -3640
rect 23320 -3760 23375 -3640
rect 23495 -3760 23540 -3640
rect 23660 -3760 23705 -3640
rect 23825 -3760 23870 -3640
rect 23990 -3760 24000 -3640
rect 18500 -3805 24000 -3760
rect 18500 -3925 18510 -3805
rect 18630 -3925 18685 -3805
rect 18805 -3925 18850 -3805
rect 18970 -3925 19015 -3805
rect 19135 -3925 19180 -3805
rect 19300 -3925 19355 -3805
rect 19475 -3925 19520 -3805
rect 19640 -3925 19685 -3805
rect 19805 -3925 19850 -3805
rect 19970 -3925 20025 -3805
rect 20145 -3925 20190 -3805
rect 20310 -3925 20355 -3805
rect 20475 -3925 20520 -3805
rect 20640 -3925 20695 -3805
rect 20815 -3925 20860 -3805
rect 20980 -3925 21025 -3805
rect 21145 -3925 21190 -3805
rect 21310 -3925 21365 -3805
rect 21485 -3925 21530 -3805
rect 21650 -3925 21695 -3805
rect 21815 -3925 21860 -3805
rect 21980 -3925 22035 -3805
rect 22155 -3925 22200 -3805
rect 22320 -3925 22365 -3805
rect 22485 -3925 22530 -3805
rect 22650 -3925 22705 -3805
rect 22825 -3925 22870 -3805
rect 22990 -3925 23035 -3805
rect 23155 -3925 23200 -3805
rect 23320 -3925 23375 -3805
rect 23495 -3925 23540 -3805
rect 23660 -3925 23705 -3805
rect 23825 -3925 23870 -3805
rect 23990 -3925 24000 -3805
rect 18500 -3980 24000 -3925
rect 18500 -4100 18510 -3980
rect 18630 -4100 18685 -3980
rect 18805 -4100 18850 -3980
rect 18970 -4100 19015 -3980
rect 19135 -4100 19180 -3980
rect 19300 -4100 19355 -3980
rect 19475 -4100 19520 -3980
rect 19640 -4100 19685 -3980
rect 19805 -4100 19850 -3980
rect 19970 -4100 20025 -3980
rect 20145 -4100 20190 -3980
rect 20310 -4100 20355 -3980
rect 20475 -4100 20520 -3980
rect 20640 -4100 20695 -3980
rect 20815 -4100 20860 -3980
rect 20980 -4100 21025 -3980
rect 21145 -4100 21190 -3980
rect 21310 -4100 21365 -3980
rect 21485 -4100 21530 -3980
rect 21650 -4100 21695 -3980
rect 21815 -4100 21860 -3980
rect 21980 -4100 22035 -3980
rect 22155 -4100 22200 -3980
rect 22320 -4100 22365 -3980
rect 22485 -4100 22530 -3980
rect 22650 -4100 22705 -3980
rect 22825 -4100 22870 -3980
rect 22990 -4100 23035 -3980
rect 23155 -4100 23200 -3980
rect 23320 -4100 23375 -3980
rect 23495 -4100 23540 -3980
rect 23660 -4100 23705 -3980
rect 23825 -4100 23870 -3980
rect 23990 -4100 24000 -3980
rect 18500 -4110 24000 -4100
rect 24190 1380 29690 1390
rect 24190 1260 24200 1380
rect 24320 1260 24375 1380
rect 24495 1260 24540 1380
rect 24660 1260 24705 1380
rect 24825 1260 24870 1380
rect 24990 1260 25045 1380
rect 25165 1260 25210 1380
rect 25330 1260 25375 1380
rect 25495 1260 25540 1380
rect 25660 1260 25715 1380
rect 25835 1260 25880 1380
rect 26000 1260 26045 1380
rect 26165 1260 26210 1380
rect 26330 1260 26385 1380
rect 26505 1260 26550 1380
rect 26670 1260 26715 1380
rect 26835 1260 26880 1380
rect 27000 1260 27055 1380
rect 27175 1260 27220 1380
rect 27340 1260 27385 1380
rect 27505 1260 27550 1380
rect 27670 1260 27725 1380
rect 27845 1260 27890 1380
rect 28010 1260 28055 1380
rect 28175 1260 28220 1380
rect 28340 1260 28395 1380
rect 28515 1260 28560 1380
rect 28680 1260 28725 1380
rect 28845 1260 28890 1380
rect 29010 1260 29065 1380
rect 29185 1260 29230 1380
rect 29350 1260 29395 1380
rect 29515 1260 29560 1380
rect 29680 1260 29690 1380
rect 24190 1215 29690 1260
rect 24190 1095 24200 1215
rect 24320 1095 24375 1215
rect 24495 1095 24540 1215
rect 24660 1095 24705 1215
rect 24825 1095 24870 1215
rect 24990 1095 25045 1215
rect 25165 1095 25210 1215
rect 25330 1095 25375 1215
rect 25495 1095 25540 1215
rect 25660 1095 25715 1215
rect 25835 1095 25880 1215
rect 26000 1095 26045 1215
rect 26165 1095 26210 1215
rect 26330 1095 26385 1215
rect 26505 1095 26550 1215
rect 26670 1095 26715 1215
rect 26835 1095 26880 1215
rect 27000 1095 27055 1215
rect 27175 1095 27220 1215
rect 27340 1095 27385 1215
rect 27505 1095 27550 1215
rect 27670 1095 27725 1215
rect 27845 1095 27890 1215
rect 28010 1095 28055 1215
rect 28175 1095 28220 1215
rect 28340 1095 28395 1215
rect 28515 1095 28560 1215
rect 28680 1095 28725 1215
rect 28845 1095 28890 1215
rect 29010 1095 29065 1215
rect 29185 1095 29230 1215
rect 29350 1095 29395 1215
rect 29515 1095 29560 1215
rect 29680 1095 29690 1215
rect 24190 1050 29690 1095
rect 24190 930 24200 1050
rect 24320 930 24375 1050
rect 24495 930 24540 1050
rect 24660 930 24705 1050
rect 24825 930 24870 1050
rect 24990 930 25045 1050
rect 25165 930 25210 1050
rect 25330 930 25375 1050
rect 25495 930 25540 1050
rect 25660 930 25715 1050
rect 25835 930 25880 1050
rect 26000 930 26045 1050
rect 26165 930 26210 1050
rect 26330 930 26385 1050
rect 26505 930 26550 1050
rect 26670 930 26715 1050
rect 26835 930 26880 1050
rect 27000 930 27055 1050
rect 27175 930 27220 1050
rect 27340 930 27385 1050
rect 27505 930 27550 1050
rect 27670 930 27725 1050
rect 27845 930 27890 1050
rect 28010 930 28055 1050
rect 28175 930 28220 1050
rect 28340 930 28395 1050
rect 28515 930 28560 1050
rect 28680 930 28725 1050
rect 28845 930 28890 1050
rect 29010 930 29065 1050
rect 29185 930 29230 1050
rect 29350 930 29395 1050
rect 29515 930 29560 1050
rect 29680 930 29690 1050
rect 24190 885 29690 930
rect 24190 765 24200 885
rect 24320 765 24375 885
rect 24495 765 24540 885
rect 24660 765 24705 885
rect 24825 765 24870 885
rect 24990 765 25045 885
rect 25165 765 25210 885
rect 25330 765 25375 885
rect 25495 765 25540 885
rect 25660 765 25715 885
rect 25835 765 25880 885
rect 26000 765 26045 885
rect 26165 765 26210 885
rect 26330 765 26385 885
rect 26505 765 26550 885
rect 26670 765 26715 885
rect 26835 765 26880 885
rect 27000 765 27055 885
rect 27175 765 27220 885
rect 27340 765 27385 885
rect 27505 765 27550 885
rect 27670 765 27725 885
rect 27845 765 27890 885
rect 28010 765 28055 885
rect 28175 765 28220 885
rect 28340 765 28395 885
rect 28515 765 28560 885
rect 28680 765 28725 885
rect 28845 765 28890 885
rect 29010 765 29065 885
rect 29185 765 29230 885
rect 29350 765 29395 885
rect 29515 765 29560 885
rect 29680 765 29690 885
rect 24190 710 29690 765
rect 24190 590 24200 710
rect 24320 590 24375 710
rect 24495 590 24540 710
rect 24660 590 24705 710
rect 24825 590 24870 710
rect 24990 590 25045 710
rect 25165 590 25210 710
rect 25330 590 25375 710
rect 25495 590 25540 710
rect 25660 590 25715 710
rect 25835 590 25880 710
rect 26000 590 26045 710
rect 26165 590 26210 710
rect 26330 590 26385 710
rect 26505 590 26550 710
rect 26670 590 26715 710
rect 26835 590 26880 710
rect 27000 590 27055 710
rect 27175 590 27220 710
rect 27340 590 27385 710
rect 27505 590 27550 710
rect 27670 590 27725 710
rect 27845 590 27890 710
rect 28010 590 28055 710
rect 28175 590 28220 710
rect 28340 590 28395 710
rect 28515 590 28560 710
rect 28680 590 28725 710
rect 28845 590 28890 710
rect 29010 590 29065 710
rect 29185 590 29230 710
rect 29350 590 29395 710
rect 29515 590 29560 710
rect 29680 590 29690 710
rect 24190 545 29690 590
rect 24190 425 24200 545
rect 24320 425 24375 545
rect 24495 425 24540 545
rect 24660 425 24705 545
rect 24825 425 24870 545
rect 24990 425 25045 545
rect 25165 425 25210 545
rect 25330 425 25375 545
rect 25495 425 25540 545
rect 25660 425 25715 545
rect 25835 425 25880 545
rect 26000 425 26045 545
rect 26165 425 26210 545
rect 26330 425 26385 545
rect 26505 425 26550 545
rect 26670 425 26715 545
rect 26835 425 26880 545
rect 27000 425 27055 545
rect 27175 425 27220 545
rect 27340 425 27385 545
rect 27505 425 27550 545
rect 27670 425 27725 545
rect 27845 425 27890 545
rect 28010 425 28055 545
rect 28175 425 28220 545
rect 28340 425 28395 545
rect 28515 425 28560 545
rect 28680 425 28725 545
rect 28845 425 28890 545
rect 29010 425 29065 545
rect 29185 425 29230 545
rect 29350 425 29395 545
rect 29515 425 29560 545
rect 29680 425 29690 545
rect 24190 380 29690 425
rect 24190 260 24200 380
rect 24320 260 24375 380
rect 24495 260 24540 380
rect 24660 260 24705 380
rect 24825 260 24870 380
rect 24990 260 25045 380
rect 25165 260 25210 380
rect 25330 260 25375 380
rect 25495 260 25540 380
rect 25660 260 25715 380
rect 25835 260 25880 380
rect 26000 260 26045 380
rect 26165 260 26210 380
rect 26330 260 26385 380
rect 26505 260 26550 380
rect 26670 260 26715 380
rect 26835 260 26880 380
rect 27000 260 27055 380
rect 27175 260 27220 380
rect 27340 260 27385 380
rect 27505 260 27550 380
rect 27670 260 27725 380
rect 27845 260 27890 380
rect 28010 260 28055 380
rect 28175 260 28220 380
rect 28340 260 28395 380
rect 28515 260 28560 380
rect 28680 260 28725 380
rect 28845 260 28890 380
rect 29010 260 29065 380
rect 29185 260 29230 380
rect 29350 260 29395 380
rect 29515 260 29560 380
rect 29680 260 29690 380
rect 24190 215 29690 260
rect 24190 95 24200 215
rect 24320 95 24375 215
rect 24495 95 24540 215
rect 24660 95 24705 215
rect 24825 95 24870 215
rect 24990 95 25045 215
rect 25165 95 25210 215
rect 25330 95 25375 215
rect 25495 95 25540 215
rect 25660 95 25715 215
rect 25835 95 25880 215
rect 26000 95 26045 215
rect 26165 95 26210 215
rect 26330 95 26385 215
rect 26505 95 26550 215
rect 26670 95 26715 215
rect 26835 95 26880 215
rect 27000 95 27055 215
rect 27175 95 27220 215
rect 27340 95 27385 215
rect 27505 95 27550 215
rect 27670 95 27725 215
rect 27845 95 27890 215
rect 28010 95 28055 215
rect 28175 95 28220 215
rect 28340 95 28395 215
rect 28515 95 28560 215
rect 28680 95 28725 215
rect 28845 95 28890 215
rect 29010 95 29065 215
rect 29185 95 29230 215
rect 29350 95 29395 215
rect 29515 95 29560 215
rect 29680 95 29690 215
rect 24190 40 29690 95
rect 24190 -80 24200 40
rect 24320 -80 24375 40
rect 24495 -80 24540 40
rect 24660 -80 24705 40
rect 24825 -80 24870 40
rect 24990 -80 25045 40
rect 25165 -80 25210 40
rect 25330 -80 25375 40
rect 25495 -80 25540 40
rect 25660 -80 25715 40
rect 25835 -80 25880 40
rect 26000 -80 26045 40
rect 26165 -80 26210 40
rect 26330 -80 26385 40
rect 26505 -80 26550 40
rect 26670 -80 26715 40
rect 26835 -80 26880 40
rect 27000 -80 27055 40
rect 27175 -80 27220 40
rect 27340 -80 27385 40
rect 27505 -80 27550 40
rect 27670 -80 27725 40
rect 27845 -80 27890 40
rect 28010 -80 28055 40
rect 28175 -80 28220 40
rect 28340 -80 28395 40
rect 28515 -80 28560 40
rect 28680 -80 28725 40
rect 28845 -80 28890 40
rect 29010 -80 29065 40
rect 29185 -80 29230 40
rect 29350 -80 29395 40
rect 29515 -80 29560 40
rect 29680 -80 29690 40
rect 24190 -125 29690 -80
rect 24190 -245 24200 -125
rect 24320 -245 24375 -125
rect 24495 -245 24540 -125
rect 24660 -245 24705 -125
rect 24825 -245 24870 -125
rect 24990 -245 25045 -125
rect 25165 -245 25210 -125
rect 25330 -245 25375 -125
rect 25495 -245 25540 -125
rect 25660 -245 25715 -125
rect 25835 -245 25880 -125
rect 26000 -245 26045 -125
rect 26165 -245 26210 -125
rect 26330 -245 26385 -125
rect 26505 -245 26550 -125
rect 26670 -245 26715 -125
rect 26835 -245 26880 -125
rect 27000 -245 27055 -125
rect 27175 -245 27220 -125
rect 27340 -245 27385 -125
rect 27505 -245 27550 -125
rect 27670 -245 27725 -125
rect 27845 -245 27890 -125
rect 28010 -245 28055 -125
rect 28175 -245 28220 -125
rect 28340 -245 28395 -125
rect 28515 -245 28560 -125
rect 28680 -245 28725 -125
rect 28845 -245 28890 -125
rect 29010 -245 29065 -125
rect 29185 -245 29230 -125
rect 29350 -245 29395 -125
rect 29515 -245 29560 -125
rect 29680 -245 29690 -125
rect 24190 -290 29690 -245
rect 24190 -410 24200 -290
rect 24320 -410 24375 -290
rect 24495 -410 24540 -290
rect 24660 -410 24705 -290
rect 24825 -410 24870 -290
rect 24990 -410 25045 -290
rect 25165 -410 25210 -290
rect 25330 -410 25375 -290
rect 25495 -410 25540 -290
rect 25660 -410 25715 -290
rect 25835 -410 25880 -290
rect 26000 -410 26045 -290
rect 26165 -410 26210 -290
rect 26330 -410 26385 -290
rect 26505 -410 26550 -290
rect 26670 -410 26715 -290
rect 26835 -410 26880 -290
rect 27000 -410 27055 -290
rect 27175 -410 27220 -290
rect 27340 -410 27385 -290
rect 27505 -410 27550 -290
rect 27670 -410 27725 -290
rect 27845 -410 27890 -290
rect 28010 -410 28055 -290
rect 28175 -410 28220 -290
rect 28340 -410 28395 -290
rect 28515 -410 28560 -290
rect 28680 -410 28725 -290
rect 28845 -410 28890 -290
rect 29010 -410 29065 -290
rect 29185 -410 29230 -290
rect 29350 -410 29395 -290
rect 29515 -410 29560 -290
rect 29680 -410 29690 -290
rect 24190 -455 29690 -410
rect 24190 -575 24200 -455
rect 24320 -575 24375 -455
rect 24495 -575 24540 -455
rect 24660 -575 24705 -455
rect 24825 -575 24870 -455
rect 24990 -575 25045 -455
rect 25165 -575 25210 -455
rect 25330 -575 25375 -455
rect 25495 -575 25540 -455
rect 25660 -575 25715 -455
rect 25835 -575 25880 -455
rect 26000 -575 26045 -455
rect 26165 -575 26210 -455
rect 26330 -575 26385 -455
rect 26505 -575 26550 -455
rect 26670 -575 26715 -455
rect 26835 -575 26880 -455
rect 27000 -575 27055 -455
rect 27175 -575 27220 -455
rect 27340 -575 27385 -455
rect 27505 -575 27550 -455
rect 27670 -575 27725 -455
rect 27845 -575 27890 -455
rect 28010 -575 28055 -455
rect 28175 -575 28220 -455
rect 28340 -575 28395 -455
rect 28515 -575 28560 -455
rect 28680 -575 28725 -455
rect 28845 -575 28890 -455
rect 29010 -575 29065 -455
rect 29185 -575 29230 -455
rect 29350 -575 29395 -455
rect 29515 -575 29560 -455
rect 29680 -575 29690 -455
rect 24190 -630 29690 -575
rect 24190 -750 24200 -630
rect 24320 -750 24375 -630
rect 24495 -750 24540 -630
rect 24660 -750 24705 -630
rect 24825 -750 24870 -630
rect 24990 -750 25045 -630
rect 25165 -750 25210 -630
rect 25330 -750 25375 -630
rect 25495 -750 25540 -630
rect 25660 -750 25715 -630
rect 25835 -750 25880 -630
rect 26000 -750 26045 -630
rect 26165 -750 26210 -630
rect 26330 -750 26385 -630
rect 26505 -750 26550 -630
rect 26670 -750 26715 -630
rect 26835 -750 26880 -630
rect 27000 -750 27055 -630
rect 27175 -750 27220 -630
rect 27340 -750 27385 -630
rect 27505 -750 27550 -630
rect 27670 -750 27725 -630
rect 27845 -750 27890 -630
rect 28010 -750 28055 -630
rect 28175 -750 28220 -630
rect 28340 -750 28395 -630
rect 28515 -750 28560 -630
rect 28680 -750 28725 -630
rect 28845 -750 28890 -630
rect 29010 -750 29065 -630
rect 29185 -750 29230 -630
rect 29350 -750 29395 -630
rect 29515 -750 29560 -630
rect 29680 -750 29690 -630
rect 24190 -795 29690 -750
rect 24190 -915 24200 -795
rect 24320 -915 24375 -795
rect 24495 -915 24540 -795
rect 24660 -915 24705 -795
rect 24825 -915 24870 -795
rect 24990 -915 25045 -795
rect 25165 -915 25210 -795
rect 25330 -915 25375 -795
rect 25495 -915 25540 -795
rect 25660 -915 25715 -795
rect 25835 -915 25880 -795
rect 26000 -915 26045 -795
rect 26165 -915 26210 -795
rect 26330 -915 26385 -795
rect 26505 -915 26550 -795
rect 26670 -915 26715 -795
rect 26835 -915 26880 -795
rect 27000 -915 27055 -795
rect 27175 -915 27220 -795
rect 27340 -915 27385 -795
rect 27505 -915 27550 -795
rect 27670 -915 27725 -795
rect 27845 -915 27890 -795
rect 28010 -915 28055 -795
rect 28175 -915 28220 -795
rect 28340 -915 28395 -795
rect 28515 -915 28560 -795
rect 28680 -915 28725 -795
rect 28845 -915 28890 -795
rect 29010 -915 29065 -795
rect 29185 -915 29230 -795
rect 29350 -915 29395 -795
rect 29515 -915 29560 -795
rect 29680 -915 29690 -795
rect 24190 -960 29690 -915
rect 24190 -1080 24200 -960
rect 24320 -1080 24375 -960
rect 24495 -1080 24540 -960
rect 24660 -1080 24705 -960
rect 24825 -1080 24870 -960
rect 24990 -1080 25045 -960
rect 25165 -1080 25210 -960
rect 25330 -1080 25375 -960
rect 25495 -1080 25540 -960
rect 25660 -1080 25715 -960
rect 25835 -1080 25880 -960
rect 26000 -1080 26045 -960
rect 26165 -1080 26210 -960
rect 26330 -1080 26385 -960
rect 26505 -1080 26550 -960
rect 26670 -1080 26715 -960
rect 26835 -1080 26880 -960
rect 27000 -1080 27055 -960
rect 27175 -1080 27220 -960
rect 27340 -1080 27385 -960
rect 27505 -1080 27550 -960
rect 27670 -1080 27725 -960
rect 27845 -1080 27890 -960
rect 28010 -1080 28055 -960
rect 28175 -1080 28220 -960
rect 28340 -1080 28395 -960
rect 28515 -1080 28560 -960
rect 28680 -1080 28725 -960
rect 28845 -1080 28890 -960
rect 29010 -1080 29065 -960
rect 29185 -1080 29230 -960
rect 29350 -1080 29395 -960
rect 29515 -1080 29560 -960
rect 29680 -1080 29690 -960
rect 24190 -1125 29690 -1080
rect 24190 -1245 24200 -1125
rect 24320 -1245 24375 -1125
rect 24495 -1245 24540 -1125
rect 24660 -1245 24705 -1125
rect 24825 -1245 24870 -1125
rect 24990 -1245 25045 -1125
rect 25165 -1245 25210 -1125
rect 25330 -1245 25375 -1125
rect 25495 -1245 25540 -1125
rect 25660 -1245 25715 -1125
rect 25835 -1245 25880 -1125
rect 26000 -1245 26045 -1125
rect 26165 -1245 26210 -1125
rect 26330 -1245 26385 -1125
rect 26505 -1245 26550 -1125
rect 26670 -1245 26715 -1125
rect 26835 -1245 26880 -1125
rect 27000 -1245 27055 -1125
rect 27175 -1245 27220 -1125
rect 27340 -1245 27385 -1125
rect 27505 -1245 27550 -1125
rect 27670 -1245 27725 -1125
rect 27845 -1245 27890 -1125
rect 28010 -1245 28055 -1125
rect 28175 -1245 28220 -1125
rect 28340 -1245 28395 -1125
rect 28515 -1245 28560 -1125
rect 28680 -1245 28725 -1125
rect 28845 -1245 28890 -1125
rect 29010 -1245 29065 -1125
rect 29185 -1245 29230 -1125
rect 29350 -1245 29395 -1125
rect 29515 -1245 29560 -1125
rect 29680 -1245 29690 -1125
rect 24190 -1300 29690 -1245
rect 24190 -1420 24200 -1300
rect 24320 -1420 24375 -1300
rect 24495 -1420 24540 -1300
rect 24660 -1420 24705 -1300
rect 24825 -1420 24870 -1300
rect 24990 -1420 25045 -1300
rect 25165 -1420 25210 -1300
rect 25330 -1420 25375 -1300
rect 25495 -1420 25540 -1300
rect 25660 -1420 25715 -1300
rect 25835 -1420 25880 -1300
rect 26000 -1420 26045 -1300
rect 26165 -1420 26210 -1300
rect 26330 -1420 26385 -1300
rect 26505 -1420 26550 -1300
rect 26670 -1420 26715 -1300
rect 26835 -1420 26880 -1300
rect 27000 -1420 27055 -1300
rect 27175 -1420 27220 -1300
rect 27340 -1420 27385 -1300
rect 27505 -1420 27550 -1300
rect 27670 -1420 27725 -1300
rect 27845 -1420 27890 -1300
rect 28010 -1420 28055 -1300
rect 28175 -1420 28220 -1300
rect 28340 -1420 28395 -1300
rect 28515 -1420 28560 -1300
rect 28680 -1420 28725 -1300
rect 28845 -1420 28890 -1300
rect 29010 -1420 29065 -1300
rect 29185 -1420 29230 -1300
rect 29350 -1420 29395 -1300
rect 29515 -1420 29560 -1300
rect 29680 -1420 29690 -1300
rect 24190 -1465 29690 -1420
rect 24190 -1585 24200 -1465
rect 24320 -1585 24375 -1465
rect 24495 -1585 24540 -1465
rect 24660 -1585 24705 -1465
rect 24825 -1585 24870 -1465
rect 24990 -1585 25045 -1465
rect 25165 -1585 25210 -1465
rect 25330 -1585 25375 -1465
rect 25495 -1585 25540 -1465
rect 25660 -1585 25715 -1465
rect 25835 -1585 25880 -1465
rect 26000 -1585 26045 -1465
rect 26165 -1585 26210 -1465
rect 26330 -1585 26385 -1465
rect 26505 -1585 26550 -1465
rect 26670 -1585 26715 -1465
rect 26835 -1585 26880 -1465
rect 27000 -1585 27055 -1465
rect 27175 -1585 27220 -1465
rect 27340 -1585 27385 -1465
rect 27505 -1585 27550 -1465
rect 27670 -1585 27725 -1465
rect 27845 -1585 27890 -1465
rect 28010 -1585 28055 -1465
rect 28175 -1585 28220 -1465
rect 28340 -1585 28395 -1465
rect 28515 -1585 28560 -1465
rect 28680 -1585 28725 -1465
rect 28845 -1585 28890 -1465
rect 29010 -1585 29065 -1465
rect 29185 -1585 29230 -1465
rect 29350 -1585 29395 -1465
rect 29515 -1585 29560 -1465
rect 29680 -1585 29690 -1465
rect 24190 -1630 29690 -1585
rect 24190 -1750 24200 -1630
rect 24320 -1750 24375 -1630
rect 24495 -1750 24540 -1630
rect 24660 -1750 24705 -1630
rect 24825 -1750 24870 -1630
rect 24990 -1750 25045 -1630
rect 25165 -1750 25210 -1630
rect 25330 -1750 25375 -1630
rect 25495 -1750 25540 -1630
rect 25660 -1750 25715 -1630
rect 25835 -1750 25880 -1630
rect 26000 -1750 26045 -1630
rect 26165 -1750 26210 -1630
rect 26330 -1750 26385 -1630
rect 26505 -1750 26550 -1630
rect 26670 -1750 26715 -1630
rect 26835 -1750 26880 -1630
rect 27000 -1750 27055 -1630
rect 27175 -1750 27220 -1630
rect 27340 -1750 27385 -1630
rect 27505 -1750 27550 -1630
rect 27670 -1750 27725 -1630
rect 27845 -1750 27890 -1630
rect 28010 -1750 28055 -1630
rect 28175 -1750 28220 -1630
rect 28340 -1750 28395 -1630
rect 28515 -1750 28560 -1630
rect 28680 -1750 28725 -1630
rect 28845 -1750 28890 -1630
rect 29010 -1750 29065 -1630
rect 29185 -1750 29230 -1630
rect 29350 -1750 29395 -1630
rect 29515 -1750 29560 -1630
rect 29680 -1750 29690 -1630
rect 24190 -1795 29690 -1750
rect 24190 -1915 24200 -1795
rect 24320 -1915 24375 -1795
rect 24495 -1915 24540 -1795
rect 24660 -1915 24705 -1795
rect 24825 -1915 24870 -1795
rect 24990 -1915 25045 -1795
rect 25165 -1915 25210 -1795
rect 25330 -1915 25375 -1795
rect 25495 -1915 25540 -1795
rect 25660 -1915 25715 -1795
rect 25835 -1915 25880 -1795
rect 26000 -1915 26045 -1795
rect 26165 -1915 26210 -1795
rect 26330 -1915 26385 -1795
rect 26505 -1915 26550 -1795
rect 26670 -1915 26715 -1795
rect 26835 -1915 26880 -1795
rect 27000 -1915 27055 -1795
rect 27175 -1915 27220 -1795
rect 27340 -1915 27385 -1795
rect 27505 -1915 27550 -1795
rect 27670 -1915 27725 -1795
rect 27845 -1915 27890 -1795
rect 28010 -1915 28055 -1795
rect 28175 -1915 28220 -1795
rect 28340 -1915 28395 -1795
rect 28515 -1915 28560 -1795
rect 28680 -1915 28725 -1795
rect 28845 -1915 28890 -1795
rect 29010 -1915 29065 -1795
rect 29185 -1915 29230 -1795
rect 29350 -1915 29395 -1795
rect 29515 -1915 29560 -1795
rect 29680 -1915 29690 -1795
rect 24190 -1970 29690 -1915
rect 24190 -2090 24200 -1970
rect 24320 -2090 24375 -1970
rect 24495 -2090 24540 -1970
rect 24660 -2090 24705 -1970
rect 24825 -2090 24870 -1970
rect 24990 -2090 25045 -1970
rect 25165 -2090 25210 -1970
rect 25330 -2090 25375 -1970
rect 25495 -2090 25540 -1970
rect 25660 -2090 25715 -1970
rect 25835 -2090 25880 -1970
rect 26000 -2090 26045 -1970
rect 26165 -2090 26210 -1970
rect 26330 -2090 26385 -1970
rect 26505 -2090 26550 -1970
rect 26670 -2090 26715 -1970
rect 26835 -2090 26880 -1970
rect 27000 -2090 27055 -1970
rect 27175 -2090 27220 -1970
rect 27340 -2090 27385 -1970
rect 27505 -2090 27550 -1970
rect 27670 -2090 27725 -1970
rect 27845 -2090 27890 -1970
rect 28010 -2090 28055 -1970
rect 28175 -2090 28220 -1970
rect 28340 -2090 28395 -1970
rect 28515 -2090 28560 -1970
rect 28680 -2090 28725 -1970
rect 28845 -2090 28890 -1970
rect 29010 -2090 29065 -1970
rect 29185 -2090 29230 -1970
rect 29350 -2090 29395 -1970
rect 29515 -2090 29560 -1970
rect 29680 -2090 29690 -1970
rect 24190 -2135 29690 -2090
rect 24190 -2255 24200 -2135
rect 24320 -2255 24375 -2135
rect 24495 -2255 24540 -2135
rect 24660 -2255 24705 -2135
rect 24825 -2255 24870 -2135
rect 24990 -2255 25045 -2135
rect 25165 -2255 25210 -2135
rect 25330 -2255 25375 -2135
rect 25495 -2255 25540 -2135
rect 25660 -2255 25715 -2135
rect 25835 -2255 25880 -2135
rect 26000 -2255 26045 -2135
rect 26165 -2255 26210 -2135
rect 26330 -2255 26385 -2135
rect 26505 -2255 26550 -2135
rect 26670 -2255 26715 -2135
rect 26835 -2255 26880 -2135
rect 27000 -2255 27055 -2135
rect 27175 -2255 27220 -2135
rect 27340 -2255 27385 -2135
rect 27505 -2255 27550 -2135
rect 27670 -2255 27725 -2135
rect 27845 -2255 27890 -2135
rect 28010 -2255 28055 -2135
rect 28175 -2255 28220 -2135
rect 28340 -2255 28395 -2135
rect 28515 -2255 28560 -2135
rect 28680 -2255 28725 -2135
rect 28845 -2255 28890 -2135
rect 29010 -2255 29065 -2135
rect 29185 -2255 29230 -2135
rect 29350 -2255 29395 -2135
rect 29515 -2255 29560 -2135
rect 29680 -2255 29690 -2135
rect 24190 -2300 29690 -2255
rect 24190 -2420 24200 -2300
rect 24320 -2420 24375 -2300
rect 24495 -2420 24540 -2300
rect 24660 -2420 24705 -2300
rect 24825 -2420 24870 -2300
rect 24990 -2420 25045 -2300
rect 25165 -2420 25210 -2300
rect 25330 -2420 25375 -2300
rect 25495 -2420 25540 -2300
rect 25660 -2420 25715 -2300
rect 25835 -2420 25880 -2300
rect 26000 -2420 26045 -2300
rect 26165 -2420 26210 -2300
rect 26330 -2420 26385 -2300
rect 26505 -2420 26550 -2300
rect 26670 -2420 26715 -2300
rect 26835 -2420 26880 -2300
rect 27000 -2420 27055 -2300
rect 27175 -2420 27220 -2300
rect 27340 -2420 27385 -2300
rect 27505 -2420 27550 -2300
rect 27670 -2420 27725 -2300
rect 27845 -2420 27890 -2300
rect 28010 -2420 28055 -2300
rect 28175 -2420 28220 -2300
rect 28340 -2420 28395 -2300
rect 28515 -2420 28560 -2300
rect 28680 -2420 28725 -2300
rect 28845 -2420 28890 -2300
rect 29010 -2420 29065 -2300
rect 29185 -2420 29230 -2300
rect 29350 -2420 29395 -2300
rect 29515 -2420 29560 -2300
rect 29680 -2420 29690 -2300
rect 24190 -2465 29690 -2420
rect 24190 -2585 24200 -2465
rect 24320 -2585 24375 -2465
rect 24495 -2585 24540 -2465
rect 24660 -2585 24705 -2465
rect 24825 -2585 24870 -2465
rect 24990 -2585 25045 -2465
rect 25165 -2585 25210 -2465
rect 25330 -2585 25375 -2465
rect 25495 -2585 25540 -2465
rect 25660 -2585 25715 -2465
rect 25835 -2585 25880 -2465
rect 26000 -2585 26045 -2465
rect 26165 -2585 26210 -2465
rect 26330 -2585 26385 -2465
rect 26505 -2585 26550 -2465
rect 26670 -2585 26715 -2465
rect 26835 -2585 26880 -2465
rect 27000 -2585 27055 -2465
rect 27175 -2585 27220 -2465
rect 27340 -2585 27385 -2465
rect 27505 -2585 27550 -2465
rect 27670 -2585 27725 -2465
rect 27845 -2585 27890 -2465
rect 28010 -2585 28055 -2465
rect 28175 -2585 28220 -2465
rect 28340 -2585 28395 -2465
rect 28515 -2585 28560 -2465
rect 28680 -2585 28725 -2465
rect 28845 -2585 28890 -2465
rect 29010 -2585 29065 -2465
rect 29185 -2585 29230 -2465
rect 29350 -2585 29395 -2465
rect 29515 -2585 29560 -2465
rect 29680 -2585 29690 -2465
rect 24190 -2640 29690 -2585
rect 24190 -2760 24200 -2640
rect 24320 -2760 24375 -2640
rect 24495 -2760 24540 -2640
rect 24660 -2760 24705 -2640
rect 24825 -2760 24870 -2640
rect 24990 -2760 25045 -2640
rect 25165 -2760 25210 -2640
rect 25330 -2760 25375 -2640
rect 25495 -2760 25540 -2640
rect 25660 -2760 25715 -2640
rect 25835 -2760 25880 -2640
rect 26000 -2760 26045 -2640
rect 26165 -2760 26210 -2640
rect 26330 -2760 26385 -2640
rect 26505 -2760 26550 -2640
rect 26670 -2760 26715 -2640
rect 26835 -2760 26880 -2640
rect 27000 -2760 27055 -2640
rect 27175 -2760 27220 -2640
rect 27340 -2760 27385 -2640
rect 27505 -2760 27550 -2640
rect 27670 -2760 27725 -2640
rect 27845 -2760 27890 -2640
rect 28010 -2760 28055 -2640
rect 28175 -2760 28220 -2640
rect 28340 -2760 28395 -2640
rect 28515 -2760 28560 -2640
rect 28680 -2760 28725 -2640
rect 28845 -2760 28890 -2640
rect 29010 -2760 29065 -2640
rect 29185 -2760 29230 -2640
rect 29350 -2760 29395 -2640
rect 29515 -2760 29560 -2640
rect 29680 -2760 29690 -2640
rect 24190 -2805 29690 -2760
rect 24190 -2925 24200 -2805
rect 24320 -2925 24375 -2805
rect 24495 -2925 24540 -2805
rect 24660 -2925 24705 -2805
rect 24825 -2925 24870 -2805
rect 24990 -2925 25045 -2805
rect 25165 -2925 25210 -2805
rect 25330 -2925 25375 -2805
rect 25495 -2925 25540 -2805
rect 25660 -2925 25715 -2805
rect 25835 -2925 25880 -2805
rect 26000 -2925 26045 -2805
rect 26165 -2925 26210 -2805
rect 26330 -2925 26385 -2805
rect 26505 -2925 26550 -2805
rect 26670 -2925 26715 -2805
rect 26835 -2925 26880 -2805
rect 27000 -2925 27055 -2805
rect 27175 -2925 27220 -2805
rect 27340 -2925 27385 -2805
rect 27505 -2925 27550 -2805
rect 27670 -2925 27725 -2805
rect 27845 -2925 27890 -2805
rect 28010 -2925 28055 -2805
rect 28175 -2925 28220 -2805
rect 28340 -2925 28395 -2805
rect 28515 -2925 28560 -2805
rect 28680 -2925 28725 -2805
rect 28845 -2925 28890 -2805
rect 29010 -2925 29065 -2805
rect 29185 -2925 29230 -2805
rect 29350 -2925 29395 -2805
rect 29515 -2925 29560 -2805
rect 29680 -2925 29690 -2805
rect 24190 -2970 29690 -2925
rect 24190 -3090 24200 -2970
rect 24320 -3090 24375 -2970
rect 24495 -3090 24540 -2970
rect 24660 -3090 24705 -2970
rect 24825 -3090 24870 -2970
rect 24990 -3090 25045 -2970
rect 25165 -3090 25210 -2970
rect 25330 -3090 25375 -2970
rect 25495 -3090 25540 -2970
rect 25660 -3090 25715 -2970
rect 25835 -3090 25880 -2970
rect 26000 -3090 26045 -2970
rect 26165 -3090 26210 -2970
rect 26330 -3090 26385 -2970
rect 26505 -3090 26550 -2970
rect 26670 -3090 26715 -2970
rect 26835 -3090 26880 -2970
rect 27000 -3090 27055 -2970
rect 27175 -3090 27220 -2970
rect 27340 -3090 27385 -2970
rect 27505 -3090 27550 -2970
rect 27670 -3090 27725 -2970
rect 27845 -3090 27890 -2970
rect 28010 -3090 28055 -2970
rect 28175 -3090 28220 -2970
rect 28340 -3090 28395 -2970
rect 28515 -3090 28560 -2970
rect 28680 -3090 28725 -2970
rect 28845 -3090 28890 -2970
rect 29010 -3090 29065 -2970
rect 29185 -3090 29230 -2970
rect 29350 -3090 29395 -2970
rect 29515 -3090 29560 -2970
rect 29680 -3090 29690 -2970
rect 24190 -3135 29690 -3090
rect 24190 -3255 24200 -3135
rect 24320 -3255 24375 -3135
rect 24495 -3255 24540 -3135
rect 24660 -3255 24705 -3135
rect 24825 -3255 24870 -3135
rect 24990 -3255 25045 -3135
rect 25165 -3255 25210 -3135
rect 25330 -3255 25375 -3135
rect 25495 -3255 25540 -3135
rect 25660 -3255 25715 -3135
rect 25835 -3255 25880 -3135
rect 26000 -3255 26045 -3135
rect 26165 -3255 26210 -3135
rect 26330 -3255 26385 -3135
rect 26505 -3255 26550 -3135
rect 26670 -3255 26715 -3135
rect 26835 -3255 26880 -3135
rect 27000 -3255 27055 -3135
rect 27175 -3255 27220 -3135
rect 27340 -3255 27385 -3135
rect 27505 -3255 27550 -3135
rect 27670 -3255 27725 -3135
rect 27845 -3255 27890 -3135
rect 28010 -3255 28055 -3135
rect 28175 -3255 28220 -3135
rect 28340 -3255 28395 -3135
rect 28515 -3255 28560 -3135
rect 28680 -3255 28725 -3135
rect 28845 -3255 28890 -3135
rect 29010 -3255 29065 -3135
rect 29185 -3255 29230 -3135
rect 29350 -3255 29395 -3135
rect 29515 -3255 29560 -3135
rect 29680 -3255 29690 -3135
rect 24190 -3310 29690 -3255
rect 24190 -3430 24200 -3310
rect 24320 -3430 24375 -3310
rect 24495 -3430 24540 -3310
rect 24660 -3430 24705 -3310
rect 24825 -3430 24870 -3310
rect 24990 -3430 25045 -3310
rect 25165 -3430 25210 -3310
rect 25330 -3430 25375 -3310
rect 25495 -3430 25540 -3310
rect 25660 -3430 25715 -3310
rect 25835 -3430 25880 -3310
rect 26000 -3430 26045 -3310
rect 26165 -3430 26210 -3310
rect 26330 -3430 26385 -3310
rect 26505 -3430 26550 -3310
rect 26670 -3430 26715 -3310
rect 26835 -3430 26880 -3310
rect 27000 -3430 27055 -3310
rect 27175 -3430 27220 -3310
rect 27340 -3430 27385 -3310
rect 27505 -3430 27550 -3310
rect 27670 -3430 27725 -3310
rect 27845 -3430 27890 -3310
rect 28010 -3430 28055 -3310
rect 28175 -3430 28220 -3310
rect 28340 -3430 28395 -3310
rect 28515 -3430 28560 -3310
rect 28680 -3430 28725 -3310
rect 28845 -3430 28890 -3310
rect 29010 -3430 29065 -3310
rect 29185 -3430 29230 -3310
rect 29350 -3430 29395 -3310
rect 29515 -3430 29560 -3310
rect 29680 -3430 29690 -3310
rect 24190 -3475 29690 -3430
rect 24190 -3595 24200 -3475
rect 24320 -3595 24375 -3475
rect 24495 -3595 24540 -3475
rect 24660 -3595 24705 -3475
rect 24825 -3595 24870 -3475
rect 24990 -3595 25045 -3475
rect 25165 -3595 25210 -3475
rect 25330 -3595 25375 -3475
rect 25495 -3595 25540 -3475
rect 25660 -3595 25715 -3475
rect 25835 -3595 25880 -3475
rect 26000 -3595 26045 -3475
rect 26165 -3595 26210 -3475
rect 26330 -3595 26385 -3475
rect 26505 -3595 26550 -3475
rect 26670 -3595 26715 -3475
rect 26835 -3595 26880 -3475
rect 27000 -3595 27055 -3475
rect 27175 -3595 27220 -3475
rect 27340 -3595 27385 -3475
rect 27505 -3595 27550 -3475
rect 27670 -3595 27725 -3475
rect 27845 -3595 27890 -3475
rect 28010 -3595 28055 -3475
rect 28175 -3595 28220 -3475
rect 28340 -3595 28395 -3475
rect 28515 -3595 28560 -3475
rect 28680 -3595 28725 -3475
rect 28845 -3595 28890 -3475
rect 29010 -3595 29065 -3475
rect 29185 -3595 29230 -3475
rect 29350 -3595 29395 -3475
rect 29515 -3595 29560 -3475
rect 29680 -3595 29690 -3475
rect 24190 -3640 29690 -3595
rect 24190 -3760 24200 -3640
rect 24320 -3760 24375 -3640
rect 24495 -3760 24540 -3640
rect 24660 -3760 24705 -3640
rect 24825 -3760 24870 -3640
rect 24990 -3760 25045 -3640
rect 25165 -3760 25210 -3640
rect 25330 -3760 25375 -3640
rect 25495 -3760 25540 -3640
rect 25660 -3760 25715 -3640
rect 25835 -3760 25880 -3640
rect 26000 -3760 26045 -3640
rect 26165 -3760 26210 -3640
rect 26330 -3760 26385 -3640
rect 26505 -3760 26550 -3640
rect 26670 -3760 26715 -3640
rect 26835 -3760 26880 -3640
rect 27000 -3760 27055 -3640
rect 27175 -3760 27220 -3640
rect 27340 -3760 27385 -3640
rect 27505 -3760 27550 -3640
rect 27670 -3760 27725 -3640
rect 27845 -3760 27890 -3640
rect 28010 -3760 28055 -3640
rect 28175 -3760 28220 -3640
rect 28340 -3760 28395 -3640
rect 28515 -3760 28560 -3640
rect 28680 -3760 28725 -3640
rect 28845 -3760 28890 -3640
rect 29010 -3760 29065 -3640
rect 29185 -3760 29230 -3640
rect 29350 -3760 29395 -3640
rect 29515 -3760 29560 -3640
rect 29680 -3760 29690 -3640
rect 24190 -3805 29690 -3760
rect 24190 -3925 24200 -3805
rect 24320 -3925 24375 -3805
rect 24495 -3925 24540 -3805
rect 24660 -3925 24705 -3805
rect 24825 -3925 24870 -3805
rect 24990 -3925 25045 -3805
rect 25165 -3925 25210 -3805
rect 25330 -3925 25375 -3805
rect 25495 -3925 25540 -3805
rect 25660 -3925 25715 -3805
rect 25835 -3925 25880 -3805
rect 26000 -3925 26045 -3805
rect 26165 -3925 26210 -3805
rect 26330 -3925 26385 -3805
rect 26505 -3925 26550 -3805
rect 26670 -3925 26715 -3805
rect 26835 -3925 26880 -3805
rect 27000 -3925 27055 -3805
rect 27175 -3925 27220 -3805
rect 27340 -3925 27385 -3805
rect 27505 -3925 27550 -3805
rect 27670 -3925 27725 -3805
rect 27845 -3925 27890 -3805
rect 28010 -3925 28055 -3805
rect 28175 -3925 28220 -3805
rect 28340 -3925 28395 -3805
rect 28515 -3925 28560 -3805
rect 28680 -3925 28725 -3805
rect 28845 -3925 28890 -3805
rect 29010 -3925 29065 -3805
rect 29185 -3925 29230 -3805
rect 29350 -3925 29395 -3805
rect 29515 -3925 29560 -3805
rect 29680 -3925 29690 -3805
rect 24190 -3980 29690 -3925
rect 24190 -4100 24200 -3980
rect 24320 -4100 24375 -3980
rect 24495 -4100 24540 -3980
rect 24660 -4100 24705 -3980
rect 24825 -4100 24870 -3980
rect 24990 -4100 25045 -3980
rect 25165 -4100 25210 -3980
rect 25330 -4100 25375 -3980
rect 25495 -4100 25540 -3980
rect 25660 -4100 25715 -3980
rect 25835 -4100 25880 -3980
rect 26000 -4100 26045 -3980
rect 26165 -4100 26210 -3980
rect 26330 -4100 26385 -3980
rect 26505 -4100 26550 -3980
rect 26670 -4100 26715 -3980
rect 26835 -4100 26880 -3980
rect 27000 -4100 27055 -3980
rect 27175 -4100 27220 -3980
rect 27340 -4100 27385 -3980
rect 27505 -4100 27550 -3980
rect 27670 -4100 27725 -3980
rect 27845 -4100 27890 -3980
rect 28010 -4100 28055 -3980
rect 28175 -4100 28220 -3980
rect 28340 -4100 28395 -3980
rect 28515 -4100 28560 -3980
rect 28680 -4100 28725 -3980
rect 28845 -4100 28890 -3980
rect 29010 -4100 29065 -3980
rect 29185 -4100 29230 -3980
rect 29350 -4100 29395 -3980
rect 29515 -4100 29560 -3980
rect 29680 -4100 29690 -3980
rect 24190 -4110 29690 -4100
rect 7120 -4310 12620 -4300
rect 7120 -4430 7130 -4310
rect 7250 -4430 7295 -4310
rect 7415 -4430 7460 -4310
rect 7580 -4430 7625 -4310
rect 7745 -4430 7800 -4310
rect 7920 -4430 7965 -4310
rect 8085 -4430 8130 -4310
rect 8250 -4430 8295 -4310
rect 8415 -4430 8470 -4310
rect 8590 -4430 8635 -4310
rect 8755 -4430 8800 -4310
rect 8920 -4430 8965 -4310
rect 9085 -4430 9140 -4310
rect 9260 -4430 9305 -4310
rect 9425 -4430 9470 -4310
rect 9590 -4430 9635 -4310
rect 9755 -4430 9810 -4310
rect 9930 -4430 9975 -4310
rect 10095 -4430 10140 -4310
rect 10260 -4430 10305 -4310
rect 10425 -4430 10480 -4310
rect 10600 -4430 10645 -4310
rect 10765 -4430 10810 -4310
rect 10930 -4430 10975 -4310
rect 11095 -4430 11150 -4310
rect 11270 -4430 11315 -4310
rect 11435 -4430 11480 -4310
rect 11600 -4430 11645 -4310
rect 11765 -4430 11820 -4310
rect 11940 -4430 11985 -4310
rect 12105 -4430 12150 -4310
rect 12270 -4430 12315 -4310
rect 12435 -4430 12490 -4310
rect 12610 -4430 12620 -4310
rect 7120 -4485 12620 -4430
rect 7120 -4605 7130 -4485
rect 7250 -4605 7295 -4485
rect 7415 -4605 7460 -4485
rect 7580 -4605 7625 -4485
rect 7745 -4605 7800 -4485
rect 7920 -4605 7965 -4485
rect 8085 -4605 8130 -4485
rect 8250 -4605 8295 -4485
rect 8415 -4605 8470 -4485
rect 8590 -4605 8635 -4485
rect 8755 -4605 8800 -4485
rect 8920 -4605 8965 -4485
rect 9085 -4605 9140 -4485
rect 9260 -4605 9305 -4485
rect 9425 -4605 9470 -4485
rect 9590 -4605 9635 -4485
rect 9755 -4605 9810 -4485
rect 9930 -4605 9975 -4485
rect 10095 -4605 10140 -4485
rect 10260 -4605 10305 -4485
rect 10425 -4605 10480 -4485
rect 10600 -4605 10645 -4485
rect 10765 -4605 10810 -4485
rect 10930 -4605 10975 -4485
rect 11095 -4605 11150 -4485
rect 11270 -4605 11315 -4485
rect 11435 -4605 11480 -4485
rect 11600 -4605 11645 -4485
rect 11765 -4605 11820 -4485
rect 11940 -4605 11985 -4485
rect 12105 -4605 12150 -4485
rect 12270 -4605 12315 -4485
rect 12435 -4605 12490 -4485
rect 12610 -4605 12620 -4485
rect 7120 -4650 12620 -4605
rect 7120 -4770 7130 -4650
rect 7250 -4770 7295 -4650
rect 7415 -4770 7460 -4650
rect 7580 -4770 7625 -4650
rect 7745 -4770 7800 -4650
rect 7920 -4770 7965 -4650
rect 8085 -4770 8130 -4650
rect 8250 -4770 8295 -4650
rect 8415 -4770 8470 -4650
rect 8590 -4770 8635 -4650
rect 8755 -4770 8800 -4650
rect 8920 -4770 8965 -4650
rect 9085 -4770 9140 -4650
rect 9260 -4770 9305 -4650
rect 9425 -4770 9470 -4650
rect 9590 -4770 9635 -4650
rect 9755 -4770 9810 -4650
rect 9930 -4770 9975 -4650
rect 10095 -4770 10140 -4650
rect 10260 -4770 10305 -4650
rect 10425 -4770 10480 -4650
rect 10600 -4770 10645 -4650
rect 10765 -4770 10810 -4650
rect 10930 -4770 10975 -4650
rect 11095 -4770 11150 -4650
rect 11270 -4770 11315 -4650
rect 11435 -4770 11480 -4650
rect 11600 -4770 11645 -4650
rect 11765 -4770 11820 -4650
rect 11940 -4770 11985 -4650
rect 12105 -4770 12150 -4650
rect 12270 -4770 12315 -4650
rect 12435 -4770 12490 -4650
rect 12610 -4770 12620 -4650
rect 7120 -4815 12620 -4770
rect 7120 -4935 7130 -4815
rect 7250 -4935 7295 -4815
rect 7415 -4935 7460 -4815
rect 7580 -4935 7625 -4815
rect 7745 -4935 7800 -4815
rect 7920 -4935 7965 -4815
rect 8085 -4935 8130 -4815
rect 8250 -4935 8295 -4815
rect 8415 -4935 8470 -4815
rect 8590 -4935 8635 -4815
rect 8755 -4935 8800 -4815
rect 8920 -4935 8965 -4815
rect 9085 -4935 9140 -4815
rect 9260 -4935 9305 -4815
rect 9425 -4935 9470 -4815
rect 9590 -4935 9635 -4815
rect 9755 -4935 9810 -4815
rect 9930 -4935 9975 -4815
rect 10095 -4935 10140 -4815
rect 10260 -4935 10305 -4815
rect 10425 -4935 10480 -4815
rect 10600 -4935 10645 -4815
rect 10765 -4935 10810 -4815
rect 10930 -4935 10975 -4815
rect 11095 -4935 11150 -4815
rect 11270 -4935 11315 -4815
rect 11435 -4935 11480 -4815
rect 11600 -4935 11645 -4815
rect 11765 -4935 11820 -4815
rect 11940 -4935 11985 -4815
rect 12105 -4935 12150 -4815
rect 12270 -4935 12315 -4815
rect 12435 -4935 12490 -4815
rect 12610 -4935 12620 -4815
rect 7120 -4980 12620 -4935
rect 7120 -5100 7130 -4980
rect 7250 -5100 7295 -4980
rect 7415 -5100 7460 -4980
rect 7580 -5100 7625 -4980
rect 7745 -5100 7800 -4980
rect 7920 -5100 7965 -4980
rect 8085 -5100 8130 -4980
rect 8250 -5100 8295 -4980
rect 8415 -5100 8470 -4980
rect 8590 -5100 8635 -4980
rect 8755 -5100 8800 -4980
rect 8920 -5100 8965 -4980
rect 9085 -5100 9140 -4980
rect 9260 -5100 9305 -4980
rect 9425 -5100 9470 -4980
rect 9590 -5100 9635 -4980
rect 9755 -5100 9810 -4980
rect 9930 -5100 9975 -4980
rect 10095 -5100 10140 -4980
rect 10260 -5100 10305 -4980
rect 10425 -5100 10480 -4980
rect 10600 -5100 10645 -4980
rect 10765 -5100 10810 -4980
rect 10930 -5100 10975 -4980
rect 11095 -5100 11150 -4980
rect 11270 -5100 11315 -4980
rect 11435 -5100 11480 -4980
rect 11600 -5100 11645 -4980
rect 11765 -5100 11820 -4980
rect 11940 -5100 11985 -4980
rect 12105 -5100 12150 -4980
rect 12270 -5100 12315 -4980
rect 12435 -5100 12490 -4980
rect 12610 -5100 12620 -4980
rect 7120 -5155 12620 -5100
rect 7120 -5275 7130 -5155
rect 7250 -5275 7295 -5155
rect 7415 -5275 7460 -5155
rect 7580 -5275 7625 -5155
rect 7745 -5275 7800 -5155
rect 7920 -5275 7965 -5155
rect 8085 -5275 8130 -5155
rect 8250 -5275 8295 -5155
rect 8415 -5275 8470 -5155
rect 8590 -5275 8635 -5155
rect 8755 -5275 8800 -5155
rect 8920 -5275 8965 -5155
rect 9085 -5275 9140 -5155
rect 9260 -5275 9305 -5155
rect 9425 -5275 9470 -5155
rect 9590 -5275 9635 -5155
rect 9755 -5275 9810 -5155
rect 9930 -5275 9975 -5155
rect 10095 -5275 10140 -5155
rect 10260 -5275 10305 -5155
rect 10425 -5275 10480 -5155
rect 10600 -5275 10645 -5155
rect 10765 -5275 10810 -5155
rect 10930 -5275 10975 -5155
rect 11095 -5275 11150 -5155
rect 11270 -5275 11315 -5155
rect 11435 -5275 11480 -5155
rect 11600 -5275 11645 -5155
rect 11765 -5275 11820 -5155
rect 11940 -5275 11985 -5155
rect 12105 -5275 12150 -5155
rect 12270 -5275 12315 -5155
rect 12435 -5275 12490 -5155
rect 12610 -5275 12620 -5155
rect 7120 -5320 12620 -5275
rect 7120 -5440 7130 -5320
rect 7250 -5440 7295 -5320
rect 7415 -5440 7460 -5320
rect 7580 -5440 7625 -5320
rect 7745 -5440 7800 -5320
rect 7920 -5440 7965 -5320
rect 8085 -5440 8130 -5320
rect 8250 -5440 8295 -5320
rect 8415 -5440 8470 -5320
rect 8590 -5440 8635 -5320
rect 8755 -5440 8800 -5320
rect 8920 -5440 8965 -5320
rect 9085 -5440 9140 -5320
rect 9260 -5440 9305 -5320
rect 9425 -5440 9470 -5320
rect 9590 -5440 9635 -5320
rect 9755 -5440 9810 -5320
rect 9930 -5440 9975 -5320
rect 10095 -5440 10140 -5320
rect 10260 -5440 10305 -5320
rect 10425 -5440 10480 -5320
rect 10600 -5440 10645 -5320
rect 10765 -5440 10810 -5320
rect 10930 -5440 10975 -5320
rect 11095 -5440 11150 -5320
rect 11270 -5440 11315 -5320
rect 11435 -5440 11480 -5320
rect 11600 -5440 11645 -5320
rect 11765 -5440 11820 -5320
rect 11940 -5440 11985 -5320
rect 12105 -5440 12150 -5320
rect 12270 -5440 12315 -5320
rect 12435 -5440 12490 -5320
rect 12610 -5440 12620 -5320
rect 7120 -5485 12620 -5440
rect 7120 -5605 7130 -5485
rect 7250 -5605 7295 -5485
rect 7415 -5605 7460 -5485
rect 7580 -5605 7625 -5485
rect 7745 -5605 7800 -5485
rect 7920 -5605 7965 -5485
rect 8085 -5605 8130 -5485
rect 8250 -5605 8295 -5485
rect 8415 -5605 8470 -5485
rect 8590 -5605 8635 -5485
rect 8755 -5605 8800 -5485
rect 8920 -5605 8965 -5485
rect 9085 -5605 9140 -5485
rect 9260 -5605 9305 -5485
rect 9425 -5605 9470 -5485
rect 9590 -5605 9635 -5485
rect 9755 -5605 9810 -5485
rect 9930 -5605 9975 -5485
rect 10095 -5605 10140 -5485
rect 10260 -5605 10305 -5485
rect 10425 -5605 10480 -5485
rect 10600 -5605 10645 -5485
rect 10765 -5605 10810 -5485
rect 10930 -5605 10975 -5485
rect 11095 -5605 11150 -5485
rect 11270 -5605 11315 -5485
rect 11435 -5605 11480 -5485
rect 11600 -5605 11645 -5485
rect 11765 -5605 11820 -5485
rect 11940 -5605 11985 -5485
rect 12105 -5605 12150 -5485
rect 12270 -5605 12315 -5485
rect 12435 -5605 12490 -5485
rect 12610 -5605 12620 -5485
rect 7120 -5650 12620 -5605
rect 7120 -5770 7130 -5650
rect 7250 -5770 7295 -5650
rect 7415 -5770 7460 -5650
rect 7580 -5770 7625 -5650
rect 7745 -5770 7800 -5650
rect 7920 -5770 7965 -5650
rect 8085 -5770 8130 -5650
rect 8250 -5770 8295 -5650
rect 8415 -5770 8470 -5650
rect 8590 -5770 8635 -5650
rect 8755 -5770 8800 -5650
rect 8920 -5770 8965 -5650
rect 9085 -5770 9140 -5650
rect 9260 -5770 9305 -5650
rect 9425 -5770 9470 -5650
rect 9590 -5770 9635 -5650
rect 9755 -5770 9810 -5650
rect 9930 -5770 9975 -5650
rect 10095 -5770 10140 -5650
rect 10260 -5770 10305 -5650
rect 10425 -5770 10480 -5650
rect 10600 -5770 10645 -5650
rect 10765 -5770 10810 -5650
rect 10930 -5770 10975 -5650
rect 11095 -5770 11150 -5650
rect 11270 -5770 11315 -5650
rect 11435 -5770 11480 -5650
rect 11600 -5770 11645 -5650
rect 11765 -5770 11820 -5650
rect 11940 -5770 11985 -5650
rect 12105 -5770 12150 -5650
rect 12270 -5770 12315 -5650
rect 12435 -5770 12490 -5650
rect 12610 -5770 12620 -5650
rect 7120 -5825 12620 -5770
rect 7120 -5945 7130 -5825
rect 7250 -5945 7295 -5825
rect 7415 -5945 7460 -5825
rect 7580 -5945 7625 -5825
rect 7745 -5945 7800 -5825
rect 7920 -5945 7965 -5825
rect 8085 -5945 8130 -5825
rect 8250 -5945 8295 -5825
rect 8415 -5945 8470 -5825
rect 8590 -5945 8635 -5825
rect 8755 -5945 8800 -5825
rect 8920 -5945 8965 -5825
rect 9085 -5945 9140 -5825
rect 9260 -5945 9305 -5825
rect 9425 -5945 9470 -5825
rect 9590 -5945 9635 -5825
rect 9755 -5945 9810 -5825
rect 9930 -5945 9975 -5825
rect 10095 -5945 10140 -5825
rect 10260 -5945 10305 -5825
rect 10425 -5945 10480 -5825
rect 10600 -5945 10645 -5825
rect 10765 -5945 10810 -5825
rect 10930 -5945 10975 -5825
rect 11095 -5945 11150 -5825
rect 11270 -5945 11315 -5825
rect 11435 -5945 11480 -5825
rect 11600 -5945 11645 -5825
rect 11765 -5945 11820 -5825
rect 11940 -5945 11985 -5825
rect 12105 -5945 12150 -5825
rect 12270 -5945 12315 -5825
rect 12435 -5945 12490 -5825
rect 12610 -5945 12620 -5825
rect 7120 -5990 12620 -5945
rect 7120 -6110 7130 -5990
rect 7250 -6110 7295 -5990
rect 7415 -6110 7460 -5990
rect 7580 -6110 7625 -5990
rect 7745 -6110 7800 -5990
rect 7920 -6110 7965 -5990
rect 8085 -6110 8130 -5990
rect 8250 -6110 8295 -5990
rect 8415 -6110 8470 -5990
rect 8590 -6110 8635 -5990
rect 8755 -6110 8800 -5990
rect 8920 -6110 8965 -5990
rect 9085 -6110 9140 -5990
rect 9260 -6110 9305 -5990
rect 9425 -6110 9470 -5990
rect 9590 -6110 9635 -5990
rect 9755 -6110 9810 -5990
rect 9930 -6110 9975 -5990
rect 10095 -6110 10140 -5990
rect 10260 -6110 10305 -5990
rect 10425 -6110 10480 -5990
rect 10600 -6110 10645 -5990
rect 10765 -6110 10810 -5990
rect 10930 -6110 10975 -5990
rect 11095 -6110 11150 -5990
rect 11270 -6110 11315 -5990
rect 11435 -6110 11480 -5990
rect 11600 -6110 11645 -5990
rect 11765 -6110 11820 -5990
rect 11940 -6110 11985 -5990
rect 12105 -6110 12150 -5990
rect 12270 -6110 12315 -5990
rect 12435 -6110 12490 -5990
rect 12610 -6110 12620 -5990
rect 7120 -6155 12620 -6110
rect 7120 -6275 7130 -6155
rect 7250 -6275 7295 -6155
rect 7415 -6275 7460 -6155
rect 7580 -6275 7625 -6155
rect 7745 -6275 7800 -6155
rect 7920 -6275 7965 -6155
rect 8085 -6275 8130 -6155
rect 8250 -6275 8295 -6155
rect 8415 -6275 8470 -6155
rect 8590 -6275 8635 -6155
rect 8755 -6275 8800 -6155
rect 8920 -6275 8965 -6155
rect 9085 -6275 9140 -6155
rect 9260 -6275 9305 -6155
rect 9425 -6275 9470 -6155
rect 9590 -6275 9635 -6155
rect 9755 -6275 9810 -6155
rect 9930 -6275 9975 -6155
rect 10095 -6275 10140 -6155
rect 10260 -6275 10305 -6155
rect 10425 -6275 10480 -6155
rect 10600 -6275 10645 -6155
rect 10765 -6275 10810 -6155
rect 10930 -6275 10975 -6155
rect 11095 -6275 11150 -6155
rect 11270 -6275 11315 -6155
rect 11435 -6275 11480 -6155
rect 11600 -6275 11645 -6155
rect 11765 -6275 11820 -6155
rect 11940 -6275 11985 -6155
rect 12105 -6275 12150 -6155
rect 12270 -6275 12315 -6155
rect 12435 -6275 12490 -6155
rect 12610 -6275 12620 -6155
rect 7120 -6320 12620 -6275
rect 7120 -6440 7130 -6320
rect 7250 -6440 7295 -6320
rect 7415 -6440 7460 -6320
rect 7580 -6440 7625 -6320
rect 7745 -6440 7800 -6320
rect 7920 -6440 7965 -6320
rect 8085 -6440 8130 -6320
rect 8250 -6440 8295 -6320
rect 8415 -6440 8470 -6320
rect 8590 -6440 8635 -6320
rect 8755 -6440 8800 -6320
rect 8920 -6440 8965 -6320
rect 9085 -6440 9140 -6320
rect 9260 -6440 9305 -6320
rect 9425 -6440 9470 -6320
rect 9590 -6440 9635 -6320
rect 9755 -6440 9810 -6320
rect 9930 -6440 9975 -6320
rect 10095 -6440 10140 -6320
rect 10260 -6440 10305 -6320
rect 10425 -6440 10480 -6320
rect 10600 -6440 10645 -6320
rect 10765 -6440 10810 -6320
rect 10930 -6440 10975 -6320
rect 11095 -6440 11150 -6320
rect 11270 -6440 11315 -6320
rect 11435 -6440 11480 -6320
rect 11600 -6440 11645 -6320
rect 11765 -6440 11820 -6320
rect 11940 -6440 11985 -6320
rect 12105 -6440 12150 -6320
rect 12270 -6440 12315 -6320
rect 12435 -6440 12490 -6320
rect 12610 -6440 12620 -6320
rect 7120 -6495 12620 -6440
rect 7120 -6615 7130 -6495
rect 7250 -6615 7295 -6495
rect 7415 -6615 7460 -6495
rect 7580 -6615 7625 -6495
rect 7745 -6615 7800 -6495
rect 7920 -6615 7965 -6495
rect 8085 -6615 8130 -6495
rect 8250 -6615 8295 -6495
rect 8415 -6615 8470 -6495
rect 8590 -6615 8635 -6495
rect 8755 -6615 8800 -6495
rect 8920 -6615 8965 -6495
rect 9085 -6615 9140 -6495
rect 9260 -6615 9305 -6495
rect 9425 -6615 9470 -6495
rect 9590 -6615 9635 -6495
rect 9755 -6615 9810 -6495
rect 9930 -6615 9975 -6495
rect 10095 -6615 10140 -6495
rect 10260 -6615 10305 -6495
rect 10425 -6615 10480 -6495
rect 10600 -6615 10645 -6495
rect 10765 -6615 10810 -6495
rect 10930 -6615 10975 -6495
rect 11095 -6615 11150 -6495
rect 11270 -6615 11315 -6495
rect 11435 -6615 11480 -6495
rect 11600 -6615 11645 -6495
rect 11765 -6615 11820 -6495
rect 11940 -6615 11985 -6495
rect 12105 -6615 12150 -6495
rect 12270 -6615 12315 -6495
rect 12435 -6615 12490 -6495
rect 12610 -6615 12620 -6495
rect 7120 -6660 12620 -6615
rect 7120 -6780 7130 -6660
rect 7250 -6780 7295 -6660
rect 7415 -6780 7460 -6660
rect 7580 -6780 7625 -6660
rect 7745 -6780 7800 -6660
rect 7920 -6780 7965 -6660
rect 8085 -6780 8130 -6660
rect 8250 -6780 8295 -6660
rect 8415 -6780 8470 -6660
rect 8590 -6780 8635 -6660
rect 8755 -6780 8800 -6660
rect 8920 -6780 8965 -6660
rect 9085 -6780 9140 -6660
rect 9260 -6780 9305 -6660
rect 9425 -6780 9470 -6660
rect 9590 -6780 9635 -6660
rect 9755 -6780 9810 -6660
rect 9930 -6780 9975 -6660
rect 10095 -6780 10140 -6660
rect 10260 -6780 10305 -6660
rect 10425 -6780 10480 -6660
rect 10600 -6780 10645 -6660
rect 10765 -6780 10810 -6660
rect 10930 -6780 10975 -6660
rect 11095 -6780 11150 -6660
rect 11270 -6780 11315 -6660
rect 11435 -6780 11480 -6660
rect 11600 -6780 11645 -6660
rect 11765 -6780 11820 -6660
rect 11940 -6780 11985 -6660
rect 12105 -6780 12150 -6660
rect 12270 -6780 12315 -6660
rect 12435 -6780 12490 -6660
rect 12610 -6780 12620 -6660
rect 7120 -6825 12620 -6780
rect 7120 -6945 7130 -6825
rect 7250 -6945 7295 -6825
rect 7415 -6945 7460 -6825
rect 7580 -6945 7625 -6825
rect 7745 -6945 7800 -6825
rect 7920 -6945 7965 -6825
rect 8085 -6945 8130 -6825
rect 8250 -6945 8295 -6825
rect 8415 -6945 8470 -6825
rect 8590 -6945 8635 -6825
rect 8755 -6945 8800 -6825
rect 8920 -6945 8965 -6825
rect 9085 -6945 9140 -6825
rect 9260 -6945 9305 -6825
rect 9425 -6945 9470 -6825
rect 9590 -6945 9635 -6825
rect 9755 -6945 9810 -6825
rect 9930 -6945 9975 -6825
rect 10095 -6945 10140 -6825
rect 10260 -6945 10305 -6825
rect 10425 -6945 10480 -6825
rect 10600 -6945 10645 -6825
rect 10765 -6945 10810 -6825
rect 10930 -6945 10975 -6825
rect 11095 -6945 11150 -6825
rect 11270 -6945 11315 -6825
rect 11435 -6945 11480 -6825
rect 11600 -6945 11645 -6825
rect 11765 -6945 11820 -6825
rect 11940 -6945 11985 -6825
rect 12105 -6945 12150 -6825
rect 12270 -6945 12315 -6825
rect 12435 -6945 12490 -6825
rect 12610 -6945 12620 -6825
rect 7120 -6990 12620 -6945
rect 7120 -7110 7130 -6990
rect 7250 -7110 7295 -6990
rect 7415 -7110 7460 -6990
rect 7580 -7110 7625 -6990
rect 7745 -7110 7800 -6990
rect 7920 -7110 7965 -6990
rect 8085 -7110 8130 -6990
rect 8250 -7110 8295 -6990
rect 8415 -7110 8470 -6990
rect 8590 -7110 8635 -6990
rect 8755 -7110 8800 -6990
rect 8920 -7110 8965 -6990
rect 9085 -7110 9140 -6990
rect 9260 -7110 9305 -6990
rect 9425 -7110 9470 -6990
rect 9590 -7110 9635 -6990
rect 9755 -7110 9810 -6990
rect 9930 -7110 9975 -6990
rect 10095 -7110 10140 -6990
rect 10260 -7110 10305 -6990
rect 10425 -7110 10480 -6990
rect 10600 -7110 10645 -6990
rect 10765 -7110 10810 -6990
rect 10930 -7110 10975 -6990
rect 11095 -7110 11150 -6990
rect 11270 -7110 11315 -6990
rect 11435 -7110 11480 -6990
rect 11600 -7110 11645 -6990
rect 11765 -7110 11820 -6990
rect 11940 -7110 11985 -6990
rect 12105 -7110 12150 -6990
rect 12270 -7110 12315 -6990
rect 12435 -7110 12490 -6990
rect 12610 -7110 12620 -6990
rect 7120 -7165 12620 -7110
rect 7120 -7285 7130 -7165
rect 7250 -7285 7295 -7165
rect 7415 -7285 7460 -7165
rect 7580 -7285 7625 -7165
rect 7745 -7285 7800 -7165
rect 7920 -7285 7965 -7165
rect 8085 -7285 8130 -7165
rect 8250 -7285 8295 -7165
rect 8415 -7285 8470 -7165
rect 8590 -7285 8635 -7165
rect 8755 -7285 8800 -7165
rect 8920 -7285 8965 -7165
rect 9085 -7285 9140 -7165
rect 9260 -7285 9305 -7165
rect 9425 -7285 9470 -7165
rect 9590 -7285 9635 -7165
rect 9755 -7285 9810 -7165
rect 9930 -7285 9975 -7165
rect 10095 -7285 10140 -7165
rect 10260 -7285 10305 -7165
rect 10425 -7285 10480 -7165
rect 10600 -7285 10645 -7165
rect 10765 -7285 10810 -7165
rect 10930 -7285 10975 -7165
rect 11095 -7285 11150 -7165
rect 11270 -7285 11315 -7165
rect 11435 -7285 11480 -7165
rect 11600 -7285 11645 -7165
rect 11765 -7285 11820 -7165
rect 11940 -7285 11985 -7165
rect 12105 -7285 12150 -7165
rect 12270 -7285 12315 -7165
rect 12435 -7285 12490 -7165
rect 12610 -7285 12620 -7165
rect 7120 -7330 12620 -7285
rect 7120 -7450 7130 -7330
rect 7250 -7450 7295 -7330
rect 7415 -7450 7460 -7330
rect 7580 -7450 7625 -7330
rect 7745 -7450 7800 -7330
rect 7920 -7450 7965 -7330
rect 8085 -7450 8130 -7330
rect 8250 -7450 8295 -7330
rect 8415 -7450 8470 -7330
rect 8590 -7450 8635 -7330
rect 8755 -7450 8800 -7330
rect 8920 -7450 8965 -7330
rect 9085 -7450 9140 -7330
rect 9260 -7450 9305 -7330
rect 9425 -7450 9470 -7330
rect 9590 -7450 9635 -7330
rect 9755 -7450 9810 -7330
rect 9930 -7450 9975 -7330
rect 10095 -7450 10140 -7330
rect 10260 -7450 10305 -7330
rect 10425 -7450 10480 -7330
rect 10600 -7450 10645 -7330
rect 10765 -7450 10810 -7330
rect 10930 -7450 10975 -7330
rect 11095 -7450 11150 -7330
rect 11270 -7450 11315 -7330
rect 11435 -7450 11480 -7330
rect 11600 -7450 11645 -7330
rect 11765 -7450 11820 -7330
rect 11940 -7450 11985 -7330
rect 12105 -7450 12150 -7330
rect 12270 -7450 12315 -7330
rect 12435 -7450 12490 -7330
rect 12610 -7450 12620 -7330
rect 7120 -7495 12620 -7450
rect 7120 -7615 7130 -7495
rect 7250 -7615 7295 -7495
rect 7415 -7615 7460 -7495
rect 7580 -7615 7625 -7495
rect 7745 -7615 7800 -7495
rect 7920 -7615 7965 -7495
rect 8085 -7615 8130 -7495
rect 8250 -7615 8295 -7495
rect 8415 -7615 8470 -7495
rect 8590 -7615 8635 -7495
rect 8755 -7615 8800 -7495
rect 8920 -7615 8965 -7495
rect 9085 -7615 9140 -7495
rect 9260 -7615 9305 -7495
rect 9425 -7615 9470 -7495
rect 9590 -7615 9635 -7495
rect 9755 -7615 9810 -7495
rect 9930 -7615 9975 -7495
rect 10095 -7615 10140 -7495
rect 10260 -7615 10305 -7495
rect 10425 -7615 10480 -7495
rect 10600 -7615 10645 -7495
rect 10765 -7615 10810 -7495
rect 10930 -7615 10975 -7495
rect 11095 -7615 11150 -7495
rect 11270 -7615 11315 -7495
rect 11435 -7615 11480 -7495
rect 11600 -7615 11645 -7495
rect 11765 -7615 11820 -7495
rect 11940 -7615 11985 -7495
rect 12105 -7615 12150 -7495
rect 12270 -7615 12315 -7495
rect 12435 -7615 12490 -7495
rect 12610 -7615 12620 -7495
rect 7120 -7660 12620 -7615
rect 7120 -7780 7130 -7660
rect 7250 -7780 7295 -7660
rect 7415 -7780 7460 -7660
rect 7580 -7780 7625 -7660
rect 7745 -7780 7800 -7660
rect 7920 -7780 7965 -7660
rect 8085 -7780 8130 -7660
rect 8250 -7780 8295 -7660
rect 8415 -7780 8470 -7660
rect 8590 -7780 8635 -7660
rect 8755 -7780 8800 -7660
rect 8920 -7780 8965 -7660
rect 9085 -7780 9140 -7660
rect 9260 -7780 9305 -7660
rect 9425 -7780 9470 -7660
rect 9590 -7780 9635 -7660
rect 9755 -7780 9810 -7660
rect 9930 -7780 9975 -7660
rect 10095 -7780 10140 -7660
rect 10260 -7780 10305 -7660
rect 10425 -7780 10480 -7660
rect 10600 -7780 10645 -7660
rect 10765 -7780 10810 -7660
rect 10930 -7780 10975 -7660
rect 11095 -7780 11150 -7660
rect 11270 -7780 11315 -7660
rect 11435 -7780 11480 -7660
rect 11600 -7780 11645 -7660
rect 11765 -7780 11820 -7660
rect 11940 -7780 11985 -7660
rect 12105 -7780 12150 -7660
rect 12270 -7780 12315 -7660
rect 12435 -7780 12490 -7660
rect 12610 -7780 12620 -7660
rect 7120 -7835 12620 -7780
rect 7120 -7955 7130 -7835
rect 7250 -7955 7295 -7835
rect 7415 -7955 7460 -7835
rect 7580 -7955 7625 -7835
rect 7745 -7955 7800 -7835
rect 7920 -7955 7965 -7835
rect 8085 -7955 8130 -7835
rect 8250 -7955 8295 -7835
rect 8415 -7955 8470 -7835
rect 8590 -7955 8635 -7835
rect 8755 -7955 8800 -7835
rect 8920 -7955 8965 -7835
rect 9085 -7955 9140 -7835
rect 9260 -7955 9305 -7835
rect 9425 -7955 9470 -7835
rect 9590 -7955 9635 -7835
rect 9755 -7955 9810 -7835
rect 9930 -7955 9975 -7835
rect 10095 -7955 10140 -7835
rect 10260 -7955 10305 -7835
rect 10425 -7955 10480 -7835
rect 10600 -7955 10645 -7835
rect 10765 -7955 10810 -7835
rect 10930 -7955 10975 -7835
rect 11095 -7955 11150 -7835
rect 11270 -7955 11315 -7835
rect 11435 -7955 11480 -7835
rect 11600 -7955 11645 -7835
rect 11765 -7955 11820 -7835
rect 11940 -7955 11985 -7835
rect 12105 -7955 12150 -7835
rect 12270 -7955 12315 -7835
rect 12435 -7955 12490 -7835
rect 12610 -7955 12620 -7835
rect 7120 -8000 12620 -7955
rect 7120 -8120 7130 -8000
rect 7250 -8120 7295 -8000
rect 7415 -8120 7460 -8000
rect 7580 -8120 7625 -8000
rect 7745 -8120 7800 -8000
rect 7920 -8120 7965 -8000
rect 8085 -8120 8130 -8000
rect 8250 -8120 8295 -8000
rect 8415 -8120 8470 -8000
rect 8590 -8120 8635 -8000
rect 8755 -8120 8800 -8000
rect 8920 -8120 8965 -8000
rect 9085 -8120 9140 -8000
rect 9260 -8120 9305 -8000
rect 9425 -8120 9470 -8000
rect 9590 -8120 9635 -8000
rect 9755 -8120 9810 -8000
rect 9930 -8120 9975 -8000
rect 10095 -8120 10140 -8000
rect 10260 -8120 10305 -8000
rect 10425 -8120 10480 -8000
rect 10600 -8120 10645 -8000
rect 10765 -8120 10810 -8000
rect 10930 -8120 10975 -8000
rect 11095 -8120 11150 -8000
rect 11270 -8120 11315 -8000
rect 11435 -8120 11480 -8000
rect 11600 -8120 11645 -8000
rect 11765 -8120 11820 -8000
rect 11940 -8120 11985 -8000
rect 12105 -8120 12150 -8000
rect 12270 -8120 12315 -8000
rect 12435 -8120 12490 -8000
rect 12610 -8120 12620 -8000
rect 7120 -8165 12620 -8120
rect 7120 -8285 7130 -8165
rect 7250 -8285 7295 -8165
rect 7415 -8285 7460 -8165
rect 7580 -8285 7625 -8165
rect 7745 -8285 7800 -8165
rect 7920 -8285 7965 -8165
rect 8085 -8285 8130 -8165
rect 8250 -8285 8295 -8165
rect 8415 -8285 8470 -8165
rect 8590 -8285 8635 -8165
rect 8755 -8285 8800 -8165
rect 8920 -8285 8965 -8165
rect 9085 -8285 9140 -8165
rect 9260 -8285 9305 -8165
rect 9425 -8285 9470 -8165
rect 9590 -8285 9635 -8165
rect 9755 -8285 9810 -8165
rect 9930 -8285 9975 -8165
rect 10095 -8285 10140 -8165
rect 10260 -8285 10305 -8165
rect 10425 -8285 10480 -8165
rect 10600 -8285 10645 -8165
rect 10765 -8285 10810 -8165
rect 10930 -8285 10975 -8165
rect 11095 -8285 11150 -8165
rect 11270 -8285 11315 -8165
rect 11435 -8285 11480 -8165
rect 11600 -8285 11645 -8165
rect 11765 -8285 11820 -8165
rect 11940 -8285 11985 -8165
rect 12105 -8285 12150 -8165
rect 12270 -8285 12315 -8165
rect 12435 -8285 12490 -8165
rect 12610 -8285 12620 -8165
rect 7120 -8330 12620 -8285
rect 7120 -8450 7130 -8330
rect 7250 -8450 7295 -8330
rect 7415 -8450 7460 -8330
rect 7580 -8450 7625 -8330
rect 7745 -8450 7800 -8330
rect 7920 -8450 7965 -8330
rect 8085 -8450 8130 -8330
rect 8250 -8450 8295 -8330
rect 8415 -8450 8470 -8330
rect 8590 -8450 8635 -8330
rect 8755 -8450 8800 -8330
rect 8920 -8450 8965 -8330
rect 9085 -8450 9140 -8330
rect 9260 -8450 9305 -8330
rect 9425 -8450 9470 -8330
rect 9590 -8450 9635 -8330
rect 9755 -8450 9810 -8330
rect 9930 -8450 9975 -8330
rect 10095 -8450 10140 -8330
rect 10260 -8450 10305 -8330
rect 10425 -8450 10480 -8330
rect 10600 -8450 10645 -8330
rect 10765 -8450 10810 -8330
rect 10930 -8450 10975 -8330
rect 11095 -8450 11150 -8330
rect 11270 -8450 11315 -8330
rect 11435 -8450 11480 -8330
rect 11600 -8450 11645 -8330
rect 11765 -8450 11820 -8330
rect 11940 -8450 11985 -8330
rect 12105 -8450 12150 -8330
rect 12270 -8450 12315 -8330
rect 12435 -8450 12490 -8330
rect 12610 -8450 12620 -8330
rect 7120 -8505 12620 -8450
rect 7120 -8625 7130 -8505
rect 7250 -8625 7295 -8505
rect 7415 -8625 7460 -8505
rect 7580 -8625 7625 -8505
rect 7745 -8625 7800 -8505
rect 7920 -8625 7965 -8505
rect 8085 -8625 8130 -8505
rect 8250 -8625 8295 -8505
rect 8415 -8625 8470 -8505
rect 8590 -8625 8635 -8505
rect 8755 -8625 8800 -8505
rect 8920 -8625 8965 -8505
rect 9085 -8625 9140 -8505
rect 9260 -8625 9305 -8505
rect 9425 -8625 9470 -8505
rect 9590 -8625 9635 -8505
rect 9755 -8625 9810 -8505
rect 9930 -8625 9975 -8505
rect 10095 -8625 10140 -8505
rect 10260 -8625 10305 -8505
rect 10425 -8625 10480 -8505
rect 10600 -8625 10645 -8505
rect 10765 -8625 10810 -8505
rect 10930 -8625 10975 -8505
rect 11095 -8625 11150 -8505
rect 11270 -8625 11315 -8505
rect 11435 -8625 11480 -8505
rect 11600 -8625 11645 -8505
rect 11765 -8625 11820 -8505
rect 11940 -8625 11985 -8505
rect 12105 -8625 12150 -8505
rect 12270 -8625 12315 -8505
rect 12435 -8625 12490 -8505
rect 12610 -8625 12620 -8505
rect 7120 -8670 12620 -8625
rect 7120 -8790 7130 -8670
rect 7250 -8790 7295 -8670
rect 7415 -8790 7460 -8670
rect 7580 -8790 7625 -8670
rect 7745 -8790 7800 -8670
rect 7920 -8790 7965 -8670
rect 8085 -8790 8130 -8670
rect 8250 -8790 8295 -8670
rect 8415 -8790 8470 -8670
rect 8590 -8790 8635 -8670
rect 8755 -8790 8800 -8670
rect 8920 -8790 8965 -8670
rect 9085 -8790 9140 -8670
rect 9260 -8790 9305 -8670
rect 9425 -8790 9470 -8670
rect 9590 -8790 9635 -8670
rect 9755 -8790 9810 -8670
rect 9930 -8790 9975 -8670
rect 10095 -8790 10140 -8670
rect 10260 -8790 10305 -8670
rect 10425 -8790 10480 -8670
rect 10600 -8790 10645 -8670
rect 10765 -8790 10810 -8670
rect 10930 -8790 10975 -8670
rect 11095 -8790 11150 -8670
rect 11270 -8790 11315 -8670
rect 11435 -8790 11480 -8670
rect 11600 -8790 11645 -8670
rect 11765 -8790 11820 -8670
rect 11940 -8790 11985 -8670
rect 12105 -8790 12150 -8670
rect 12270 -8790 12315 -8670
rect 12435 -8790 12490 -8670
rect 12610 -8790 12620 -8670
rect 7120 -8835 12620 -8790
rect 7120 -8955 7130 -8835
rect 7250 -8955 7295 -8835
rect 7415 -8955 7460 -8835
rect 7580 -8955 7625 -8835
rect 7745 -8955 7800 -8835
rect 7920 -8955 7965 -8835
rect 8085 -8955 8130 -8835
rect 8250 -8955 8295 -8835
rect 8415 -8955 8470 -8835
rect 8590 -8955 8635 -8835
rect 8755 -8955 8800 -8835
rect 8920 -8955 8965 -8835
rect 9085 -8955 9140 -8835
rect 9260 -8955 9305 -8835
rect 9425 -8955 9470 -8835
rect 9590 -8955 9635 -8835
rect 9755 -8955 9810 -8835
rect 9930 -8955 9975 -8835
rect 10095 -8955 10140 -8835
rect 10260 -8955 10305 -8835
rect 10425 -8955 10480 -8835
rect 10600 -8955 10645 -8835
rect 10765 -8955 10810 -8835
rect 10930 -8955 10975 -8835
rect 11095 -8955 11150 -8835
rect 11270 -8955 11315 -8835
rect 11435 -8955 11480 -8835
rect 11600 -8955 11645 -8835
rect 11765 -8955 11820 -8835
rect 11940 -8955 11985 -8835
rect 12105 -8955 12150 -8835
rect 12270 -8955 12315 -8835
rect 12435 -8955 12490 -8835
rect 12610 -8955 12620 -8835
rect 7120 -9000 12620 -8955
rect 7120 -9120 7130 -9000
rect 7250 -9120 7295 -9000
rect 7415 -9120 7460 -9000
rect 7580 -9120 7625 -9000
rect 7745 -9120 7800 -9000
rect 7920 -9120 7965 -9000
rect 8085 -9120 8130 -9000
rect 8250 -9120 8295 -9000
rect 8415 -9120 8470 -9000
rect 8590 -9120 8635 -9000
rect 8755 -9120 8800 -9000
rect 8920 -9120 8965 -9000
rect 9085 -9120 9140 -9000
rect 9260 -9120 9305 -9000
rect 9425 -9120 9470 -9000
rect 9590 -9120 9635 -9000
rect 9755 -9120 9810 -9000
rect 9930 -9120 9975 -9000
rect 10095 -9120 10140 -9000
rect 10260 -9120 10305 -9000
rect 10425 -9120 10480 -9000
rect 10600 -9120 10645 -9000
rect 10765 -9120 10810 -9000
rect 10930 -9120 10975 -9000
rect 11095 -9120 11150 -9000
rect 11270 -9120 11315 -9000
rect 11435 -9120 11480 -9000
rect 11600 -9120 11645 -9000
rect 11765 -9120 11820 -9000
rect 11940 -9120 11985 -9000
rect 12105 -9120 12150 -9000
rect 12270 -9120 12315 -9000
rect 12435 -9120 12490 -9000
rect 12610 -9120 12620 -9000
rect 7120 -9175 12620 -9120
rect 7120 -9295 7130 -9175
rect 7250 -9295 7295 -9175
rect 7415 -9295 7460 -9175
rect 7580 -9295 7625 -9175
rect 7745 -9295 7800 -9175
rect 7920 -9295 7965 -9175
rect 8085 -9295 8130 -9175
rect 8250 -9295 8295 -9175
rect 8415 -9295 8470 -9175
rect 8590 -9295 8635 -9175
rect 8755 -9295 8800 -9175
rect 8920 -9295 8965 -9175
rect 9085 -9295 9140 -9175
rect 9260 -9295 9305 -9175
rect 9425 -9295 9470 -9175
rect 9590 -9295 9635 -9175
rect 9755 -9295 9810 -9175
rect 9930 -9295 9975 -9175
rect 10095 -9295 10140 -9175
rect 10260 -9295 10305 -9175
rect 10425 -9295 10480 -9175
rect 10600 -9295 10645 -9175
rect 10765 -9295 10810 -9175
rect 10930 -9295 10975 -9175
rect 11095 -9295 11150 -9175
rect 11270 -9295 11315 -9175
rect 11435 -9295 11480 -9175
rect 11600 -9295 11645 -9175
rect 11765 -9295 11820 -9175
rect 11940 -9295 11985 -9175
rect 12105 -9295 12150 -9175
rect 12270 -9295 12315 -9175
rect 12435 -9295 12490 -9175
rect 12610 -9295 12620 -9175
rect 7120 -9340 12620 -9295
rect 7120 -9460 7130 -9340
rect 7250 -9460 7295 -9340
rect 7415 -9460 7460 -9340
rect 7580 -9460 7625 -9340
rect 7745 -9460 7800 -9340
rect 7920 -9460 7965 -9340
rect 8085 -9460 8130 -9340
rect 8250 -9460 8295 -9340
rect 8415 -9460 8470 -9340
rect 8590 -9460 8635 -9340
rect 8755 -9460 8800 -9340
rect 8920 -9460 8965 -9340
rect 9085 -9460 9140 -9340
rect 9260 -9460 9305 -9340
rect 9425 -9460 9470 -9340
rect 9590 -9460 9635 -9340
rect 9755 -9460 9810 -9340
rect 9930 -9460 9975 -9340
rect 10095 -9460 10140 -9340
rect 10260 -9460 10305 -9340
rect 10425 -9460 10480 -9340
rect 10600 -9460 10645 -9340
rect 10765 -9460 10810 -9340
rect 10930 -9460 10975 -9340
rect 11095 -9460 11150 -9340
rect 11270 -9460 11315 -9340
rect 11435 -9460 11480 -9340
rect 11600 -9460 11645 -9340
rect 11765 -9460 11820 -9340
rect 11940 -9460 11985 -9340
rect 12105 -9460 12150 -9340
rect 12270 -9460 12315 -9340
rect 12435 -9460 12490 -9340
rect 12610 -9460 12620 -9340
rect 7120 -9505 12620 -9460
rect 7120 -9625 7130 -9505
rect 7250 -9625 7295 -9505
rect 7415 -9625 7460 -9505
rect 7580 -9625 7625 -9505
rect 7745 -9625 7800 -9505
rect 7920 -9625 7965 -9505
rect 8085 -9625 8130 -9505
rect 8250 -9625 8295 -9505
rect 8415 -9625 8470 -9505
rect 8590 -9625 8635 -9505
rect 8755 -9625 8800 -9505
rect 8920 -9625 8965 -9505
rect 9085 -9625 9140 -9505
rect 9260 -9625 9305 -9505
rect 9425 -9625 9470 -9505
rect 9590 -9625 9635 -9505
rect 9755 -9625 9810 -9505
rect 9930 -9625 9975 -9505
rect 10095 -9625 10140 -9505
rect 10260 -9625 10305 -9505
rect 10425 -9625 10480 -9505
rect 10600 -9625 10645 -9505
rect 10765 -9625 10810 -9505
rect 10930 -9625 10975 -9505
rect 11095 -9625 11150 -9505
rect 11270 -9625 11315 -9505
rect 11435 -9625 11480 -9505
rect 11600 -9625 11645 -9505
rect 11765 -9625 11820 -9505
rect 11940 -9625 11985 -9505
rect 12105 -9625 12150 -9505
rect 12270 -9625 12315 -9505
rect 12435 -9625 12490 -9505
rect 12610 -9625 12620 -9505
rect 7120 -9670 12620 -9625
rect 7120 -9790 7130 -9670
rect 7250 -9790 7295 -9670
rect 7415 -9790 7460 -9670
rect 7580 -9790 7625 -9670
rect 7745 -9790 7800 -9670
rect 7920 -9790 7965 -9670
rect 8085 -9790 8130 -9670
rect 8250 -9790 8295 -9670
rect 8415 -9790 8470 -9670
rect 8590 -9790 8635 -9670
rect 8755 -9790 8800 -9670
rect 8920 -9790 8965 -9670
rect 9085 -9790 9140 -9670
rect 9260 -9790 9305 -9670
rect 9425 -9790 9470 -9670
rect 9590 -9790 9635 -9670
rect 9755 -9790 9810 -9670
rect 9930 -9790 9975 -9670
rect 10095 -9790 10140 -9670
rect 10260 -9790 10305 -9670
rect 10425 -9790 10480 -9670
rect 10600 -9790 10645 -9670
rect 10765 -9790 10810 -9670
rect 10930 -9790 10975 -9670
rect 11095 -9790 11150 -9670
rect 11270 -9790 11315 -9670
rect 11435 -9790 11480 -9670
rect 11600 -9790 11645 -9670
rect 11765 -9790 11820 -9670
rect 11940 -9790 11985 -9670
rect 12105 -9790 12150 -9670
rect 12270 -9790 12315 -9670
rect 12435 -9790 12490 -9670
rect 12610 -9790 12620 -9670
rect 7120 -9800 12620 -9790
rect 12810 -4310 18310 -4300
rect 12810 -4430 12820 -4310
rect 12940 -4430 12985 -4310
rect 13105 -4430 13150 -4310
rect 13270 -4430 13315 -4310
rect 13435 -4430 13490 -4310
rect 13610 -4430 13655 -4310
rect 13775 -4430 13820 -4310
rect 13940 -4430 13985 -4310
rect 14105 -4430 14160 -4310
rect 14280 -4430 14325 -4310
rect 14445 -4430 14490 -4310
rect 14610 -4430 14655 -4310
rect 14775 -4430 14830 -4310
rect 14950 -4430 14995 -4310
rect 15115 -4430 15160 -4310
rect 15280 -4430 15325 -4310
rect 15445 -4430 15500 -4310
rect 15620 -4430 15665 -4310
rect 15785 -4430 15830 -4310
rect 15950 -4430 15995 -4310
rect 16115 -4430 16170 -4310
rect 16290 -4430 16335 -4310
rect 16455 -4430 16500 -4310
rect 16620 -4430 16665 -4310
rect 16785 -4430 16840 -4310
rect 16960 -4430 17005 -4310
rect 17125 -4430 17170 -4310
rect 17290 -4430 17335 -4310
rect 17455 -4430 17510 -4310
rect 17630 -4430 17675 -4310
rect 17795 -4430 17840 -4310
rect 17960 -4430 18005 -4310
rect 18125 -4430 18180 -4310
rect 18300 -4430 18310 -4310
rect 12810 -4485 18310 -4430
rect 12810 -4605 12820 -4485
rect 12940 -4605 12985 -4485
rect 13105 -4605 13150 -4485
rect 13270 -4605 13315 -4485
rect 13435 -4605 13490 -4485
rect 13610 -4605 13655 -4485
rect 13775 -4605 13820 -4485
rect 13940 -4605 13985 -4485
rect 14105 -4605 14160 -4485
rect 14280 -4605 14325 -4485
rect 14445 -4605 14490 -4485
rect 14610 -4605 14655 -4485
rect 14775 -4605 14830 -4485
rect 14950 -4605 14995 -4485
rect 15115 -4605 15160 -4485
rect 15280 -4605 15325 -4485
rect 15445 -4605 15500 -4485
rect 15620 -4605 15665 -4485
rect 15785 -4605 15830 -4485
rect 15950 -4605 15995 -4485
rect 16115 -4605 16170 -4485
rect 16290 -4605 16335 -4485
rect 16455 -4605 16500 -4485
rect 16620 -4605 16665 -4485
rect 16785 -4605 16840 -4485
rect 16960 -4605 17005 -4485
rect 17125 -4605 17170 -4485
rect 17290 -4605 17335 -4485
rect 17455 -4605 17510 -4485
rect 17630 -4605 17675 -4485
rect 17795 -4605 17840 -4485
rect 17960 -4605 18005 -4485
rect 18125 -4605 18180 -4485
rect 18300 -4605 18310 -4485
rect 12810 -4650 18310 -4605
rect 12810 -4770 12820 -4650
rect 12940 -4770 12985 -4650
rect 13105 -4770 13150 -4650
rect 13270 -4770 13315 -4650
rect 13435 -4770 13490 -4650
rect 13610 -4770 13655 -4650
rect 13775 -4770 13820 -4650
rect 13940 -4770 13985 -4650
rect 14105 -4770 14160 -4650
rect 14280 -4770 14325 -4650
rect 14445 -4770 14490 -4650
rect 14610 -4770 14655 -4650
rect 14775 -4770 14830 -4650
rect 14950 -4770 14995 -4650
rect 15115 -4770 15160 -4650
rect 15280 -4770 15325 -4650
rect 15445 -4770 15500 -4650
rect 15620 -4770 15665 -4650
rect 15785 -4770 15830 -4650
rect 15950 -4770 15995 -4650
rect 16115 -4770 16170 -4650
rect 16290 -4770 16335 -4650
rect 16455 -4770 16500 -4650
rect 16620 -4770 16665 -4650
rect 16785 -4770 16840 -4650
rect 16960 -4770 17005 -4650
rect 17125 -4770 17170 -4650
rect 17290 -4770 17335 -4650
rect 17455 -4770 17510 -4650
rect 17630 -4770 17675 -4650
rect 17795 -4770 17840 -4650
rect 17960 -4770 18005 -4650
rect 18125 -4770 18180 -4650
rect 18300 -4770 18310 -4650
rect 12810 -4815 18310 -4770
rect 12810 -4935 12820 -4815
rect 12940 -4935 12985 -4815
rect 13105 -4935 13150 -4815
rect 13270 -4935 13315 -4815
rect 13435 -4935 13490 -4815
rect 13610 -4935 13655 -4815
rect 13775 -4935 13820 -4815
rect 13940 -4935 13985 -4815
rect 14105 -4935 14160 -4815
rect 14280 -4935 14325 -4815
rect 14445 -4935 14490 -4815
rect 14610 -4935 14655 -4815
rect 14775 -4935 14830 -4815
rect 14950 -4935 14995 -4815
rect 15115 -4935 15160 -4815
rect 15280 -4935 15325 -4815
rect 15445 -4935 15500 -4815
rect 15620 -4935 15665 -4815
rect 15785 -4935 15830 -4815
rect 15950 -4935 15995 -4815
rect 16115 -4935 16170 -4815
rect 16290 -4935 16335 -4815
rect 16455 -4935 16500 -4815
rect 16620 -4935 16665 -4815
rect 16785 -4935 16840 -4815
rect 16960 -4935 17005 -4815
rect 17125 -4935 17170 -4815
rect 17290 -4935 17335 -4815
rect 17455 -4935 17510 -4815
rect 17630 -4935 17675 -4815
rect 17795 -4935 17840 -4815
rect 17960 -4935 18005 -4815
rect 18125 -4935 18180 -4815
rect 18300 -4935 18310 -4815
rect 12810 -4980 18310 -4935
rect 12810 -5100 12820 -4980
rect 12940 -5100 12985 -4980
rect 13105 -5100 13150 -4980
rect 13270 -5100 13315 -4980
rect 13435 -5100 13490 -4980
rect 13610 -5100 13655 -4980
rect 13775 -5100 13820 -4980
rect 13940 -5100 13985 -4980
rect 14105 -5100 14160 -4980
rect 14280 -5100 14325 -4980
rect 14445 -5100 14490 -4980
rect 14610 -5100 14655 -4980
rect 14775 -5100 14830 -4980
rect 14950 -5100 14995 -4980
rect 15115 -5100 15160 -4980
rect 15280 -5100 15325 -4980
rect 15445 -5100 15500 -4980
rect 15620 -5100 15665 -4980
rect 15785 -5100 15830 -4980
rect 15950 -5100 15995 -4980
rect 16115 -5100 16170 -4980
rect 16290 -5100 16335 -4980
rect 16455 -5100 16500 -4980
rect 16620 -5100 16665 -4980
rect 16785 -5100 16840 -4980
rect 16960 -5100 17005 -4980
rect 17125 -5100 17170 -4980
rect 17290 -5100 17335 -4980
rect 17455 -5100 17510 -4980
rect 17630 -5100 17675 -4980
rect 17795 -5100 17840 -4980
rect 17960 -5100 18005 -4980
rect 18125 -5100 18180 -4980
rect 18300 -5100 18310 -4980
rect 12810 -5155 18310 -5100
rect 12810 -5275 12820 -5155
rect 12940 -5275 12985 -5155
rect 13105 -5275 13150 -5155
rect 13270 -5275 13315 -5155
rect 13435 -5275 13490 -5155
rect 13610 -5275 13655 -5155
rect 13775 -5275 13820 -5155
rect 13940 -5275 13985 -5155
rect 14105 -5275 14160 -5155
rect 14280 -5275 14325 -5155
rect 14445 -5275 14490 -5155
rect 14610 -5275 14655 -5155
rect 14775 -5275 14830 -5155
rect 14950 -5275 14995 -5155
rect 15115 -5275 15160 -5155
rect 15280 -5275 15325 -5155
rect 15445 -5275 15500 -5155
rect 15620 -5275 15665 -5155
rect 15785 -5275 15830 -5155
rect 15950 -5275 15995 -5155
rect 16115 -5275 16170 -5155
rect 16290 -5275 16335 -5155
rect 16455 -5275 16500 -5155
rect 16620 -5275 16665 -5155
rect 16785 -5275 16840 -5155
rect 16960 -5275 17005 -5155
rect 17125 -5275 17170 -5155
rect 17290 -5275 17335 -5155
rect 17455 -5275 17510 -5155
rect 17630 -5275 17675 -5155
rect 17795 -5275 17840 -5155
rect 17960 -5275 18005 -5155
rect 18125 -5275 18180 -5155
rect 18300 -5275 18310 -5155
rect 12810 -5320 18310 -5275
rect 12810 -5440 12820 -5320
rect 12940 -5440 12985 -5320
rect 13105 -5440 13150 -5320
rect 13270 -5440 13315 -5320
rect 13435 -5440 13490 -5320
rect 13610 -5440 13655 -5320
rect 13775 -5440 13820 -5320
rect 13940 -5440 13985 -5320
rect 14105 -5440 14160 -5320
rect 14280 -5440 14325 -5320
rect 14445 -5440 14490 -5320
rect 14610 -5440 14655 -5320
rect 14775 -5440 14830 -5320
rect 14950 -5440 14995 -5320
rect 15115 -5440 15160 -5320
rect 15280 -5440 15325 -5320
rect 15445 -5440 15500 -5320
rect 15620 -5440 15665 -5320
rect 15785 -5440 15830 -5320
rect 15950 -5440 15995 -5320
rect 16115 -5440 16170 -5320
rect 16290 -5440 16335 -5320
rect 16455 -5440 16500 -5320
rect 16620 -5440 16665 -5320
rect 16785 -5440 16840 -5320
rect 16960 -5440 17005 -5320
rect 17125 -5440 17170 -5320
rect 17290 -5440 17335 -5320
rect 17455 -5440 17510 -5320
rect 17630 -5440 17675 -5320
rect 17795 -5440 17840 -5320
rect 17960 -5440 18005 -5320
rect 18125 -5440 18180 -5320
rect 18300 -5440 18310 -5320
rect 12810 -5485 18310 -5440
rect 12810 -5605 12820 -5485
rect 12940 -5605 12985 -5485
rect 13105 -5605 13150 -5485
rect 13270 -5605 13315 -5485
rect 13435 -5605 13490 -5485
rect 13610 -5605 13655 -5485
rect 13775 -5605 13820 -5485
rect 13940 -5605 13985 -5485
rect 14105 -5605 14160 -5485
rect 14280 -5605 14325 -5485
rect 14445 -5605 14490 -5485
rect 14610 -5605 14655 -5485
rect 14775 -5605 14830 -5485
rect 14950 -5605 14995 -5485
rect 15115 -5605 15160 -5485
rect 15280 -5605 15325 -5485
rect 15445 -5605 15500 -5485
rect 15620 -5605 15665 -5485
rect 15785 -5605 15830 -5485
rect 15950 -5605 15995 -5485
rect 16115 -5605 16170 -5485
rect 16290 -5605 16335 -5485
rect 16455 -5605 16500 -5485
rect 16620 -5605 16665 -5485
rect 16785 -5605 16840 -5485
rect 16960 -5605 17005 -5485
rect 17125 -5605 17170 -5485
rect 17290 -5605 17335 -5485
rect 17455 -5605 17510 -5485
rect 17630 -5605 17675 -5485
rect 17795 -5605 17840 -5485
rect 17960 -5605 18005 -5485
rect 18125 -5605 18180 -5485
rect 18300 -5605 18310 -5485
rect 12810 -5650 18310 -5605
rect 12810 -5770 12820 -5650
rect 12940 -5770 12985 -5650
rect 13105 -5770 13150 -5650
rect 13270 -5770 13315 -5650
rect 13435 -5770 13490 -5650
rect 13610 -5770 13655 -5650
rect 13775 -5770 13820 -5650
rect 13940 -5770 13985 -5650
rect 14105 -5770 14160 -5650
rect 14280 -5770 14325 -5650
rect 14445 -5770 14490 -5650
rect 14610 -5770 14655 -5650
rect 14775 -5770 14830 -5650
rect 14950 -5770 14995 -5650
rect 15115 -5770 15160 -5650
rect 15280 -5770 15325 -5650
rect 15445 -5770 15500 -5650
rect 15620 -5770 15665 -5650
rect 15785 -5770 15830 -5650
rect 15950 -5770 15995 -5650
rect 16115 -5770 16170 -5650
rect 16290 -5770 16335 -5650
rect 16455 -5770 16500 -5650
rect 16620 -5770 16665 -5650
rect 16785 -5770 16840 -5650
rect 16960 -5770 17005 -5650
rect 17125 -5770 17170 -5650
rect 17290 -5770 17335 -5650
rect 17455 -5770 17510 -5650
rect 17630 -5770 17675 -5650
rect 17795 -5770 17840 -5650
rect 17960 -5770 18005 -5650
rect 18125 -5770 18180 -5650
rect 18300 -5770 18310 -5650
rect 12810 -5825 18310 -5770
rect 12810 -5945 12820 -5825
rect 12940 -5945 12985 -5825
rect 13105 -5945 13150 -5825
rect 13270 -5945 13315 -5825
rect 13435 -5945 13490 -5825
rect 13610 -5945 13655 -5825
rect 13775 -5945 13820 -5825
rect 13940 -5945 13985 -5825
rect 14105 -5945 14160 -5825
rect 14280 -5945 14325 -5825
rect 14445 -5945 14490 -5825
rect 14610 -5945 14655 -5825
rect 14775 -5945 14830 -5825
rect 14950 -5945 14995 -5825
rect 15115 -5945 15160 -5825
rect 15280 -5945 15325 -5825
rect 15445 -5945 15500 -5825
rect 15620 -5945 15665 -5825
rect 15785 -5945 15830 -5825
rect 15950 -5945 15995 -5825
rect 16115 -5945 16170 -5825
rect 16290 -5945 16335 -5825
rect 16455 -5945 16500 -5825
rect 16620 -5945 16665 -5825
rect 16785 -5945 16840 -5825
rect 16960 -5945 17005 -5825
rect 17125 -5945 17170 -5825
rect 17290 -5945 17335 -5825
rect 17455 -5945 17510 -5825
rect 17630 -5945 17675 -5825
rect 17795 -5945 17840 -5825
rect 17960 -5945 18005 -5825
rect 18125 -5945 18180 -5825
rect 18300 -5945 18310 -5825
rect 12810 -5990 18310 -5945
rect 12810 -6110 12820 -5990
rect 12940 -6110 12985 -5990
rect 13105 -6110 13150 -5990
rect 13270 -6110 13315 -5990
rect 13435 -6110 13490 -5990
rect 13610 -6110 13655 -5990
rect 13775 -6110 13820 -5990
rect 13940 -6110 13985 -5990
rect 14105 -6110 14160 -5990
rect 14280 -6110 14325 -5990
rect 14445 -6110 14490 -5990
rect 14610 -6110 14655 -5990
rect 14775 -6110 14830 -5990
rect 14950 -6110 14995 -5990
rect 15115 -6110 15160 -5990
rect 15280 -6110 15325 -5990
rect 15445 -6110 15500 -5990
rect 15620 -6110 15665 -5990
rect 15785 -6110 15830 -5990
rect 15950 -6110 15995 -5990
rect 16115 -6110 16170 -5990
rect 16290 -6110 16335 -5990
rect 16455 -6110 16500 -5990
rect 16620 -6110 16665 -5990
rect 16785 -6110 16840 -5990
rect 16960 -6110 17005 -5990
rect 17125 -6110 17170 -5990
rect 17290 -6110 17335 -5990
rect 17455 -6110 17510 -5990
rect 17630 -6110 17675 -5990
rect 17795 -6110 17840 -5990
rect 17960 -6110 18005 -5990
rect 18125 -6110 18180 -5990
rect 18300 -6110 18310 -5990
rect 12810 -6155 18310 -6110
rect 12810 -6275 12820 -6155
rect 12940 -6275 12985 -6155
rect 13105 -6275 13150 -6155
rect 13270 -6275 13315 -6155
rect 13435 -6275 13490 -6155
rect 13610 -6275 13655 -6155
rect 13775 -6275 13820 -6155
rect 13940 -6275 13985 -6155
rect 14105 -6275 14160 -6155
rect 14280 -6275 14325 -6155
rect 14445 -6275 14490 -6155
rect 14610 -6275 14655 -6155
rect 14775 -6275 14830 -6155
rect 14950 -6275 14995 -6155
rect 15115 -6275 15160 -6155
rect 15280 -6275 15325 -6155
rect 15445 -6275 15500 -6155
rect 15620 -6275 15665 -6155
rect 15785 -6275 15830 -6155
rect 15950 -6275 15995 -6155
rect 16115 -6275 16170 -6155
rect 16290 -6275 16335 -6155
rect 16455 -6275 16500 -6155
rect 16620 -6275 16665 -6155
rect 16785 -6275 16840 -6155
rect 16960 -6275 17005 -6155
rect 17125 -6275 17170 -6155
rect 17290 -6275 17335 -6155
rect 17455 -6275 17510 -6155
rect 17630 -6275 17675 -6155
rect 17795 -6275 17840 -6155
rect 17960 -6275 18005 -6155
rect 18125 -6275 18180 -6155
rect 18300 -6275 18310 -6155
rect 12810 -6320 18310 -6275
rect 12810 -6440 12820 -6320
rect 12940 -6440 12985 -6320
rect 13105 -6440 13150 -6320
rect 13270 -6440 13315 -6320
rect 13435 -6440 13490 -6320
rect 13610 -6440 13655 -6320
rect 13775 -6440 13820 -6320
rect 13940 -6440 13985 -6320
rect 14105 -6440 14160 -6320
rect 14280 -6440 14325 -6320
rect 14445 -6440 14490 -6320
rect 14610 -6440 14655 -6320
rect 14775 -6440 14830 -6320
rect 14950 -6440 14995 -6320
rect 15115 -6440 15160 -6320
rect 15280 -6440 15325 -6320
rect 15445 -6440 15500 -6320
rect 15620 -6440 15665 -6320
rect 15785 -6440 15830 -6320
rect 15950 -6440 15995 -6320
rect 16115 -6440 16170 -6320
rect 16290 -6440 16335 -6320
rect 16455 -6440 16500 -6320
rect 16620 -6440 16665 -6320
rect 16785 -6440 16840 -6320
rect 16960 -6440 17005 -6320
rect 17125 -6440 17170 -6320
rect 17290 -6440 17335 -6320
rect 17455 -6440 17510 -6320
rect 17630 -6440 17675 -6320
rect 17795 -6440 17840 -6320
rect 17960 -6440 18005 -6320
rect 18125 -6440 18180 -6320
rect 18300 -6440 18310 -6320
rect 12810 -6495 18310 -6440
rect 12810 -6615 12820 -6495
rect 12940 -6615 12985 -6495
rect 13105 -6615 13150 -6495
rect 13270 -6615 13315 -6495
rect 13435 -6615 13490 -6495
rect 13610 -6615 13655 -6495
rect 13775 -6615 13820 -6495
rect 13940 -6615 13985 -6495
rect 14105 -6615 14160 -6495
rect 14280 -6615 14325 -6495
rect 14445 -6615 14490 -6495
rect 14610 -6615 14655 -6495
rect 14775 -6615 14830 -6495
rect 14950 -6615 14995 -6495
rect 15115 -6615 15160 -6495
rect 15280 -6615 15325 -6495
rect 15445 -6615 15500 -6495
rect 15620 -6615 15665 -6495
rect 15785 -6615 15830 -6495
rect 15950 -6615 15995 -6495
rect 16115 -6615 16170 -6495
rect 16290 -6615 16335 -6495
rect 16455 -6615 16500 -6495
rect 16620 -6615 16665 -6495
rect 16785 -6615 16840 -6495
rect 16960 -6615 17005 -6495
rect 17125 -6615 17170 -6495
rect 17290 -6615 17335 -6495
rect 17455 -6615 17510 -6495
rect 17630 -6615 17675 -6495
rect 17795 -6615 17840 -6495
rect 17960 -6615 18005 -6495
rect 18125 -6615 18180 -6495
rect 18300 -6615 18310 -6495
rect 12810 -6660 18310 -6615
rect 12810 -6780 12820 -6660
rect 12940 -6780 12985 -6660
rect 13105 -6780 13150 -6660
rect 13270 -6780 13315 -6660
rect 13435 -6780 13490 -6660
rect 13610 -6780 13655 -6660
rect 13775 -6780 13820 -6660
rect 13940 -6780 13985 -6660
rect 14105 -6780 14160 -6660
rect 14280 -6780 14325 -6660
rect 14445 -6780 14490 -6660
rect 14610 -6780 14655 -6660
rect 14775 -6780 14830 -6660
rect 14950 -6780 14995 -6660
rect 15115 -6780 15160 -6660
rect 15280 -6780 15325 -6660
rect 15445 -6780 15500 -6660
rect 15620 -6780 15665 -6660
rect 15785 -6780 15830 -6660
rect 15950 -6780 15995 -6660
rect 16115 -6780 16170 -6660
rect 16290 -6780 16335 -6660
rect 16455 -6780 16500 -6660
rect 16620 -6780 16665 -6660
rect 16785 -6780 16840 -6660
rect 16960 -6780 17005 -6660
rect 17125 -6780 17170 -6660
rect 17290 -6780 17335 -6660
rect 17455 -6780 17510 -6660
rect 17630 -6780 17675 -6660
rect 17795 -6780 17840 -6660
rect 17960 -6780 18005 -6660
rect 18125 -6780 18180 -6660
rect 18300 -6780 18310 -6660
rect 12810 -6825 18310 -6780
rect 12810 -6945 12820 -6825
rect 12940 -6945 12985 -6825
rect 13105 -6945 13150 -6825
rect 13270 -6945 13315 -6825
rect 13435 -6945 13490 -6825
rect 13610 -6945 13655 -6825
rect 13775 -6945 13820 -6825
rect 13940 -6945 13985 -6825
rect 14105 -6945 14160 -6825
rect 14280 -6945 14325 -6825
rect 14445 -6945 14490 -6825
rect 14610 -6945 14655 -6825
rect 14775 -6945 14830 -6825
rect 14950 -6945 14995 -6825
rect 15115 -6945 15160 -6825
rect 15280 -6945 15325 -6825
rect 15445 -6945 15500 -6825
rect 15620 -6945 15665 -6825
rect 15785 -6945 15830 -6825
rect 15950 -6945 15995 -6825
rect 16115 -6945 16170 -6825
rect 16290 -6945 16335 -6825
rect 16455 -6945 16500 -6825
rect 16620 -6945 16665 -6825
rect 16785 -6945 16840 -6825
rect 16960 -6945 17005 -6825
rect 17125 -6945 17170 -6825
rect 17290 -6945 17335 -6825
rect 17455 -6945 17510 -6825
rect 17630 -6945 17675 -6825
rect 17795 -6945 17840 -6825
rect 17960 -6945 18005 -6825
rect 18125 -6945 18180 -6825
rect 18300 -6945 18310 -6825
rect 12810 -6990 18310 -6945
rect 12810 -7110 12820 -6990
rect 12940 -7110 12985 -6990
rect 13105 -7110 13150 -6990
rect 13270 -7110 13315 -6990
rect 13435 -7110 13490 -6990
rect 13610 -7110 13655 -6990
rect 13775 -7110 13820 -6990
rect 13940 -7110 13985 -6990
rect 14105 -7110 14160 -6990
rect 14280 -7110 14325 -6990
rect 14445 -7110 14490 -6990
rect 14610 -7110 14655 -6990
rect 14775 -7110 14830 -6990
rect 14950 -7110 14995 -6990
rect 15115 -7110 15160 -6990
rect 15280 -7110 15325 -6990
rect 15445 -7110 15500 -6990
rect 15620 -7110 15665 -6990
rect 15785 -7110 15830 -6990
rect 15950 -7110 15995 -6990
rect 16115 -7110 16170 -6990
rect 16290 -7110 16335 -6990
rect 16455 -7110 16500 -6990
rect 16620 -7110 16665 -6990
rect 16785 -7110 16840 -6990
rect 16960 -7110 17005 -6990
rect 17125 -7110 17170 -6990
rect 17290 -7110 17335 -6990
rect 17455 -7110 17510 -6990
rect 17630 -7110 17675 -6990
rect 17795 -7110 17840 -6990
rect 17960 -7110 18005 -6990
rect 18125 -7110 18180 -6990
rect 18300 -7110 18310 -6990
rect 12810 -7165 18310 -7110
rect 12810 -7285 12820 -7165
rect 12940 -7285 12985 -7165
rect 13105 -7285 13150 -7165
rect 13270 -7285 13315 -7165
rect 13435 -7285 13490 -7165
rect 13610 -7285 13655 -7165
rect 13775 -7285 13820 -7165
rect 13940 -7285 13985 -7165
rect 14105 -7285 14160 -7165
rect 14280 -7285 14325 -7165
rect 14445 -7285 14490 -7165
rect 14610 -7285 14655 -7165
rect 14775 -7285 14830 -7165
rect 14950 -7285 14995 -7165
rect 15115 -7285 15160 -7165
rect 15280 -7285 15325 -7165
rect 15445 -7285 15500 -7165
rect 15620 -7285 15665 -7165
rect 15785 -7285 15830 -7165
rect 15950 -7285 15995 -7165
rect 16115 -7285 16170 -7165
rect 16290 -7285 16335 -7165
rect 16455 -7285 16500 -7165
rect 16620 -7285 16665 -7165
rect 16785 -7285 16840 -7165
rect 16960 -7285 17005 -7165
rect 17125 -7285 17170 -7165
rect 17290 -7285 17335 -7165
rect 17455 -7285 17510 -7165
rect 17630 -7285 17675 -7165
rect 17795 -7285 17840 -7165
rect 17960 -7285 18005 -7165
rect 18125 -7285 18180 -7165
rect 18300 -7285 18310 -7165
rect 12810 -7330 18310 -7285
rect 12810 -7450 12820 -7330
rect 12940 -7450 12985 -7330
rect 13105 -7450 13150 -7330
rect 13270 -7450 13315 -7330
rect 13435 -7450 13490 -7330
rect 13610 -7450 13655 -7330
rect 13775 -7450 13820 -7330
rect 13940 -7450 13985 -7330
rect 14105 -7450 14160 -7330
rect 14280 -7450 14325 -7330
rect 14445 -7450 14490 -7330
rect 14610 -7450 14655 -7330
rect 14775 -7450 14830 -7330
rect 14950 -7450 14995 -7330
rect 15115 -7450 15160 -7330
rect 15280 -7450 15325 -7330
rect 15445 -7450 15500 -7330
rect 15620 -7450 15665 -7330
rect 15785 -7450 15830 -7330
rect 15950 -7450 15995 -7330
rect 16115 -7450 16170 -7330
rect 16290 -7450 16335 -7330
rect 16455 -7450 16500 -7330
rect 16620 -7450 16665 -7330
rect 16785 -7450 16840 -7330
rect 16960 -7450 17005 -7330
rect 17125 -7450 17170 -7330
rect 17290 -7450 17335 -7330
rect 17455 -7450 17510 -7330
rect 17630 -7450 17675 -7330
rect 17795 -7450 17840 -7330
rect 17960 -7450 18005 -7330
rect 18125 -7450 18180 -7330
rect 18300 -7450 18310 -7330
rect 12810 -7495 18310 -7450
rect 12810 -7615 12820 -7495
rect 12940 -7615 12985 -7495
rect 13105 -7615 13150 -7495
rect 13270 -7615 13315 -7495
rect 13435 -7615 13490 -7495
rect 13610 -7615 13655 -7495
rect 13775 -7615 13820 -7495
rect 13940 -7615 13985 -7495
rect 14105 -7615 14160 -7495
rect 14280 -7615 14325 -7495
rect 14445 -7615 14490 -7495
rect 14610 -7615 14655 -7495
rect 14775 -7615 14830 -7495
rect 14950 -7615 14995 -7495
rect 15115 -7615 15160 -7495
rect 15280 -7615 15325 -7495
rect 15445 -7615 15500 -7495
rect 15620 -7615 15665 -7495
rect 15785 -7615 15830 -7495
rect 15950 -7615 15995 -7495
rect 16115 -7615 16170 -7495
rect 16290 -7615 16335 -7495
rect 16455 -7615 16500 -7495
rect 16620 -7615 16665 -7495
rect 16785 -7615 16840 -7495
rect 16960 -7615 17005 -7495
rect 17125 -7615 17170 -7495
rect 17290 -7615 17335 -7495
rect 17455 -7615 17510 -7495
rect 17630 -7615 17675 -7495
rect 17795 -7615 17840 -7495
rect 17960 -7615 18005 -7495
rect 18125 -7615 18180 -7495
rect 18300 -7615 18310 -7495
rect 12810 -7660 18310 -7615
rect 12810 -7780 12820 -7660
rect 12940 -7780 12985 -7660
rect 13105 -7780 13150 -7660
rect 13270 -7780 13315 -7660
rect 13435 -7780 13490 -7660
rect 13610 -7780 13655 -7660
rect 13775 -7780 13820 -7660
rect 13940 -7780 13985 -7660
rect 14105 -7780 14160 -7660
rect 14280 -7780 14325 -7660
rect 14445 -7780 14490 -7660
rect 14610 -7780 14655 -7660
rect 14775 -7780 14830 -7660
rect 14950 -7780 14995 -7660
rect 15115 -7780 15160 -7660
rect 15280 -7780 15325 -7660
rect 15445 -7780 15500 -7660
rect 15620 -7780 15665 -7660
rect 15785 -7780 15830 -7660
rect 15950 -7780 15995 -7660
rect 16115 -7780 16170 -7660
rect 16290 -7780 16335 -7660
rect 16455 -7780 16500 -7660
rect 16620 -7780 16665 -7660
rect 16785 -7780 16840 -7660
rect 16960 -7780 17005 -7660
rect 17125 -7780 17170 -7660
rect 17290 -7780 17335 -7660
rect 17455 -7780 17510 -7660
rect 17630 -7780 17675 -7660
rect 17795 -7780 17840 -7660
rect 17960 -7780 18005 -7660
rect 18125 -7780 18180 -7660
rect 18300 -7780 18310 -7660
rect 12810 -7835 18310 -7780
rect 12810 -7955 12820 -7835
rect 12940 -7955 12985 -7835
rect 13105 -7955 13150 -7835
rect 13270 -7955 13315 -7835
rect 13435 -7955 13490 -7835
rect 13610 -7955 13655 -7835
rect 13775 -7955 13820 -7835
rect 13940 -7955 13985 -7835
rect 14105 -7955 14160 -7835
rect 14280 -7955 14325 -7835
rect 14445 -7955 14490 -7835
rect 14610 -7955 14655 -7835
rect 14775 -7955 14830 -7835
rect 14950 -7955 14995 -7835
rect 15115 -7955 15160 -7835
rect 15280 -7955 15325 -7835
rect 15445 -7955 15500 -7835
rect 15620 -7955 15665 -7835
rect 15785 -7955 15830 -7835
rect 15950 -7955 15995 -7835
rect 16115 -7955 16170 -7835
rect 16290 -7955 16335 -7835
rect 16455 -7955 16500 -7835
rect 16620 -7955 16665 -7835
rect 16785 -7955 16840 -7835
rect 16960 -7955 17005 -7835
rect 17125 -7955 17170 -7835
rect 17290 -7955 17335 -7835
rect 17455 -7955 17510 -7835
rect 17630 -7955 17675 -7835
rect 17795 -7955 17840 -7835
rect 17960 -7955 18005 -7835
rect 18125 -7955 18180 -7835
rect 18300 -7955 18310 -7835
rect 12810 -8000 18310 -7955
rect 12810 -8120 12820 -8000
rect 12940 -8120 12985 -8000
rect 13105 -8120 13150 -8000
rect 13270 -8120 13315 -8000
rect 13435 -8120 13490 -8000
rect 13610 -8120 13655 -8000
rect 13775 -8120 13820 -8000
rect 13940 -8120 13985 -8000
rect 14105 -8120 14160 -8000
rect 14280 -8120 14325 -8000
rect 14445 -8120 14490 -8000
rect 14610 -8120 14655 -8000
rect 14775 -8120 14830 -8000
rect 14950 -8120 14995 -8000
rect 15115 -8120 15160 -8000
rect 15280 -8120 15325 -8000
rect 15445 -8120 15500 -8000
rect 15620 -8120 15665 -8000
rect 15785 -8120 15830 -8000
rect 15950 -8120 15995 -8000
rect 16115 -8120 16170 -8000
rect 16290 -8120 16335 -8000
rect 16455 -8120 16500 -8000
rect 16620 -8120 16665 -8000
rect 16785 -8120 16840 -8000
rect 16960 -8120 17005 -8000
rect 17125 -8120 17170 -8000
rect 17290 -8120 17335 -8000
rect 17455 -8120 17510 -8000
rect 17630 -8120 17675 -8000
rect 17795 -8120 17840 -8000
rect 17960 -8120 18005 -8000
rect 18125 -8120 18180 -8000
rect 18300 -8120 18310 -8000
rect 12810 -8165 18310 -8120
rect 12810 -8285 12820 -8165
rect 12940 -8285 12985 -8165
rect 13105 -8285 13150 -8165
rect 13270 -8285 13315 -8165
rect 13435 -8285 13490 -8165
rect 13610 -8285 13655 -8165
rect 13775 -8285 13820 -8165
rect 13940 -8285 13985 -8165
rect 14105 -8285 14160 -8165
rect 14280 -8285 14325 -8165
rect 14445 -8285 14490 -8165
rect 14610 -8285 14655 -8165
rect 14775 -8285 14830 -8165
rect 14950 -8285 14995 -8165
rect 15115 -8285 15160 -8165
rect 15280 -8285 15325 -8165
rect 15445 -8285 15500 -8165
rect 15620 -8285 15665 -8165
rect 15785 -8285 15830 -8165
rect 15950 -8285 15995 -8165
rect 16115 -8285 16170 -8165
rect 16290 -8285 16335 -8165
rect 16455 -8285 16500 -8165
rect 16620 -8285 16665 -8165
rect 16785 -8285 16840 -8165
rect 16960 -8285 17005 -8165
rect 17125 -8285 17170 -8165
rect 17290 -8285 17335 -8165
rect 17455 -8285 17510 -8165
rect 17630 -8285 17675 -8165
rect 17795 -8285 17840 -8165
rect 17960 -8285 18005 -8165
rect 18125 -8285 18180 -8165
rect 18300 -8285 18310 -8165
rect 12810 -8330 18310 -8285
rect 12810 -8450 12820 -8330
rect 12940 -8450 12985 -8330
rect 13105 -8450 13150 -8330
rect 13270 -8450 13315 -8330
rect 13435 -8450 13490 -8330
rect 13610 -8450 13655 -8330
rect 13775 -8450 13820 -8330
rect 13940 -8450 13985 -8330
rect 14105 -8450 14160 -8330
rect 14280 -8450 14325 -8330
rect 14445 -8450 14490 -8330
rect 14610 -8450 14655 -8330
rect 14775 -8450 14830 -8330
rect 14950 -8450 14995 -8330
rect 15115 -8450 15160 -8330
rect 15280 -8450 15325 -8330
rect 15445 -8450 15500 -8330
rect 15620 -8450 15665 -8330
rect 15785 -8450 15830 -8330
rect 15950 -8450 15995 -8330
rect 16115 -8450 16170 -8330
rect 16290 -8450 16335 -8330
rect 16455 -8450 16500 -8330
rect 16620 -8450 16665 -8330
rect 16785 -8450 16840 -8330
rect 16960 -8450 17005 -8330
rect 17125 -8450 17170 -8330
rect 17290 -8450 17335 -8330
rect 17455 -8450 17510 -8330
rect 17630 -8450 17675 -8330
rect 17795 -8450 17840 -8330
rect 17960 -8450 18005 -8330
rect 18125 -8450 18180 -8330
rect 18300 -8450 18310 -8330
rect 12810 -8505 18310 -8450
rect 12810 -8625 12820 -8505
rect 12940 -8625 12985 -8505
rect 13105 -8625 13150 -8505
rect 13270 -8625 13315 -8505
rect 13435 -8625 13490 -8505
rect 13610 -8625 13655 -8505
rect 13775 -8625 13820 -8505
rect 13940 -8625 13985 -8505
rect 14105 -8625 14160 -8505
rect 14280 -8625 14325 -8505
rect 14445 -8625 14490 -8505
rect 14610 -8625 14655 -8505
rect 14775 -8625 14830 -8505
rect 14950 -8625 14995 -8505
rect 15115 -8625 15160 -8505
rect 15280 -8625 15325 -8505
rect 15445 -8625 15500 -8505
rect 15620 -8625 15665 -8505
rect 15785 -8625 15830 -8505
rect 15950 -8625 15995 -8505
rect 16115 -8625 16170 -8505
rect 16290 -8625 16335 -8505
rect 16455 -8625 16500 -8505
rect 16620 -8625 16665 -8505
rect 16785 -8625 16840 -8505
rect 16960 -8625 17005 -8505
rect 17125 -8625 17170 -8505
rect 17290 -8625 17335 -8505
rect 17455 -8625 17510 -8505
rect 17630 -8625 17675 -8505
rect 17795 -8625 17840 -8505
rect 17960 -8625 18005 -8505
rect 18125 -8625 18180 -8505
rect 18300 -8625 18310 -8505
rect 12810 -8670 18310 -8625
rect 12810 -8790 12820 -8670
rect 12940 -8790 12985 -8670
rect 13105 -8790 13150 -8670
rect 13270 -8790 13315 -8670
rect 13435 -8790 13490 -8670
rect 13610 -8790 13655 -8670
rect 13775 -8790 13820 -8670
rect 13940 -8790 13985 -8670
rect 14105 -8790 14160 -8670
rect 14280 -8790 14325 -8670
rect 14445 -8790 14490 -8670
rect 14610 -8790 14655 -8670
rect 14775 -8790 14830 -8670
rect 14950 -8790 14995 -8670
rect 15115 -8790 15160 -8670
rect 15280 -8790 15325 -8670
rect 15445 -8790 15500 -8670
rect 15620 -8790 15665 -8670
rect 15785 -8790 15830 -8670
rect 15950 -8790 15995 -8670
rect 16115 -8790 16170 -8670
rect 16290 -8790 16335 -8670
rect 16455 -8790 16500 -8670
rect 16620 -8790 16665 -8670
rect 16785 -8790 16840 -8670
rect 16960 -8790 17005 -8670
rect 17125 -8790 17170 -8670
rect 17290 -8790 17335 -8670
rect 17455 -8790 17510 -8670
rect 17630 -8790 17675 -8670
rect 17795 -8790 17840 -8670
rect 17960 -8790 18005 -8670
rect 18125 -8790 18180 -8670
rect 18300 -8790 18310 -8670
rect 12810 -8835 18310 -8790
rect 12810 -8955 12820 -8835
rect 12940 -8955 12985 -8835
rect 13105 -8955 13150 -8835
rect 13270 -8955 13315 -8835
rect 13435 -8955 13490 -8835
rect 13610 -8955 13655 -8835
rect 13775 -8955 13820 -8835
rect 13940 -8955 13985 -8835
rect 14105 -8955 14160 -8835
rect 14280 -8955 14325 -8835
rect 14445 -8955 14490 -8835
rect 14610 -8955 14655 -8835
rect 14775 -8955 14830 -8835
rect 14950 -8955 14995 -8835
rect 15115 -8955 15160 -8835
rect 15280 -8955 15325 -8835
rect 15445 -8955 15500 -8835
rect 15620 -8955 15665 -8835
rect 15785 -8955 15830 -8835
rect 15950 -8955 15995 -8835
rect 16115 -8955 16170 -8835
rect 16290 -8955 16335 -8835
rect 16455 -8955 16500 -8835
rect 16620 -8955 16665 -8835
rect 16785 -8955 16840 -8835
rect 16960 -8955 17005 -8835
rect 17125 -8955 17170 -8835
rect 17290 -8955 17335 -8835
rect 17455 -8955 17510 -8835
rect 17630 -8955 17675 -8835
rect 17795 -8955 17840 -8835
rect 17960 -8955 18005 -8835
rect 18125 -8955 18180 -8835
rect 18300 -8955 18310 -8835
rect 12810 -9000 18310 -8955
rect 12810 -9120 12820 -9000
rect 12940 -9120 12985 -9000
rect 13105 -9120 13150 -9000
rect 13270 -9120 13315 -9000
rect 13435 -9120 13490 -9000
rect 13610 -9120 13655 -9000
rect 13775 -9120 13820 -9000
rect 13940 -9120 13985 -9000
rect 14105 -9120 14160 -9000
rect 14280 -9120 14325 -9000
rect 14445 -9120 14490 -9000
rect 14610 -9120 14655 -9000
rect 14775 -9120 14830 -9000
rect 14950 -9120 14995 -9000
rect 15115 -9120 15160 -9000
rect 15280 -9120 15325 -9000
rect 15445 -9120 15500 -9000
rect 15620 -9120 15665 -9000
rect 15785 -9120 15830 -9000
rect 15950 -9120 15995 -9000
rect 16115 -9120 16170 -9000
rect 16290 -9120 16335 -9000
rect 16455 -9120 16500 -9000
rect 16620 -9120 16665 -9000
rect 16785 -9120 16840 -9000
rect 16960 -9120 17005 -9000
rect 17125 -9120 17170 -9000
rect 17290 -9120 17335 -9000
rect 17455 -9120 17510 -9000
rect 17630 -9120 17675 -9000
rect 17795 -9120 17840 -9000
rect 17960 -9120 18005 -9000
rect 18125 -9120 18180 -9000
rect 18300 -9120 18310 -9000
rect 12810 -9175 18310 -9120
rect 12810 -9295 12820 -9175
rect 12940 -9295 12985 -9175
rect 13105 -9295 13150 -9175
rect 13270 -9295 13315 -9175
rect 13435 -9295 13490 -9175
rect 13610 -9295 13655 -9175
rect 13775 -9295 13820 -9175
rect 13940 -9295 13985 -9175
rect 14105 -9295 14160 -9175
rect 14280 -9295 14325 -9175
rect 14445 -9295 14490 -9175
rect 14610 -9295 14655 -9175
rect 14775 -9295 14830 -9175
rect 14950 -9295 14995 -9175
rect 15115 -9295 15160 -9175
rect 15280 -9295 15325 -9175
rect 15445 -9295 15500 -9175
rect 15620 -9295 15665 -9175
rect 15785 -9295 15830 -9175
rect 15950 -9295 15995 -9175
rect 16115 -9295 16170 -9175
rect 16290 -9295 16335 -9175
rect 16455 -9295 16500 -9175
rect 16620 -9295 16665 -9175
rect 16785 -9295 16840 -9175
rect 16960 -9295 17005 -9175
rect 17125 -9295 17170 -9175
rect 17290 -9295 17335 -9175
rect 17455 -9295 17510 -9175
rect 17630 -9295 17675 -9175
rect 17795 -9295 17840 -9175
rect 17960 -9295 18005 -9175
rect 18125 -9295 18180 -9175
rect 18300 -9295 18310 -9175
rect 12810 -9340 18310 -9295
rect 12810 -9460 12820 -9340
rect 12940 -9460 12985 -9340
rect 13105 -9460 13150 -9340
rect 13270 -9460 13315 -9340
rect 13435 -9460 13490 -9340
rect 13610 -9460 13655 -9340
rect 13775 -9460 13820 -9340
rect 13940 -9460 13985 -9340
rect 14105 -9460 14160 -9340
rect 14280 -9460 14325 -9340
rect 14445 -9460 14490 -9340
rect 14610 -9460 14655 -9340
rect 14775 -9460 14830 -9340
rect 14950 -9460 14995 -9340
rect 15115 -9460 15160 -9340
rect 15280 -9460 15325 -9340
rect 15445 -9460 15500 -9340
rect 15620 -9460 15665 -9340
rect 15785 -9460 15830 -9340
rect 15950 -9460 15995 -9340
rect 16115 -9460 16170 -9340
rect 16290 -9460 16335 -9340
rect 16455 -9460 16500 -9340
rect 16620 -9460 16665 -9340
rect 16785 -9460 16840 -9340
rect 16960 -9460 17005 -9340
rect 17125 -9460 17170 -9340
rect 17290 -9460 17335 -9340
rect 17455 -9460 17510 -9340
rect 17630 -9460 17675 -9340
rect 17795 -9460 17840 -9340
rect 17960 -9460 18005 -9340
rect 18125 -9460 18180 -9340
rect 18300 -9460 18310 -9340
rect 12810 -9505 18310 -9460
rect 12810 -9625 12820 -9505
rect 12940 -9625 12985 -9505
rect 13105 -9625 13150 -9505
rect 13270 -9625 13315 -9505
rect 13435 -9625 13490 -9505
rect 13610 -9625 13655 -9505
rect 13775 -9625 13820 -9505
rect 13940 -9625 13985 -9505
rect 14105 -9625 14160 -9505
rect 14280 -9625 14325 -9505
rect 14445 -9625 14490 -9505
rect 14610 -9625 14655 -9505
rect 14775 -9625 14830 -9505
rect 14950 -9625 14995 -9505
rect 15115 -9625 15160 -9505
rect 15280 -9625 15325 -9505
rect 15445 -9625 15500 -9505
rect 15620 -9625 15665 -9505
rect 15785 -9625 15830 -9505
rect 15950 -9625 15995 -9505
rect 16115 -9625 16170 -9505
rect 16290 -9625 16335 -9505
rect 16455 -9625 16500 -9505
rect 16620 -9625 16665 -9505
rect 16785 -9625 16840 -9505
rect 16960 -9625 17005 -9505
rect 17125 -9625 17170 -9505
rect 17290 -9625 17335 -9505
rect 17455 -9625 17510 -9505
rect 17630 -9625 17675 -9505
rect 17795 -9625 17840 -9505
rect 17960 -9625 18005 -9505
rect 18125 -9625 18180 -9505
rect 18300 -9625 18310 -9505
rect 12810 -9670 18310 -9625
rect 12810 -9790 12820 -9670
rect 12940 -9790 12985 -9670
rect 13105 -9790 13150 -9670
rect 13270 -9790 13315 -9670
rect 13435 -9790 13490 -9670
rect 13610 -9790 13655 -9670
rect 13775 -9790 13820 -9670
rect 13940 -9790 13985 -9670
rect 14105 -9790 14160 -9670
rect 14280 -9790 14325 -9670
rect 14445 -9790 14490 -9670
rect 14610 -9790 14655 -9670
rect 14775 -9790 14830 -9670
rect 14950 -9790 14995 -9670
rect 15115 -9790 15160 -9670
rect 15280 -9790 15325 -9670
rect 15445 -9790 15500 -9670
rect 15620 -9790 15665 -9670
rect 15785 -9790 15830 -9670
rect 15950 -9790 15995 -9670
rect 16115 -9790 16170 -9670
rect 16290 -9790 16335 -9670
rect 16455 -9790 16500 -9670
rect 16620 -9790 16665 -9670
rect 16785 -9790 16840 -9670
rect 16960 -9790 17005 -9670
rect 17125 -9790 17170 -9670
rect 17290 -9790 17335 -9670
rect 17455 -9790 17510 -9670
rect 17630 -9790 17675 -9670
rect 17795 -9790 17840 -9670
rect 17960 -9790 18005 -9670
rect 18125 -9790 18180 -9670
rect 18300 -9790 18310 -9670
rect 12810 -9800 18310 -9790
rect 18500 -4310 24000 -4300
rect 18500 -4430 18510 -4310
rect 18630 -4430 18675 -4310
rect 18795 -4430 18840 -4310
rect 18960 -4430 19005 -4310
rect 19125 -4430 19180 -4310
rect 19300 -4430 19345 -4310
rect 19465 -4430 19510 -4310
rect 19630 -4430 19675 -4310
rect 19795 -4430 19850 -4310
rect 19970 -4430 20015 -4310
rect 20135 -4430 20180 -4310
rect 20300 -4430 20345 -4310
rect 20465 -4430 20520 -4310
rect 20640 -4430 20685 -4310
rect 20805 -4430 20850 -4310
rect 20970 -4430 21015 -4310
rect 21135 -4430 21190 -4310
rect 21310 -4430 21355 -4310
rect 21475 -4430 21520 -4310
rect 21640 -4430 21685 -4310
rect 21805 -4430 21860 -4310
rect 21980 -4430 22025 -4310
rect 22145 -4430 22190 -4310
rect 22310 -4430 22355 -4310
rect 22475 -4430 22530 -4310
rect 22650 -4430 22695 -4310
rect 22815 -4430 22860 -4310
rect 22980 -4430 23025 -4310
rect 23145 -4430 23200 -4310
rect 23320 -4430 23365 -4310
rect 23485 -4430 23530 -4310
rect 23650 -4430 23695 -4310
rect 23815 -4430 23870 -4310
rect 23990 -4430 24000 -4310
rect 18500 -4485 24000 -4430
rect 18500 -4605 18510 -4485
rect 18630 -4605 18675 -4485
rect 18795 -4605 18840 -4485
rect 18960 -4605 19005 -4485
rect 19125 -4605 19180 -4485
rect 19300 -4605 19345 -4485
rect 19465 -4605 19510 -4485
rect 19630 -4605 19675 -4485
rect 19795 -4605 19850 -4485
rect 19970 -4605 20015 -4485
rect 20135 -4605 20180 -4485
rect 20300 -4605 20345 -4485
rect 20465 -4605 20520 -4485
rect 20640 -4605 20685 -4485
rect 20805 -4605 20850 -4485
rect 20970 -4605 21015 -4485
rect 21135 -4605 21190 -4485
rect 21310 -4605 21355 -4485
rect 21475 -4605 21520 -4485
rect 21640 -4605 21685 -4485
rect 21805 -4605 21860 -4485
rect 21980 -4605 22025 -4485
rect 22145 -4605 22190 -4485
rect 22310 -4605 22355 -4485
rect 22475 -4605 22530 -4485
rect 22650 -4605 22695 -4485
rect 22815 -4605 22860 -4485
rect 22980 -4605 23025 -4485
rect 23145 -4605 23200 -4485
rect 23320 -4605 23365 -4485
rect 23485 -4605 23530 -4485
rect 23650 -4605 23695 -4485
rect 23815 -4605 23870 -4485
rect 23990 -4605 24000 -4485
rect 18500 -4650 24000 -4605
rect 18500 -4770 18510 -4650
rect 18630 -4770 18675 -4650
rect 18795 -4770 18840 -4650
rect 18960 -4770 19005 -4650
rect 19125 -4770 19180 -4650
rect 19300 -4770 19345 -4650
rect 19465 -4770 19510 -4650
rect 19630 -4770 19675 -4650
rect 19795 -4770 19850 -4650
rect 19970 -4770 20015 -4650
rect 20135 -4770 20180 -4650
rect 20300 -4770 20345 -4650
rect 20465 -4770 20520 -4650
rect 20640 -4770 20685 -4650
rect 20805 -4770 20850 -4650
rect 20970 -4770 21015 -4650
rect 21135 -4770 21190 -4650
rect 21310 -4770 21355 -4650
rect 21475 -4770 21520 -4650
rect 21640 -4770 21685 -4650
rect 21805 -4770 21860 -4650
rect 21980 -4770 22025 -4650
rect 22145 -4770 22190 -4650
rect 22310 -4770 22355 -4650
rect 22475 -4770 22530 -4650
rect 22650 -4770 22695 -4650
rect 22815 -4770 22860 -4650
rect 22980 -4770 23025 -4650
rect 23145 -4770 23200 -4650
rect 23320 -4770 23365 -4650
rect 23485 -4770 23530 -4650
rect 23650 -4770 23695 -4650
rect 23815 -4770 23870 -4650
rect 23990 -4770 24000 -4650
rect 18500 -4815 24000 -4770
rect 18500 -4935 18510 -4815
rect 18630 -4935 18675 -4815
rect 18795 -4935 18840 -4815
rect 18960 -4935 19005 -4815
rect 19125 -4935 19180 -4815
rect 19300 -4935 19345 -4815
rect 19465 -4935 19510 -4815
rect 19630 -4935 19675 -4815
rect 19795 -4935 19850 -4815
rect 19970 -4935 20015 -4815
rect 20135 -4935 20180 -4815
rect 20300 -4935 20345 -4815
rect 20465 -4935 20520 -4815
rect 20640 -4935 20685 -4815
rect 20805 -4935 20850 -4815
rect 20970 -4935 21015 -4815
rect 21135 -4935 21190 -4815
rect 21310 -4935 21355 -4815
rect 21475 -4935 21520 -4815
rect 21640 -4935 21685 -4815
rect 21805 -4935 21860 -4815
rect 21980 -4935 22025 -4815
rect 22145 -4935 22190 -4815
rect 22310 -4935 22355 -4815
rect 22475 -4935 22530 -4815
rect 22650 -4935 22695 -4815
rect 22815 -4935 22860 -4815
rect 22980 -4935 23025 -4815
rect 23145 -4935 23200 -4815
rect 23320 -4935 23365 -4815
rect 23485 -4935 23530 -4815
rect 23650 -4935 23695 -4815
rect 23815 -4935 23870 -4815
rect 23990 -4935 24000 -4815
rect 18500 -4980 24000 -4935
rect 18500 -5100 18510 -4980
rect 18630 -5100 18675 -4980
rect 18795 -5100 18840 -4980
rect 18960 -5100 19005 -4980
rect 19125 -5100 19180 -4980
rect 19300 -5100 19345 -4980
rect 19465 -5100 19510 -4980
rect 19630 -5100 19675 -4980
rect 19795 -5100 19850 -4980
rect 19970 -5100 20015 -4980
rect 20135 -5100 20180 -4980
rect 20300 -5100 20345 -4980
rect 20465 -5100 20520 -4980
rect 20640 -5100 20685 -4980
rect 20805 -5100 20850 -4980
rect 20970 -5100 21015 -4980
rect 21135 -5100 21190 -4980
rect 21310 -5100 21355 -4980
rect 21475 -5100 21520 -4980
rect 21640 -5100 21685 -4980
rect 21805 -5100 21860 -4980
rect 21980 -5100 22025 -4980
rect 22145 -5100 22190 -4980
rect 22310 -5100 22355 -4980
rect 22475 -5100 22530 -4980
rect 22650 -5100 22695 -4980
rect 22815 -5100 22860 -4980
rect 22980 -5100 23025 -4980
rect 23145 -5100 23200 -4980
rect 23320 -5100 23365 -4980
rect 23485 -5100 23530 -4980
rect 23650 -5100 23695 -4980
rect 23815 -5100 23870 -4980
rect 23990 -5100 24000 -4980
rect 18500 -5155 24000 -5100
rect 18500 -5275 18510 -5155
rect 18630 -5275 18675 -5155
rect 18795 -5275 18840 -5155
rect 18960 -5275 19005 -5155
rect 19125 -5275 19180 -5155
rect 19300 -5275 19345 -5155
rect 19465 -5275 19510 -5155
rect 19630 -5275 19675 -5155
rect 19795 -5275 19850 -5155
rect 19970 -5275 20015 -5155
rect 20135 -5275 20180 -5155
rect 20300 -5275 20345 -5155
rect 20465 -5275 20520 -5155
rect 20640 -5275 20685 -5155
rect 20805 -5275 20850 -5155
rect 20970 -5275 21015 -5155
rect 21135 -5275 21190 -5155
rect 21310 -5275 21355 -5155
rect 21475 -5275 21520 -5155
rect 21640 -5275 21685 -5155
rect 21805 -5275 21860 -5155
rect 21980 -5275 22025 -5155
rect 22145 -5275 22190 -5155
rect 22310 -5275 22355 -5155
rect 22475 -5275 22530 -5155
rect 22650 -5275 22695 -5155
rect 22815 -5275 22860 -5155
rect 22980 -5275 23025 -5155
rect 23145 -5275 23200 -5155
rect 23320 -5275 23365 -5155
rect 23485 -5275 23530 -5155
rect 23650 -5275 23695 -5155
rect 23815 -5275 23870 -5155
rect 23990 -5275 24000 -5155
rect 18500 -5320 24000 -5275
rect 18500 -5440 18510 -5320
rect 18630 -5440 18675 -5320
rect 18795 -5440 18840 -5320
rect 18960 -5440 19005 -5320
rect 19125 -5440 19180 -5320
rect 19300 -5440 19345 -5320
rect 19465 -5440 19510 -5320
rect 19630 -5440 19675 -5320
rect 19795 -5440 19850 -5320
rect 19970 -5440 20015 -5320
rect 20135 -5440 20180 -5320
rect 20300 -5440 20345 -5320
rect 20465 -5440 20520 -5320
rect 20640 -5440 20685 -5320
rect 20805 -5440 20850 -5320
rect 20970 -5440 21015 -5320
rect 21135 -5440 21190 -5320
rect 21310 -5440 21355 -5320
rect 21475 -5440 21520 -5320
rect 21640 -5440 21685 -5320
rect 21805 -5440 21860 -5320
rect 21980 -5440 22025 -5320
rect 22145 -5440 22190 -5320
rect 22310 -5440 22355 -5320
rect 22475 -5440 22530 -5320
rect 22650 -5440 22695 -5320
rect 22815 -5440 22860 -5320
rect 22980 -5440 23025 -5320
rect 23145 -5440 23200 -5320
rect 23320 -5440 23365 -5320
rect 23485 -5440 23530 -5320
rect 23650 -5440 23695 -5320
rect 23815 -5440 23870 -5320
rect 23990 -5440 24000 -5320
rect 18500 -5485 24000 -5440
rect 18500 -5605 18510 -5485
rect 18630 -5605 18675 -5485
rect 18795 -5605 18840 -5485
rect 18960 -5605 19005 -5485
rect 19125 -5605 19180 -5485
rect 19300 -5605 19345 -5485
rect 19465 -5605 19510 -5485
rect 19630 -5605 19675 -5485
rect 19795 -5605 19850 -5485
rect 19970 -5605 20015 -5485
rect 20135 -5605 20180 -5485
rect 20300 -5605 20345 -5485
rect 20465 -5605 20520 -5485
rect 20640 -5605 20685 -5485
rect 20805 -5605 20850 -5485
rect 20970 -5605 21015 -5485
rect 21135 -5605 21190 -5485
rect 21310 -5605 21355 -5485
rect 21475 -5605 21520 -5485
rect 21640 -5605 21685 -5485
rect 21805 -5605 21860 -5485
rect 21980 -5605 22025 -5485
rect 22145 -5605 22190 -5485
rect 22310 -5605 22355 -5485
rect 22475 -5605 22530 -5485
rect 22650 -5605 22695 -5485
rect 22815 -5605 22860 -5485
rect 22980 -5605 23025 -5485
rect 23145 -5605 23200 -5485
rect 23320 -5605 23365 -5485
rect 23485 -5605 23530 -5485
rect 23650 -5605 23695 -5485
rect 23815 -5605 23870 -5485
rect 23990 -5605 24000 -5485
rect 18500 -5650 24000 -5605
rect 18500 -5770 18510 -5650
rect 18630 -5770 18675 -5650
rect 18795 -5770 18840 -5650
rect 18960 -5770 19005 -5650
rect 19125 -5770 19180 -5650
rect 19300 -5770 19345 -5650
rect 19465 -5770 19510 -5650
rect 19630 -5770 19675 -5650
rect 19795 -5770 19850 -5650
rect 19970 -5770 20015 -5650
rect 20135 -5770 20180 -5650
rect 20300 -5770 20345 -5650
rect 20465 -5770 20520 -5650
rect 20640 -5770 20685 -5650
rect 20805 -5770 20850 -5650
rect 20970 -5770 21015 -5650
rect 21135 -5770 21190 -5650
rect 21310 -5770 21355 -5650
rect 21475 -5770 21520 -5650
rect 21640 -5770 21685 -5650
rect 21805 -5770 21860 -5650
rect 21980 -5770 22025 -5650
rect 22145 -5770 22190 -5650
rect 22310 -5770 22355 -5650
rect 22475 -5770 22530 -5650
rect 22650 -5770 22695 -5650
rect 22815 -5770 22860 -5650
rect 22980 -5770 23025 -5650
rect 23145 -5770 23200 -5650
rect 23320 -5770 23365 -5650
rect 23485 -5770 23530 -5650
rect 23650 -5770 23695 -5650
rect 23815 -5770 23870 -5650
rect 23990 -5770 24000 -5650
rect 18500 -5825 24000 -5770
rect 18500 -5945 18510 -5825
rect 18630 -5945 18675 -5825
rect 18795 -5945 18840 -5825
rect 18960 -5945 19005 -5825
rect 19125 -5945 19180 -5825
rect 19300 -5945 19345 -5825
rect 19465 -5945 19510 -5825
rect 19630 -5945 19675 -5825
rect 19795 -5945 19850 -5825
rect 19970 -5945 20015 -5825
rect 20135 -5945 20180 -5825
rect 20300 -5945 20345 -5825
rect 20465 -5945 20520 -5825
rect 20640 -5945 20685 -5825
rect 20805 -5945 20850 -5825
rect 20970 -5945 21015 -5825
rect 21135 -5945 21190 -5825
rect 21310 -5945 21355 -5825
rect 21475 -5945 21520 -5825
rect 21640 -5945 21685 -5825
rect 21805 -5945 21860 -5825
rect 21980 -5945 22025 -5825
rect 22145 -5945 22190 -5825
rect 22310 -5945 22355 -5825
rect 22475 -5945 22530 -5825
rect 22650 -5945 22695 -5825
rect 22815 -5945 22860 -5825
rect 22980 -5945 23025 -5825
rect 23145 -5945 23200 -5825
rect 23320 -5945 23365 -5825
rect 23485 -5945 23530 -5825
rect 23650 -5945 23695 -5825
rect 23815 -5945 23870 -5825
rect 23990 -5945 24000 -5825
rect 18500 -5990 24000 -5945
rect 18500 -6110 18510 -5990
rect 18630 -6110 18675 -5990
rect 18795 -6110 18840 -5990
rect 18960 -6110 19005 -5990
rect 19125 -6110 19180 -5990
rect 19300 -6110 19345 -5990
rect 19465 -6110 19510 -5990
rect 19630 -6110 19675 -5990
rect 19795 -6110 19850 -5990
rect 19970 -6110 20015 -5990
rect 20135 -6110 20180 -5990
rect 20300 -6110 20345 -5990
rect 20465 -6110 20520 -5990
rect 20640 -6110 20685 -5990
rect 20805 -6110 20850 -5990
rect 20970 -6110 21015 -5990
rect 21135 -6110 21190 -5990
rect 21310 -6110 21355 -5990
rect 21475 -6110 21520 -5990
rect 21640 -6110 21685 -5990
rect 21805 -6110 21860 -5990
rect 21980 -6110 22025 -5990
rect 22145 -6110 22190 -5990
rect 22310 -6110 22355 -5990
rect 22475 -6110 22530 -5990
rect 22650 -6110 22695 -5990
rect 22815 -6110 22860 -5990
rect 22980 -6110 23025 -5990
rect 23145 -6110 23200 -5990
rect 23320 -6110 23365 -5990
rect 23485 -6110 23530 -5990
rect 23650 -6110 23695 -5990
rect 23815 -6110 23870 -5990
rect 23990 -6110 24000 -5990
rect 18500 -6155 24000 -6110
rect 18500 -6275 18510 -6155
rect 18630 -6275 18675 -6155
rect 18795 -6275 18840 -6155
rect 18960 -6275 19005 -6155
rect 19125 -6275 19180 -6155
rect 19300 -6275 19345 -6155
rect 19465 -6275 19510 -6155
rect 19630 -6275 19675 -6155
rect 19795 -6275 19850 -6155
rect 19970 -6275 20015 -6155
rect 20135 -6275 20180 -6155
rect 20300 -6275 20345 -6155
rect 20465 -6275 20520 -6155
rect 20640 -6275 20685 -6155
rect 20805 -6275 20850 -6155
rect 20970 -6275 21015 -6155
rect 21135 -6275 21190 -6155
rect 21310 -6275 21355 -6155
rect 21475 -6275 21520 -6155
rect 21640 -6275 21685 -6155
rect 21805 -6275 21860 -6155
rect 21980 -6275 22025 -6155
rect 22145 -6275 22190 -6155
rect 22310 -6275 22355 -6155
rect 22475 -6275 22530 -6155
rect 22650 -6275 22695 -6155
rect 22815 -6275 22860 -6155
rect 22980 -6275 23025 -6155
rect 23145 -6275 23200 -6155
rect 23320 -6275 23365 -6155
rect 23485 -6275 23530 -6155
rect 23650 -6275 23695 -6155
rect 23815 -6275 23870 -6155
rect 23990 -6275 24000 -6155
rect 18500 -6320 24000 -6275
rect 18500 -6440 18510 -6320
rect 18630 -6440 18675 -6320
rect 18795 -6440 18840 -6320
rect 18960 -6440 19005 -6320
rect 19125 -6440 19180 -6320
rect 19300 -6440 19345 -6320
rect 19465 -6440 19510 -6320
rect 19630 -6440 19675 -6320
rect 19795 -6440 19850 -6320
rect 19970 -6440 20015 -6320
rect 20135 -6440 20180 -6320
rect 20300 -6440 20345 -6320
rect 20465 -6440 20520 -6320
rect 20640 -6440 20685 -6320
rect 20805 -6440 20850 -6320
rect 20970 -6440 21015 -6320
rect 21135 -6440 21190 -6320
rect 21310 -6440 21355 -6320
rect 21475 -6440 21520 -6320
rect 21640 -6440 21685 -6320
rect 21805 -6440 21860 -6320
rect 21980 -6440 22025 -6320
rect 22145 -6440 22190 -6320
rect 22310 -6440 22355 -6320
rect 22475 -6440 22530 -6320
rect 22650 -6440 22695 -6320
rect 22815 -6440 22860 -6320
rect 22980 -6440 23025 -6320
rect 23145 -6440 23200 -6320
rect 23320 -6440 23365 -6320
rect 23485 -6440 23530 -6320
rect 23650 -6440 23695 -6320
rect 23815 -6440 23870 -6320
rect 23990 -6440 24000 -6320
rect 18500 -6495 24000 -6440
rect 18500 -6615 18510 -6495
rect 18630 -6615 18675 -6495
rect 18795 -6615 18840 -6495
rect 18960 -6615 19005 -6495
rect 19125 -6615 19180 -6495
rect 19300 -6615 19345 -6495
rect 19465 -6615 19510 -6495
rect 19630 -6615 19675 -6495
rect 19795 -6615 19850 -6495
rect 19970 -6615 20015 -6495
rect 20135 -6615 20180 -6495
rect 20300 -6615 20345 -6495
rect 20465 -6615 20520 -6495
rect 20640 -6615 20685 -6495
rect 20805 -6615 20850 -6495
rect 20970 -6615 21015 -6495
rect 21135 -6615 21190 -6495
rect 21310 -6615 21355 -6495
rect 21475 -6615 21520 -6495
rect 21640 -6615 21685 -6495
rect 21805 -6615 21860 -6495
rect 21980 -6615 22025 -6495
rect 22145 -6615 22190 -6495
rect 22310 -6615 22355 -6495
rect 22475 -6615 22530 -6495
rect 22650 -6615 22695 -6495
rect 22815 -6615 22860 -6495
rect 22980 -6615 23025 -6495
rect 23145 -6615 23200 -6495
rect 23320 -6615 23365 -6495
rect 23485 -6615 23530 -6495
rect 23650 -6615 23695 -6495
rect 23815 -6615 23870 -6495
rect 23990 -6615 24000 -6495
rect 18500 -6660 24000 -6615
rect 18500 -6780 18510 -6660
rect 18630 -6780 18675 -6660
rect 18795 -6780 18840 -6660
rect 18960 -6780 19005 -6660
rect 19125 -6780 19180 -6660
rect 19300 -6780 19345 -6660
rect 19465 -6780 19510 -6660
rect 19630 -6780 19675 -6660
rect 19795 -6780 19850 -6660
rect 19970 -6780 20015 -6660
rect 20135 -6780 20180 -6660
rect 20300 -6780 20345 -6660
rect 20465 -6780 20520 -6660
rect 20640 -6780 20685 -6660
rect 20805 -6780 20850 -6660
rect 20970 -6780 21015 -6660
rect 21135 -6780 21190 -6660
rect 21310 -6780 21355 -6660
rect 21475 -6780 21520 -6660
rect 21640 -6780 21685 -6660
rect 21805 -6780 21860 -6660
rect 21980 -6780 22025 -6660
rect 22145 -6780 22190 -6660
rect 22310 -6780 22355 -6660
rect 22475 -6780 22530 -6660
rect 22650 -6780 22695 -6660
rect 22815 -6780 22860 -6660
rect 22980 -6780 23025 -6660
rect 23145 -6780 23200 -6660
rect 23320 -6780 23365 -6660
rect 23485 -6780 23530 -6660
rect 23650 -6780 23695 -6660
rect 23815 -6780 23870 -6660
rect 23990 -6780 24000 -6660
rect 18500 -6825 24000 -6780
rect 18500 -6945 18510 -6825
rect 18630 -6945 18675 -6825
rect 18795 -6945 18840 -6825
rect 18960 -6945 19005 -6825
rect 19125 -6945 19180 -6825
rect 19300 -6945 19345 -6825
rect 19465 -6945 19510 -6825
rect 19630 -6945 19675 -6825
rect 19795 -6945 19850 -6825
rect 19970 -6945 20015 -6825
rect 20135 -6945 20180 -6825
rect 20300 -6945 20345 -6825
rect 20465 -6945 20520 -6825
rect 20640 -6945 20685 -6825
rect 20805 -6945 20850 -6825
rect 20970 -6945 21015 -6825
rect 21135 -6945 21190 -6825
rect 21310 -6945 21355 -6825
rect 21475 -6945 21520 -6825
rect 21640 -6945 21685 -6825
rect 21805 -6945 21860 -6825
rect 21980 -6945 22025 -6825
rect 22145 -6945 22190 -6825
rect 22310 -6945 22355 -6825
rect 22475 -6945 22530 -6825
rect 22650 -6945 22695 -6825
rect 22815 -6945 22860 -6825
rect 22980 -6945 23025 -6825
rect 23145 -6945 23200 -6825
rect 23320 -6945 23365 -6825
rect 23485 -6945 23530 -6825
rect 23650 -6945 23695 -6825
rect 23815 -6945 23870 -6825
rect 23990 -6945 24000 -6825
rect 18500 -6990 24000 -6945
rect 18500 -7110 18510 -6990
rect 18630 -7110 18675 -6990
rect 18795 -7110 18840 -6990
rect 18960 -7110 19005 -6990
rect 19125 -7110 19180 -6990
rect 19300 -7110 19345 -6990
rect 19465 -7110 19510 -6990
rect 19630 -7110 19675 -6990
rect 19795 -7110 19850 -6990
rect 19970 -7110 20015 -6990
rect 20135 -7110 20180 -6990
rect 20300 -7110 20345 -6990
rect 20465 -7110 20520 -6990
rect 20640 -7110 20685 -6990
rect 20805 -7110 20850 -6990
rect 20970 -7110 21015 -6990
rect 21135 -7110 21190 -6990
rect 21310 -7110 21355 -6990
rect 21475 -7110 21520 -6990
rect 21640 -7110 21685 -6990
rect 21805 -7110 21860 -6990
rect 21980 -7110 22025 -6990
rect 22145 -7110 22190 -6990
rect 22310 -7110 22355 -6990
rect 22475 -7110 22530 -6990
rect 22650 -7110 22695 -6990
rect 22815 -7110 22860 -6990
rect 22980 -7110 23025 -6990
rect 23145 -7110 23200 -6990
rect 23320 -7110 23365 -6990
rect 23485 -7110 23530 -6990
rect 23650 -7110 23695 -6990
rect 23815 -7110 23870 -6990
rect 23990 -7110 24000 -6990
rect 18500 -7165 24000 -7110
rect 18500 -7285 18510 -7165
rect 18630 -7285 18675 -7165
rect 18795 -7285 18840 -7165
rect 18960 -7285 19005 -7165
rect 19125 -7285 19180 -7165
rect 19300 -7285 19345 -7165
rect 19465 -7285 19510 -7165
rect 19630 -7285 19675 -7165
rect 19795 -7285 19850 -7165
rect 19970 -7285 20015 -7165
rect 20135 -7285 20180 -7165
rect 20300 -7285 20345 -7165
rect 20465 -7285 20520 -7165
rect 20640 -7285 20685 -7165
rect 20805 -7285 20850 -7165
rect 20970 -7285 21015 -7165
rect 21135 -7285 21190 -7165
rect 21310 -7285 21355 -7165
rect 21475 -7285 21520 -7165
rect 21640 -7285 21685 -7165
rect 21805 -7285 21860 -7165
rect 21980 -7285 22025 -7165
rect 22145 -7285 22190 -7165
rect 22310 -7285 22355 -7165
rect 22475 -7285 22530 -7165
rect 22650 -7285 22695 -7165
rect 22815 -7285 22860 -7165
rect 22980 -7285 23025 -7165
rect 23145 -7285 23200 -7165
rect 23320 -7285 23365 -7165
rect 23485 -7285 23530 -7165
rect 23650 -7285 23695 -7165
rect 23815 -7285 23870 -7165
rect 23990 -7285 24000 -7165
rect 18500 -7330 24000 -7285
rect 18500 -7450 18510 -7330
rect 18630 -7450 18675 -7330
rect 18795 -7450 18840 -7330
rect 18960 -7450 19005 -7330
rect 19125 -7450 19180 -7330
rect 19300 -7450 19345 -7330
rect 19465 -7450 19510 -7330
rect 19630 -7450 19675 -7330
rect 19795 -7450 19850 -7330
rect 19970 -7450 20015 -7330
rect 20135 -7450 20180 -7330
rect 20300 -7450 20345 -7330
rect 20465 -7450 20520 -7330
rect 20640 -7450 20685 -7330
rect 20805 -7450 20850 -7330
rect 20970 -7450 21015 -7330
rect 21135 -7450 21190 -7330
rect 21310 -7450 21355 -7330
rect 21475 -7450 21520 -7330
rect 21640 -7450 21685 -7330
rect 21805 -7450 21860 -7330
rect 21980 -7450 22025 -7330
rect 22145 -7450 22190 -7330
rect 22310 -7450 22355 -7330
rect 22475 -7450 22530 -7330
rect 22650 -7450 22695 -7330
rect 22815 -7450 22860 -7330
rect 22980 -7450 23025 -7330
rect 23145 -7450 23200 -7330
rect 23320 -7450 23365 -7330
rect 23485 -7450 23530 -7330
rect 23650 -7450 23695 -7330
rect 23815 -7450 23870 -7330
rect 23990 -7450 24000 -7330
rect 18500 -7495 24000 -7450
rect 18500 -7615 18510 -7495
rect 18630 -7615 18675 -7495
rect 18795 -7615 18840 -7495
rect 18960 -7615 19005 -7495
rect 19125 -7615 19180 -7495
rect 19300 -7615 19345 -7495
rect 19465 -7615 19510 -7495
rect 19630 -7615 19675 -7495
rect 19795 -7615 19850 -7495
rect 19970 -7615 20015 -7495
rect 20135 -7615 20180 -7495
rect 20300 -7615 20345 -7495
rect 20465 -7615 20520 -7495
rect 20640 -7615 20685 -7495
rect 20805 -7615 20850 -7495
rect 20970 -7615 21015 -7495
rect 21135 -7615 21190 -7495
rect 21310 -7615 21355 -7495
rect 21475 -7615 21520 -7495
rect 21640 -7615 21685 -7495
rect 21805 -7615 21860 -7495
rect 21980 -7615 22025 -7495
rect 22145 -7615 22190 -7495
rect 22310 -7615 22355 -7495
rect 22475 -7615 22530 -7495
rect 22650 -7615 22695 -7495
rect 22815 -7615 22860 -7495
rect 22980 -7615 23025 -7495
rect 23145 -7615 23200 -7495
rect 23320 -7615 23365 -7495
rect 23485 -7615 23530 -7495
rect 23650 -7615 23695 -7495
rect 23815 -7615 23870 -7495
rect 23990 -7615 24000 -7495
rect 18500 -7660 24000 -7615
rect 18500 -7780 18510 -7660
rect 18630 -7780 18675 -7660
rect 18795 -7780 18840 -7660
rect 18960 -7780 19005 -7660
rect 19125 -7780 19180 -7660
rect 19300 -7780 19345 -7660
rect 19465 -7780 19510 -7660
rect 19630 -7780 19675 -7660
rect 19795 -7780 19850 -7660
rect 19970 -7780 20015 -7660
rect 20135 -7780 20180 -7660
rect 20300 -7780 20345 -7660
rect 20465 -7780 20520 -7660
rect 20640 -7780 20685 -7660
rect 20805 -7780 20850 -7660
rect 20970 -7780 21015 -7660
rect 21135 -7780 21190 -7660
rect 21310 -7780 21355 -7660
rect 21475 -7780 21520 -7660
rect 21640 -7780 21685 -7660
rect 21805 -7780 21860 -7660
rect 21980 -7780 22025 -7660
rect 22145 -7780 22190 -7660
rect 22310 -7780 22355 -7660
rect 22475 -7780 22530 -7660
rect 22650 -7780 22695 -7660
rect 22815 -7780 22860 -7660
rect 22980 -7780 23025 -7660
rect 23145 -7780 23200 -7660
rect 23320 -7780 23365 -7660
rect 23485 -7780 23530 -7660
rect 23650 -7780 23695 -7660
rect 23815 -7780 23870 -7660
rect 23990 -7780 24000 -7660
rect 18500 -7835 24000 -7780
rect 18500 -7955 18510 -7835
rect 18630 -7955 18675 -7835
rect 18795 -7955 18840 -7835
rect 18960 -7955 19005 -7835
rect 19125 -7955 19180 -7835
rect 19300 -7955 19345 -7835
rect 19465 -7955 19510 -7835
rect 19630 -7955 19675 -7835
rect 19795 -7955 19850 -7835
rect 19970 -7955 20015 -7835
rect 20135 -7955 20180 -7835
rect 20300 -7955 20345 -7835
rect 20465 -7955 20520 -7835
rect 20640 -7955 20685 -7835
rect 20805 -7955 20850 -7835
rect 20970 -7955 21015 -7835
rect 21135 -7955 21190 -7835
rect 21310 -7955 21355 -7835
rect 21475 -7955 21520 -7835
rect 21640 -7955 21685 -7835
rect 21805 -7955 21860 -7835
rect 21980 -7955 22025 -7835
rect 22145 -7955 22190 -7835
rect 22310 -7955 22355 -7835
rect 22475 -7955 22530 -7835
rect 22650 -7955 22695 -7835
rect 22815 -7955 22860 -7835
rect 22980 -7955 23025 -7835
rect 23145 -7955 23200 -7835
rect 23320 -7955 23365 -7835
rect 23485 -7955 23530 -7835
rect 23650 -7955 23695 -7835
rect 23815 -7955 23870 -7835
rect 23990 -7955 24000 -7835
rect 18500 -8000 24000 -7955
rect 18500 -8120 18510 -8000
rect 18630 -8120 18675 -8000
rect 18795 -8120 18840 -8000
rect 18960 -8120 19005 -8000
rect 19125 -8120 19180 -8000
rect 19300 -8120 19345 -8000
rect 19465 -8120 19510 -8000
rect 19630 -8120 19675 -8000
rect 19795 -8120 19850 -8000
rect 19970 -8120 20015 -8000
rect 20135 -8120 20180 -8000
rect 20300 -8120 20345 -8000
rect 20465 -8120 20520 -8000
rect 20640 -8120 20685 -8000
rect 20805 -8120 20850 -8000
rect 20970 -8120 21015 -8000
rect 21135 -8120 21190 -8000
rect 21310 -8120 21355 -8000
rect 21475 -8120 21520 -8000
rect 21640 -8120 21685 -8000
rect 21805 -8120 21860 -8000
rect 21980 -8120 22025 -8000
rect 22145 -8120 22190 -8000
rect 22310 -8120 22355 -8000
rect 22475 -8120 22530 -8000
rect 22650 -8120 22695 -8000
rect 22815 -8120 22860 -8000
rect 22980 -8120 23025 -8000
rect 23145 -8120 23200 -8000
rect 23320 -8120 23365 -8000
rect 23485 -8120 23530 -8000
rect 23650 -8120 23695 -8000
rect 23815 -8120 23870 -8000
rect 23990 -8120 24000 -8000
rect 18500 -8165 24000 -8120
rect 18500 -8285 18510 -8165
rect 18630 -8285 18675 -8165
rect 18795 -8285 18840 -8165
rect 18960 -8285 19005 -8165
rect 19125 -8285 19180 -8165
rect 19300 -8285 19345 -8165
rect 19465 -8285 19510 -8165
rect 19630 -8285 19675 -8165
rect 19795 -8285 19850 -8165
rect 19970 -8285 20015 -8165
rect 20135 -8285 20180 -8165
rect 20300 -8285 20345 -8165
rect 20465 -8285 20520 -8165
rect 20640 -8285 20685 -8165
rect 20805 -8285 20850 -8165
rect 20970 -8285 21015 -8165
rect 21135 -8285 21190 -8165
rect 21310 -8285 21355 -8165
rect 21475 -8285 21520 -8165
rect 21640 -8285 21685 -8165
rect 21805 -8285 21860 -8165
rect 21980 -8285 22025 -8165
rect 22145 -8285 22190 -8165
rect 22310 -8285 22355 -8165
rect 22475 -8285 22530 -8165
rect 22650 -8285 22695 -8165
rect 22815 -8285 22860 -8165
rect 22980 -8285 23025 -8165
rect 23145 -8285 23200 -8165
rect 23320 -8285 23365 -8165
rect 23485 -8285 23530 -8165
rect 23650 -8285 23695 -8165
rect 23815 -8285 23870 -8165
rect 23990 -8285 24000 -8165
rect 18500 -8330 24000 -8285
rect 18500 -8450 18510 -8330
rect 18630 -8450 18675 -8330
rect 18795 -8450 18840 -8330
rect 18960 -8450 19005 -8330
rect 19125 -8450 19180 -8330
rect 19300 -8450 19345 -8330
rect 19465 -8450 19510 -8330
rect 19630 -8450 19675 -8330
rect 19795 -8450 19850 -8330
rect 19970 -8450 20015 -8330
rect 20135 -8450 20180 -8330
rect 20300 -8450 20345 -8330
rect 20465 -8450 20520 -8330
rect 20640 -8450 20685 -8330
rect 20805 -8450 20850 -8330
rect 20970 -8450 21015 -8330
rect 21135 -8450 21190 -8330
rect 21310 -8450 21355 -8330
rect 21475 -8450 21520 -8330
rect 21640 -8450 21685 -8330
rect 21805 -8450 21860 -8330
rect 21980 -8450 22025 -8330
rect 22145 -8450 22190 -8330
rect 22310 -8450 22355 -8330
rect 22475 -8450 22530 -8330
rect 22650 -8450 22695 -8330
rect 22815 -8450 22860 -8330
rect 22980 -8450 23025 -8330
rect 23145 -8450 23200 -8330
rect 23320 -8450 23365 -8330
rect 23485 -8450 23530 -8330
rect 23650 -8450 23695 -8330
rect 23815 -8450 23870 -8330
rect 23990 -8450 24000 -8330
rect 18500 -8505 24000 -8450
rect 18500 -8625 18510 -8505
rect 18630 -8625 18675 -8505
rect 18795 -8625 18840 -8505
rect 18960 -8625 19005 -8505
rect 19125 -8625 19180 -8505
rect 19300 -8625 19345 -8505
rect 19465 -8625 19510 -8505
rect 19630 -8625 19675 -8505
rect 19795 -8625 19850 -8505
rect 19970 -8625 20015 -8505
rect 20135 -8625 20180 -8505
rect 20300 -8625 20345 -8505
rect 20465 -8625 20520 -8505
rect 20640 -8625 20685 -8505
rect 20805 -8625 20850 -8505
rect 20970 -8625 21015 -8505
rect 21135 -8625 21190 -8505
rect 21310 -8625 21355 -8505
rect 21475 -8625 21520 -8505
rect 21640 -8625 21685 -8505
rect 21805 -8625 21860 -8505
rect 21980 -8625 22025 -8505
rect 22145 -8625 22190 -8505
rect 22310 -8625 22355 -8505
rect 22475 -8625 22530 -8505
rect 22650 -8625 22695 -8505
rect 22815 -8625 22860 -8505
rect 22980 -8625 23025 -8505
rect 23145 -8625 23200 -8505
rect 23320 -8625 23365 -8505
rect 23485 -8625 23530 -8505
rect 23650 -8625 23695 -8505
rect 23815 -8625 23870 -8505
rect 23990 -8625 24000 -8505
rect 18500 -8670 24000 -8625
rect 18500 -8790 18510 -8670
rect 18630 -8790 18675 -8670
rect 18795 -8790 18840 -8670
rect 18960 -8790 19005 -8670
rect 19125 -8790 19180 -8670
rect 19300 -8790 19345 -8670
rect 19465 -8790 19510 -8670
rect 19630 -8790 19675 -8670
rect 19795 -8790 19850 -8670
rect 19970 -8790 20015 -8670
rect 20135 -8790 20180 -8670
rect 20300 -8790 20345 -8670
rect 20465 -8790 20520 -8670
rect 20640 -8790 20685 -8670
rect 20805 -8790 20850 -8670
rect 20970 -8790 21015 -8670
rect 21135 -8790 21190 -8670
rect 21310 -8790 21355 -8670
rect 21475 -8790 21520 -8670
rect 21640 -8790 21685 -8670
rect 21805 -8790 21860 -8670
rect 21980 -8790 22025 -8670
rect 22145 -8790 22190 -8670
rect 22310 -8790 22355 -8670
rect 22475 -8790 22530 -8670
rect 22650 -8790 22695 -8670
rect 22815 -8790 22860 -8670
rect 22980 -8790 23025 -8670
rect 23145 -8790 23200 -8670
rect 23320 -8790 23365 -8670
rect 23485 -8790 23530 -8670
rect 23650 -8790 23695 -8670
rect 23815 -8790 23870 -8670
rect 23990 -8790 24000 -8670
rect 18500 -8835 24000 -8790
rect 18500 -8955 18510 -8835
rect 18630 -8955 18675 -8835
rect 18795 -8955 18840 -8835
rect 18960 -8955 19005 -8835
rect 19125 -8955 19180 -8835
rect 19300 -8955 19345 -8835
rect 19465 -8955 19510 -8835
rect 19630 -8955 19675 -8835
rect 19795 -8955 19850 -8835
rect 19970 -8955 20015 -8835
rect 20135 -8955 20180 -8835
rect 20300 -8955 20345 -8835
rect 20465 -8955 20520 -8835
rect 20640 -8955 20685 -8835
rect 20805 -8955 20850 -8835
rect 20970 -8955 21015 -8835
rect 21135 -8955 21190 -8835
rect 21310 -8955 21355 -8835
rect 21475 -8955 21520 -8835
rect 21640 -8955 21685 -8835
rect 21805 -8955 21860 -8835
rect 21980 -8955 22025 -8835
rect 22145 -8955 22190 -8835
rect 22310 -8955 22355 -8835
rect 22475 -8955 22530 -8835
rect 22650 -8955 22695 -8835
rect 22815 -8955 22860 -8835
rect 22980 -8955 23025 -8835
rect 23145 -8955 23200 -8835
rect 23320 -8955 23365 -8835
rect 23485 -8955 23530 -8835
rect 23650 -8955 23695 -8835
rect 23815 -8955 23870 -8835
rect 23990 -8955 24000 -8835
rect 18500 -9000 24000 -8955
rect 18500 -9120 18510 -9000
rect 18630 -9120 18675 -9000
rect 18795 -9120 18840 -9000
rect 18960 -9120 19005 -9000
rect 19125 -9120 19180 -9000
rect 19300 -9120 19345 -9000
rect 19465 -9120 19510 -9000
rect 19630 -9120 19675 -9000
rect 19795 -9120 19850 -9000
rect 19970 -9120 20015 -9000
rect 20135 -9120 20180 -9000
rect 20300 -9120 20345 -9000
rect 20465 -9120 20520 -9000
rect 20640 -9120 20685 -9000
rect 20805 -9120 20850 -9000
rect 20970 -9120 21015 -9000
rect 21135 -9120 21190 -9000
rect 21310 -9120 21355 -9000
rect 21475 -9120 21520 -9000
rect 21640 -9120 21685 -9000
rect 21805 -9120 21860 -9000
rect 21980 -9120 22025 -9000
rect 22145 -9120 22190 -9000
rect 22310 -9120 22355 -9000
rect 22475 -9120 22530 -9000
rect 22650 -9120 22695 -9000
rect 22815 -9120 22860 -9000
rect 22980 -9120 23025 -9000
rect 23145 -9120 23200 -9000
rect 23320 -9120 23365 -9000
rect 23485 -9120 23530 -9000
rect 23650 -9120 23695 -9000
rect 23815 -9120 23870 -9000
rect 23990 -9120 24000 -9000
rect 18500 -9175 24000 -9120
rect 18500 -9295 18510 -9175
rect 18630 -9295 18675 -9175
rect 18795 -9295 18840 -9175
rect 18960 -9295 19005 -9175
rect 19125 -9295 19180 -9175
rect 19300 -9295 19345 -9175
rect 19465 -9295 19510 -9175
rect 19630 -9295 19675 -9175
rect 19795 -9295 19850 -9175
rect 19970 -9295 20015 -9175
rect 20135 -9295 20180 -9175
rect 20300 -9295 20345 -9175
rect 20465 -9295 20520 -9175
rect 20640 -9295 20685 -9175
rect 20805 -9295 20850 -9175
rect 20970 -9295 21015 -9175
rect 21135 -9295 21190 -9175
rect 21310 -9295 21355 -9175
rect 21475 -9295 21520 -9175
rect 21640 -9295 21685 -9175
rect 21805 -9295 21860 -9175
rect 21980 -9295 22025 -9175
rect 22145 -9295 22190 -9175
rect 22310 -9295 22355 -9175
rect 22475 -9295 22530 -9175
rect 22650 -9295 22695 -9175
rect 22815 -9295 22860 -9175
rect 22980 -9295 23025 -9175
rect 23145 -9295 23200 -9175
rect 23320 -9295 23365 -9175
rect 23485 -9295 23530 -9175
rect 23650 -9295 23695 -9175
rect 23815 -9295 23870 -9175
rect 23990 -9295 24000 -9175
rect 18500 -9340 24000 -9295
rect 18500 -9460 18510 -9340
rect 18630 -9460 18675 -9340
rect 18795 -9460 18840 -9340
rect 18960 -9460 19005 -9340
rect 19125 -9460 19180 -9340
rect 19300 -9460 19345 -9340
rect 19465 -9460 19510 -9340
rect 19630 -9460 19675 -9340
rect 19795 -9460 19850 -9340
rect 19970 -9460 20015 -9340
rect 20135 -9460 20180 -9340
rect 20300 -9460 20345 -9340
rect 20465 -9460 20520 -9340
rect 20640 -9460 20685 -9340
rect 20805 -9460 20850 -9340
rect 20970 -9460 21015 -9340
rect 21135 -9460 21190 -9340
rect 21310 -9460 21355 -9340
rect 21475 -9460 21520 -9340
rect 21640 -9460 21685 -9340
rect 21805 -9460 21860 -9340
rect 21980 -9460 22025 -9340
rect 22145 -9460 22190 -9340
rect 22310 -9460 22355 -9340
rect 22475 -9460 22530 -9340
rect 22650 -9460 22695 -9340
rect 22815 -9460 22860 -9340
rect 22980 -9460 23025 -9340
rect 23145 -9460 23200 -9340
rect 23320 -9460 23365 -9340
rect 23485 -9460 23530 -9340
rect 23650 -9460 23695 -9340
rect 23815 -9460 23870 -9340
rect 23990 -9460 24000 -9340
rect 18500 -9505 24000 -9460
rect 18500 -9625 18510 -9505
rect 18630 -9625 18675 -9505
rect 18795 -9625 18840 -9505
rect 18960 -9625 19005 -9505
rect 19125 -9625 19180 -9505
rect 19300 -9625 19345 -9505
rect 19465 -9625 19510 -9505
rect 19630 -9625 19675 -9505
rect 19795 -9625 19850 -9505
rect 19970 -9625 20015 -9505
rect 20135 -9625 20180 -9505
rect 20300 -9625 20345 -9505
rect 20465 -9625 20520 -9505
rect 20640 -9625 20685 -9505
rect 20805 -9625 20850 -9505
rect 20970 -9625 21015 -9505
rect 21135 -9625 21190 -9505
rect 21310 -9625 21355 -9505
rect 21475 -9625 21520 -9505
rect 21640 -9625 21685 -9505
rect 21805 -9625 21860 -9505
rect 21980 -9625 22025 -9505
rect 22145 -9625 22190 -9505
rect 22310 -9625 22355 -9505
rect 22475 -9625 22530 -9505
rect 22650 -9625 22695 -9505
rect 22815 -9625 22860 -9505
rect 22980 -9625 23025 -9505
rect 23145 -9625 23200 -9505
rect 23320 -9625 23365 -9505
rect 23485 -9625 23530 -9505
rect 23650 -9625 23695 -9505
rect 23815 -9625 23870 -9505
rect 23990 -9625 24000 -9505
rect 18500 -9670 24000 -9625
rect 18500 -9790 18510 -9670
rect 18630 -9790 18675 -9670
rect 18795 -9790 18840 -9670
rect 18960 -9790 19005 -9670
rect 19125 -9790 19180 -9670
rect 19300 -9790 19345 -9670
rect 19465 -9790 19510 -9670
rect 19630 -9790 19675 -9670
rect 19795 -9790 19850 -9670
rect 19970 -9790 20015 -9670
rect 20135 -9790 20180 -9670
rect 20300 -9790 20345 -9670
rect 20465 -9790 20520 -9670
rect 20640 -9790 20685 -9670
rect 20805 -9790 20850 -9670
rect 20970 -9790 21015 -9670
rect 21135 -9790 21190 -9670
rect 21310 -9790 21355 -9670
rect 21475 -9790 21520 -9670
rect 21640 -9790 21685 -9670
rect 21805 -9790 21860 -9670
rect 21980 -9790 22025 -9670
rect 22145 -9790 22190 -9670
rect 22310 -9790 22355 -9670
rect 22475 -9790 22530 -9670
rect 22650 -9790 22695 -9670
rect 22815 -9790 22860 -9670
rect 22980 -9790 23025 -9670
rect 23145 -9790 23200 -9670
rect 23320 -9790 23365 -9670
rect 23485 -9790 23530 -9670
rect 23650 -9790 23695 -9670
rect 23815 -9790 23870 -9670
rect 23990 -9790 24000 -9670
rect 18500 -9800 24000 -9790
rect 24190 -4310 29690 -4300
rect 24190 -4430 24200 -4310
rect 24320 -4430 24365 -4310
rect 24485 -4430 24530 -4310
rect 24650 -4430 24695 -4310
rect 24815 -4430 24870 -4310
rect 24990 -4430 25035 -4310
rect 25155 -4430 25200 -4310
rect 25320 -4430 25365 -4310
rect 25485 -4430 25540 -4310
rect 25660 -4430 25705 -4310
rect 25825 -4430 25870 -4310
rect 25990 -4430 26035 -4310
rect 26155 -4430 26210 -4310
rect 26330 -4430 26375 -4310
rect 26495 -4430 26540 -4310
rect 26660 -4430 26705 -4310
rect 26825 -4430 26880 -4310
rect 27000 -4430 27045 -4310
rect 27165 -4430 27210 -4310
rect 27330 -4430 27375 -4310
rect 27495 -4430 27550 -4310
rect 27670 -4430 27715 -4310
rect 27835 -4430 27880 -4310
rect 28000 -4430 28045 -4310
rect 28165 -4430 28220 -4310
rect 28340 -4430 28385 -4310
rect 28505 -4430 28550 -4310
rect 28670 -4430 28715 -4310
rect 28835 -4430 28890 -4310
rect 29010 -4430 29055 -4310
rect 29175 -4430 29220 -4310
rect 29340 -4430 29385 -4310
rect 29505 -4430 29560 -4310
rect 29680 -4430 29690 -4310
rect 24190 -4485 29690 -4430
rect 24190 -4605 24200 -4485
rect 24320 -4605 24365 -4485
rect 24485 -4605 24530 -4485
rect 24650 -4605 24695 -4485
rect 24815 -4605 24870 -4485
rect 24990 -4605 25035 -4485
rect 25155 -4605 25200 -4485
rect 25320 -4605 25365 -4485
rect 25485 -4605 25540 -4485
rect 25660 -4605 25705 -4485
rect 25825 -4605 25870 -4485
rect 25990 -4605 26035 -4485
rect 26155 -4605 26210 -4485
rect 26330 -4605 26375 -4485
rect 26495 -4605 26540 -4485
rect 26660 -4605 26705 -4485
rect 26825 -4605 26880 -4485
rect 27000 -4605 27045 -4485
rect 27165 -4605 27210 -4485
rect 27330 -4605 27375 -4485
rect 27495 -4605 27550 -4485
rect 27670 -4605 27715 -4485
rect 27835 -4605 27880 -4485
rect 28000 -4605 28045 -4485
rect 28165 -4605 28220 -4485
rect 28340 -4605 28385 -4485
rect 28505 -4605 28550 -4485
rect 28670 -4605 28715 -4485
rect 28835 -4605 28890 -4485
rect 29010 -4605 29055 -4485
rect 29175 -4605 29220 -4485
rect 29340 -4605 29385 -4485
rect 29505 -4605 29560 -4485
rect 29680 -4605 29690 -4485
rect 24190 -4650 29690 -4605
rect 24190 -4770 24200 -4650
rect 24320 -4770 24365 -4650
rect 24485 -4770 24530 -4650
rect 24650 -4770 24695 -4650
rect 24815 -4770 24870 -4650
rect 24990 -4770 25035 -4650
rect 25155 -4770 25200 -4650
rect 25320 -4770 25365 -4650
rect 25485 -4770 25540 -4650
rect 25660 -4770 25705 -4650
rect 25825 -4770 25870 -4650
rect 25990 -4770 26035 -4650
rect 26155 -4770 26210 -4650
rect 26330 -4770 26375 -4650
rect 26495 -4770 26540 -4650
rect 26660 -4770 26705 -4650
rect 26825 -4770 26880 -4650
rect 27000 -4770 27045 -4650
rect 27165 -4770 27210 -4650
rect 27330 -4770 27375 -4650
rect 27495 -4770 27550 -4650
rect 27670 -4770 27715 -4650
rect 27835 -4770 27880 -4650
rect 28000 -4770 28045 -4650
rect 28165 -4770 28220 -4650
rect 28340 -4770 28385 -4650
rect 28505 -4770 28550 -4650
rect 28670 -4770 28715 -4650
rect 28835 -4770 28890 -4650
rect 29010 -4770 29055 -4650
rect 29175 -4770 29220 -4650
rect 29340 -4770 29385 -4650
rect 29505 -4770 29560 -4650
rect 29680 -4770 29690 -4650
rect 24190 -4815 29690 -4770
rect 24190 -4935 24200 -4815
rect 24320 -4935 24365 -4815
rect 24485 -4935 24530 -4815
rect 24650 -4935 24695 -4815
rect 24815 -4935 24870 -4815
rect 24990 -4935 25035 -4815
rect 25155 -4935 25200 -4815
rect 25320 -4935 25365 -4815
rect 25485 -4935 25540 -4815
rect 25660 -4935 25705 -4815
rect 25825 -4935 25870 -4815
rect 25990 -4935 26035 -4815
rect 26155 -4935 26210 -4815
rect 26330 -4935 26375 -4815
rect 26495 -4935 26540 -4815
rect 26660 -4935 26705 -4815
rect 26825 -4935 26880 -4815
rect 27000 -4935 27045 -4815
rect 27165 -4935 27210 -4815
rect 27330 -4935 27375 -4815
rect 27495 -4935 27550 -4815
rect 27670 -4935 27715 -4815
rect 27835 -4935 27880 -4815
rect 28000 -4935 28045 -4815
rect 28165 -4935 28220 -4815
rect 28340 -4935 28385 -4815
rect 28505 -4935 28550 -4815
rect 28670 -4935 28715 -4815
rect 28835 -4935 28890 -4815
rect 29010 -4935 29055 -4815
rect 29175 -4935 29220 -4815
rect 29340 -4935 29385 -4815
rect 29505 -4935 29560 -4815
rect 29680 -4935 29690 -4815
rect 24190 -4980 29690 -4935
rect 24190 -5100 24200 -4980
rect 24320 -5100 24365 -4980
rect 24485 -5100 24530 -4980
rect 24650 -5100 24695 -4980
rect 24815 -5100 24870 -4980
rect 24990 -5100 25035 -4980
rect 25155 -5100 25200 -4980
rect 25320 -5100 25365 -4980
rect 25485 -5100 25540 -4980
rect 25660 -5100 25705 -4980
rect 25825 -5100 25870 -4980
rect 25990 -5100 26035 -4980
rect 26155 -5100 26210 -4980
rect 26330 -5100 26375 -4980
rect 26495 -5100 26540 -4980
rect 26660 -5100 26705 -4980
rect 26825 -5100 26880 -4980
rect 27000 -5100 27045 -4980
rect 27165 -5100 27210 -4980
rect 27330 -5100 27375 -4980
rect 27495 -5100 27550 -4980
rect 27670 -5100 27715 -4980
rect 27835 -5100 27880 -4980
rect 28000 -5100 28045 -4980
rect 28165 -5100 28220 -4980
rect 28340 -5100 28385 -4980
rect 28505 -5100 28550 -4980
rect 28670 -5100 28715 -4980
rect 28835 -5100 28890 -4980
rect 29010 -5100 29055 -4980
rect 29175 -5100 29220 -4980
rect 29340 -5100 29385 -4980
rect 29505 -5100 29560 -4980
rect 29680 -5100 29690 -4980
rect 24190 -5155 29690 -5100
rect 24190 -5275 24200 -5155
rect 24320 -5275 24365 -5155
rect 24485 -5275 24530 -5155
rect 24650 -5275 24695 -5155
rect 24815 -5275 24870 -5155
rect 24990 -5275 25035 -5155
rect 25155 -5275 25200 -5155
rect 25320 -5275 25365 -5155
rect 25485 -5275 25540 -5155
rect 25660 -5275 25705 -5155
rect 25825 -5275 25870 -5155
rect 25990 -5275 26035 -5155
rect 26155 -5275 26210 -5155
rect 26330 -5275 26375 -5155
rect 26495 -5275 26540 -5155
rect 26660 -5275 26705 -5155
rect 26825 -5275 26880 -5155
rect 27000 -5275 27045 -5155
rect 27165 -5275 27210 -5155
rect 27330 -5275 27375 -5155
rect 27495 -5275 27550 -5155
rect 27670 -5275 27715 -5155
rect 27835 -5275 27880 -5155
rect 28000 -5275 28045 -5155
rect 28165 -5275 28220 -5155
rect 28340 -5275 28385 -5155
rect 28505 -5275 28550 -5155
rect 28670 -5275 28715 -5155
rect 28835 -5275 28890 -5155
rect 29010 -5275 29055 -5155
rect 29175 -5275 29220 -5155
rect 29340 -5275 29385 -5155
rect 29505 -5275 29560 -5155
rect 29680 -5275 29690 -5155
rect 24190 -5320 29690 -5275
rect 24190 -5440 24200 -5320
rect 24320 -5440 24365 -5320
rect 24485 -5440 24530 -5320
rect 24650 -5440 24695 -5320
rect 24815 -5440 24870 -5320
rect 24990 -5440 25035 -5320
rect 25155 -5440 25200 -5320
rect 25320 -5440 25365 -5320
rect 25485 -5440 25540 -5320
rect 25660 -5440 25705 -5320
rect 25825 -5440 25870 -5320
rect 25990 -5440 26035 -5320
rect 26155 -5440 26210 -5320
rect 26330 -5440 26375 -5320
rect 26495 -5440 26540 -5320
rect 26660 -5440 26705 -5320
rect 26825 -5440 26880 -5320
rect 27000 -5440 27045 -5320
rect 27165 -5440 27210 -5320
rect 27330 -5440 27375 -5320
rect 27495 -5440 27550 -5320
rect 27670 -5440 27715 -5320
rect 27835 -5440 27880 -5320
rect 28000 -5440 28045 -5320
rect 28165 -5440 28220 -5320
rect 28340 -5440 28385 -5320
rect 28505 -5440 28550 -5320
rect 28670 -5440 28715 -5320
rect 28835 -5440 28890 -5320
rect 29010 -5440 29055 -5320
rect 29175 -5440 29220 -5320
rect 29340 -5440 29385 -5320
rect 29505 -5440 29560 -5320
rect 29680 -5440 29690 -5320
rect 24190 -5485 29690 -5440
rect 24190 -5605 24200 -5485
rect 24320 -5605 24365 -5485
rect 24485 -5605 24530 -5485
rect 24650 -5605 24695 -5485
rect 24815 -5605 24870 -5485
rect 24990 -5605 25035 -5485
rect 25155 -5605 25200 -5485
rect 25320 -5605 25365 -5485
rect 25485 -5605 25540 -5485
rect 25660 -5605 25705 -5485
rect 25825 -5605 25870 -5485
rect 25990 -5605 26035 -5485
rect 26155 -5605 26210 -5485
rect 26330 -5605 26375 -5485
rect 26495 -5605 26540 -5485
rect 26660 -5605 26705 -5485
rect 26825 -5605 26880 -5485
rect 27000 -5605 27045 -5485
rect 27165 -5605 27210 -5485
rect 27330 -5605 27375 -5485
rect 27495 -5605 27550 -5485
rect 27670 -5605 27715 -5485
rect 27835 -5605 27880 -5485
rect 28000 -5605 28045 -5485
rect 28165 -5605 28220 -5485
rect 28340 -5605 28385 -5485
rect 28505 -5605 28550 -5485
rect 28670 -5605 28715 -5485
rect 28835 -5605 28890 -5485
rect 29010 -5605 29055 -5485
rect 29175 -5605 29220 -5485
rect 29340 -5605 29385 -5485
rect 29505 -5605 29560 -5485
rect 29680 -5605 29690 -5485
rect 24190 -5650 29690 -5605
rect 24190 -5770 24200 -5650
rect 24320 -5770 24365 -5650
rect 24485 -5770 24530 -5650
rect 24650 -5770 24695 -5650
rect 24815 -5770 24870 -5650
rect 24990 -5770 25035 -5650
rect 25155 -5770 25200 -5650
rect 25320 -5770 25365 -5650
rect 25485 -5770 25540 -5650
rect 25660 -5770 25705 -5650
rect 25825 -5770 25870 -5650
rect 25990 -5770 26035 -5650
rect 26155 -5770 26210 -5650
rect 26330 -5770 26375 -5650
rect 26495 -5770 26540 -5650
rect 26660 -5770 26705 -5650
rect 26825 -5770 26880 -5650
rect 27000 -5770 27045 -5650
rect 27165 -5770 27210 -5650
rect 27330 -5770 27375 -5650
rect 27495 -5770 27550 -5650
rect 27670 -5770 27715 -5650
rect 27835 -5770 27880 -5650
rect 28000 -5770 28045 -5650
rect 28165 -5770 28220 -5650
rect 28340 -5770 28385 -5650
rect 28505 -5770 28550 -5650
rect 28670 -5770 28715 -5650
rect 28835 -5770 28890 -5650
rect 29010 -5770 29055 -5650
rect 29175 -5770 29220 -5650
rect 29340 -5770 29385 -5650
rect 29505 -5770 29560 -5650
rect 29680 -5770 29690 -5650
rect 24190 -5825 29690 -5770
rect 24190 -5945 24200 -5825
rect 24320 -5945 24365 -5825
rect 24485 -5945 24530 -5825
rect 24650 -5945 24695 -5825
rect 24815 -5945 24870 -5825
rect 24990 -5945 25035 -5825
rect 25155 -5945 25200 -5825
rect 25320 -5945 25365 -5825
rect 25485 -5945 25540 -5825
rect 25660 -5945 25705 -5825
rect 25825 -5945 25870 -5825
rect 25990 -5945 26035 -5825
rect 26155 -5945 26210 -5825
rect 26330 -5945 26375 -5825
rect 26495 -5945 26540 -5825
rect 26660 -5945 26705 -5825
rect 26825 -5945 26880 -5825
rect 27000 -5945 27045 -5825
rect 27165 -5945 27210 -5825
rect 27330 -5945 27375 -5825
rect 27495 -5945 27550 -5825
rect 27670 -5945 27715 -5825
rect 27835 -5945 27880 -5825
rect 28000 -5945 28045 -5825
rect 28165 -5945 28220 -5825
rect 28340 -5945 28385 -5825
rect 28505 -5945 28550 -5825
rect 28670 -5945 28715 -5825
rect 28835 -5945 28890 -5825
rect 29010 -5945 29055 -5825
rect 29175 -5945 29220 -5825
rect 29340 -5945 29385 -5825
rect 29505 -5945 29560 -5825
rect 29680 -5945 29690 -5825
rect 24190 -5990 29690 -5945
rect 24190 -6110 24200 -5990
rect 24320 -6110 24365 -5990
rect 24485 -6110 24530 -5990
rect 24650 -6110 24695 -5990
rect 24815 -6110 24870 -5990
rect 24990 -6110 25035 -5990
rect 25155 -6110 25200 -5990
rect 25320 -6110 25365 -5990
rect 25485 -6110 25540 -5990
rect 25660 -6110 25705 -5990
rect 25825 -6110 25870 -5990
rect 25990 -6110 26035 -5990
rect 26155 -6110 26210 -5990
rect 26330 -6110 26375 -5990
rect 26495 -6110 26540 -5990
rect 26660 -6110 26705 -5990
rect 26825 -6110 26880 -5990
rect 27000 -6110 27045 -5990
rect 27165 -6110 27210 -5990
rect 27330 -6110 27375 -5990
rect 27495 -6110 27550 -5990
rect 27670 -6110 27715 -5990
rect 27835 -6110 27880 -5990
rect 28000 -6110 28045 -5990
rect 28165 -6110 28220 -5990
rect 28340 -6110 28385 -5990
rect 28505 -6110 28550 -5990
rect 28670 -6110 28715 -5990
rect 28835 -6110 28890 -5990
rect 29010 -6110 29055 -5990
rect 29175 -6110 29220 -5990
rect 29340 -6110 29385 -5990
rect 29505 -6110 29560 -5990
rect 29680 -6110 29690 -5990
rect 24190 -6155 29690 -6110
rect 24190 -6275 24200 -6155
rect 24320 -6275 24365 -6155
rect 24485 -6275 24530 -6155
rect 24650 -6275 24695 -6155
rect 24815 -6275 24870 -6155
rect 24990 -6275 25035 -6155
rect 25155 -6275 25200 -6155
rect 25320 -6275 25365 -6155
rect 25485 -6275 25540 -6155
rect 25660 -6275 25705 -6155
rect 25825 -6275 25870 -6155
rect 25990 -6275 26035 -6155
rect 26155 -6275 26210 -6155
rect 26330 -6275 26375 -6155
rect 26495 -6275 26540 -6155
rect 26660 -6275 26705 -6155
rect 26825 -6275 26880 -6155
rect 27000 -6275 27045 -6155
rect 27165 -6275 27210 -6155
rect 27330 -6275 27375 -6155
rect 27495 -6275 27550 -6155
rect 27670 -6275 27715 -6155
rect 27835 -6275 27880 -6155
rect 28000 -6275 28045 -6155
rect 28165 -6275 28220 -6155
rect 28340 -6275 28385 -6155
rect 28505 -6275 28550 -6155
rect 28670 -6275 28715 -6155
rect 28835 -6275 28890 -6155
rect 29010 -6275 29055 -6155
rect 29175 -6275 29220 -6155
rect 29340 -6275 29385 -6155
rect 29505 -6275 29560 -6155
rect 29680 -6275 29690 -6155
rect 24190 -6320 29690 -6275
rect 24190 -6440 24200 -6320
rect 24320 -6440 24365 -6320
rect 24485 -6440 24530 -6320
rect 24650 -6440 24695 -6320
rect 24815 -6440 24870 -6320
rect 24990 -6440 25035 -6320
rect 25155 -6440 25200 -6320
rect 25320 -6440 25365 -6320
rect 25485 -6440 25540 -6320
rect 25660 -6440 25705 -6320
rect 25825 -6440 25870 -6320
rect 25990 -6440 26035 -6320
rect 26155 -6440 26210 -6320
rect 26330 -6440 26375 -6320
rect 26495 -6440 26540 -6320
rect 26660 -6440 26705 -6320
rect 26825 -6440 26880 -6320
rect 27000 -6440 27045 -6320
rect 27165 -6440 27210 -6320
rect 27330 -6440 27375 -6320
rect 27495 -6440 27550 -6320
rect 27670 -6440 27715 -6320
rect 27835 -6440 27880 -6320
rect 28000 -6440 28045 -6320
rect 28165 -6440 28220 -6320
rect 28340 -6440 28385 -6320
rect 28505 -6440 28550 -6320
rect 28670 -6440 28715 -6320
rect 28835 -6440 28890 -6320
rect 29010 -6440 29055 -6320
rect 29175 -6440 29220 -6320
rect 29340 -6440 29385 -6320
rect 29505 -6440 29560 -6320
rect 29680 -6440 29690 -6320
rect 24190 -6495 29690 -6440
rect 24190 -6615 24200 -6495
rect 24320 -6615 24365 -6495
rect 24485 -6615 24530 -6495
rect 24650 -6615 24695 -6495
rect 24815 -6615 24870 -6495
rect 24990 -6615 25035 -6495
rect 25155 -6615 25200 -6495
rect 25320 -6615 25365 -6495
rect 25485 -6615 25540 -6495
rect 25660 -6615 25705 -6495
rect 25825 -6615 25870 -6495
rect 25990 -6615 26035 -6495
rect 26155 -6615 26210 -6495
rect 26330 -6615 26375 -6495
rect 26495 -6615 26540 -6495
rect 26660 -6615 26705 -6495
rect 26825 -6615 26880 -6495
rect 27000 -6615 27045 -6495
rect 27165 -6615 27210 -6495
rect 27330 -6615 27375 -6495
rect 27495 -6615 27550 -6495
rect 27670 -6615 27715 -6495
rect 27835 -6615 27880 -6495
rect 28000 -6615 28045 -6495
rect 28165 -6615 28220 -6495
rect 28340 -6615 28385 -6495
rect 28505 -6615 28550 -6495
rect 28670 -6615 28715 -6495
rect 28835 -6615 28890 -6495
rect 29010 -6615 29055 -6495
rect 29175 -6615 29220 -6495
rect 29340 -6615 29385 -6495
rect 29505 -6615 29560 -6495
rect 29680 -6615 29690 -6495
rect 24190 -6660 29690 -6615
rect 24190 -6780 24200 -6660
rect 24320 -6780 24365 -6660
rect 24485 -6780 24530 -6660
rect 24650 -6780 24695 -6660
rect 24815 -6780 24870 -6660
rect 24990 -6780 25035 -6660
rect 25155 -6780 25200 -6660
rect 25320 -6780 25365 -6660
rect 25485 -6780 25540 -6660
rect 25660 -6780 25705 -6660
rect 25825 -6780 25870 -6660
rect 25990 -6780 26035 -6660
rect 26155 -6780 26210 -6660
rect 26330 -6780 26375 -6660
rect 26495 -6780 26540 -6660
rect 26660 -6780 26705 -6660
rect 26825 -6780 26880 -6660
rect 27000 -6780 27045 -6660
rect 27165 -6780 27210 -6660
rect 27330 -6780 27375 -6660
rect 27495 -6780 27550 -6660
rect 27670 -6780 27715 -6660
rect 27835 -6780 27880 -6660
rect 28000 -6780 28045 -6660
rect 28165 -6780 28220 -6660
rect 28340 -6780 28385 -6660
rect 28505 -6780 28550 -6660
rect 28670 -6780 28715 -6660
rect 28835 -6780 28890 -6660
rect 29010 -6780 29055 -6660
rect 29175 -6780 29220 -6660
rect 29340 -6780 29385 -6660
rect 29505 -6780 29560 -6660
rect 29680 -6780 29690 -6660
rect 24190 -6825 29690 -6780
rect 24190 -6945 24200 -6825
rect 24320 -6945 24365 -6825
rect 24485 -6945 24530 -6825
rect 24650 -6945 24695 -6825
rect 24815 -6945 24870 -6825
rect 24990 -6945 25035 -6825
rect 25155 -6945 25200 -6825
rect 25320 -6945 25365 -6825
rect 25485 -6945 25540 -6825
rect 25660 -6945 25705 -6825
rect 25825 -6945 25870 -6825
rect 25990 -6945 26035 -6825
rect 26155 -6945 26210 -6825
rect 26330 -6945 26375 -6825
rect 26495 -6945 26540 -6825
rect 26660 -6945 26705 -6825
rect 26825 -6945 26880 -6825
rect 27000 -6945 27045 -6825
rect 27165 -6945 27210 -6825
rect 27330 -6945 27375 -6825
rect 27495 -6945 27550 -6825
rect 27670 -6945 27715 -6825
rect 27835 -6945 27880 -6825
rect 28000 -6945 28045 -6825
rect 28165 -6945 28220 -6825
rect 28340 -6945 28385 -6825
rect 28505 -6945 28550 -6825
rect 28670 -6945 28715 -6825
rect 28835 -6945 28890 -6825
rect 29010 -6945 29055 -6825
rect 29175 -6945 29220 -6825
rect 29340 -6945 29385 -6825
rect 29505 -6945 29560 -6825
rect 29680 -6945 29690 -6825
rect 24190 -6990 29690 -6945
rect 24190 -7110 24200 -6990
rect 24320 -7110 24365 -6990
rect 24485 -7110 24530 -6990
rect 24650 -7110 24695 -6990
rect 24815 -7110 24870 -6990
rect 24990 -7110 25035 -6990
rect 25155 -7110 25200 -6990
rect 25320 -7110 25365 -6990
rect 25485 -7110 25540 -6990
rect 25660 -7110 25705 -6990
rect 25825 -7110 25870 -6990
rect 25990 -7110 26035 -6990
rect 26155 -7110 26210 -6990
rect 26330 -7110 26375 -6990
rect 26495 -7110 26540 -6990
rect 26660 -7110 26705 -6990
rect 26825 -7110 26880 -6990
rect 27000 -7110 27045 -6990
rect 27165 -7110 27210 -6990
rect 27330 -7110 27375 -6990
rect 27495 -7110 27550 -6990
rect 27670 -7110 27715 -6990
rect 27835 -7110 27880 -6990
rect 28000 -7110 28045 -6990
rect 28165 -7110 28220 -6990
rect 28340 -7110 28385 -6990
rect 28505 -7110 28550 -6990
rect 28670 -7110 28715 -6990
rect 28835 -7110 28890 -6990
rect 29010 -7110 29055 -6990
rect 29175 -7110 29220 -6990
rect 29340 -7110 29385 -6990
rect 29505 -7110 29560 -6990
rect 29680 -7110 29690 -6990
rect 24190 -7165 29690 -7110
rect 24190 -7285 24200 -7165
rect 24320 -7285 24365 -7165
rect 24485 -7285 24530 -7165
rect 24650 -7285 24695 -7165
rect 24815 -7285 24870 -7165
rect 24990 -7285 25035 -7165
rect 25155 -7285 25200 -7165
rect 25320 -7285 25365 -7165
rect 25485 -7285 25540 -7165
rect 25660 -7285 25705 -7165
rect 25825 -7285 25870 -7165
rect 25990 -7285 26035 -7165
rect 26155 -7285 26210 -7165
rect 26330 -7285 26375 -7165
rect 26495 -7285 26540 -7165
rect 26660 -7285 26705 -7165
rect 26825 -7285 26880 -7165
rect 27000 -7285 27045 -7165
rect 27165 -7285 27210 -7165
rect 27330 -7285 27375 -7165
rect 27495 -7285 27550 -7165
rect 27670 -7285 27715 -7165
rect 27835 -7285 27880 -7165
rect 28000 -7285 28045 -7165
rect 28165 -7285 28220 -7165
rect 28340 -7285 28385 -7165
rect 28505 -7285 28550 -7165
rect 28670 -7285 28715 -7165
rect 28835 -7285 28890 -7165
rect 29010 -7285 29055 -7165
rect 29175 -7285 29220 -7165
rect 29340 -7285 29385 -7165
rect 29505 -7285 29560 -7165
rect 29680 -7285 29690 -7165
rect 24190 -7330 29690 -7285
rect 24190 -7450 24200 -7330
rect 24320 -7450 24365 -7330
rect 24485 -7450 24530 -7330
rect 24650 -7450 24695 -7330
rect 24815 -7450 24870 -7330
rect 24990 -7450 25035 -7330
rect 25155 -7450 25200 -7330
rect 25320 -7450 25365 -7330
rect 25485 -7450 25540 -7330
rect 25660 -7450 25705 -7330
rect 25825 -7450 25870 -7330
rect 25990 -7450 26035 -7330
rect 26155 -7450 26210 -7330
rect 26330 -7450 26375 -7330
rect 26495 -7450 26540 -7330
rect 26660 -7450 26705 -7330
rect 26825 -7450 26880 -7330
rect 27000 -7450 27045 -7330
rect 27165 -7450 27210 -7330
rect 27330 -7450 27375 -7330
rect 27495 -7450 27550 -7330
rect 27670 -7450 27715 -7330
rect 27835 -7450 27880 -7330
rect 28000 -7450 28045 -7330
rect 28165 -7450 28220 -7330
rect 28340 -7450 28385 -7330
rect 28505 -7450 28550 -7330
rect 28670 -7450 28715 -7330
rect 28835 -7450 28890 -7330
rect 29010 -7450 29055 -7330
rect 29175 -7450 29220 -7330
rect 29340 -7450 29385 -7330
rect 29505 -7450 29560 -7330
rect 29680 -7450 29690 -7330
rect 24190 -7495 29690 -7450
rect 24190 -7615 24200 -7495
rect 24320 -7615 24365 -7495
rect 24485 -7615 24530 -7495
rect 24650 -7615 24695 -7495
rect 24815 -7615 24870 -7495
rect 24990 -7615 25035 -7495
rect 25155 -7615 25200 -7495
rect 25320 -7615 25365 -7495
rect 25485 -7615 25540 -7495
rect 25660 -7615 25705 -7495
rect 25825 -7615 25870 -7495
rect 25990 -7615 26035 -7495
rect 26155 -7615 26210 -7495
rect 26330 -7615 26375 -7495
rect 26495 -7615 26540 -7495
rect 26660 -7615 26705 -7495
rect 26825 -7615 26880 -7495
rect 27000 -7615 27045 -7495
rect 27165 -7615 27210 -7495
rect 27330 -7615 27375 -7495
rect 27495 -7615 27550 -7495
rect 27670 -7615 27715 -7495
rect 27835 -7615 27880 -7495
rect 28000 -7615 28045 -7495
rect 28165 -7615 28220 -7495
rect 28340 -7615 28385 -7495
rect 28505 -7615 28550 -7495
rect 28670 -7615 28715 -7495
rect 28835 -7615 28890 -7495
rect 29010 -7615 29055 -7495
rect 29175 -7615 29220 -7495
rect 29340 -7615 29385 -7495
rect 29505 -7615 29560 -7495
rect 29680 -7615 29690 -7495
rect 24190 -7660 29690 -7615
rect 24190 -7780 24200 -7660
rect 24320 -7780 24365 -7660
rect 24485 -7780 24530 -7660
rect 24650 -7780 24695 -7660
rect 24815 -7780 24870 -7660
rect 24990 -7780 25035 -7660
rect 25155 -7780 25200 -7660
rect 25320 -7780 25365 -7660
rect 25485 -7780 25540 -7660
rect 25660 -7780 25705 -7660
rect 25825 -7780 25870 -7660
rect 25990 -7780 26035 -7660
rect 26155 -7780 26210 -7660
rect 26330 -7780 26375 -7660
rect 26495 -7780 26540 -7660
rect 26660 -7780 26705 -7660
rect 26825 -7780 26880 -7660
rect 27000 -7780 27045 -7660
rect 27165 -7780 27210 -7660
rect 27330 -7780 27375 -7660
rect 27495 -7780 27550 -7660
rect 27670 -7780 27715 -7660
rect 27835 -7780 27880 -7660
rect 28000 -7780 28045 -7660
rect 28165 -7780 28220 -7660
rect 28340 -7780 28385 -7660
rect 28505 -7780 28550 -7660
rect 28670 -7780 28715 -7660
rect 28835 -7780 28890 -7660
rect 29010 -7780 29055 -7660
rect 29175 -7780 29220 -7660
rect 29340 -7780 29385 -7660
rect 29505 -7780 29560 -7660
rect 29680 -7780 29690 -7660
rect 24190 -7835 29690 -7780
rect 24190 -7955 24200 -7835
rect 24320 -7955 24365 -7835
rect 24485 -7955 24530 -7835
rect 24650 -7955 24695 -7835
rect 24815 -7955 24870 -7835
rect 24990 -7955 25035 -7835
rect 25155 -7955 25200 -7835
rect 25320 -7955 25365 -7835
rect 25485 -7955 25540 -7835
rect 25660 -7955 25705 -7835
rect 25825 -7955 25870 -7835
rect 25990 -7955 26035 -7835
rect 26155 -7955 26210 -7835
rect 26330 -7955 26375 -7835
rect 26495 -7955 26540 -7835
rect 26660 -7955 26705 -7835
rect 26825 -7955 26880 -7835
rect 27000 -7955 27045 -7835
rect 27165 -7955 27210 -7835
rect 27330 -7955 27375 -7835
rect 27495 -7955 27550 -7835
rect 27670 -7955 27715 -7835
rect 27835 -7955 27880 -7835
rect 28000 -7955 28045 -7835
rect 28165 -7955 28220 -7835
rect 28340 -7955 28385 -7835
rect 28505 -7955 28550 -7835
rect 28670 -7955 28715 -7835
rect 28835 -7955 28890 -7835
rect 29010 -7955 29055 -7835
rect 29175 -7955 29220 -7835
rect 29340 -7955 29385 -7835
rect 29505 -7955 29560 -7835
rect 29680 -7955 29690 -7835
rect 24190 -8000 29690 -7955
rect 24190 -8120 24200 -8000
rect 24320 -8120 24365 -8000
rect 24485 -8120 24530 -8000
rect 24650 -8120 24695 -8000
rect 24815 -8120 24870 -8000
rect 24990 -8120 25035 -8000
rect 25155 -8120 25200 -8000
rect 25320 -8120 25365 -8000
rect 25485 -8120 25540 -8000
rect 25660 -8120 25705 -8000
rect 25825 -8120 25870 -8000
rect 25990 -8120 26035 -8000
rect 26155 -8120 26210 -8000
rect 26330 -8120 26375 -8000
rect 26495 -8120 26540 -8000
rect 26660 -8120 26705 -8000
rect 26825 -8120 26880 -8000
rect 27000 -8120 27045 -8000
rect 27165 -8120 27210 -8000
rect 27330 -8120 27375 -8000
rect 27495 -8120 27550 -8000
rect 27670 -8120 27715 -8000
rect 27835 -8120 27880 -8000
rect 28000 -8120 28045 -8000
rect 28165 -8120 28220 -8000
rect 28340 -8120 28385 -8000
rect 28505 -8120 28550 -8000
rect 28670 -8120 28715 -8000
rect 28835 -8120 28890 -8000
rect 29010 -8120 29055 -8000
rect 29175 -8120 29220 -8000
rect 29340 -8120 29385 -8000
rect 29505 -8120 29560 -8000
rect 29680 -8120 29690 -8000
rect 24190 -8165 29690 -8120
rect 24190 -8285 24200 -8165
rect 24320 -8285 24365 -8165
rect 24485 -8285 24530 -8165
rect 24650 -8285 24695 -8165
rect 24815 -8285 24870 -8165
rect 24990 -8285 25035 -8165
rect 25155 -8285 25200 -8165
rect 25320 -8285 25365 -8165
rect 25485 -8285 25540 -8165
rect 25660 -8285 25705 -8165
rect 25825 -8285 25870 -8165
rect 25990 -8285 26035 -8165
rect 26155 -8285 26210 -8165
rect 26330 -8285 26375 -8165
rect 26495 -8285 26540 -8165
rect 26660 -8285 26705 -8165
rect 26825 -8285 26880 -8165
rect 27000 -8285 27045 -8165
rect 27165 -8285 27210 -8165
rect 27330 -8285 27375 -8165
rect 27495 -8285 27550 -8165
rect 27670 -8285 27715 -8165
rect 27835 -8285 27880 -8165
rect 28000 -8285 28045 -8165
rect 28165 -8285 28220 -8165
rect 28340 -8285 28385 -8165
rect 28505 -8285 28550 -8165
rect 28670 -8285 28715 -8165
rect 28835 -8285 28890 -8165
rect 29010 -8285 29055 -8165
rect 29175 -8285 29220 -8165
rect 29340 -8285 29385 -8165
rect 29505 -8285 29560 -8165
rect 29680 -8285 29690 -8165
rect 24190 -8330 29690 -8285
rect 24190 -8450 24200 -8330
rect 24320 -8450 24365 -8330
rect 24485 -8450 24530 -8330
rect 24650 -8450 24695 -8330
rect 24815 -8450 24870 -8330
rect 24990 -8450 25035 -8330
rect 25155 -8450 25200 -8330
rect 25320 -8450 25365 -8330
rect 25485 -8450 25540 -8330
rect 25660 -8450 25705 -8330
rect 25825 -8450 25870 -8330
rect 25990 -8450 26035 -8330
rect 26155 -8450 26210 -8330
rect 26330 -8450 26375 -8330
rect 26495 -8450 26540 -8330
rect 26660 -8450 26705 -8330
rect 26825 -8450 26880 -8330
rect 27000 -8450 27045 -8330
rect 27165 -8450 27210 -8330
rect 27330 -8450 27375 -8330
rect 27495 -8450 27550 -8330
rect 27670 -8450 27715 -8330
rect 27835 -8450 27880 -8330
rect 28000 -8450 28045 -8330
rect 28165 -8450 28220 -8330
rect 28340 -8450 28385 -8330
rect 28505 -8450 28550 -8330
rect 28670 -8450 28715 -8330
rect 28835 -8450 28890 -8330
rect 29010 -8450 29055 -8330
rect 29175 -8450 29220 -8330
rect 29340 -8450 29385 -8330
rect 29505 -8450 29560 -8330
rect 29680 -8450 29690 -8330
rect 24190 -8505 29690 -8450
rect 24190 -8625 24200 -8505
rect 24320 -8625 24365 -8505
rect 24485 -8625 24530 -8505
rect 24650 -8625 24695 -8505
rect 24815 -8625 24870 -8505
rect 24990 -8625 25035 -8505
rect 25155 -8625 25200 -8505
rect 25320 -8625 25365 -8505
rect 25485 -8625 25540 -8505
rect 25660 -8625 25705 -8505
rect 25825 -8625 25870 -8505
rect 25990 -8625 26035 -8505
rect 26155 -8625 26210 -8505
rect 26330 -8625 26375 -8505
rect 26495 -8625 26540 -8505
rect 26660 -8625 26705 -8505
rect 26825 -8625 26880 -8505
rect 27000 -8625 27045 -8505
rect 27165 -8625 27210 -8505
rect 27330 -8625 27375 -8505
rect 27495 -8625 27550 -8505
rect 27670 -8625 27715 -8505
rect 27835 -8625 27880 -8505
rect 28000 -8625 28045 -8505
rect 28165 -8625 28220 -8505
rect 28340 -8625 28385 -8505
rect 28505 -8625 28550 -8505
rect 28670 -8625 28715 -8505
rect 28835 -8625 28890 -8505
rect 29010 -8625 29055 -8505
rect 29175 -8625 29220 -8505
rect 29340 -8625 29385 -8505
rect 29505 -8625 29560 -8505
rect 29680 -8625 29690 -8505
rect 24190 -8670 29690 -8625
rect 24190 -8790 24200 -8670
rect 24320 -8790 24365 -8670
rect 24485 -8790 24530 -8670
rect 24650 -8790 24695 -8670
rect 24815 -8790 24870 -8670
rect 24990 -8790 25035 -8670
rect 25155 -8790 25200 -8670
rect 25320 -8790 25365 -8670
rect 25485 -8790 25540 -8670
rect 25660 -8790 25705 -8670
rect 25825 -8790 25870 -8670
rect 25990 -8790 26035 -8670
rect 26155 -8790 26210 -8670
rect 26330 -8790 26375 -8670
rect 26495 -8790 26540 -8670
rect 26660 -8790 26705 -8670
rect 26825 -8790 26880 -8670
rect 27000 -8790 27045 -8670
rect 27165 -8790 27210 -8670
rect 27330 -8790 27375 -8670
rect 27495 -8790 27550 -8670
rect 27670 -8790 27715 -8670
rect 27835 -8790 27880 -8670
rect 28000 -8790 28045 -8670
rect 28165 -8790 28220 -8670
rect 28340 -8790 28385 -8670
rect 28505 -8790 28550 -8670
rect 28670 -8790 28715 -8670
rect 28835 -8790 28890 -8670
rect 29010 -8790 29055 -8670
rect 29175 -8790 29220 -8670
rect 29340 -8790 29385 -8670
rect 29505 -8790 29560 -8670
rect 29680 -8790 29690 -8670
rect 24190 -8835 29690 -8790
rect 24190 -8955 24200 -8835
rect 24320 -8955 24365 -8835
rect 24485 -8955 24530 -8835
rect 24650 -8955 24695 -8835
rect 24815 -8955 24870 -8835
rect 24990 -8955 25035 -8835
rect 25155 -8955 25200 -8835
rect 25320 -8955 25365 -8835
rect 25485 -8955 25540 -8835
rect 25660 -8955 25705 -8835
rect 25825 -8955 25870 -8835
rect 25990 -8955 26035 -8835
rect 26155 -8955 26210 -8835
rect 26330 -8955 26375 -8835
rect 26495 -8955 26540 -8835
rect 26660 -8955 26705 -8835
rect 26825 -8955 26880 -8835
rect 27000 -8955 27045 -8835
rect 27165 -8955 27210 -8835
rect 27330 -8955 27375 -8835
rect 27495 -8955 27550 -8835
rect 27670 -8955 27715 -8835
rect 27835 -8955 27880 -8835
rect 28000 -8955 28045 -8835
rect 28165 -8955 28220 -8835
rect 28340 -8955 28385 -8835
rect 28505 -8955 28550 -8835
rect 28670 -8955 28715 -8835
rect 28835 -8955 28890 -8835
rect 29010 -8955 29055 -8835
rect 29175 -8955 29220 -8835
rect 29340 -8955 29385 -8835
rect 29505 -8955 29560 -8835
rect 29680 -8955 29690 -8835
rect 24190 -9000 29690 -8955
rect 24190 -9120 24200 -9000
rect 24320 -9120 24365 -9000
rect 24485 -9120 24530 -9000
rect 24650 -9120 24695 -9000
rect 24815 -9120 24870 -9000
rect 24990 -9120 25035 -9000
rect 25155 -9120 25200 -9000
rect 25320 -9120 25365 -9000
rect 25485 -9120 25540 -9000
rect 25660 -9120 25705 -9000
rect 25825 -9120 25870 -9000
rect 25990 -9120 26035 -9000
rect 26155 -9120 26210 -9000
rect 26330 -9120 26375 -9000
rect 26495 -9120 26540 -9000
rect 26660 -9120 26705 -9000
rect 26825 -9120 26880 -9000
rect 27000 -9120 27045 -9000
rect 27165 -9120 27210 -9000
rect 27330 -9120 27375 -9000
rect 27495 -9120 27550 -9000
rect 27670 -9120 27715 -9000
rect 27835 -9120 27880 -9000
rect 28000 -9120 28045 -9000
rect 28165 -9120 28220 -9000
rect 28340 -9120 28385 -9000
rect 28505 -9120 28550 -9000
rect 28670 -9120 28715 -9000
rect 28835 -9120 28890 -9000
rect 29010 -9120 29055 -9000
rect 29175 -9120 29220 -9000
rect 29340 -9120 29385 -9000
rect 29505 -9120 29560 -9000
rect 29680 -9120 29690 -9000
rect 24190 -9175 29690 -9120
rect 24190 -9295 24200 -9175
rect 24320 -9295 24365 -9175
rect 24485 -9295 24530 -9175
rect 24650 -9295 24695 -9175
rect 24815 -9295 24870 -9175
rect 24990 -9295 25035 -9175
rect 25155 -9295 25200 -9175
rect 25320 -9295 25365 -9175
rect 25485 -9295 25540 -9175
rect 25660 -9295 25705 -9175
rect 25825 -9295 25870 -9175
rect 25990 -9295 26035 -9175
rect 26155 -9295 26210 -9175
rect 26330 -9295 26375 -9175
rect 26495 -9295 26540 -9175
rect 26660 -9295 26705 -9175
rect 26825 -9295 26880 -9175
rect 27000 -9295 27045 -9175
rect 27165 -9295 27210 -9175
rect 27330 -9295 27375 -9175
rect 27495 -9295 27550 -9175
rect 27670 -9295 27715 -9175
rect 27835 -9295 27880 -9175
rect 28000 -9295 28045 -9175
rect 28165 -9295 28220 -9175
rect 28340 -9295 28385 -9175
rect 28505 -9295 28550 -9175
rect 28670 -9295 28715 -9175
rect 28835 -9295 28890 -9175
rect 29010 -9295 29055 -9175
rect 29175 -9295 29220 -9175
rect 29340 -9295 29385 -9175
rect 29505 -9295 29560 -9175
rect 29680 -9295 29690 -9175
rect 24190 -9340 29690 -9295
rect 24190 -9460 24200 -9340
rect 24320 -9460 24365 -9340
rect 24485 -9460 24530 -9340
rect 24650 -9460 24695 -9340
rect 24815 -9460 24870 -9340
rect 24990 -9460 25035 -9340
rect 25155 -9460 25200 -9340
rect 25320 -9460 25365 -9340
rect 25485 -9460 25540 -9340
rect 25660 -9460 25705 -9340
rect 25825 -9460 25870 -9340
rect 25990 -9460 26035 -9340
rect 26155 -9460 26210 -9340
rect 26330 -9460 26375 -9340
rect 26495 -9460 26540 -9340
rect 26660 -9460 26705 -9340
rect 26825 -9460 26880 -9340
rect 27000 -9460 27045 -9340
rect 27165 -9460 27210 -9340
rect 27330 -9460 27375 -9340
rect 27495 -9460 27550 -9340
rect 27670 -9460 27715 -9340
rect 27835 -9460 27880 -9340
rect 28000 -9460 28045 -9340
rect 28165 -9460 28220 -9340
rect 28340 -9460 28385 -9340
rect 28505 -9460 28550 -9340
rect 28670 -9460 28715 -9340
rect 28835 -9460 28890 -9340
rect 29010 -9460 29055 -9340
rect 29175 -9460 29220 -9340
rect 29340 -9460 29385 -9340
rect 29505 -9460 29560 -9340
rect 29680 -9460 29690 -9340
rect 24190 -9505 29690 -9460
rect 24190 -9625 24200 -9505
rect 24320 -9625 24365 -9505
rect 24485 -9625 24530 -9505
rect 24650 -9625 24695 -9505
rect 24815 -9625 24870 -9505
rect 24990 -9625 25035 -9505
rect 25155 -9625 25200 -9505
rect 25320 -9625 25365 -9505
rect 25485 -9625 25540 -9505
rect 25660 -9625 25705 -9505
rect 25825 -9625 25870 -9505
rect 25990 -9625 26035 -9505
rect 26155 -9625 26210 -9505
rect 26330 -9625 26375 -9505
rect 26495 -9625 26540 -9505
rect 26660 -9625 26705 -9505
rect 26825 -9625 26880 -9505
rect 27000 -9625 27045 -9505
rect 27165 -9625 27210 -9505
rect 27330 -9625 27375 -9505
rect 27495 -9625 27550 -9505
rect 27670 -9625 27715 -9505
rect 27835 -9625 27880 -9505
rect 28000 -9625 28045 -9505
rect 28165 -9625 28220 -9505
rect 28340 -9625 28385 -9505
rect 28505 -9625 28550 -9505
rect 28670 -9625 28715 -9505
rect 28835 -9625 28890 -9505
rect 29010 -9625 29055 -9505
rect 29175 -9625 29220 -9505
rect 29340 -9625 29385 -9505
rect 29505 -9625 29560 -9505
rect 29680 -9625 29690 -9505
rect 24190 -9670 29690 -9625
rect 24190 -9790 24200 -9670
rect 24320 -9790 24365 -9670
rect 24485 -9790 24530 -9670
rect 24650 -9790 24695 -9670
rect 24815 -9790 24870 -9670
rect 24990 -9790 25035 -9670
rect 25155 -9790 25200 -9670
rect 25320 -9790 25365 -9670
rect 25485 -9790 25540 -9670
rect 25660 -9790 25705 -9670
rect 25825 -9790 25870 -9670
rect 25990 -9790 26035 -9670
rect 26155 -9790 26210 -9670
rect 26330 -9790 26375 -9670
rect 26495 -9790 26540 -9670
rect 26660 -9790 26705 -9670
rect 26825 -9790 26880 -9670
rect 27000 -9790 27045 -9670
rect 27165 -9790 27210 -9670
rect 27330 -9790 27375 -9670
rect 27495 -9790 27550 -9670
rect 27670 -9790 27715 -9670
rect 27835 -9790 27880 -9670
rect 28000 -9790 28045 -9670
rect 28165 -9790 28220 -9670
rect 28340 -9790 28385 -9670
rect 28505 -9790 28550 -9670
rect 28670 -9790 28715 -9670
rect 28835 -9790 28890 -9670
rect 29010 -9790 29055 -9670
rect 29175 -9790 29220 -9670
rect 29340 -9790 29385 -9670
rect 29505 -9790 29560 -9670
rect 29680 -9790 29690 -9670
rect 24190 -9800 29690 -9790
rect 7120 -10090 12620 -10080
rect 7120 -10210 7130 -10090
rect 7250 -10210 7305 -10090
rect 7425 -10210 7470 -10090
rect 7590 -10210 7635 -10090
rect 7755 -10210 7800 -10090
rect 7920 -10210 7975 -10090
rect 8095 -10210 8140 -10090
rect 8260 -10210 8305 -10090
rect 8425 -10210 8470 -10090
rect 8590 -10210 8645 -10090
rect 8765 -10210 8810 -10090
rect 8930 -10210 8975 -10090
rect 9095 -10210 9140 -10090
rect 9260 -10210 9315 -10090
rect 9435 -10210 9480 -10090
rect 9600 -10210 9645 -10090
rect 9765 -10210 9810 -10090
rect 9930 -10210 9985 -10090
rect 10105 -10210 10150 -10090
rect 10270 -10210 10315 -10090
rect 10435 -10210 10480 -10090
rect 10600 -10210 10655 -10090
rect 10775 -10210 10820 -10090
rect 10940 -10210 10985 -10090
rect 11105 -10210 11150 -10090
rect 11270 -10210 11325 -10090
rect 11445 -10210 11490 -10090
rect 11610 -10210 11655 -10090
rect 11775 -10210 11820 -10090
rect 11940 -10210 11995 -10090
rect 12115 -10210 12160 -10090
rect 12280 -10210 12325 -10090
rect 12445 -10210 12490 -10090
rect 12610 -10210 12620 -10090
rect 7120 -10255 12620 -10210
rect 7120 -10375 7130 -10255
rect 7250 -10375 7305 -10255
rect 7425 -10375 7470 -10255
rect 7590 -10375 7635 -10255
rect 7755 -10375 7800 -10255
rect 7920 -10375 7975 -10255
rect 8095 -10375 8140 -10255
rect 8260 -10375 8305 -10255
rect 8425 -10375 8470 -10255
rect 8590 -10375 8645 -10255
rect 8765 -10375 8810 -10255
rect 8930 -10375 8975 -10255
rect 9095 -10375 9140 -10255
rect 9260 -10375 9315 -10255
rect 9435 -10375 9480 -10255
rect 9600 -10375 9645 -10255
rect 9765 -10375 9810 -10255
rect 9930 -10375 9985 -10255
rect 10105 -10375 10150 -10255
rect 10270 -10375 10315 -10255
rect 10435 -10375 10480 -10255
rect 10600 -10375 10655 -10255
rect 10775 -10375 10820 -10255
rect 10940 -10375 10985 -10255
rect 11105 -10375 11150 -10255
rect 11270 -10375 11325 -10255
rect 11445 -10375 11490 -10255
rect 11610 -10375 11655 -10255
rect 11775 -10375 11820 -10255
rect 11940 -10375 11995 -10255
rect 12115 -10375 12160 -10255
rect 12280 -10375 12325 -10255
rect 12445 -10375 12490 -10255
rect 12610 -10375 12620 -10255
rect 7120 -10420 12620 -10375
rect 7120 -10540 7130 -10420
rect 7250 -10540 7305 -10420
rect 7425 -10540 7470 -10420
rect 7590 -10540 7635 -10420
rect 7755 -10540 7800 -10420
rect 7920 -10540 7975 -10420
rect 8095 -10540 8140 -10420
rect 8260 -10540 8305 -10420
rect 8425 -10540 8470 -10420
rect 8590 -10540 8645 -10420
rect 8765 -10540 8810 -10420
rect 8930 -10540 8975 -10420
rect 9095 -10540 9140 -10420
rect 9260 -10540 9315 -10420
rect 9435 -10540 9480 -10420
rect 9600 -10540 9645 -10420
rect 9765 -10540 9810 -10420
rect 9930 -10540 9985 -10420
rect 10105 -10540 10150 -10420
rect 10270 -10540 10315 -10420
rect 10435 -10540 10480 -10420
rect 10600 -10540 10655 -10420
rect 10775 -10540 10820 -10420
rect 10940 -10540 10985 -10420
rect 11105 -10540 11150 -10420
rect 11270 -10540 11325 -10420
rect 11445 -10540 11490 -10420
rect 11610 -10540 11655 -10420
rect 11775 -10540 11820 -10420
rect 11940 -10540 11995 -10420
rect 12115 -10540 12160 -10420
rect 12280 -10540 12325 -10420
rect 12445 -10540 12490 -10420
rect 12610 -10540 12620 -10420
rect 7120 -10585 12620 -10540
rect 7120 -10705 7130 -10585
rect 7250 -10705 7305 -10585
rect 7425 -10705 7470 -10585
rect 7590 -10705 7635 -10585
rect 7755 -10705 7800 -10585
rect 7920 -10705 7975 -10585
rect 8095 -10705 8140 -10585
rect 8260 -10705 8305 -10585
rect 8425 -10705 8470 -10585
rect 8590 -10705 8645 -10585
rect 8765 -10705 8810 -10585
rect 8930 -10705 8975 -10585
rect 9095 -10705 9140 -10585
rect 9260 -10705 9315 -10585
rect 9435 -10705 9480 -10585
rect 9600 -10705 9645 -10585
rect 9765 -10705 9810 -10585
rect 9930 -10705 9985 -10585
rect 10105 -10705 10150 -10585
rect 10270 -10705 10315 -10585
rect 10435 -10705 10480 -10585
rect 10600 -10705 10655 -10585
rect 10775 -10705 10820 -10585
rect 10940 -10705 10985 -10585
rect 11105 -10705 11150 -10585
rect 11270 -10705 11325 -10585
rect 11445 -10705 11490 -10585
rect 11610 -10705 11655 -10585
rect 11775 -10705 11820 -10585
rect 11940 -10705 11995 -10585
rect 12115 -10705 12160 -10585
rect 12280 -10705 12325 -10585
rect 12445 -10705 12490 -10585
rect 12610 -10705 12620 -10585
rect 7120 -10760 12620 -10705
rect 7120 -10880 7130 -10760
rect 7250 -10880 7305 -10760
rect 7425 -10880 7470 -10760
rect 7590 -10880 7635 -10760
rect 7755 -10880 7800 -10760
rect 7920 -10880 7975 -10760
rect 8095 -10880 8140 -10760
rect 8260 -10880 8305 -10760
rect 8425 -10880 8470 -10760
rect 8590 -10880 8645 -10760
rect 8765 -10880 8810 -10760
rect 8930 -10880 8975 -10760
rect 9095 -10880 9140 -10760
rect 9260 -10880 9315 -10760
rect 9435 -10880 9480 -10760
rect 9600 -10880 9645 -10760
rect 9765 -10880 9810 -10760
rect 9930 -10880 9985 -10760
rect 10105 -10880 10150 -10760
rect 10270 -10880 10315 -10760
rect 10435 -10880 10480 -10760
rect 10600 -10880 10655 -10760
rect 10775 -10880 10820 -10760
rect 10940 -10880 10985 -10760
rect 11105 -10880 11150 -10760
rect 11270 -10880 11325 -10760
rect 11445 -10880 11490 -10760
rect 11610 -10880 11655 -10760
rect 11775 -10880 11820 -10760
rect 11940 -10880 11995 -10760
rect 12115 -10880 12160 -10760
rect 12280 -10880 12325 -10760
rect 12445 -10880 12490 -10760
rect 12610 -10880 12620 -10760
rect 7120 -10925 12620 -10880
rect 7120 -11045 7130 -10925
rect 7250 -11045 7305 -10925
rect 7425 -11045 7470 -10925
rect 7590 -11045 7635 -10925
rect 7755 -11045 7800 -10925
rect 7920 -11045 7975 -10925
rect 8095 -11045 8140 -10925
rect 8260 -11045 8305 -10925
rect 8425 -11045 8470 -10925
rect 8590 -11045 8645 -10925
rect 8765 -11045 8810 -10925
rect 8930 -11045 8975 -10925
rect 9095 -11045 9140 -10925
rect 9260 -11045 9315 -10925
rect 9435 -11045 9480 -10925
rect 9600 -11045 9645 -10925
rect 9765 -11045 9810 -10925
rect 9930 -11045 9985 -10925
rect 10105 -11045 10150 -10925
rect 10270 -11045 10315 -10925
rect 10435 -11045 10480 -10925
rect 10600 -11045 10655 -10925
rect 10775 -11045 10820 -10925
rect 10940 -11045 10985 -10925
rect 11105 -11045 11150 -10925
rect 11270 -11045 11325 -10925
rect 11445 -11045 11490 -10925
rect 11610 -11045 11655 -10925
rect 11775 -11045 11820 -10925
rect 11940 -11045 11995 -10925
rect 12115 -11045 12160 -10925
rect 12280 -11045 12325 -10925
rect 12445 -11045 12490 -10925
rect 12610 -11045 12620 -10925
rect 7120 -11090 12620 -11045
rect 7120 -11210 7130 -11090
rect 7250 -11210 7305 -11090
rect 7425 -11210 7470 -11090
rect 7590 -11210 7635 -11090
rect 7755 -11210 7800 -11090
rect 7920 -11210 7975 -11090
rect 8095 -11210 8140 -11090
rect 8260 -11210 8305 -11090
rect 8425 -11210 8470 -11090
rect 8590 -11210 8645 -11090
rect 8765 -11210 8810 -11090
rect 8930 -11210 8975 -11090
rect 9095 -11210 9140 -11090
rect 9260 -11210 9315 -11090
rect 9435 -11210 9480 -11090
rect 9600 -11210 9645 -11090
rect 9765 -11210 9810 -11090
rect 9930 -11210 9985 -11090
rect 10105 -11210 10150 -11090
rect 10270 -11210 10315 -11090
rect 10435 -11210 10480 -11090
rect 10600 -11210 10655 -11090
rect 10775 -11210 10820 -11090
rect 10940 -11210 10985 -11090
rect 11105 -11210 11150 -11090
rect 11270 -11210 11325 -11090
rect 11445 -11210 11490 -11090
rect 11610 -11210 11655 -11090
rect 11775 -11210 11820 -11090
rect 11940 -11210 11995 -11090
rect 12115 -11210 12160 -11090
rect 12280 -11210 12325 -11090
rect 12445 -11210 12490 -11090
rect 12610 -11210 12620 -11090
rect 7120 -11255 12620 -11210
rect 7120 -11375 7130 -11255
rect 7250 -11375 7305 -11255
rect 7425 -11375 7470 -11255
rect 7590 -11375 7635 -11255
rect 7755 -11375 7800 -11255
rect 7920 -11375 7975 -11255
rect 8095 -11375 8140 -11255
rect 8260 -11375 8305 -11255
rect 8425 -11375 8470 -11255
rect 8590 -11375 8645 -11255
rect 8765 -11375 8810 -11255
rect 8930 -11375 8975 -11255
rect 9095 -11375 9140 -11255
rect 9260 -11375 9315 -11255
rect 9435 -11375 9480 -11255
rect 9600 -11375 9645 -11255
rect 9765 -11375 9810 -11255
rect 9930 -11375 9985 -11255
rect 10105 -11375 10150 -11255
rect 10270 -11375 10315 -11255
rect 10435 -11375 10480 -11255
rect 10600 -11375 10655 -11255
rect 10775 -11375 10820 -11255
rect 10940 -11375 10985 -11255
rect 11105 -11375 11150 -11255
rect 11270 -11375 11325 -11255
rect 11445 -11375 11490 -11255
rect 11610 -11375 11655 -11255
rect 11775 -11375 11820 -11255
rect 11940 -11375 11995 -11255
rect 12115 -11375 12160 -11255
rect 12280 -11375 12325 -11255
rect 12445 -11375 12490 -11255
rect 12610 -11375 12620 -11255
rect 7120 -11430 12620 -11375
rect 7120 -11550 7130 -11430
rect 7250 -11550 7305 -11430
rect 7425 -11550 7470 -11430
rect 7590 -11550 7635 -11430
rect 7755 -11550 7800 -11430
rect 7920 -11550 7975 -11430
rect 8095 -11550 8140 -11430
rect 8260 -11550 8305 -11430
rect 8425 -11550 8470 -11430
rect 8590 -11550 8645 -11430
rect 8765 -11550 8810 -11430
rect 8930 -11550 8975 -11430
rect 9095 -11550 9140 -11430
rect 9260 -11550 9315 -11430
rect 9435 -11550 9480 -11430
rect 9600 -11550 9645 -11430
rect 9765 -11550 9810 -11430
rect 9930 -11550 9985 -11430
rect 10105 -11550 10150 -11430
rect 10270 -11550 10315 -11430
rect 10435 -11550 10480 -11430
rect 10600 -11550 10655 -11430
rect 10775 -11550 10820 -11430
rect 10940 -11550 10985 -11430
rect 11105 -11550 11150 -11430
rect 11270 -11550 11325 -11430
rect 11445 -11550 11490 -11430
rect 11610 -11550 11655 -11430
rect 11775 -11550 11820 -11430
rect 11940 -11550 11995 -11430
rect 12115 -11550 12160 -11430
rect 12280 -11550 12325 -11430
rect 12445 -11550 12490 -11430
rect 12610 -11550 12620 -11430
rect 7120 -11595 12620 -11550
rect 7120 -11715 7130 -11595
rect 7250 -11715 7305 -11595
rect 7425 -11715 7470 -11595
rect 7590 -11715 7635 -11595
rect 7755 -11715 7800 -11595
rect 7920 -11715 7975 -11595
rect 8095 -11715 8140 -11595
rect 8260 -11715 8305 -11595
rect 8425 -11715 8470 -11595
rect 8590 -11715 8645 -11595
rect 8765 -11715 8810 -11595
rect 8930 -11715 8975 -11595
rect 9095 -11715 9140 -11595
rect 9260 -11715 9315 -11595
rect 9435 -11715 9480 -11595
rect 9600 -11715 9645 -11595
rect 9765 -11715 9810 -11595
rect 9930 -11715 9985 -11595
rect 10105 -11715 10150 -11595
rect 10270 -11715 10315 -11595
rect 10435 -11715 10480 -11595
rect 10600 -11715 10655 -11595
rect 10775 -11715 10820 -11595
rect 10940 -11715 10985 -11595
rect 11105 -11715 11150 -11595
rect 11270 -11715 11325 -11595
rect 11445 -11715 11490 -11595
rect 11610 -11715 11655 -11595
rect 11775 -11715 11820 -11595
rect 11940 -11715 11995 -11595
rect 12115 -11715 12160 -11595
rect 12280 -11715 12325 -11595
rect 12445 -11715 12490 -11595
rect 12610 -11715 12620 -11595
rect 7120 -11760 12620 -11715
rect 7120 -11880 7130 -11760
rect 7250 -11880 7305 -11760
rect 7425 -11880 7470 -11760
rect 7590 -11880 7635 -11760
rect 7755 -11880 7800 -11760
rect 7920 -11880 7975 -11760
rect 8095 -11880 8140 -11760
rect 8260 -11880 8305 -11760
rect 8425 -11880 8470 -11760
rect 8590 -11880 8645 -11760
rect 8765 -11880 8810 -11760
rect 8930 -11880 8975 -11760
rect 9095 -11880 9140 -11760
rect 9260 -11880 9315 -11760
rect 9435 -11880 9480 -11760
rect 9600 -11880 9645 -11760
rect 9765 -11880 9810 -11760
rect 9930 -11880 9985 -11760
rect 10105 -11880 10150 -11760
rect 10270 -11880 10315 -11760
rect 10435 -11880 10480 -11760
rect 10600 -11880 10655 -11760
rect 10775 -11880 10820 -11760
rect 10940 -11880 10985 -11760
rect 11105 -11880 11150 -11760
rect 11270 -11880 11325 -11760
rect 11445 -11880 11490 -11760
rect 11610 -11880 11655 -11760
rect 11775 -11880 11820 -11760
rect 11940 -11880 11995 -11760
rect 12115 -11880 12160 -11760
rect 12280 -11880 12325 -11760
rect 12445 -11880 12490 -11760
rect 12610 -11880 12620 -11760
rect 7120 -11925 12620 -11880
rect 7120 -12045 7130 -11925
rect 7250 -12045 7305 -11925
rect 7425 -12045 7470 -11925
rect 7590 -12045 7635 -11925
rect 7755 -12045 7800 -11925
rect 7920 -12045 7975 -11925
rect 8095 -12045 8140 -11925
rect 8260 -12045 8305 -11925
rect 8425 -12045 8470 -11925
rect 8590 -12045 8645 -11925
rect 8765 -12045 8810 -11925
rect 8930 -12045 8975 -11925
rect 9095 -12045 9140 -11925
rect 9260 -12045 9315 -11925
rect 9435 -12045 9480 -11925
rect 9600 -12045 9645 -11925
rect 9765 -12045 9810 -11925
rect 9930 -12045 9985 -11925
rect 10105 -12045 10150 -11925
rect 10270 -12045 10315 -11925
rect 10435 -12045 10480 -11925
rect 10600 -12045 10655 -11925
rect 10775 -12045 10820 -11925
rect 10940 -12045 10985 -11925
rect 11105 -12045 11150 -11925
rect 11270 -12045 11325 -11925
rect 11445 -12045 11490 -11925
rect 11610 -12045 11655 -11925
rect 11775 -12045 11820 -11925
rect 11940 -12045 11995 -11925
rect 12115 -12045 12160 -11925
rect 12280 -12045 12325 -11925
rect 12445 -12045 12490 -11925
rect 12610 -12045 12620 -11925
rect 7120 -12100 12620 -12045
rect 7120 -12220 7130 -12100
rect 7250 -12220 7305 -12100
rect 7425 -12220 7470 -12100
rect 7590 -12220 7635 -12100
rect 7755 -12220 7800 -12100
rect 7920 -12220 7975 -12100
rect 8095 -12220 8140 -12100
rect 8260 -12220 8305 -12100
rect 8425 -12220 8470 -12100
rect 8590 -12220 8645 -12100
rect 8765 -12220 8810 -12100
rect 8930 -12220 8975 -12100
rect 9095 -12220 9140 -12100
rect 9260 -12220 9315 -12100
rect 9435 -12220 9480 -12100
rect 9600 -12220 9645 -12100
rect 9765 -12220 9810 -12100
rect 9930 -12220 9985 -12100
rect 10105 -12220 10150 -12100
rect 10270 -12220 10315 -12100
rect 10435 -12220 10480 -12100
rect 10600 -12220 10655 -12100
rect 10775 -12220 10820 -12100
rect 10940 -12220 10985 -12100
rect 11105 -12220 11150 -12100
rect 11270 -12220 11325 -12100
rect 11445 -12220 11490 -12100
rect 11610 -12220 11655 -12100
rect 11775 -12220 11820 -12100
rect 11940 -12220 11995 -12100
rect 12115 -12220 12160 -12100
rect 12280 -12220 12325 -12100
rect 12445 -12220 12490 -12100
rect 12610 -12220 12620 -12100
rect 7120 -12265 12620 -12220
rect 7120 -12385 7130 -12265
rect 7250 -12385 7305 -12265
rect 7425 -12385 7470 -12265
rect 7590 -12385 7635 -12265
rect 7755 -12385 7800 -12265
rect 7920 -12385 7975 -12265
rect 8095 -12385 8140 -12265
rect 8260 -12385 8305 -12265
rect 8425 -12385 8470 -12265
rect 8590 -12385 8645 -12265
rect 8765 -12385 8810 -12265
rect 8930 -12385 8975 -12265
rect 9095 -12385 9140 -12265
rect 9260 -12385 9315 -12265
rect 9435 -12385 9480 -12265
rect 9600 -12385 9645 -12265
rect 9765 -12385 9810 -12265
rect 9930 -12385 9985 -12265
rect 10105 -12385 10150 -12265
rect 10270 -12385 10315 -12265
rect 10435 -12385 10480 -12265
rect 10600 -12385 10655 -12265
rect 10775 -12385 10820 -12265
rect 10940 -12385 10985 -12265
rect 11105 -12385 11150 -12265
rect 11270 -12385 11325 -12265
rect 11445 -12385 11490 -12265
rect 11610 -12385 11655 -12265
rect 11775 -12385 11820 -12265
rect 11940 -12385 11995 -12265
rect 12115 -12385 12160 -12265
rect 12280 -12385 12325 -12265
rect 12445 -12385 12490 -12265
rect 12610 -12385 12620 -12265
rect 7120 -12430 12620 -12385
rect 7120 -12550 7130 -12430
rect 7250 -12550 7305 -12430
rect 7425 -12550 7470 -12430
rect 7590 -12550 7635 -12430
rect 7755 -12550 7800 -12430
rect 7920 -12550 7975 -12430
rect 8095 -12550 8140 -12430
rect 8260 -12550 8305 -12430
rect 8425 -12550 8470 -12430
rect 8590 -12550 8645 -12430
rect 8765 -12550 8810 -12430
rect 8930 -12550 8975 -12430
rect 9095 -12550 9140 -12430
rect 9260 -12550 9315 -12430
rect 9435 -12550 9480 -12430
rect 9600 -12550 9645 -12430
rect 9765 -12550 9810 -12430
rect 9930 -12550 9985 -12430
rect 10105 -12550 10150 -12430
rect 10270 -12550 10315 -12430
rect 10435 -12550 10480 -12430
rect 10600 -12550 10655 -12430
rect 10775 -12550 10820 -12430
rect 10940 -12550 10985 -12430
rect 11105 -12550 11150 -12430
rect 11270 -12550 11325 -12430
rect 11445 -12550 11490 -12430
rect 11610 -12550 11655 -12430
rect 11775 -12550 11820 -12430
rect 11940 -12550 11995 -12430
rect 12115 -12550 12160 -12430
rect 12280 -12550 12325 -12430
rect 12445 -12550 12490 -12430
rect 12610 -12550 12620 -12430
rect 7120 -12595 12620 -12550
rect 7120 -12715 7130 -12595
rect 7250 -12715 7305 -12595
rect 7425 -12715 7470 -12595
rect 7590 -12715 7635 -12595
rect 7755 -12715 7800 -12595
rect 7920 -12715 7975 -12595
rect 8095 -12715 8140 -12595
rect 8260 -12715 8305 -12595
rect 8425 -12715 8470 -12595
rect 8590 -12715 8645 -12595
rect 8765 -12715 8810 -12595
rect 8930 -12715 8975 -12595
rect 9095 -12715 9140 -12595
rect 9260 -12715 9315 -12595
rect 9435 -12715 9480 -12595
rect 9600 -12715 9645 -12595
rect 9765 -12715 9810 -12595
rect 9930 -12715 9985 -12595
rect 10105 -12715 10150 -12595
rect 10270 -12715 10315 -12595
rect 10435 -12715 10480 -12595
rect 10600 -12715 10655 -12595
rect 10775 -12715 10820 -12595
rect 10940 -12715 10985 -12595
rect 11105 -12715 11150 -12595
rect 11270 -12715 11325 -12595
rect 11445 -12715 11490 -12595
rect 11610 -12715 11655 -12595
rect 11775 -12715 11820 -12595
rect 11940 -12715 11995 -12595
rect 12115 -12715 12160 -12595
rect 12280 -12715 12325 -12595
rect 12445 -12715 12490 -12595
rect 12610 -12715 12620 -12595
rect 7120 -12770 12620 -12715
rect 7120 -12890 7130 -12770
rect 7250 -12890 7305 -12770
rect 7425 -12890 7470 -12770
rect 7590 -12890 7635 -12770
rect 7755 -12890 7800 -12770
rect 7920 -12890 7975 -12770
rect 8095 -12890 8140 -12770
rect 8260 -12890 8305 -12770
rect 8425 -12890 8470 -12770
rect 8590 -12890 8645 -12770
rect 8765 -12890 8810 -12770
rect 8930 -12890 8975 -12770
rect 9095 -12890 9140 -12770
rect 9260 -12890 9315 -12770
rect 9435 -12890 9480 -12770
rect 9600 -12890 9645 -12770
rect 9765 -12890 9810 -12770
rect 9930 -12890 9985 -12770
rect 10105 -12890 10150 -12770
rect 10270 -12890 10315 -12770
rect 10435 -12890 10480 -12770
rect 10600 -12890 10655 -12770
rect 10775 -12890 10820 -12770
rect 10940 -12890 10985 -12770
rect 11105 -12890 11150 -12770
rect 11270 -12890 11325 -12770
rect 11445 -12890 11490 -12770
rect 11610 -12890 11655 -12770
rect 11775 -12890 11820 -12770
rect 11940 -12890 11995 -12770
rect 12115 -12890 12160 -12770
rect 12280 -12890 12325 -12770
rect 12445 -12890 12490 -12770
rect 12610 -12890 12620 -12770
rect 7120 -12935 12620 -12890
rect 7120 -13055 7130 -12935
rect 7250 -13055 7305 -12935
rect 7425 -13055 7470 -12935
rect 7590 -13055 7635 -12935
rect 7755 -13055 7800 -12935
rect 7920 -13055 7975 -12935
rect 8095 -13055 8140 -12935
rect 8260 -13055 8305 -12935
rect 8425 -13055 8470 -12935
rect 8590 -13055 8645 -12935
rect 8765 -13055 8810 -12935
rect 8930 -13055 8975 -12935
rect 9095 -13055 9140 -12935
rect 9260 -13055 9315 -12935
rect 9435 -13055 9480 -12935
rect 9600 -13055 9645 -12935
rect 9765 -13055 9810 -12935
rect 9930 -13055 9985 -12935
rect 10105 -13055 10150 -12935
rect 10270 -13055 10315 -12935
rect 10435 -13055 10480 -12935
rect 10600 -13055 10655 -12935
rect 10775 -13055 10820 -12935
rect 10940 -13055 10985 -12935
rect 11105 -13055 11150 -12935
rect 11270 -13055 11325 -12935
rect 11445 -13055 11490 -12935
rect 11610 -13055 11655 -12935
rect 11775 -13055 11820 -12935
rect 11940 -13055 11995 -12935
rect 12115 -13055 12160 -12935
rect 12280 -13055 12325 -12935
rect 12445 -13055 12490 -12935
rect 12610 -13055 12620 -12935
rect 7120 -13100 12620 -13055
rect 7120 -13220 7130 -13100
rect 7250 -13220 7305 -13100
rect 7425 -13220 7470 -13100
rect 7590 -13220 7635 -13100
rect 7755 -13220 7800 -13100
rect 7920 -13220 7975 -13100
rect 8095 -13220 8140 -13100
rect 8260 -13220 8305 -13100
rect 8425 -13220 8470 -13100
rect 8590 -13220 8645 -13100
rect 8765 -13220 8810 -13100
rect 8930 -13220 8975 -13100
rect 9095 -13220 9140 -13100
rect 9260 -13220 9315 -13100
rect 9435 -13220 9480 -13100
rect 9600 -13220 9645 -13100
rect 9765 -13220 9810 -13100
rect 9930 -13220 9985 -13100
rect 10105 -13220 10150 -13100
rect 10270 -13220 10315 -13100
rect 10435 -13220 10480 -13100
rect 10600 -13220 10655 -13100
rect 10775 -13220 10820 -13100
rect 10940 -13220 10985 -13100
rect 11105 -13220 11150 -13100
rect 11270 -13220 11325 -13100
rect 11445 -13220 11490 -13100
rect 11610 -13220 11655 -13100
rect 11775 -13220 11820 -13100
rect 11940 -13220 11995 -13100
rect 12115 -13220 12160 -13100
rect 12280 -13220 12325 -13100
rect 12445 -13220 12490 -13100
rect 12610 -13220 12620 -13100
rect 7120 -13265 12620 -13220
rect 7120 -13385 7130 -13265
rect 7250 -13385 7305 -13265
rect 7425 -13385 7470 -13265
rect 7590 -13385 7635 -13265
rect 7755 -13385 7800 -13265
rect 7920 -13385 7975 -13265
rect 8095 -13385 8140 -13265
rect 8260 -13385 8305 -13265
rect 8425 -13385 8470 -13265
rect 8590 -13385 8645 -13265
rect 8765 -13385 8810 -13265
rect 8930 -13385 8975 -13265
rect 9095 -13385 9140 -13265
rect 9260 -13385 9315 -13265
rect 9435 -13385 9480 -13265
rect 9600 -13385 9645 -13265
rect 9765 -13385 9810 -13265
rect 9930 -13385 9985 -13265
rect 10105 -13385 10150 -13265
rect 10270 -13385 10315 -13265
rect 10435 -13385 10480 -13265
rect 10600 -13385 10655 -13265
rect 10775 -13385 10820 -13265
rect 10940 -13385 10985 -13265
rect 11105 -13385 11150 -13265
rect 11270 -13385 11325 -13265
rect 11445 -13385 11490 -13265
rect 11610 -13385 11655 -13265
rect 11775 -13385 11820 -13265
rect 11940 -13385 11995 -13265
rect 12115 -13385 12160 -13265
rect 12280 -13385 12325 -13265
rect 12445 -13385 12490 -13265
rect 12610 -13385 12620 -13265
rect 7120 -13440 12620 -13385
rect 7120 -13560 7130 -13440
rect 7250 -13560 7305 -13440
rect 7425 -13560 7470 -13440
rect 7590 -13560 7635 -13440
rect 7755 -13560 7800 -13440
rect 7920 -13560 7975 -13440
rect 8095 -13560 8140 -13440
rect 8260 -13560 8305 -13440
rect 8425 -13560 8470 -13440
rect 8590 -13560 8645 -13440
rect 8765 -13560 8810 -13440
rect 8930 -13560 8975 -13440
rect 9095 -13560 9140 -13440
rect 9260 -13560 9315 -13440
rect 9435 -13560 9480 -13440
rect 9600 -13560 9645 -13440
rect 9765 -13560 9810 -13440
rect 9930 -13560 9985 -13440
rect 10105 -13560 10150 -13440
rect 10270 -13560 10315 -13440
rect 10435 -13560 10480 -13440
rect 10600 -13560 10655 -13440
rect 10775 -13560 10820 -13440
rect 10940 -13560 10985 -13440
rect 11105 -13560 11150 -13440
rect 11270 -13560 11325 -13440
rect 11445 -13560 11490 -13440
rect 11610 -13560 11655 -13440
rect 11775 -13560 11820 -13440
rect 11940 -13560 11995 -13440
rect 12115 -13560 12160 -13440
rect 12280 -13560 12325 -13440
rect 12445 -13560 12490 -13440
rect 12610 -13560 12620 -13440
rect 7120 -13605 12620 -13560
rect 7120 -13725 7130 -13605
rect 7250 -13725 7305 -13605
rect 7425 -13725 7470 -13605
rect 7590 -13725 7635 -13605
rect 7755 -13725 7800 -13605
rect 7920 -13725 7975 -13605
rect 8095 -13725 8140 -13605
rect 8260 -13725 8305 -13605
rect 8425 -13725 8470 -13605
rect 8590 -13725 8645 -13605
rect 8765 -13725 8810 -13605
rect 8930 -13725 8975 -13605
rect 9095 -13725 9140 -13605
rect 9260 -13725 9315 -13605
rect 9435 -13725 9480 -13605
rect 9600 -13725 9645 -13605
rect 9765 -13725 9810 -13605
rect 9930 -13725 9985 -13605
rect 10105 -13725 10150 -13605
rect 10270 -13725 10315 -13605
rect 10435 -13725 10480 -13605
rect 10600 -13725 10655 -13605
rect 10775 -13725 10820 -13605
rect 10940 -13725 10985 -13605
rect 11105 -13725 11150 -13605
rect 11270 -13725 11325 -13605
rect 11445 -13725 11490 -13605
rect 11610 -13725 11655 -13605
rect 11775 -13725 11820 -13605
rect 11940 -13725 11995 -13605
rect 12115 -13725 12160 -13605
rect 12280 -13725 12325 -13605
rect 12445 -13725 12490 -13605
rect 12610 -13725 12620 -13605
rect 7120 -13770 12620 -13725
rect 7120 -13890 7130 -13770
rect 7250 -13890 7305 -13770
rect 7425 -13890 7470 -13770
rect 7590 -13890 7635 -13770
rect 7755 -13890 7800 -13770
rect 7920 -13890 7975 -13770
rect 8095 -13890 8140 -13770
rect 8260 -13890 8305 -13770
rect 8425 -13890 8470 -13770
rect 8590 -13890 8645 -13770
rect 8765 -13890 8810 -13770
rect 8930 -13890 8975 -13770
rect 9095 -13890 9140 -13770
rect 9260 -13890 9315 -13770
rect 9435 -13890 9480 -13770
rect 9600 -13890 9645 -13770
rect 9765 -13890 9810 -13770
rect 9930 -13890 9985 -13770
rect 10105 -13890 10150 -13770
rect 10270 -13890 10315 -13770
rect 10435 -13890 10480 -13770
rect 10600 -13890 10655 -13770
rect 10775 -13890 10820 -13770
rect 10940 -13890 10985 -13770
rect 11105 -13890 11150 -13770
rect 11270 -13890 11325 -13770
rect 11445 -13890 11490 -13770
rect 11610 -13890 11655 -13770
rect 11775 -13890 11820 -13770
rect 11940 -13890 11995 -13770
rect 12115 -13890 12160 -13770
rect 12280 -13890 12325 -13770
rect 12445 -13890 12490 -13770
rect 12610 -13890 12620 -13770
rect 7120 -13935 12620 -13890
rect 7120 -14055 7130 -13935
rect 7250 -14055 7305 -13935
rect 7425 -14055 7470 -13935
rect 7590 -14055 7635 -13935
rect 7755 -14055 7800 -13935
rect 7920 -14055 7975 -13935
rect 8095 -14055 8140 -13935
rect 8260 -14055 8305 -13935
rect 8425 -14055 8470 -13935
rect 8590 -14055 8645 -13935
rect 8765 -14055 8810 -13935
rect 8930 -14055 8975 -13935
rect 9095 -14055 9140 -13935
rect 9260 -14055 9315 -13935
rect 9435 -14055 9480 -13935
rect 9600 -14055 9645 -13935
rect 9765 -14055 9810 -13935
rect 9930 -14055 9985 -13935
rect 10105 -14055 10150 -13935
rect 10270 -14055 10315 -13935
rect 10435 -14055 10480 -13935
rect 10600 -14055 10655 -13935
rect 10775 -14055 10820 -13935
rect 10940 -14055 10985 -13935
rect 11105 -14055 11150 -13935
rect 11270 -14055 11325 -13935
rect 11445 -14055 11490 -13935
rect 11610 -14055 11655 -13935
rect 11775 -14055 11820 -13935
rect 11940 -14055 11995 -13935
rect 12115 -14055 12160 -13935
rect 12280 -14055 12325 -13935
rect 12445 -14055 12490 -13935
rect 12610 -14055 12620 -13935
rect 7120 -14110 12620 -14055
rect 7120 -14230 7130 -14110
rect 7250 -14230 7305 -14110
rect 7425 -14230 7470 -14110
rect 7590 -14230 7635 -14110
rect 7755 -14230 7800 -14110
rect 7920 -14230 7975 -14110
rect 8095 -14230 8140 -14110
rect 8260 -14230 8305 -14110
rect 8425 -14230 8470 -14110
rect 8590 -14230 8645 -14110
rect 8765 -14230 8810 -14110
rect 8930 -14230 8975 -14110
rect 9095 -14230 9140 -14110
rect 9260 -14230 9315 -14110
rect 9435 -14230 9480 -14110
rect 9600 -14230 9645 -14110
rect 9765 -14230 9810 -14110
rect 9930 -14230 9985 -14110
rect 10105 -14230 10150 -14110
rect 10270 -14230 10315 -14110
rect 10435 -14230 10480 -14110
rect 10600 -14230 10655 -14110
rect 10775 -14230 10820 -14110
rect 10940 -14230 10985 -14110
rect 11105 -14230 11150 -14110
rect 11270 -14230 11325 -14110
rect 11445 -14230 11490 -14110
rect 11610 -14230 11655 -14110
rect 11775 -14230 11820 -14110
rect 11940 -14230 11995 -14110
rect 12115 -14230 12160 -14110
rect 12280 -14230 12325 -14110
rect 12445 -14230 12490 -14110
rect 12610 -14230 12620 -14110
rect 7120 -14275 12620 -14230
rect 7120 -14395 7130 -14275
rect 7250 -14395 7305 -14275
rect 7425 -14395 7470 -14275
rect 7590 -14395 7635 -14275
rect 7755 -14395 7800 -14275
rect 7920 -14395 7975 -14275
rect 8095 -14395 8140 -14275
rect 8260 -14395 8305 -14275
rect 8425 -14395 8470 -14275
rect 8590 -14395 8645 -14275
rect 8765 -14395 8810 -14275
rect 8930 -14395 8975 -14275
rect 9095 -14395 9140 -14275
rect 9260 -14395 9315 -14275
rect 9435 -14395 9480 -14275
rect 9600 -14395 9645 -14275
rect 9765 -14395 9810 -14275
rect 9930 -14395 9985 -14275
rect 10105 -14395 10150 -14275
rect 10270 -14395 10315 -14275
rect 10435 -14395 10480 -14275
rect 10600 -14395 10655 -14275
rect 10775 -14395 10820 -14275
rect 10940 -14395 10985 -14275
rect 11105 -14395 11150 -14275
rect 11270 -14395 11325 -14275
rect 11445 -14395 11490 -14275
rect 11610 -14395 11655 -14275
rect 11775 -14395 11820 -14275
rect 11940 -14395 11995 -14275
rect 12115 -14395 12160 -14275
rect 12280 -14395 12325 -14275
rect 12445 -14395 12490 -14275
rect 12610 -14395 12620 -14275
rect 7120 -14440 12620 -14395
rect 7120 -14560 7130 -14440
rect 7250 -14560 7305 -14440
rect 7425 -14560 7470 -14440
rect 7590 -14560 7635 -14440
rect 7755 -14560 7800 -14440
rect 7920 -14560 7975 -14440
rect 8095 -14560 8140 -14440
rect 8260 -14560 8305 -14440
rect 8425 -14560 8470 -14440
rect 8590 -14560 8645 -14440
rect 8765 -14560 8810 -14440
rect 8930 -14560 8975 -14440
rect 9095 -14560 9140 -14440
rect 9260 -14560 9315 -14440
rect 9435 -14560 9480 -14440
rect 9600 -14560 9645 -14440
rect 9765 -14560 9810 -14440
rect 9930 -14560 9985 -14440
rect 10105 -14560 10150 -14440
rect 10270 -14560 10315 -14440
rect 10435 -14560 10480 -14440
rect 10600 -14560 10655 -14440
rect 10775 -14560 10820 -14440
rect 10940 -14560 10985 -14440
rect 11105 -14560 11150 -14440
rect 11270 -14560 11325 -14440
rect 11445 -14560 11490 -14440
rect 11610 -14560 11655 -14440
rect 11775 -14560 11820 -14440
rect 11940 -14560 11995 -14440
rect 12115 -14560 12160 -14440
rect 12280 -14560 12325 -14440
rect 12445 -14560 12490 -14440
rect 12610 -14560 12620 -14440
rect 7120 -14605 12620 -14560
rect 7120 -14725 7130 -14605
rect 7250 -14725 7305 -14605
rect 7425 -14725 7470 -14605
rect 7590 -14725 7635 -14605
rect 7755 -14725 7800 -14605
rect 7920 -14725 7975 -14605
rect 8095 -14725 8140 -14605
rect 8260 -14725 8305 -14605
rect 8425 -14725 8470 -14605
rect 8590 -14725 8645 -14605
rect 8765 -14725 8810 -14605
rect 8930 -14725 8975 -14605
rect 9095 -14725 9140 -14605
rect 9260 -14725 9315 -14605
rect 9435 -14725 9480 -14605
rect 9600 -14725 9645 -14605
rect 9765 -14725 9810 -14605
rect 9930 -14725 9985 -14605
rect 10105 -14725 10150 -14605
rect 10270 -14725 10315 -14605
rect 10435 -14725 10480 -14605
rect 10600 -14725 10655 -14605
rect 10775 -14725 10820 -14605
rect 10940 -14725 10985 -14605
rect 11105 -14725 11150 -14605
rect 11270 -14725 11325 -14605
rect 11445 -14725 11490 -14605
rect 11610 -14725 11655 -14605
rect 11775 -14725 11820 -14605
rect 11940 -14725 11995 -14605
rect 12115 -14725 12160 -14605
rect 12280 -14725 12325 -14605
rect 12445 -14725 12490 -14605
rect 12610 -14725 12620 -14605
rect 7120 -14780 12620 -14725
rect 7120 -14900 7130 -14780
rect 7250 -14900 7305 -14780
rect 7425 -14900 7470 -14780
rect 7590 -14900 7635 -14780
rect 7755 -14900 7800 -14780
rect 7920 -14900 7975 -14780
rect 8095 -14900 8140 -14780
rect 8260 -14900 8305 -14780
rect 8425 -14900 8470 -14780
rect 8590 -14900 8645 -14780
rect 8765 -14900 8810 -14780
rect 8930 -14900 8975 -14780
rect 9095 -14900 9140 -14780
rect 9260 -14900 9315 -14780
rect 9435 -14900 9480 -14780
rect 9600 -14900 9645 -14780
rect 9765 -14900 9810 -14780
rect 9930 -14900 9985 -14780
rect 10105 -14900 10150 -14780
rect 10270 -14900 10315 -14780
rect 10435 -14900 10480 -14780
rect 10600 -14900 10655 -14780
rect 10775 -14900 10820 -14780
rect 10940 -14900 10985 -14780
rect 11105 -14900 11150 -14780
rect 11270 -14900 11325 -14780
rect 11445 -14900 11490 -14780
rect 11610 -14900 11655 -14780
rect 11775 -14900 11820 -14780
rect 11940 -14900 11995 -14780
rect 12115 -14900 12160 -14780
rect 12280 -14900 12325 -14780
rect 12445 -14900 12490 -14780
rect 12610 -14900 12620 -14780
rect 7120 -14945 12620 -14900
rect 7120 -15065 7130 -14945
rect 7250 -15065 7305 -14945
rect 7425 -15065 7470 -14945
rect 7590 -15065 7635 -14945
rect 7755 -15065 7800 -14945
rect 7920 -15065 7975 -14945
rect 8095 -15065 8140 -14945
rect 8260 -15065 8305 -14945
rect 8425 -15065 8470 -14945
rect 8590 -15065 8645 -14945
rect 8765 -15065 8810 -14945
rect 8930 -15065 8975 -14945
rect 9095 -15065 9140 -14945
rect 9260 -15065 9315 -14945
rect 9435 -15065 9480 -14945
rect 9600 -15065 9645 -14945
rect 9765 -15065 9810 -14945
rect 9930 -15065 9985 -14945
rect 10105 -15065 10150 -14945
rect 10270 -15065 10315 -14945
rect 10435 -15065 10480 -14945
rect 10600 -15065 10655 -14945
rect 10775 -15065 10820 -14945
rect 10940 -15065 10985 -14945
rect 11105 -15065 11150 -14945
rect 11270 -15065 11325 -14945
rect 11445 -15065 11490 -14945
rect 11610 -15065 11655 -14945
rect 11775 -15065 11820 -14945
rect 11940 -15065 11995 -14945
rect 12115 -15065 12160 -14945
rect 12280 -15065 12325 -14945
rect 12445 -15065 12490 -14945
rect 12610 -15065 12620 -14945
rect 7120 -15110 12620 -15065
rect 7120 -15230 7130 -15110
rect 7250 -15230 7305 -15110
rect 7425 -15230 7470 -15110
rect 7590 -15230 7635 -15110
rect 7755 -15230 7800 -15110
rect 7920 -15230 7975 -15110
rect 8095 -15230 8140 -15110
rect 8260 -15230 8305 -15110
rect 8425 -15230 8470 -15110
rect 8590 -15230 8645 -15110
rect 8765 -15230 8810 -15110
rect 8930 -15230 8975 -15110
rect 9095 -15230 9140 -15110
rect 9260 -15230 9315 -15110
rect 9435 -15230 9480 -15110
rect 9600 -15230 9645 -15110
rect 9765 -15230 9810 -15110
rect 9930 -15230 9985 -15110
rect 10105 -15230 10150 -15110
rect 10270 -15230 10315 -15110
rect 10435 -15230 10480 -15110
rect 10600 -15230 10655 -15110
rect 10775 -15230 10820 -15110
rect 10940 -15230 10985 -15110
rect 11105 -15230 11150 -15110
rect 11270 -15230 11325 -15110
rect 11445 -15230 11490 -15110
rect 11610 -15230 11655 -15110
rect 11775 -15230 11820 -15110
rect 11940 -15230 11995 -15110
rect 12115 -15230 12160 -15110
rect 12280 -15230 12325 -15110
rect 12445 -15230 12490 -15110
rect 12610 -15230 12620 -15110
rect 7120 -15275 12620 -15230
rect 7120 -15395 7130 -15275
rect 7250 -15395 7305 -15275
rect 7425 -15395 7470 -15275
rect 7590 -15395 7635 -15275
rect 7755 -15395 7800 -15275
rect 7920 -15395 7975 -15275
rect 8095 -15395 8140 -15275
rect 8260 -15395 8305 -15275
rect 8425 -15395 8470 -15275
rect 8590 -15395 8645 -15275
rect 8765 -15395 8810 -15275
rect 8930 -15395 8975 -15275
rect 9095 -15395 9140 -15275
rect 9260 -15395 9315 -15275
rect 9435 -15395 9480 -15275
rect 9600 -15395 9645 -15275
rect 9765 -15395 9810 -15275
rect 9930 -15395 9985 -15275
rect 10105 -15395 10150 -15275
rect 10270 -15395 10315 -15275
rect 10435 -15395 10480 -15275
rect 10600 -15395 10655 -15275
rect 10775 -15395 10820 -15275
rect 10940 -15395 10985 -15275
rect 11105 -15395 11150 -15275
rect 11270 -15395 11325 -15275
rect 11445 -15395 11490 -15275
rect 11610 -15395 11655 -15275
rect 11775 -15395 11820 -15275
rect 11940 -15395 11995 -15275
rect 12115 -15395 12160 -15275
rect 12280 -15395 12325 -15275
rect 12445 -15395 12490 -15275
rect 12610 -15395 12620 -15275
rect 7120 -15450 12620 -15395
rect 7120 -15570 7130 -15450
rect 7250 -15570 7305 -15450
rect 7425 -15570 7470 -15450
rect 7590 -15570 7635 -15450
rect 7755 -15570 7800 -15450
rect 7920 -15570 7975 -15450
rect 8095 -15570 8140 -15450
rect 8260 -15570 8305 -15450
rect 8425 -15570 8470 -15450
rect 8590 -15570 8645 -15450
rect 8765 -15570 8810 -15450
rect 8930 -15570 8975 -15450
rect 9095 -15570 9140 -15450
rect 9260 -15570 9315 -15450
rect 9435 -15570 9480 -15450
rect 9600 -15570 9645 -15450
rect 9765 -15570 9810 -15450
rect 9930 -15570 9985 -15450
rect 10105 -15570 10150 -15450
rect 10270 -15570 10315 -15450
rect 10435 -15570 10480 -15450
rect 10600 -15570 10655 -15450
rect 10775 -15570 10820 -15450
rect 10940 -15570 10985 -15450
rect 11105 -15570 11150 -15450
rect 11270 -15570 11325 -15450
rect 11445 -15570 11490 -15450
rect 11610 -15570 11655 -15450
rect 11775 -15570 11820 -15450
rect 11940 -15570 11995 -15450
rect 12115 -15570 12160 -15450
rect 12280 -15570 12325 -15450
rect 12445 -15570 12490 -15450
rect 12610 -15570 12620 -15450
rect 7120 -15580 12620 -15570
rect 12810 -10090 18310 -10080
rect 12810 -10210 12820 -10090
rect 12940 -10210 12995 -10090
rect 13115 -10210 13160 -10090
rect 13280 -10210 13325 -10090
rect 13445 -10210 13490 -10090
rect 13610 -10210 13665 -10090
rect 13785 -10210 13830 -10090
rect 13950 -10210 13995 -10090
rect 14115 -10210 14160 -10090
rect 14280 -10210 14335 -10090
rect 14455 -10210 14500 -10090
rect 14620 -10210 14665 -10090
rect 14785 -10210 14830 -10090
rect 14950 -10210 15005 -10090
rect 15125 -10210 15170 -10090
rect 15290 -10210 15335 -10090
rect 15455 -10210 15500 -10090
rect 15620 -10210 15675 -10090
rect 15795 -10210 15840 -10090
rect 15960 -10210 16005 -10090
rect 16125 -10210 16170 -10090
rect 16290 -10210 16345 -10090
rect 16465 -10210 16510 -10090
rect 16630 -10210 16675 -10090
rect 16795 -10210 16840 -10090
rect 16960 -10210 17015 -10090
rect 17135 -10210 17180 -10090
rect 17300 -10210 17345 -10090
rect 17465 -10210 17510 -10090
rect 17630 -10210 17685 -10090
rect 17805 -10210 17850 -10090
rect 17970 -10210 18015 -10090
rect 18135 -10210 18180 -10090
rect 18300 -10210 18310 -10090
rect 12810 -10255 18310 -10210
rect 12810 -10375 12820 -10255
rect 12940 -10375 12995 -10255
rect 13115 -10375 13160 -10255
rect 13280 -10375 13325 -10255
rect 13445 -10375 13490 -10255
rect 13610 -10375 13665 -10255
rect 13785 -10375 13830 -10255
rect 13950 -10375 13995 -10255
rect 14115 -10375 14160 -10255
rect 14280 -10375 14335 -10255
rect 14455 -10375 14500 -10255
rect 14620 -10375 14665 -10255
rect 14785 -10375 14830 -10255
rect 14950 -10375 15005 -10255
rect 15125 -10375 15170 -10255
rect 15290 -10375 15335 -10255
rect 15455 -10375 15500 -10255
rect 15620 -10375 15675 -10255
rect 15795 -10375 15840 -10255
rect 15960 -10375 16005 -10255
rect 16125 -10375 16170 -10255
rect 16290 -10375 16345 -10255
rect 16465 -10375 16510 -10255
rect 16630 -10375 16675 -10255
rect 16795 -10375 16840 -10255
rect 16960 -10375 17015 -10255
rect 17135 -10375 17180 -10255
rect 17300 -10375 17345 -10255
rect 17465 -10375 17510 -10255
rect 17630 -10375 17685 -10255
rect 17805 -10375 17850 -10255
rect 17970 -10375 18015 -10255
rect 18135 -10375 18180 -10255
rect 18300 -10375 18310 -10255
rect 12810 -10420 18310 -10375
rect 12810 -10540 12820 -10420
rect 12940 -10540 12995 -10420
rect 13115 -10540 13160 -10420
rect 13280 -10540 13325 -10420
rect 13445 -10540 13490 -10420
rect 13610 -10540 13665 -10420
rect 13785 -10540 13830 -10420
rect 13950 -10540 13995 -10420
rect 14115 -10540 14160 -10420
rect 14280 -10540 14335 -10420
rect 14455 -10540 14500 -10420
rect 14620 -10540 14665 -10420
rect 14785 -10540 14830 -10420
rect 14950 -10540 15005 -10420
rect 15125 -10540 15170 -10420
rect 15290 -10540 15335 -10420
rect 15455 -10540 15500 -10420
rect 15620 -10540 15675 -10420
rect 15795 -10540 15840 -10420
rect 15960 -10540 16005 -10420
rect 16125 -10540 16170 -10420
rect 16290 -10540 16345 -10420
rect 16465 -10540 16510 -10420
rect 16630 -10540 16675 -10420
rect 16795 -10540 16840 -10420
rect 16960 -10540 17015 -10420
rect 17135 -10540 17180 -10420
rect 17300 -10540 17345 -10420
rect 17465 -10540 17510 -10420
rect 17630 -10540 17685 -10420
rect 17805 -10540 17850 -10420
rect 17970 -10540 18015 -10420
rect 18135 -10540 18180 -10420
rect 18300 -10540 18310 -10420
rect 12810 -10585 18310 -10540
rect 12810 -10705 12820 -10585
rect 12940 -10705 12995 -10585
rect 13115 -10705 13160 -10585
rect 13280 -10705 13325 -10585
rect 13445 -10705 13490 -10585
rect 13610 -10705 13665 -10585
rect 13785 -10705 13830 -10585
rect 13950 -10705 13995 -10585
rect 14115 -10705 14160 -10585
rect 14280 -10705 14335 -10585
rect 14455 -10705 14500 -10585
rect 14620 -10705 14665 -10585
rect 14785 -10705 14830 -10585
rect 14950 -10705 15005 -10585
rect 15125 -10705 15170 -10585
rect 15290 -10705 15335 -10585
rect 15455 -10705 15500 -10585
rect 15620 -10705 15675 -10585
rect 15795 -10705 15840 -10585
rect 15960 -10705 16005 -10585
rect 16125 -10705 16170 -10585
rect 16290 -10705 16345 -10585
rect 16465 -10705 16510 -10585
rect 16630 -10705 16675 -10585
rect 16795 -10705 16840 -10585
rect 16960 -10705 17015 -10585
rect 17135 -10705 17180 -10585
rect 17300 -10705 17345 -10585
rect 17465 -10705 17510 -10585
rect 17630 -10705 17685 -10585
rect 17805 -10705 17850 -10585
rect 17970 -10705 18015 -10585
rect 18135 -10705 18180 -10585
rect 18300 -10705 18310 -10585
rect 12810 -10760 18310 -10705
rect 12810 -10880 12820 -10760
rect 12940 -10880 12995 -10760
rect 13115 -10880 13160 -10760
rect 13280 -10880 13325 -10760
rect 13445 -10880 13490 -10760
rect 13610 -10880 13665 -10760
rect 13785 -10880 13830 -10760
rect 13950 -10880 13995 -10760
rect 14115 -10880 14160 -10760
rect 14280 -10880 14335 -10760
rect 14455 -10880 14500 -10760
rect 14620 -10880 14665 -10760
rect 14785 -10880 14830 -10760
rect 14950 -10880 15005 -10760
rect 15125 -10880 15170 -10760
rect 15290 -10880 15335 -10760
rect 15455 -10880 15500 -10760
rect 15620 -10880 15675 -10760
rect 15795 -10880 15840 -10760
rect 15960 -10880 16005 -10760
rect 16125 -10880 16170 -10760
rect 16290 -10880 16345 -10760
rect 16465 -10880 16510 -10760
rect 16630 -10880 16675 -10760
rect 16795 -10880 16840 -10760
rect 16960 -10880 17015 -10760
rect 17135 -10880 17180 -10760
rect 17300 -10880 17345 -10760
rect 17465 -10880 17510 -10760
rect 17630 -10880 17685 -10760
rect 17805 -10880 17850 -10760
rect 17970 -10880 18015 -10760
rect 18135 -10880 18180 -10760
rect 18300 -10880 18310 -10760
rect 12810 -10925 18310 -10880
rect 12810 -11045 12820 -10925
rect 12940 -11045 12995 -10925
rect 13115 -11045 13160 -10925
rect 13280 -11045 13325 -10925
rect 13445 -11045 13490 -10925
rect 13610 -11045 13665 -10925
rect 13785 -11045 13830 -10925
rect 13950 -11045 13995 -10925
rect 14115 -11045 14160 -10925
rect 14280 -11045 14335 -10925
rect 14455 -11045 14500 -10925
rect 14620 -11045 14665 -10925
rect 14785 -11045 14830 -10925
rect 14950 -11045 15005 -10925
rect 15125 -11045 15170 -10925
rect 15290 -11045 15335 -10925
rect 15455 -11045 15500 -10925
rect 15620 -11045 15675 -10925
rect 15795 -11045 15840 -10925
rect 15960 -11045 16005 -10925
rect 16125 -11045 16170 -10925
rect 16290 -11045 16345 -10925
rect 16465 -11045 16510 -10925
rect 16630 -11045 16675 -10925
rect 16795 -11045 16840 -10925
rect 16960 -11045 17015 -10925
rect 17135 -11045 17180 -10925
rect 17300 -11045 17345 -10925
rect 17465 -11045 17510 -10925
rect 17630 -11045 17685 -10925
rect 17805 -11045 17850 -10925
rect 17970 -11045 18015 -10925
rect 18135 -11045 18180 -10925
rect 18300 -11045 18310 -10925
rect 12810 -11090 18310 -11045
rect 12810 -11210 12820 -11090
rect 12940 -11210 12995 -11090
rect 13115 -11210 13160 -11090
rect 13280 -11210 13325 -11090
rect 13445 -11210 13490 -11090
rect 13610 -11210 13665 -11090
rect 13785 -11210 13830 -11090
rect 13950 -11210 13995 -11090
rect 14115 -11210 14160 -11090
rect 14280 -11210 14335 -11090
rect 14455 -11210 14500 -11090
rect 14620 -11210 14665 -11090
rect 14785 -11210 14830 -11090
rect 14950 -11210 15005 -11090
rect 15125 -11210 15170 -11090
rect 15290 -11210 15335 -11090
rect 15455 -11210 15500 -11090
rect 15620 -11210 15675 -11090
rect 15795 -11210 15840 -11090
rect 15960 -11210 16005 -11090
rect 16125 -11210 16170 -11090
rect 16290 -11210 16345 -11090
rect 16465 -11210 16510 -11090
rect 16630 -11210 16675 -11090
rect 16795 -11210 16840 -11090
rect 16960 -11210 17015 -11090
rect 17135 -11210 17180 -11090
rect 17300 -11210 17345 -11090
rect 17465 -11210 17510 -11090
rect 17630 -11210 17685 -11090
rect 17805 -11210 17850 -11090
rect 17970 -11210 18015 -11090
rect 18135 -11210 18180 -11090
rect 18300 -11210 18310 -11090
rect 12810 -11255 18310 -11210
rect 12810 -11375 12820 -11255
rect 12940 -11375 12995 -11255
rect 13115 -11375 13160 -11255
rect 13280 -11375 13325 -11255
rect 13445 -11375 13490 -11255
rect 13610 -11375 13665 -11255
rect 13785 -11375 13830 -11255
rect 13950 -11375 13995 -11255
rect 14115 -11375 14160 -11255
rect 14280 -11375 14335 -11255
rect 14455 -11375 14500 -11255
rect 14620 -11375 14665 -11255
rect 14785 -11375 14830 -11255
rect 14950 -11375 15005 -11255
rect 15125 -11375 15170 -11255
rect 15290 -11375 15335 -11255
rect 15455 -11375 15500 -11255
rect 15620 -11375 15675 -11255
rect 15795 -11375 15840 -11255
rect 15960 -11375 16005 -11255
rect 16125 -11375 16170 -11255
rect 16290 -11375 16345 -11255
rect 16465 -11375 16510 -11255
rect 16630 -11375 16675 -11255
rect 16795 -11375 16840 -11255
rect 16960 -11375 17015 -11255
rect 17135 -11375 17180 -11255
rect 17300 -11375 17345 -11255
rect 17465 -11375 17510 -11255
rect 17630 -11375 17685 -11255
rect 17805 -11375 17850 -11255
rect 17970 -11375 18015 -11255
rect 18135 -11375 18180 -11255
rect 18300 -11375 18310 -11255
rect 12810 -11430 18310 -11375
rect 12810 -11550 12820 -11430
rect 12940 -11550 12995 -11430
rect 13115 -11550 13160 -11430
rect 13280 -11550 13325 -11430
rect 13445 -11550 13490 -11430
rect 13610 -11550 13665 -11430
rect 13785 -11550 13830 -11430
rect 13950 -11550 13995 -11430
rect 14115 -11550 14160 -11430
rect 14280 -11550 14335 -11430
rect 14455 -11550 14500 -11430
rect 14620 -11550 14665 -11430
rect 14785 -11550 14830 -11430
rect 14950 -11550 15005 -11430
rect 15125 -11550 15170 -11430
rect 15290 -11550 15335 -11430
rect 15455 -11550 15500 -11430
rect 15620 -11550 15675 -11430
rect 15795 -11550 15840 -11430
rect 15960 -11550 16005 -11430
rect 16125 -11550 16170 -11430
rect 16290 -11550 16345 -11430
rect 16465 -11550 16510 -11430
rect 16630 -11550 16675 -11430
rect 16795 -11550 16840 -11430
rect 16960 -11550 17015 -11430
rect 17135 -11550 17180 -11430
rect 17300 -11550 17345 -11430
rect 17465 -11550 17510 -11430
rect 17630 -11550 17685 -11430
rect 17805 -11550 17850 -11430
rect 17970 -11550 18015 -11430
rect 18135 -11550 18180 -11430
rect 18300 -11550 18310 -11430
rect 12810 -11595 18310 -11550
rect 12810 -11715 12820 -11595
rect 12940 -11715 12995 -11595
rect 13115 -11715 13160 -11595
rect 13280 -11715 13325 -11595
rect 13445 -11715 13490 -11595
rect 13610 -11715 13665 -11595
rect 13785 -11715 13830 -11595
rect 13950 -11715 13995 -11595
rect 14115 -11715 14160 -11595
rect 14280 -11715 14335 -11595
rect 14455 -11715 14500 -11595
rect 14620 -11715 14665 -11595
rect 14785 -11715 14830 -11595
rect 14950 -11715 15005 -11595
rect 15125 -11715 15170 -11595
rect 15290 -11715 15335 -11595
rect 15455 -11715 15500 -11595
rect 15620 -11715 15675 -11595
rect 15795 -11715 15840 -11595
rect 15960 -11715 16005 -11595
rect 16125 -11715 16170 -11595
rect 16290 -11715 16345 -11595
rect 16465 -11715 16510 -11595
rect 16630 -11715 16675 -11595
rect 16795 -11715 16840 -11595
rect 16960 -11715 17015 -11595
rect 17135 -11715 17180 -11595
rect 17300 -11715 17345 -11595
rect 17465 -11715 17510 -11595
rect 17630 -11715 17685 -11595
rect 17805 -11715 17850 -11595
rect 17970 -11715 18015 -11595
rect 18135 -11715 18180 -11595
rect 18300 -11715 18310 -11595
rect 12810 -11760 18310 -11715
rect 12810 -11880 12820 -11760
rect 12940 -11880 12995 -11760
rect 13115 -11880 13160 -11760
rect 13280 -11880 13325 -11760
rect 13445 -11880 13490 -11760
rect 13610 -11880 13665 -11760
rect 13785 -11880 13830 -11760
rect 13950 -11880 13995 -11760
rect 14115 -11880 14160 -11760
rect 14280 -11880 14335 -11760
rect 14455 -11880 14500 -11760
rect 14620 -11880 14665 -11760
rect 14785 -11880 14830 -11760
rect 14950 -11880 15005 -11760
rect 15125 -11880 15170 -11760
rect 15290 -11880 15335 -11760
rect 15455 -11880 15500 -11760
rect 15620 -11880 15675 -11760
rect 15795 -11880 15840 -11760
rect 15960 -11880 16005 -11760
rect 16125 -11880 16170 -11760
rect 16290 -11880 16345 -11760
rect 16465 -11880 16510 -11760
rect 16630 -11880 16675 -11760
rect 16795 -11880 16840 -11760
rect 16960 -11880 17015 -11760
rect 17135 -11880 17180 -11760
rect 17300 -11880 17345 -11760
rect 17465 -11880 17510 -11760
rect 17630 -11880 17685 -11760
rect 17805 -11880 17850 -11760
rect 17970 -11880 18015 -11760
rect 18135 -11880 18180 -11760
rect 18300 -11880 18310 -11760
rect 12810 -11925 18310 -11880
rect 12810 -12045 12820 -11925
rect 12940 -12045 12995 -11925
rect 13115 -12045 13160 -11925
rect 13280 -12045 13325 -11925
rect 13445 -12045 13490 -11925
rect 13610 -12045 13665 -11925
rect 13785 -12045 13830 -11925
rect 13950 -12045 13995 -11925
rect 14115 -12045 14160 -11925
rect 14280 -12045 14335 -11925
rect 14455 -12045 14500 -11925
rect 14620 -12045 14665 -11925
rect 14785 -12045 14830 -11925
rect 14950 -12045 15005 -11925
rect 15125 -12045 15170 -11925
rect 15290 -12045 15335 -11925
rect 15455 -12045 15500 -11925
rect 15620 -12045 15675 -11925
rect 15795 -12045 15840 -11925
rect 15960 -12045 16005 -11925
rect 16125 -12045 16170 -11925
rect 16290 -12045 16345 -11925
rect 16465 -12045 16510 -11925
rect 16630 -12045 16675 -11925
rect 16795 -12045 16840 -11925
rect 16960 -12045 17015 -11925
rect 17135 -12045 17180 -11925
rect 17300 -12045 17345 -11925
rect 17465 -12045 17510 -11925
rect 17630 -12045 17685 -11925
rect 17805 -12045 17850 -11925
rect 17970 -12045 18015 -11925
rect 18135 -12045 18180 -11925
rect 18300 -12045 18310 -11925
rect 12810 -12100 18310 -12045
rect 12810 -12220 12820 -12100
rect 12940 -12220 12995 -12100
rect 13115 -12220 13160 -12100
rect 13280 -12220 13325 -12100
rect 13445 -12220 13490 -12100
rect 13610 -12220 13665 -12100
rect 13785 -12220 13830 -12100
rect 13950 -12220 13995 -12100
rect 14115 -12220 14160 -12100
rect 14280 -12220 14335 -12100
rect 14455 -12220 14500 -12100
rect 14620 -12220 14665 -12100
rect 14785 -12220 14830 -12100
rect 14950 -12220 15005 -12100
rect 15125 -12220 15170 -12100
rect 15290 -12220 15335 -12100
rect 15455 -12220 15500 -12100
rect 15620 -12220 15675 -12100
rect 15795 -12220 15840 -12100
rect 15960 -12220 16005 -12100
rect 16125 -12220 16170 -12100
rect 16290 -12220 16345 -12100
rect 16465 -12220 16510 -12100
rect 16630 -12220 16675 -12100
rect 16795 -12220 16840 -12100
rect 16960 -12220 17015 -12100
rect 17135 -12220 17180 -12100
rect 17300 -12220 17345 -12100
rect 17465 -12220 17510 -12100
rect 17630 -12220 17685 -12100
rect 17805 -12220 17850 -12100
rect 17970 -12220 18015 -12100
rect 18135 -12220 18180 -12100
rect 18300 -12220 18310 -12100
rect 12810 -12265 18310 -12220
rect 12810 -12385 12820 -12265
rect 12940 -12385 12995 -12265
rect 13115 -12385 13160 -12265
rect 13280 -12385 13325 -12265
rect 13445 -12385 13490 -12265
rect 13610 -12385 13665 -12265
rect 13785 -12385 13830 -12265
rect 13950 -12385 13995 -12265
rect 14115 -12385 14160 -12265
rect 14280 -12385 14335 -12265
rect 14455 -12385 14500 -12265
rect 14620 -12385 14665 -12265
rect 14785 -12385 14830 -12265
rect 14950 -12385 15005 -12265
rect 15125 -12385 15170 -12265
rect 15290 -12385 15335 -12265
rect 15455 -12385 15500 -12265
rect 15620 -12385 15675 -12265
rect 15795 -12385 15840 -12265
rect 15960 -12385 16005 -12265
rect 16125 -12385 16170 -12265
rect 16290 -12385 16345 -12265
rect 16465 -12385 16510 -12265
rect 16630 -12385 16675 -12265
rect 16795 -12385 16840 -12265
rect 16960 -12385 17015 -12265
rect 17135 -12385 17180 -12265
rect 17300 -12385 17345 -12265
rect 17465 -12385 17510 -12265
rect 17630 -12385 17685 -12265
rect 17805 -12385 17850 -12265
rect 17970 -12385 18015 -12265
rect 18135 -12385 18180 -12265
rect 18300 -12385 18310 -12265
rect 12810 -12430 18310 -12385
rect 12810 -12550 12820 -12430
rect 12940 -12550 12995 -12430
rect 13115 -12550 13160 -12430
rect 13280 -12550 13325 -12430
rect 13445 -12550 13490 -12430
rect 13610 -12550 13665 -12430
rect 13785 -12550 13830 -12430
rect 13950 -12550 13995 -12430
rect 14115 -12550 14160 -12430
rect 14280 -12550 14335 -12430
rect 14455 -12550 14500 -12430
rect 14620 -12550 14665 -12430
rect 14785 -12550 14830 -12430
rect 14950 -12550 15005 -12430
rect 15125 -12550 15170 -12430
rect 15290 -12550 15335 -12430
rect 15455 -12550 15500 -12430
rect 15620 -12550 15675 -12430
rect 15795 -12550 15840 -12430
rect 15960 -12550 16005 -12430
rect 16125 -12550 16170 -12430
rect 16290 -12550 16345 -12430
rect 16465 -12550 16510 -12430
rect 16630 -12550 16675 -12430
rect 16795 -12550 16840 -12430
rect 16960 -12550 17015 -12430
rect 17135 -12550 17180 -12430
rect 17300 -12550 17345 -12430
rect 17465 -12550 17510 -12430
rect 17630 -12550 17685 -12430
rect 17805 -12550 17850 -12430
rect 17970 -12550 18015 -12430
rect 18135 -12550 18180 -12430
rect 18300 -12550 18310 -12430
rect 12810 -12595 18310 -12550
rect 12810 -12715 12820 -12595
rect 12940 -12715 12995 -12595
rect 13115 -12715 13160 -12595
rect 13280 -12715 13325 -12595
rect 13445 -12715 13490 -12595
rect 13610 -12715 13665 -12595
rect 13785 -12715 13830 -12595
rect 13950 -12715 13995 -12595
rect 14115 -12715 14160 -12595
rect 14280 -12715 14335 -12595
rect 14455 -12715 14500 -12595
rect 14620 -12715 14665 -12595
rect 14785 -12715 14830 -12595
rect 14950 -12715 15005 -12595
rect 15125 -12715 15170 -12595
rect 15290 -12715 15335 -12595
rect 15455 -12715 15500 -12595
rect 15620 -12715 15675 -12595
rect 15795 -12715 15840 -12595
rect 15960 -12715 16005 -12595
rect 16125 -12715 16170 -12595
rect 16290 -12715 16345 -12595
rect 16465 -12715 16510 -12595
rect 16630 -12715 16675 -12595
rect 16795 -12715 16840 -12595
rect 16960 -12715 17015 -12595
rect 17135 -12715 17180 -12595
rect 17300 -12715 17345 -12595
rect 17465 -12715 17510 -12595
rect 17630 -12715 17685 -12595
rect 17805 -12715 17850 -12595
rect 17970 -12715 18015 -12595
rect 18135 -12715 18180 -12595
rect 18300 -12715 18310 -12595
rect 12810 -12770 18310 -12715
rect 12810 -12890 12820 -12770
rect 12940 -12890 12995 -12770
rect 13115 -12890 13160 -12770
rect 13280 -12890 13325 -12770
rect 13445 -12890 13490 -12770
rect 13610 -12890 13665 -12770
rect 13785 -12890 13830 -12770
rect 13950 -12890 13995 -12770
rect 14115 -12890 14160 -12770
rect 14280 -12890 14335 -12770
rect 14455 -12890 14500 -12770
rect 14620 -12890 14665 -12770
rect 14785 -12890 14830 -12770
rect 14950 -12890 15005 -12770
rect 15125 -12890 15170 -12770
rect 15290 -12890 15335 -12770
rect 15455 -12890 15500 -12770
rect 15620 -12890 15675 -12770
rect 15795 -12890 15840 -12770
rect 15960 -12890 16005 -12770
rect 16125 -12890 16170 -12770
rect 16290 -12890 16345 -12770
rect 16465 -12890 16510 -12770
rect 16630 -12890 16675 -12770
rect 16795 -12890 16840 -12770
rect 16960 -12890 17015 -12770
rect 17135 -12890 17180 -12770
rect 17300 -12890 17345 -12770
rect 17465 -12890 17510 -12770
rect 17630 -12890 17685 -12770
rect 17805 -12890 17850 -12770
rect 17970 -12890 18015 -12770
rect 18135 -12890 18180 -12770
rect 18300 -12890 18310 -12770
rect 12810 -12935 18310 -12890
rect 12810 -13055 12820 -12935
rect 12940 -13055 12995 -12935
rect 13115 -13055 13160 -12935
rect 13280 -13055 13325 -12935
rect 13445 -13055 13490 -12935
rect 13610 -13055 13665 -12935
rect 13785 -13055 13830 -12935
rect 13950 -13055 13995 -12935
rect 14115 -13055 14160 -12935
rect 14280 -13055 14335 -12935
rect 14455 -13055 14500 -12935
rect 14620 -13055 14665 -12935
rect 14785 -13055 14830 -12935
rect 14950 -13055 15005 -12935
rect 15125 -13055 15170 -12935
rect 15290 -13055 15335 -12935
rect 15455 -13055 15500 -12935
rect 15620 -13055 15675 -12935
rect 15795 -13055 15840 -12935
rect 15960 -13055 16005 -12935
rect 16125 -13055 16170 -12935
rect 16290 -13055 16345 -12935
rect 16465 -13055 16510 -12935
rect 16630 -13055 16675 -12935
rect 16795 -13055 16840 -12935
rect 16960 -13055 17015 -12935
rect 17135 -13055 17180 -12935
rect 17300 -13055 17345 -12935
rect 17465 -13055 17510 -12935
rect 17630 -13055 17685 -12935
rect 17805 -13055 17850 -12935
rect 17970 -13055 18015 -12935
rect 18135 -13055 18180 -12935
rect 18300 -13055 18310 -12935
rect 12810 -13100 18310 -13055
rect 12810 -13220 12820 -13100
rect 12940 -13220 12995 -13100
rect 13115 -13220 13160 -13100
rect 13280 -13220 13325 -13100
rect 13445 -13220 13490 -13100
rect 13610 -13220 13665 -13100
rect 13785 -13220 13830 -13100
rect 13950 -13220 13995 -13100
rect 14115 -13220 14160 -13100
rect 14280 -13220 14335 -13100
rect 14455 -13220 14500 -13100
rect 14620 -13220 14665 -13100
rect 14785 -13220 14830 -13100
rect 14950 -13220 15005 -13100
rect 15125 -13220 15170 -13100
rect 15290 -13220 15335 -13100
rect 15455 -13220 15500 -13100
rect 15620 -13220 15675 -13100
rect 15795 -13220 15840 -13100
rect 15960 -13220 16005 -13100
rect 16125 -13220 16170 -13100
rect 16290 -13220 16345 -13100
rect 16465 -13220 16510 -13100
rect 16630 -13220 16675 -13100
rect 16795 -13220 16840 -13100
rect 16960 -13220 17015 -13100
rect 17135 -13220 17180 -13100
rect 17300 -13220 17345 -13100
rect 17465 -13220 17510 -13100
rect 17630 -13220 17685 -13100
rect 17805 -13220 17850 -13100
rect 17970 -13220 18015 -13100
rect 18135 -13220 18180 -13100
rect 18300 -13220 18310 -13100
rect 12810 -13265 18310 -13220
rect 12810 -13385 12820 -13265
rect 12940 -13385 12995 -13265
rect 13115 -13385 13160 -13265
rect 13280 -13385 13325 -13265
rect 13445 -13385 13490 -13265
rect 13610 -13385 13665 -13265
rect 13785 -13385 13830 -13265
rect 13950 -13385 13995 -13265
rect 14115 -13385 14160 -13265
rect 14280 -13385 14335 -13265
rect 14455 -13385 14500 -13265
rect 14620 -13385 14665 -13265
rect 14785 -13385 14830 -13265
rect 14950 -13385 15005 -13265
rect 15125 -13385 15170 -13265
rect 15290 -13385 15335 -13265
rect 15455 -13385 15500 -13265
rect 15620 -13385 15675 -13265
rect 15795 -13385 15840 -13265
rect 15960 -13385 16005 -13265
rect 16125 -13385 16170 -13265
rect 16290 -13385 16345 -13265
rect 16465 -13385 16510 -13265
rect 16630 -13385 16675 -13265
rect 16795 -13385 16840 -13265
rect 16960 -13385 17015 -13265
rect 17135 -13385 17180 -13265
rect 17300 -13385 17345 -13265
rect 17465 -13385 17510 -13265
rect 17630 -13385 17685 -13265
rect 17805 -13385 17850 -13265
rect 17970 -13385 18015 -13265
rect 18135 -13385 18180 -13265
rect 18300 -13385 18310 -13265
rect 12810 -13440 18310 -13385
rect 12810 -13560 12820 -13440
rect 12940 -13560 12995 -13440
rect 13115 -13560 13160 -13440
rect 13280 -13560 13325 -13440
rect 13445 -13560 13490 -13440
rect 13610 -13560 13665 -13440
rect 13785 -13560 13830 -13440
rect 13950 -13560 13995 -13440
rect 14115 -13560 14160 -13440
rect 14280 -13560 14335 -13440
rect 14455 -13560 14500 -13440
rect 14620 -13560 14665 -13440
rect 14785 -13560 14830 -13440
rect 14950 -13560 15005 -13440
rect 15125 -13560 15170 -13440
rect 15290 -13560 15335 -13440
rect 15455 -13560 15500 -13440
rect 15620 -13560 15675 -13440
rect 15795 -13560 15840 -13440
rect 15960 -13560 16005 -13440
rect 16125 -13560 16170 -13440
rect 16290 -13560 16345 -13440
rect 16465 -13560 16510 -13440
rect 16630 -13560 16675 -13440
rect 16795 -13560 16840 -13440
rect 16960 -13560 17015 -13440
rect 17135 -13560 17180 -13440
rect 17300 -13560 17345 -13440
rect 17465 -13560 17510 -13440
rect 17630 -13560 17685 -13440
rect 17805 -13560 17850 -13440
rect 17970 -13560 18015 -13440
rect 18135 -13560 18180 -13440
rect 18300 -13560 18310 -13440
rect 12810 -13605 18310 -13560
rect 12810 -13725 12820 -13605
rect 12940 -13725 12995 -13605
rect 13115 -13725 13160 -13605
rect 13280 -13725 13325 -13605
rect 13445 -13725 13490 -13605
rect 13610 -13725 13665 -13605
rect 13785 -13725 13830 -13605
rect 13950 -13725 13995 -13605
rect 14115 -13725 14160 -13605
rect 14280 -13725 14335 -13605
rect 14455 -13725 14500 -13605
rect 14620 -13725 14665 -13605
rect 14785 -13725 14830 -13605
rect 14950 -13725 15005 -13605
rect 15125 -13725 15170 -13605
rect 15290 -13725 15335 -13605
rect 15455 -13725 15500 -13605
rect 15620 -13725 15675 -13605
rect 15795 -13725 15840 -13605
rect 15960 -13725 16005 -13605
rect 16125 -13725 16170 -13605
rect 16290 -13725 16345 -13605
rect 16465 -13725 16510 -13605
rect 16630 -13725 16675 -13605
rect 16795 -13725 16840 -13605
rect 16960 -13725 17015 -13605
rect 17135 -13725 17180 -13605
rect 17300 -13725 17345 -13605
rect 17465 -13725 17510 -13605
rect 17630 -13725 17685 -13605
rect 17805 -13725 17850 -13605
rect 17970 -13725 18015 -13605
rect 18135 -13725 18180 -13605
rect 18300 -13725 18310 -13605
rect 12810 -13770 18310 -13725
rect 12810 -13890 12820 -13770
rect 12940 -13890 12995 -13770
rect 13115 -13890 13160 -13770
rect 13280 -13890 13325 -13770
rect 13445 -13890 13490 -13770
rect 13610 -13890 13665 -13770
rect 13785 -13890 13830 -13770
rect 13950 -13890 13995 -13770
rect 14115 -13890 14160 -13770
rect 14280 -13890 14335 -13770
rect 14455 -13890 14500 -13770
rect 14620 -13890 14665 -13770
rect 14785 -13890 14830 -13770
rect 14950 -13890 15005 -13770
rect 15125 -13890 15170 -13770
rect 15290 -13890 15335 -13770
rect 15455 -13890 15500 -13770
rect 15620 -13890 15675 -13770
rect 15795 -13890 15840 -13770
rect 15960 -13890 16005 -13770
rect 16125 -13890 16170 -13770
rect 16290 -13890 16345 -13770
rect 16465 -13890 16510 -13770
rect 16630 -13890 16675 -13770
rect 16795 -13890 16840 -13770
rect 16960 -13890 17015 -13770
rect 17135 -13890 17180 -13770
rect 17300 -13890 17345 -13770
rect 17465 -13890 17510 -13770
rect 17630 -13890 17685 -13770
rect 17805 -13890 17850 -13770
rect 17970 -13890 18015 -13770
rect 18135 -13890 18180 -13770
rect 18300 -13890 18310 -13770
rect 12810 -13935 18310 -13890
rect 12810 -14055 12820 -13935
rect 12940 -14055 12995 -13935
rect 13115 -14055 13160 -13935
rect 13280 -14055 13325 -13935
rect 13445 -14055 13490 -13935
rect 13610 -14055 13665 -13935
rect 13785 -14055 13830 -13935
rect 13950 -14055 13995 -13935
rect 14115 -14055 14160 -13935
rect 14280 -14055 14335 -13935
rect 14455 -14055 14500 -13935
rect 14620 -14055 14665 -13935
rect 14785 -14055 14830 -13935
rect 14950 -14055 15005 -13935
rect 15125 -14055 15170 -13935
rect 15290 -14055 15335 -13935
rect 15455 -14055 15500 -13935
rect 15620 -14055 15675 -13935
rect 15795 -14055 15840 -13935
rect 15960 -14055 16005 -13935
rect 16125 -14055 16170 -13935
rect 16290 -14055 16345 -13935
rect 16465 -14055 16510 -13935
rect 16630 -14055 16675 -13935
rect 16795 -14055 16840 -13935
rect 16960 -14055 17015 -13935
rect 17135 -14055 17180 -13935
rect 17300 -14055 17345 -13935
rect 17465 -14055 17510 -13935
rect 17630 -14055 17685 -13935
rect 17805 -14055 17850 -13935
rect 17970 -14055 18015 -13935
rect 18135 -14055 18180 -13935
rect 18300 -14055 18310 -13935
rect 12810 -14110 18310 -14055
rect 12810 -14230 12820 -14110
rect 12940 -14230 12995 -14110
rect 13115 -14230 13160 -14110
rect 13280 -14230 13325 -14110
rect 13445 -14230 13490 -14110
rect 13610 -14230 13665 -14110
rect 13785 -14230 13830 -14110
rect 13950 -14230 13995 -14110
rect 14115 -14230 14160 -14110
rect 14280 -14230 14335 -14110
rect 14455 -14230 14500 -14110
rect 14620 -14230 14665 -14110
rect 14785 -14230 14830 -14110
rect 14950 -14230 15005 -14110
rect 15125 -14230 15170 -14110
rect 15290 -14230 15335 -14110
rect 15455 -14230 15500 -14110
rect 15620 -14230 15675 -14110
rect 15795 -14230 15840 -14110
rect 15960 -14230 16005 -14110
rect 16125 -14230 16170 -14110
rect 16290 -14230 16345 -14110
rect 16465 -14230 16510 -14110
rect 16630 -14230 16675 -14110
rect 16795 -14230 16840 -14110
rect 16960 -14230 17015 -14110
rect 17135 -14230 17180 -14110
rect 17300 -14230 17345 -14110
rect 17465 -14230 17510 -14110
rect 17630 -14230 17685 -14110
rect 17805 -14230 17850 -14110
rect 17970 -14230 18015 -14110
rect 18135 -14230 18180 -14110
rect 18300 -14230 18310 -14110
rect 12810 -14275 18310 -14230
rect 12810 -14395 12820 -14275
rect 12940 -14395 12995 -14275
rect 13115 -14395 13160 -14275
rect 13280 -14395 13325 -14275
rect 13445 -14395 13490 -14275
rect 13610 -14395 13665 -14275
rect 13785 -14395 13830 -14275
rect 13950 -14395 13995 -14275
rect 14115 -14395 14160 -14275
rect 14280 -14395 14335 -14275
rect 14455 -14395 14500 -14275
rect 14620 -14395 14665 -14275
rect 14785 -14395 14830 -14275
rect 14950 -14395 15005 -14275
rect 15125 -14395 15170 -14275
rect 15290 -14395 15335 -14275
rect 15455 -14395 15500 -14275
rect 15620 -14395 15675 -14275
rect 15795 -14395 15840 -14275
rect 15960 -14395 16005 -14275
rect 16125 -14395 16170 -14275
rect 16290 -14395 16345 -14275
rect 16465 -14395 16510 -14275
rect 16630 -14395 16675 -14275
rect 16795 -14395 16840 -14275
rect 16960 -14395 17015 -14275
rect 17135 -14395 17180 -14275
rect 17300 -14395 17345 -14275
rect 17465 -14395 17510 -14275
rect 17630 -14395 17685 -14275
rect 17805 -14395 17850 -14275
rect 17970 -14395 18015 -14275
rect 18135 -14395 18180 -14275
rect 18300 -14395 18310 -14275
rect 12810 -14440 18310 -14395
rect 12810 -14560 12820 -14440
rect 12940 -14560 12995 -14440
rect 13115 -14560 13160 -14440
rect 13280 -14560 13325 -14440
rect 13445 -14560 13490 -14440
rect 13610 -14560 13665 -14440
rect 13785 -14560 13830 -14440
rect 13950 -14560 13995 -14440
rect 14115 -14560 14160 -14440
rect 14280 -14560 14335 -14440
rect 14455 -14560 14500 -14440
rect 14620 -14560 14665 -14440
rect 14785 -14560 14830 -14440
rect 14950 -14560 15005 -14440
rect 15125 -14560 15170 -14440
rect 15290 -14560 15335 -14440
rect 15455 -14560 15500 -14440
rect 15620 -14560 15675 -14440
rect 15795 -14560 15840 -14440
rect 15960 -14560 16005 -14440
rect 16125 -14560 16170 -14440
rect 16290 -14560 16345 -14440
rect 16465 -14560 16510 -14440
rect 16630 -14560 16675 -14440
rect 16795 -14560 16840 -14440
rect 16960 -14560 17015 -14440
rect 17135 -14560 17180 -14440
rect 17300 -14560 17345 -14440
rect 17465 -14560 17510 -14440
rect 17630 -14560 17685 -14440
rect 17805 -14560 17850 -14440
rect 17970 -14560 18015 -14440
rect 18135 -14560 18180 -14440
rect 18300 -14560 18310 -14440
rect 12810 -14605 18310 -14560
rect 12810 -14725 12820 -14605
rect 12940 -14725 12995 -14605
rect 13115 -14725 13160 -14605
rect 13280 -14725 13325 -14605
rect 13445 -14725 13490 -14605
rect 13610 -14725 13665 -14605
rect 13785 -14725 13830 -14605
rect 13950 -14725 13995 -14605
rect 14115 -14725 14160 -14605
rect 14280 -14725 14335 -14605
rect 14455 -14725 14500 -14605
rect 14620 -14725 14665 -14605
rect 14785 -14725 14830 -14605
rect 14950 -14725 15005 -14605
rect 15125 -14725 15170 -14605
rect 15290 -14725 15335 -14605
rect 15455 -14725 15500 -14605
rect 15620 -14725 15675 -14605
rect 15795 -14725 15840 -14605
rect 15960 -14725 16005 -14605
rect 16125 -14725 16170 -14605
rect 16290 -14725 16345 -14605
rect 16465 -14725 16510 -14605
rect 16630 -14725 16675 -14605
rect 16795 -14725 16840 -14605
rect 16960 -14725 17015 -14605
rect 17135 -14725 17180 -14605
rect 17300 -14725 17345 -14605
rect 17465 -14725 17510 -14605
rect 17630 -14725 17685 -14605
rect 17805 -14725 17850 -14605
rect 17970 -14725 18015 -14605
rect 18135 -14725 18180 -14605
rect 18300 -14725 18310 -14605
rect 12810 -14780 18310 -14725
rect 12810 -14900 12820 -14780
rect 12940 -14900 12995 -14780
rect 13115 -14900 13160 -14780
rect 13280 -14900 13325 -14780
rect 13445 -14900 13490 -14780
rect 13610 -14900 13665 -14780
rect 13785 -14900 13830 -14780
rect 13950 -14900 13995 -14780
rect 14115 -14900 14160 -14780
rect 14280 -14900 14335 -14780
rect 14455 -14900 14500 -14780
rect 14620 -14900 14665 -14780
rect 14785 -14900 14830 -14780
rect 14950 -14900 15005 -14780
rect 15125 -14900 15170 -14780
rect 15290 -14900 15335 -14780
rect 15455 -14900 15500 -14780
rect 15620 -14900 15675 -14780
rect 15795 -14900 15840 -14780
rect 15960 -14900 16005 -14780
rect 16125 -14900 16170 -14780
rect 16290 -14900 16345 -14780
rect 16465 -14900 16510 -14780
rect 16630 -14900 16675 -14780
rect 16795 -14900 16840 -14780
rect 16960 -14900 17015 -14780
rect 17135 -14900 17180 -14780
rect 17300 -14900 17345 -14780
rect 17465 -14900 17510 -14780
rect 17630 -14900 17685 -14780
rect 17805 -14900 17850 -14780
rect 17970 -14900 18015 -14780
rect 18135 -14900 18180 -14780
rect 18300 -14900 18310 -14780
rect 12810 -14945 18310 -14900
rect 12810 -15065 12820 -14945
rect 12940 -15065 12995 -14945
rect 13115 -15065 13160 -14945
rect 13280 -15065 13325 -14945
rect 13445 -15065 13490 -14945
rect 13610 -15065 13665 -14945
rect 13785 -15065 13830 -14945
rect 13950 -15065 13995 -14945
rect 14115 -15065 14160 -14945
rect 14280 -15065 14335 -14945
rect 14455 -15065 14500 -14945
rect 14620 -15065 14665 -14945
rect 14785 -15065 14830 -14945
rect 14950 -15065 15005 -14945
rect 15125 -15065 15170 -14945
rect 15290 -15065 15335 -14945
rect 15455 -15065 15500 -14945
rect 15620 -15065 15675 -14945
rect 15795 -15065 15840 -14945
rect 15960 -15065 16005 -14945
rect 16125 -15065 16170 -14945
rect 16290 -15065 16345 -14945
rect 16465 -15065 16510 -14945
rect 16630 -15065 16675 -14945
rect 16795 -15065 16840 -14945
rect 16960 -15065 17015 -14945
rect 17135 -15065 17180 -14945
rect 17300 -15065 17345 -14945
rect 17465 -15065 17510 -14945
rect 17630 -15065 17685 -14945
rect 17805 -15065 17850 -14945
rect 17970 -15065 18015 -14945
rect 18135 -15065 18180 -14945
rect 18300 -15065 18310 -14945
rect 12810 -15110 18310 -15065
rect 12810 -15230 12820 -15110
rect 12940 -15230 12995 -15110
rect 13115 -15230 13160 -15110
rect 13280 -15230 13325 -15110
rect 13445 -15230 13490 -15110
rect 13610 -15230 13665 -15110
rect 13785 -15230 13830 -15110
rect 13950 -15230 13995 -15110
rect 14115 -15230 14160 -15110
rect 14280 -15230 14335 -15110
rect 14455 -15230 14500 -15110
rect 14620 -15230 14665 -15110
rect 14785 -15230 14830 -15110
rect 14950 -15230 15005 -15110
rect 15125 -15230 15170 -15110
rect 15290 -15230 15335 -15110
rect 15455 -15230 15500 -15110
rect 15620 -15230 15675 -15110
rect 15795 -15230 15840 -15110
rect 15960 -15230 16005 -15110
rect 16125 -15230 16170 -15110
rect 16290 -15230 16345 -15110
rect 16465 -15230 16510 -15110
rect 16630 -15230 16675 -15110
rect 16795 -15230 16840 -15110
rect 16960 -15230 17015 -15110
rect 17135 -15230 17180 -15110
rect 17300 -15230 17345 -15110
rect 17465 -15230 17510 -15110
rect 17630 -15230 17685 -15110
rect 17805 -15230 17850 -15110
rect 17970 -15230 18015 -15110
rect 18135 -15230 18180 -15110
rect 18300 -15230 18310 -15110
rect 12810 -15275 18310 -15230
rect 12810 -15395 12820 -15275
rect 12940 -15395 12995 -15275
rect 13115 -15395 13160 -15275
rect 13280 -15395 13325 -15275
rect 13445 -15395 13490 -15275
rect 13610 -15395 13665 -15275
rect 13785 -15395 13830 -15275
rect 13950 -15395 13995 -15275
rect 14115 -15395 14160 -15275
rect 14280 -15395 14335 -15275
rect 14455 -15395 14500 -15275
rect 14620 -15395 14665 -15275
rect 14785 -15395 14830 -15275
rect 14950 -15395 15005 -15275
rect 15125 -15395 15170 -15275
rect 15290 -15395 15335 -15275
rect 15455 -15395 15500 -15275
rect 15620 -15395 15675 -15275
rect 15795 -15395 15840 -15275
rect 15960 -15395 16005 -15275
rect 16125 -15395 16170 -15275
rect 16290 -15395 16345 -15275
rect 16465 -15395 16510 -15275
rect 16630 -15395 16675 -15275
rect 16795 -15395 16840 -15275
rect 16960 -15395 17015 -15275
rect 17135 -15395 17180 -15275
rect 17300 -15395 17345 -15275
rect 17465 -15395 17510 -15275
rect 17630 -15395 17685 -15275
rect 17805 -15395 17850 -15275
rect 17970 -15395 18015 -15275
rect 18135 -15395 18180 -15275
rect 18300 -15395 18310 -15275
rect 12810 -15450 18310 -15395
rect 12810 -15570 12820 -15450
rect 12940 -15570 12995 -15450
rect 13115 -15570 13160 -15450
rect 13280 -15570 13325 -15450
rect 13445 -15570 13490 -15450
rect 13610 -15570 13665 -15450
rect 13785 -15570 13830 -15450
rect 13950 -15570 13995 -15450
rect 14115 -15570 14160 -15450
rect 14280 -15570 14335 -15450
rect 14455 -15570 14500 -15450
rect 14620 -15570 14665 -15450
rect 14785 -15570 14830 -15450
rect 14950 -15570 15005 -15450
rect 15125 -15570 15170 -15450
rect 15290 -15570 15335 -15450
rect 15455 -15570 15500 -15450
rect 15620 -15570 15675 -15450
rect 15795 -15570 15840 -15450
rect 15960 -15570 16005 -15450
rect 16125 -15570 16170 -15450
rect 16290 -15570 16345 -15450
rect 16465 -15570 16510 -15450
rect 16630 -15570 16675 -15450
rect 16795 -15570 16840 -15450
rect 16960 -15570 17015 -15450
rect 17135 -15570 17180 -15450
rect 17300 -15570 17345 -15450
rect 17465 -15570 17510 -15450
rect 17630 -15570 17685 -15450
rect 17805 -15570 17850 -15450
rect 17970 -15570 18015 -15450
rect 18135 -15570 18180 -15450
rect 18300 -15570 18310 -15450
rect 12810 -15580 18310 -15570
rect 18500 -10090 24000 -10080
rect 18500 -10210 18510 -10090
rect 18630 -10210 18685 -10090
rect 18805 -10210 18850 -10090
rect 18970 -10210 19015 -10090
rect 19135 -10210 19180 -10090
rect 19300 -10210 19355 -10090
rect 19475 -10210 19520 -10090
rect 19640 -10210 19685 -10090
rect 19805 -10210 19850 -10090
rect 19970 -10210 20025 -10090
rect 20145 -10210 20190 -10090
rect 20310 -10210 20355 -10090
rect 20475 -10210 20520 -10090
rect 20640 -10210 20695 -10090
rect 20815 -10210 20860 -10090
rect 20980 -10210 21025 -10090
rect 21145 -10210 21190 -10090
rect 21310 -10210 21365 -10090
rect 21485 -10210 21530 -10090
rect 21650 -10210 21695 -10090
rect 21815 -10210 21860 -10090
rect 21980 -10210 22035 -10090
rect 22155 -10210 22200 -10090
rect 22320 -10210 22365 -10090
rect 22485 -10210 22530 -10090
rect 22650 -10210 22705 -10090
rect 22825 -10210 22870 -10090
rect 22990 -10210 23035 -10090
rect 23155 -10210 23200 -10090
rect 23320 -10210 23375 -10090
rect 23495 -10210 23540 -10090
rect 23660 -10210 23705 -10090
rect 23825 -10210 23870 -10090
rect 23990 -10210 24000 -10090
rect 18500 -10255 24000 -10210
rect 18500 -10375 18510 -10255
rect 18630 -10375 18685 -10255
rect 18805 -10375 18850 -10255
rect 18970 -10375 19015 -10255
rect 19135 -10375 19180 -10255
rect 19300 -10375 19355 -10255
rect 19475 -10375 19520 -10255
rect 19640 -10375 19685 -10255
rect 19805 -10375 19850 -10255
rect 19970 -10375 20025 -10255
rect 20145 -10375 20190 -10255
rect 20310 -10375 20355 -10255
rect 20475 -10375 20520 -10255
rect 20640 -10375 20695 -10255
rect 20815 -10375 20860 -10255
rect 20980 -10375 21025 -10255
rect 21145 -10375 21190 -10255
rect 21310 -10375 21365 -10255
rect 21485 -10375 21530 -10255
rect 21650 -10375 21695 -10255
rect 21815 -10375 21860 -10255
rect 21980 -10375 22035 -10255
rect 22155 -10375 22200 -10255
rect 22320 -10375 22365 -10255
rect 22485 -10375 22530 -10255
rect 22650 -10375 22705 -10255
rect 22825 -10375 22870 -10255
rect 22990 -10375 23035 -10255
rect 23155 -10375 23200 -10255
rect 23320 -10375 23375 -10255
rect 23495 -10375 23540 -10255
rect 23660 -10375 23705 -10255
rect 23825 -10375 23870 -10255
rect 23990 -10375 24000 -10255
rect 18500 -10420 24000 -10375
rect 18500 -10540 18510 -10420
rect 18630 -10540 18685 -10420
rect 18805 -10540 18850 -10420
rect 18970 -10540 19015 -10420
rect 19135 -10540 19180 -10420
rect 19300 -10540 19355 -10420
rect 19475 -10540 19520 -10420
rect 19640 -10540 19685 -10420
rect 19805 -10540 19850 -10420
rect 19970 -10540 20025 -10420
rect 20145 -10540 20190 -10420
rect 20310 -10540 20355 -10420
rect 20475 -10540 20520 -10420
rect 20640 -10540 20695 -10420
rect 20815 -10540 20860 -10420
rect 20980 -10540 21025 -10420
rect 21145 -10540 21190 -10420
rect 21310 -10540 21365 -10420
rect 21485 -10540 21530 -10420
rect 21650 -10540 21695 -10420
rect 21815 -10540 21860 -10420
rect 21980 -10540 22035 -10420
rect 22155 -10540 22200 -10420
rect 22320 -10540 22365 -10420
rect 22485 -10540 22530 -10420
rect 22650 -10540 22705 -10420
rect 22825 -10540 22870 -10420
rect 22990 -10540 23035 -10420
rect 23155 -10540 23200 -10420
rect 23320 -10540 23375 -10420
rect 23495 -10540 23540 -10420
rect 23660 -10540 23705 -10420
rect 23825 -10540 23870 -10420
rect 23990 -10540 24000 -10420
rect 18500 -10585 24000 -10540
rect 18500 -10705 18510 -10585
rect 18630 -10705 18685 -10585
rect 18805 -10705 18850 -10585
rect 18970 -10705 19015 -10585
rect 19135 -10705 19180 -10585
rect 19300 -10705 19355 -10585
rect 19475 -10705 19520 -10585
rect 19640 -10705 19685 -10585
rect 19805 -10705 19850 -10585
rect 19970 -10705 20025 -10585
rect 20145 -10705 20190 -10585
rect 20310 -10705 20355 -10585
rect 20475 -10705 20520 -10585
rect 20640 -10705 20695 -10585
rect 20815 -10705 20860 -10585
rect 20980 -10705 21025 -10585
rect 21145 -10705 21190 -10585
rect 21310 -10705 21365 -10585
rect 21485 -10705 21530 -10585
rect 21650 -10705 21695 -10585
rect 21815 -10705 21860 -10585
rect 21980 -10705 22035 -10585
rect 22155 -10705 22200 -10585
rect 22320 -10705 22365 -10585
rect 22485 -10705 22530 -10585
rect 22650 -10705 22705 -10585
rect 22825 -10705 22870 -10585
rect 22990 -10705 23035 -10585
rect 23155 -10705 23200 -10585
rect 23320 -10705 23375 -10585
rect 23495 -10705 23540 -10585
rect 23660 -10705 23705 -10585
rect 23825 -10705 23870 -10585
rect 23990 -10705 24000 -10585
rect 18500 -10760 24000 -10705
rect 18500 -10880 18510 -10760
rect 18630 -10880 18685 -10760
rect 18805 -10880 18850 -10760
rect 18970 -10880 19015 -10760
rect 19135 -10880 19180 -10760
rect 19300 -10880 19355 -10760
rect 19475 -10880 19520 -10760
rect 19640 -10880 19685 -10760
rect 19805 -10880 19850 -10760
rect 19970 -10880 20025 -10760
rect 20145 -10880 20190 -10760
rect 20310 -10880 20355 -10760
rect 20475 -10880 20520 -10760
rect 20640 -10880 20695 -10760
rect 20815 -10880 20860 -10760
rect 20980 -10880 21025 -10760
rect 21145 -10880 21190 -10760
rect 21310 -10880 21365 -10760
rect 21485 -10880 21530 -10760
rect 21650 -10880 21695 -10760
rect 21815 -10880 21860 -10760
rect 21980 -10880 22035 -10760
rect 22155 -10880 22200 -10760
rect 22320 -10880 22365 -10760
rect 22485 -10880 22530 -10760
rect 22650 -10880 22705 -10760
rect 22825 -10880 22870 -10760
rect 22990 -10880 23035 -10760
rect 23155 -10880 23200 -10760
rect 23320 -10880 23375 -10760
rect 23495 -10880 23540 -10760
rect 23660 -10880 23705 -10760
rect 23825 -10880 23870 -10760
rect 23990 -10880 24000 -10760
rect 18500 -10925 24000 -10880
rect 18500 -11045 18510 -10925
rect 18630 -11045 18685 -10925
rect 18805 -11045 18850 -10925
rect 18970 -11045 19015 -10925
rect 19135 -11045 19180 -10925
rect 19300 -11045 19355 -10925
rect 19475 -11045 19520 -10925
rect 19640 -11045 19685 -10925
rect 19805 -11045 19850 -10925
rect 19970 -11045 20025 -10925
rect 20145 -11045 20190 -10925
rect 20310 -11045 20355 -10925
rect 20475 -11045 20520 -10925
rect 20640 -11045 20695 -10925
rect 20815 -11045 20860 -10925
rect 20980 -11045 21025 -10925
rect 21145 -11045 21190 -10925
rect 21310 -11045 21365 -10925
rect 21485 -11045 21530 -10925
rect 21650 -11045 21695 -10925
rect 21815 -11045 21860 -10925
rect 21980 -11045 22035 -10925
rect 22155 -11045 22200 -10925
rect 22320 -11045 22365 -10925
rect 22485 -11045 22530 -10925
rect 22650 -11045 22705 -10925
rect 22825 -11045 22870 -10925
rect 22990 -11045 23035 -10925
rect 23155 -11045 23200 -10925
rect 23320 -11045 23375 -10925
rect 23495 -11045 23540 -10925
rect 23660 -11045 23705 -10925
rect 23825 -11045 23870 -10925
rect 23990 -11045 24000 -10925
rect 18500 -11090 24000 -11045
rect 18500 -11210 18510 -11090
rect 18630 -11210 18685 -11090
rect 18805 -11210 18850 -11090
rect 18970 -11210 19015 -11090
rect 19135 -11210 19180 -11090
rect 19300 -11210 19355 -11090
rect 19475 -11210 19520 -11090
rect 19640 -11210 19685 -11090
rect 19805 -11210 19850 -11090
rect 19970 -11210 20025 -11090
rect 20145 -11210 20190 -11090
rect 20310 -11210 20355 -11090
rect 20475 -11210 20520 -11090
rect 20640 -11210 20695 -11090
rect 20815 -11210 20860 -11090
rect 20980 -11210 21025 -11090
rect 21145 -11210 21190 -11090
rect 21310 -11210 21365 -11090
rect 21485 -11210 21530 -11090
rect 21650 -11210 21695 -11090
rect 21815 -11210 21860 -11090
rect 21980 -11210 22035 -11090
rect 22155 -11210 22200 -11090
rect 22320 -11210 22365 -11090
rect 22485 -11210 22530 -11090
rect 22650 -11210 22705 -11090
rect 22825 -11210 22870 -11090
rect 22990 -11210 23035 -11090
rect 23155 -11210 23200 -11090
rect 23320 -11210 23375 -11090
rect 23495 -11210 23540 -11090
rect 23660 -11210 23705 -11090
rect 23825 -11210 23870 -11090
rect 23990 -11210 24000 -11090
rect 18500 -11255 24000 -11210
rect 18500 -11375 18510 -11255
rect 18630 -11375 18685 -11255
rect 18805 -11375 18850 -11255
rect 18970 -11375 19015 -11255
rect 19135 -11375 19180 -11255
rect 19300 -11375 19355 -11255
rect 19475 -11375 19520 -11255
rect 19640 -11375 19685 -11255
rect 19805 -11375 19850 -11255
rect 19970 -11375 20025 -11255
rect 20145 -11375 20190 -11255
rect 20310 -11375 20355 -11255
rect 20475 -11375 20520 -11255
rect 20640 -11375 20695 -11255
rect 20815 -11375 20860 -11255
rect 20980 -11375 21025 -11255
rect 21145 -11375 21190 -11255
rect 21310 -11375 21365 -11255
rect 21485 -11375 21530 -11255
rect 21650 -11375 21695 -11255
rect 21815 -11375 21860 -11255
rect 21980 -11375 22035 -11255
rect 22155 -11375 22200 -11255
rect 22320 -11375 22365 -11255
rect 22485 -11375 22530 -11255
rect 22650 -11375 22705 -11255
rect 22825 -11375 22870 -11255
rect 22990 -11375 23035 -11255
rect 23155 -11375 23200 -11255
rect 23320 -11375 23375 -11255
rect 23495 -11375 23540 -11255
rect 23660 -11375 23705 -11255
rect 23825 -11375 23870 -11255
rect 23990 -11375 24000 -11255
rect 18500 -11430 24000 -11375
rect 18500 -11550 18510 -11430
rect 18630 -11550 18685 -11430
rect 18805 -11550 18850 -11430
rect 18970 -11550 19015 -11430
rect 19135 -11550 19180 -11430
rect 19300 -11550 19355 -11430
rect 19475 -11550 19520 -11430
rect 19640 -11550 19685 -11430
rect 19805 -11550 19850 -11430
rect 19970 -11550 20025 -11430
rect 20145 -11550 20190 -11430
rect 20310 -11550 20355 -11430
rect 20475 -11550 20520 -11430
rect 20640 -11550 20695 -11430
rect 20815 -11550 20860 -11430
rect 20980 -11550 21025 -11430
rect 21145 -11550 21190 -11430
rect 21310 -11550 21365 -11430
rect 21485 -11550 21530 -11430
rect 21650 -11550 21695 -11430
rect 21815 -11550 21860 -11430
rect 21980 -11550 22035 -11430
rect 22155 -11550 22200 -11430
rect 22320 -11550 22365 -11430
rect 22485 -11550 22530 -11430
rect 22650 -11550 22705 -11430
rect 22825 -11550 22870 -11430
rect 22990 -11550 23035 -11430
rect 23155 -11550 23200 -11430
rect 23320 -11550 23375 -11430
rect 23495 -11550 23540 -11430
rect 23660 -11550 23705 -11430
rect 23825 -11550 23870 -11430
rect 23990 -11550 24000 -11430
rect 18500 -11595 24000 -11550
rect 18500 -11715 18510 -11595
rect 18630 -11715 18685 -11595
rect 18805 -11715 18850 -11595
rect 18970 -11715 19015 -11595
rect 19135 -11715 19180 -11595
rect 19300 -11715 19355 -11595
rect 19475 -11715 19520 -11595
rect 19640 -11715 19685 -11595
rect 19805 -11715 19850 -11595
rect 19970 -11715 20025 -11595
rect 20145 -11715 20190 -11595
rect 20310 -11715 20355 -11595
rect 20475 -11715 20520 -11595
rect 20640 -11715 20695 -11595
rect 20815 -11715 20860 -11595
rect 20980 -11715 21025 -11595
rect 21145 -11715 21190 -11595
rect 21310 -11715 21365 -11595
rect 21485 -11715 21530 -11595
rect 21650 -11715 21695 -11595
rect 21815 -11715 21860 -11595
rect 21980 -11715 22035 -11595
rect 22155 -11715 22200 -11595
rect 22320 -11715 22365 -11595
rect 22485 -11715 22530 -11595
rect 22650 -11715 22705 -11595
rect 22825 -11715 22870 -11595
rect 22990 -11715 23035 -11595
rect 23155 -11715 23200 -11595
rect 23320 -11715 23375 -11595
rect 23495 -11715 23540 -11595
rect 23660 -11715 23705 -11595
rect 23825 -11715 23870 -11595
rect 23990 -11715 24000 -11595
rect 18500 -11760 24000 -11715
rect 18500 -11880 18510 -11760
rect 18630 -11880 18685 -11760
rect 18805 -11880 18850 -11760
rect 18970 -11880 19015 -11760
rect 19135 -11880 19180 -11760
rect 19300 -11880 19355 -11760
rect 19475 -11880 19520 -11760
rect 19640 -11880 19685 -11760
rect 19805 -11880 19850 -11760
rect 19970 -11880 20025 -11760
rect 20145 -11880 20190 -11760
rect 20310 -11880 20355 -11760
rect 20475 -11880 20520 -11760
rect 20640 -11880 20695 -11760
rect 20815 -11880 20860 -11760
rect 20980 -11880 21025 -11760
rect 21145 -11880 21190 -11760
rect 21310 -11880 21365 -11760
rect 21485 -11880 21530 -11760
rect 21650 -11880 21695 -11760
rect 21815 -11880 21860 -11760
rect 21980 -11880 22035 -11760
rect 22155 -11880 22200 -11760
rect 22320 -11880 22365 -11760
rect 22485 -11880 22530 -11760
rect 22650 -11880 22705 -11760
rect 22825 -11880 22870 -11760
rect 22990 -11880 23035 -11760
rect 23155 -11880 23200 -11760
rect 23320 -11880 23375 -11760
rect 23495 -11880 23540 -11760
rect 23660 -11880 23705 -11760
rect 23825 -11880 23870 -11760
rect 23990 -11880 24000 -11760
rect 18500 -11925 24000 -11880
rect 18500 -12045 18510 -11925
rect 18630 -12045 18685 -11925
rect 18805 -12045 18850 -11925
rect 18970 -12045 19015 -11925
rect 19135 -12045 19180 -11925
rect 19300 -12045 19355 -11925
rect 19475 -12045 19520 -11925
rect 19640 -12045 19685 -11925
rect 19805 -12045 19850 -11925
rect 19970 -12045 20025 -11925
rect 20145 -12045 20190 -11925
rect 20310 -12045 20355 -11925
rect 20475 -12045 20520 -11925
rect 20640 -12045 20695 -11925
rect 20815 -12045 20860 -11925
rect 20980 -12045 21025 -11925
rect 21145 -12045 21190 -11925
rect 21310 -12045 21365 -11925
rect 21485 -12045 21530 -11925
rect 21650 -12045 21695 -11925
rect 21815 -12045 21860 -11925
rect 21980 -12045 22035 -11925
rect 22155 -12045 22200 -11925
rect 22320 -12045 22365 -11925
rect 22485 -12045 22530 -11925
rect 22650 -12045 22705 -11925
rect 22825 -12045 22870 -11925
rect 22990 -12045 23035 -11925
rect 23155 -12045 23200 -11925
rect 23320 -12045 23375 -11925
rect 23495 -12045 23540 -11925
rect 23660 -12045 23705 -11925
rect 23825 -12045 23870 -11925
rect 23990 -12045 24000 -11925
rect 18500 -12100 24000 -12045
rect 18500 -12220 18510 -12100
rect 18630 -12220 18685 -12100
rect 18805 -12220 18850 -12100
rect 18970 -12220 19015 -12100
rect 19135 -12220 19180 -12100
rect 19300 -12220 19355 -12100
rect 19475 -12220 19520 -12100
rect 19640 -12220 19685 -12100
rect 19805 -12220 19850 -12100
rect 19970 -12220 20025 -12100
rect 20145 -12220 20190 -12100
rect 20310 -12220 20355 -12100
rect 20475 -12220 20520 -12100
rect 20640 -12220 20695 -12100
rect 20815 -12220 20860 -12100
rect 20980 -12220 21025 -12100
rect 21145 -12220 21190 -12100
rect 21310 -12220 21365 -12100
rect 21485 -12220 21530 -12100
rect 21650 -12220 21695 -12100
rect 21815 -12220 21860 -12100
rect 21980 -12220 22035 -12100
rect 22155 -12220 22200 -12100
rect 22320 -12220 22365 -12100
rect 22485 -12220 22530 -12100
rect 22650 -12220 22705 -12100
rect 22825 -12220 22870 -12100
rect 22990 -12220 23035 -12100
rect 23155 -12220 23200 -12100
rect 23320 -12220 23375 -12100
rect 23495 -12220 23540 -12100
rect 23660 -12220 23705 -12100
rect 23825 -12220 23870 -12100
rect 23990 -12220 24000 -12100
rect 18500 -12265 24000 -12220
rect 18500 -12385 18510 -12265
rect 18630 -12385 18685 -12265
rect 18805 -12385 18850 -12265
rect 18970 -12385 19015 -12265
rect 19135 -12385 19180 -12265
rect 19300 -12385 19355 -12265
rect 19475 -12385 19520 -12265
rect 19640 -12385 19685 -12265
rect 19805 -12385 19850 -12265
rect 19970 -12385 20025 -12265
rect 20145 -12385 20190 -12265
rect 20310 -12385 20355 -12265
rect 20475 -12385 20520 -12265
rect 20640 -12385 20695 -12265
rect 20815 -12385 20860 -12265
rect 20980 -12385 21025 -12265
rect 21145 -12385 21190 -12265
rect 21310 -12385 21365 -12265
rect 21485 -12385 21530 -12265
rect 21650 -12385 21695 -12265
rect 21815 -12385 21860 -12265
rect 21980 -12385 22035 -12265
rect 22155 -12385 22200 -12265
rect 22320 -12385 22365 -12265
rect 22485 -12385 22530 -12265
rect 22650 -12385 22705 -12265
rect 22825 -12385 22870 -12265
rect 22990 -12385 23035 -12265
rect 23155 -12385 23200 -12265
rect 23320 -12385 23375 -12265
rect 23495 -12385 23540 -12265
rect 23660 -12385 23705 -12265
rect 23825 -12385 23870 -12265
rect 23990 -12385 24000 -12265
rect 18500 -12430 24000 -12385
rect 18500 -12550 18510 -12430
rect 18630 -12550 18685 -12430
rect 18805 -12550 18850 -12430
rect 18970 -12550 19015 -12430
rect 19135 -12550 19180 -12430
rect 19300 -12550 19355 -12430
rect 19475 -12550 19520 -12430
rect 19640 -12550 19685 -12430
rect 19805 -12550 19850 -12430
rect 19970 -12550 20025 -12430
rect 20145 -12550 20190 -12430
rect 20310 -12550 20355 -12430
rect 20475 -12550 20520 -12430
rect 20640 -12550 20695 -12430
rect 20815 -12550 20860 -12430
rect 20980 -12550 21025 -12430
rect 21145 -12550 21190 -12430
rect 21310 -12550 21365 -12430
rect 21485 -12550 21530 -12430
rect 21650 -12550 21695 -12430
rect 21815 -12550 21860 -12430
rect 21980 -12550 22035 -12430
rect 22155 -12550 22200 -12430
rect 22320 -12550 22365 -12430
rect 22485 -12550 22530 -12430
rect 22650 -12550 22705 -12430
rect 22825 -12550 22870 -12430
rect 22990 -12550 23035 -12430
rect 23155 -12550 23200 -12430
rect 23320 -12550 23375 -12430
rect 23495 -12550 23540 -12430
rect 23660 -12550 23705 -12430
rect 23825 -12550 23870 -12430
rect 23990 -12550 24000 -12430
rect 18500 -12595 24000 -12550
rect 18500 -12715 18510 -12595
rect 18630 -12715 18685 -12595
rect 18805 -12715 18850 -12595
rect 18970 -12715 19015 -12595
rect 19135 -12715 19180 -12595
rect 19300 -12715 19355 -12595
rect 19475 -12715 19520 -12595
rect 19640 -12715 19685 -12595
rect 19805 -12715 19850 -12595
rect 19970 -12715 20025 -12595
rect 20145 -12715 20190 -12595
rect 20310 -12715 20355 -12595
rect 20475 -12715 20520 -12595
rect 20640 -12715 20695 -12595
rect 20815 -12715 20860 -12595
rect 20980 -12715 21025 -12595
rect 21145 -12715 21190 -12595
rect 21310 -12715 21365 -12595
rect 21485 -12715 21530 -12595
rect 21650 -12715 21695 -12595
rect 21815 -12715 21860 -12595
rect 21980 -12715 22035 -12595
rect 22155 -12715 22200 -12595
rect 22320 -12715 22365 -12595
rect 22485 -12715 22530 -12595
rect 22650 -12715 22705 -12595
rect 22825 -12715 22870 -12595
rect 22990 -12715 23035 -12595
rect 23155 -12715 23200 -12595
rect 23320 -12715 23375 -12595
rect 23495 -12715 23540 -12595
rect 23660 -12715 23705 -12595
rect 23825 -12715 23870 -12595
rect 23990 -12715 24000 -12595
rect 18500 -12770 24000 -12715
rect 18500 -12890 18510 -12770
rect 18630 -12890 18685 -12770
rect 18805 -12890 18850 -12770
rect 18970 -12890 19015 -12770
rect 19135 -12890 19180 -12770
rect 19300 -12890 19355 -12770
rect 19475 -12890 19520 -12770
rect 19640 -12890 19685 -12770
rect 19805 -12890 19850 -12770
rect 19970 -12890 20025 -12770
rect 20145 -12890 20190 -12770
rect 20310 -12890 20355 -12770
rect 20475 -12890 20520 -12770
rect 20640 -12890 20695 -12770
rect 20815 -12890 20860 -12770
rect 20980 -12890 21025 -12770
rect 21145 -12890 21190 -12770
rect 21310 -12890 21365 -12770
rect 21485 -12890 21530 -12770
rect 21650 -12890 21695 -12770
rect 21815 -12890 21860 -12770
rect 21980 -12890 22035 -12770
rect 22155 -12890 22200 -12770
rect 22320 -12890 22365 -12770
rect 22485 -12890 22530 -12770
rect 22650 -12890 22705 -12770
rect 22825 -12890 22870 -12770
rect 22990 -12890 23035 -12770
rect 23155 -12890 23200 -12770
rect 23320 -12890 23375 -12770
rect 23495 -12890 23540 -12770
rect 23660 -12890 23705 -12770
rect 23825 -12890 23870 -12770
rect 23990 -12890 24000 -12770
rect 18500 -12935 24000 -12890
rect 18500 -13055 18510 -12935
rect 18630 -13055 18685 -12935
rect 18805 -13055 18850 -12935
rect 18970 -13055 19015 -12935
rect 19135 -13055 19180 -12935
rect 19300 -13055 19355 -12935
rect 19475 -13055 19520 -12935
rect 19640 -13055 19685 -12935
rect 19805 -13055 19850 -12935
rect 19970 -13055 20025 -12935
rect 20145 -13055 20190 -12935
rect 20310 -13055 20355 -12935
rect 20475 -13055 20520 -12935
rect 20640 -13055 20695 -12935
rect 20815 -13055 20860 -12935
rect 20980 -13055 21025 -12935
rect 21145 -13055 21190 -12935
rect 21310 -13055 21365 -12935
rect 21485 -13055 21530 -12935
rect 21650 -13055 21695 -12935
rect 21815 -13055 21860 -12935
rect 21980 -13055 22035 -12935
rect 22155 -13055 22200 -12935
rect 22320 -13055 22365 -12935
rect 22485 -13055 22530 -12935
rect 22650 -13055 22705 -12935
rect 22825 -13055 22870 -12935
rect 22990 -13055 23035 -12935
rect 23155 -13055 23200 -12935
rect 23320 -13055 23375 -12935
rect 23495 -13055 23540 -12935
rect 23660 -13055 23705 -12935
rect 23825 -13055 23870 -12935
rect 23990 -13055 24000 -12935
rect 18500 -13100 24000 -13055
rect 18500 -13220 18510 -13100
rect 18630 -13220 18685 -13100
rect 18805 -13220 18850 -13100
rect 18970 -13220 19015 -13100
rect 19135 -13220 19180 -13100
rect 19300 -13220 19355 -13100
rect 19475 -13220 19520 -13100
rect 19640 -13220 19685 -13100
rect 19805 -13220 19850 -13100
rect 19970 -13220 20025 -13100
rect 20145 -13220 20190 -13100
rect 20310 -13220 20355 -13100
rect 20475 -13220 20520 -13100
rect 20640 -13220 20695 -13100
rect 20815 -13220 20860 -13100
rect 20980 -13220 21025 -13100
rect 21145 -13220 21190 -13100
rect 21310 -13220 21365 -13100
rect 21485 -13220 21530 -13100
rect 21650 -13220 21695 -13100
rect 21815 -13220 21860 -13100
rect 21980 -13220 22035 -13100
rect 22155 -13220 22200 -13100
rect 22320 -13220 22365 -13100
rect 22485 -13220 22530 -13100
rect 22650 -13220 22705 -13100
rect 22825 -13220 22870 -13100
rect 22990 -13220 23035 -13100
rect 23155 -13220 23200 -13100
rect 23320 -13220 23375 -13100
rect 23495 -13220 23540 -13100
rect 23660 -13220 23705 -13100
rect 23825 -13220 23870 -13100
rect 23990 -13220 24000 -13100
rect 18500 -13265 24000 -13220
rect 18500 -13385 18510 -13265
rect 18630 -13385 18685 -13265
rect 18805 -13385 18850 -13265
rect 18970 -13385 19015 -13265
rect 19135 -13385 19180 -13265
rect 19300 -13385 19355 -13265
rect 19475 -13385 19520 -13265
rect 19640 -13385 19685 -13265
rect 19805 -13385 19850 -13265
rect 19970 -13385 20025 -13265
rect 20145 -13385 20190 -13265
rect 20310 -13385 20355 -13265
rect 20475 -13385 20520 -13265
rect 20640 -13385 20695 -13265
rect 20815 -13385 20860 -13265
rect 20980 -13385 21025 -13265
rect 21145 -13385 21190 -13265
rect 21310 -13385 21365 -13265
rect 21485 -13385 21530 -13265
rect 21650 -13385 21695 -13265
rect 21815 -13385 21860 -13265
rect 21980 -13385 22035 -13265
rect 22155 -13385 22200 -13265
rect 22320 -13385 22365 -13265
rect 22485 -13385 22530 -13265
rect 22650 -13385 22705 -13265
rect 22825 -13385 22870 -13265
rect 22990 -13385 23035 -13265
rect 23155 -13385 23200 -13265
rect 23320 -13385 23375 -13265
rect 23495 -13385 23540 -13265
rect 23660 -13385 23705 -13265
rect 23825 -13385 23870 -13265
rect 23990 -13385 24000 -13265
rect 18500 -13440 24000 -13385
rect 18500 -13560 18510 -13440
rect 18630 -13560 18685 -13440
rect 18805 -13560 18850 -13440
rect 18970 -13560 19015 -13440
rect 19135 -13560 19180 -13440
rect 19300 -13560 19355 -13440
rect 19475 -13560 19520 -13440
rect 19640 -13560 19685 -13440
rect 19805 -13560 19850 -13440
rect 19970 -13560 20025 -13440
rect 20145 -13560 20190 -13440
rect 20310 -13560 20355 -13440
rect 20475 -13560 20520 -13440
rect 20640 -13560 20695 -13440
rect 20815 -13560 20860 -13440
rect 20980 -13560 21025 -13440
rect 21145 -13560 21190 -13440
rect 21310 -13560 21365 -13440
rect 21485 -13560 21530 -13440
rect 21650 -13560 21695 -13440
rect 21815 -13560 21860 -13440
rect 21980 -13560 22035 -13440
rect 22155 -13560 22200 -13440
rect 22320 -13560 22365 -13440
rect 22485 -13560 22530 -13440
rect 22650 -13560 22705 -13440
rect 22825 -13560 22870 -13440
rect 22990 -13560 23035 -13440
rect 23155 -13560 23200 -13440
rect 23320 -13560 23375 -13440
rect 23495 -13560 23540 -13440
rect 23660 -13560 23705 -13440
rect 23825 -13560 23870 -13440
rect 23990 -13560 24000 -13440
rect 18500 -13605 24000 -13560
rect 18500 -13725 18510 -13605
rect 18630 -13725 18685 -13605
rect 18805 -13725 18850 -13605
rect 18970 -13725 19015 -13605
rect 19135 -13725 19180 -13605
rect 19300 -13725 19355 -13605
rect 19475 -13725 19520 -13605
rect 19640 -13725 19685 -13605
rect 19805 -13725 19850 -13605
rect 19970 -13725 20025 -13605
rect 20145 -13725 20190 -13605
rect 20310 -13725 20355 -13605
rect 20475 -13725 20520 -13605
rect 20640 -13725 20695 -13605
rect 20815 -13725 20860 -13605
rect 20980 -13725 21025 -13605
rect 21145 -13725 21190 -13605
rect 21310 -13725 21365 -13605
rect 21485 -13725 21530 -13605
rect 21650 -13725 21695 -13605
rect 21815 -13725 21860 -13605
rect 21980 -13725 22035 -13605
rect 22155 -13725 22200 -13605
rect 22320 -13725 22365 -13605
rect 22485 -13725 22530 -13605
rect 22650 -13725 22705 -13605
rect 22825 -13725 22870 -13605
rect 22990 -13725 23035 -13605
rect 23155 -13725 23200 -13605
rect 23320 -13725 23375 -13605
rect 23495 -13725 23540 -13605
rect 23660 -13725 23705 -13605
rect 23825 -13725 23870 -13605
rect 23990 -13725 24000 -13605
rect 18500 -13770 24000 -13725
rect 18500 -13890 18510 -13770
rect 18630 -13890 18685 -13770
rect 18805 -13890 18850 -13770
rect 18970 -13890 19015 -13770
rect 19135 -13890 19180 -13770
rect 19300 -13890 19355 -13770
rect 19475 -13890 19520 -13770
rect 19640 -13890 19685 -13770
rect 19805 -13890 19850 -13770
rect 19970 -13890 20025 -13770
rect 20145 -13890 20190 -13770
rect 20310 -13890 20355 -13770
rect 20475 -13890 20520 -13770
rect 20640 -13890 20695 -13770
rect 20815 -13890 20860 -13770
rect 20980 -13890 21025 -13770
rect 21145 -13890 21190 -13770
rect 21310 -13890 21365 -13770
rect 21485 -13890 21530 -13770
rect 21650 -13890 21695 -13770
rect 21815 -13890 21860 -13770
rect 21980 -13890 22035 -13770
rect 22155 -13890 22200 -13770
rect 22320 -13890 22365 -13770
rect 22485 -13890 22530 -13770
rect 22650 -13890 22705 -13770
rect 22825 -13890 22870 -13770
rect 22990 -13890 23035 -13770
rect 23155 -13890 23200 -13770
rect 23320 -13890 23375 -13770
rect 23495 -13890 23540 -13770
rect 23660 -13890 23705 -13770
rect 23825 -13890 23870 -13770
rect 23990 -13890 24000 -13770
rect 18500 -13935 24000 -13890
rect 18500 -14055 18510 -13935
rect 18630 -14055 18685 -13935
rect 18805 -14055 18850 -13935
rect 18970 -14055 19015 -13935
rect 19135 -14055 19180 -13935
rect 19300 -14055 19355 -13935
rect 19475 -14055 19520 -13935
rect 19640 -14055 19685 -13935
rect 19805 -14055 19850 -13935
rect 19970 -14055 20025 -13935
rect 20145 -14055 20190 -13935
rect 20310 -14055 20355 -13935
rect 20475 -14055 20520 -13935
rect 20640 -14055 20695 -13935
rect 20815 -14055 20860 -13935
rect 20980 -14055 21025 -13935
rect 21145 -14055 21190 -13935
rect 21310 -14055 21365 -13935
rect 21485 -14055 21530 -13935
rect 21650 -14055 21695 -13935
rect 21815 -14055 21860 -13935
rect 21980 -14055 22035 -13935
rect 22155 -14055 22200 -13935
rect 22320 -14055 22365 -13935
rect 22485 -14055 22530 -13935
rect 22650 -14055 22705 -13935
rect 22825 -14055 22870 -13935
rect 22990 -14055 23035 -13935
rect 23155 -14055 23200 -13935
rect 23320 -14055 23375 -13935
rect 23495 -14055 23540 -13935
rect 23660 -14055 23705 -13935
rect 23825 -14055 23870 -13935
rect 23990 -14055 24000 -13935
rect 18500 -14110 24000 -14055
rect 18500 -14230 18510 -14110
rect 18630 -14230 18685 -14110
rect 18805 -14230 18850 -14110
rect 18970 -14230 19015 -14110
rect 19135 -14230 19180 -14110
rect 19300 -14230 19355 -14110
rect 19475 -14230 19520 -14110
rect 19640 -14230 19685 -14110
rect 19805 -14230 19850 -14110
rect 19970 -14230 20025 -14110
rect 20145 -14230 20190 -14110
rect 20310 -14230 20355 -14110
rect 20475 -14230 20520 -14110
rect 20640 -14230 20695 -14110
rect 20815 -14230 20860 -14110
rect 20980 -14230 21025 -14110
rect 21145 -14230 21190 -14110
rect 21310 -14230 21365 -14110
rect 21485 -14230 21530 -14110
rect 21650 -14230 21695 -14110
rect 21815 -14230 21860 -14110
rect 21980 -14230 22035 -14110
rect 22155 -14230 22200 -14110
rect 22320 -14230 22365 -14110
rect 22485 -14230 22530 -14110
rect 22650 -14230 22705 -14110
rect 22825 -14230 22870 -14110
rect 22990 -14230 23035 -14110
rect 23155 -14230 23200 -14110
rect 23320 -14230 23375 -14110
rect 23495 -14230 23540 -14110
rect 23660 -14230 23705 -14110
rect 23825 -14230 23870 -14110
rect 23990 -14230 24000 -14110
rect 18500 -14275 24000 -14230
rect 18500 -14395 18510 -14275
rect 18630 -14395 18685 -14275
rect 18805 -14395 18850 -14275
rect 18970 -14395 19015 -14275
rect 19135 -14395 19180 -14275
rect 19300 -14395 19355 -14275
rect 19475 -14395 19520 -14275
rect 19640 -14395 19685 -14275
rect 19805 -14395 19850 -14275
rect 19970 -14395 20025 -14275
rect 20145 -14395 20190 -14275
rect 20310 -14395 20355 -14275
rect 20475 -14395 20520 -14275
rect 20640 -14395 20695 -14275
rect 20815 -14395 20860 -14275
rect 20980 -14395 21025 -14275
rect 21145 -14395 21190 -14275
rect 21310 -14395 21365 -14275
rect 21485 -14395 21530 -14275
rect 21650 -14395 21695 -14275
rect 21815 -14395 21860 -14275
rect 21980 -14395 22035 -14275
rect 22155 -14395 22200 -14275
rect 22320 -14395 22365 -14275
rect 22485 -14395 22530 -14275
rect 22650 -14395 22705 -14275
rect 22825 -14395 22870 -14275
rect 22990 -14395 23035 -14275
rect 23155 -14395 23200 -14275
rect 23320 -14395 23375 -14275
rect 23495 -14395 23540 -14275
rect 23660 -14395 23705 -14275
rect 23825 -14395 23870 -14275
rect 23990 -14395 24000 -14275
rect 18500 -14440 24000 -14395
rect 18500 -14560 18510 -14440
rect 18630 -14560 18685 -14440
rect 18805 -14560 18850 -14440
rect 18970 -14560 19015 -14440
rect 19135 -14560 19180 -14440
rect 19300 -14560 19355 -14440
rect 19475 -14560 19520 -14440
rect 19640 -14560 19685 -14440
rect 19805 -14560 19850 -14440
rect 19970 -14560 20025 -14440
rect 20145 -14560 20190 -14440
rect 20310 -14560 20355 -14440
rect 20475 -14560 20520 -14440
rect 20640 -14560 20695 -14440
rect 20815 -14560 20860 -14440
rect 20980 -14560 21025 -14440
rect 21145 -14560 21190 -14440
rect 21310 -14560 21365 -14440
rect 21485 -14560 21530 -14440
rect 21650 -14560 21695 -14440
rect 21815 -14560 21860 -14440
rect 21980 -14560 22035 -14440
rect 22155 -14560 22200 -14440
rect 22320 -14560 22365 -14440
rect 22485 -14560 22530 -14440
rect 22650 -14560 22705 -14440
rect 22825 -14560 22870 -14440
rect 22990 -14560 23035 -14440
rect 23155 -14560 23200 -14440
rect 23320 -14560 23375 -14440
rect 23495 -14560 23540 -14440
rect 23660 -14560 23705 -14440
rect 23825 -14560 23870 -14440
rect 23990 -14560 24000 -14440
rect 18500 -14605 24000 -14560
rect 18500 -14725 18510 -14605
rect 18630 -14725 18685 -14605
rect 18805 -14725 18850 -14605
rect 18970 -14725 19015 -14605
rect 19135 -14725 19180 -14605
rect 19300 -14725 19355 -14605
rect 19475 -14725 19520 -14605
rect 19640 -14725 19685 -14605
rect 19805 -14725 19850 -14605
rect 19970 -14725 20025 -14605
rect 20145 -14725 20190 -14605
rect 20310 -14725 20355 -14605
rect 20475 -14725 20520 -14605
rect 20640 -14725 20695 -14605
rect 20815 -14725 20860 -14605
rect 20980 -14725 21025 -14605
rect 21145 -14725 21190 -14605
rect 21310 -14725 21365 -14605
rect 21485 -14725 21530 -14605
rect 21650 -14725 21695 -14605
rect 21815 -14725 21860 -14605
rect 21980 -14725 22035 -14605
rect 22155 -14725 22200 -14605
rect 22320 -14725 22365 -14605
rect 22485 -14725 22530 -14605
rect 22650 -14725 22705 -14605
rect 22825 -14725 22870 -14605
rect 22990 -14725 23035 -14605
rect 23155 -14725 23200 -14605
rect 23320 -14725 23375 -14605
rect 23495 -14725 23540 -14605
rect 23660 -14725 23705 -14605
rect 23825 -14725 23870 -14605
rect 23990 -14725 24000 -14605
rect 18500 -14780 24000 -14725
rect 18500 -14900 18510 -14780
rect 18630 -14900 18685 -14780
rect 18805 -14900 18850 -14780
rect 18970 -14900 19015 -14780
rect 19135 -14900 19180 -14780
rect 19300 -14900 19355 -14780
rect 19475 -14900 19520 -14780
rect 19640 -14900 19685 -14780
rect 19805 -14900 19850 -14780
rect 19970 -14900 20025 -14780
rect 20145 -14900 20190 -14780
rect 20310 -14900 20355 -14780
rect 20475 -14900 20520 -14780
rect 20640 -14900 20695 -14780
rect 20815 -14900 20860 -14780
rect 20980 -14900 21025 -14780
rect 21145 -14900 21190 -14780
rect 21310 -14900 21365 -14780
rect 21485 -14900 21530 -14780
rect 21650 -14900 21695 -14780
rect 21815 -14900 21860 -14780
rect 21980 -14900 22035 -14780
rect 22155 -14900 22200 -14780
rect 22320 -14900 22365 -14780
rect 22485 -14900 22530 -14780
rect 22650 -14900 22705 -14780
rect 22825 -14900 22870 -14780
rect 22990 -14900 23035 -14780
rect 23155 -14900 23200 -14780
rect 23320 -14900 23375 -14780
rect 23495 -14900 23540 -14780
rect 23660 -14900 23705 -14780
rect 23825 -14900 23870 -14780
rect 23990 -14900 24000 -14780
rect 18500 -14945 24000 -14900
rect 18500 -15065 18510 -14945
rect 18630 -15065 18685 -14945
rect 18805 -15065 18850 -14945
rect 18970 -15065 19015 -14945
rect 19135 -15065 19180 -14945
rect 19300 -15065 19355 -14945
rect 19475 -15065 19520 -14945
rect 19640 -15065 19685 -14945
rect 19805 -15065 19850 -14945
rect 19970 -15065 20025 -14945
rect 20145 -15065 20190 -14945
rect 20310 -15065 20355 -14945
rect 20475 -15065 20520 -14945
rect 20640 -15065 20695 -14945
rect 20815 -15065 20860 -14945
rect 20980 -15065 21025 -14945
rect 21145 -15065 21190 -14945
rect 21310 -15065 21365 -14945
rect 21485 -15065 21530 -14945
rect 21650 -15065 21695 -14945
rect 21815 -15065 21860 -14945
rect 21980 -15065 22035 -14945
rect 22155 -15065 22200 -14945
rect 22320 -15065 22365 -14945
rect 22485 -15065 22530 -14945
rect 22650 -15065 22705 -14945
rect 22825 -15065 22870 -14945
rect 22990 -15065 23035 -14945
rect 23155 -15065 23200 -14945
rect 23320 -15065 23375 -14945
rect 23495 -15065 23540 -14945
rect 23660 -15065 23705 -14945
rect 23825 -15065 23870 -14945
rect 23990 -15065 24000 -14945
rect 18500 -15110 24000 -15065
rect 18500 -15230 18510 -15110
rect 18630 -15230 18685 -15110
rect 18805 -15230 18850 -15110
rect 18970 -15230 19015 -15110
rect 19135 -15230 19180 -15110
rect 19300 -15230 19355 -15110
rect 19475 -15230 19520 -15110
rect 19640 -15230 19685 -15110
rect 19805 -15230 19850 -15110
rect 19970 -15230 20025 -15110
rect 20145 -15230 20190 -15110
rect 20310 -15230 20355 -15110
rect 20475 -15230 20520 -15110
rect 20640 -15230 20695 -15110
rect 20815 -15230 20860 -15110
rect 20980 -15230 21025 -15110
rect 21145 -15230 21190 -15110
rect 21310 -15230 21365 -15110
rect 21485 -15230 21530 -15110
rect 21650 -15230 21695 -15110
rect 21815 -15230 21860 -15110
rect 21980 -15230 22035 -15110
rect 22155 -15230 22200 -15110
rect 22320 -15230 22365 -15110
rect 22485 -15230 22530 -15110
rect 22650 -15230 22705 -15110
rect 22825 -15230 22870 -15110
rect 22990 -15230 23035 -15110
rect 23155 -15230 23200 -15110
rect 23320 -15230 23375 -15110
rect 23495 -15230 23540 -15110
rect 23660 -15230 23705 -15110
rect 23825 -15230 23870 -15110
rect 23990 -15230 24000 -15110
rect 18500 -15275 24000 -15230
rect 18500 -15395 18510 -15275
rect 18630 -15395 18685 -15275
rect 18805 -15395 18850 -15275
rect 18970 -15395 19015 -15275
rect 19135 -15395 19180 -15275
rect 19300 -15395 19355 -15275
rect 19475 -15395 19520 -15275
rect 19640 -15395 19685 -15275
rect 19805 -15395 19850 -15275
rect 19970 -15395 20025 -15275
rect 20145 -15395 20190 -15275
rect 20310 -15395 20355 -15275
rect 20475 -15395 20520 -15275
rect 20640 -15395 20695 -15275
rect 20815 -15395 20860 -15275
rect 20980 -15395 21025 -15275
rect 21145 -15395 21190 -15275
rect 21310 -15395 21365 -15275
rect 21485 -15395 21530 -15275
rect 21650 -15395 21695 -15275
rect 21815 -15395 21860 -15275
rect 21980 -15395 22035 -15275
rect 22155 -15395 22200 -15275
rect 22320 -15395 22365 -15275
rect 22485 -15395 22530 -15275
rect 22650 -15395 22705 -15275
rect 22825 -15395 22870 -15275
rect 22990 -15395 23035 -15275
rect 23155 -15395 23200 -15275
rect 23320 -15395 23375 -15275
rect 23495 -15395 23540 -15275
rect 23660 -15395 23705 -15275
rect 23825 -15395 23870 -15275
rect 23990 -15395 24000 -15275
rect 18500 -15450 24000 -15395
rect 18500 -15570 18510 -15450
rect 18630 -15570 18685 -15450
rect 18805 -15570 18850 -15450
rect 18970 -15570 19015 -15450
rect 19135 -15570 19180 -15450
rect 19300 -15570 19355 -15450
rect 19475 -15570 19520 -15450
rect 19640 -15570 19685 -15450
rect 19805 -15570 19850 -15450
rect 19970 -15570 20025 -15450
rect 20145 -15570 20190 -15450
rect 20310 -15570 20355 -15450
rect 20475 -15570 20520 -15450
rect 20640 -15570 20695 -15450
rect 20815 -15570 20860 -15450
rect 20980 -15570 21025 -15450
rect 21145 -15570 21190 -15450
rect 21310 -15570 21365 -15450
rect 21485 -15570 21530 -15450
rect 21650 -15570 21695 -15450
rect 21815 -15570 21860 -15450
rect 21980 -15570 22035 -15450
rect 22155 -15570 22200 -15450
rect 22320 -15570 22365 -15450
rect 22485 -15570 22530 -15450
rect 22650 -15570 22705 -15450
rect 22825 -15570 22870 -15450
rect 22990 -15570 23035 -15450
rect 23155 -15570 23200 -15450
rect 23320 -15570 23375 -15450
rect 23495 -15570 23540 -15450
rect 23660 -15570 23705 -15450
rect 23825 -15570 23870 -15450
rect 23990 -15570 24000 -15450
rect 18500 -15580 24000 -15570
rect 24190 -10090 29690 -10080
rect 24190 -10210 24200 -10090
rect 24320 -10210 24375 -10090
rect 24495 -10210 24540 -10090
rect 24660 -10210 24705 -10090
rect 24825 -10210 24870 -10090
rect 24990 -10210 25045 -10090
rect 25165 -10210 25210 -10090
rect 25330 -10210 25375 -10090
rect 25495 -10210 25540 -10090
rect 25660 -10210 25715 -10090
rect 25835 -10210 25880 -10090
rect 26000 -10210 26045 -10090
rect 26165 -10210 26210 -10090
rect 26330 -10210 26385 -10090
rect 26505 -10210 26550 -10090
rect 26670 -10210 26715 -10090
rect 26835 -10210 26880 -10090
rect 27000 -10210 27055 -10090
rect 27175 -10210 27220 -10090
rect 27340 -10210 27385 -10090
rect 27505 -10210 27550 -10090
rect 27670 -10210 27725 -10090
rect 27845 -10210 27890 -10090
rect 28010 -10210 28055 -10090
rect 28175 -10210 28220 -10090
rect 28340 -10210 28395 -10090
rect 28515 -10210 28560 -10090
rect 28680 -10210 28725 -10090
rect 28845 -10210 28890 -10090
rect 29010 -10210 29065 -10090
rect 29185 -10210 29230 -10090
rect 29350 -10210 29395 -10090
rect 29515 -10210 29560 -10090
rect 29680 -10210 29690 -10090
rect 24190 -10255 29690 -10210
rect 24190 -10375 24200 -10255
rect 24320 -10375 24375 -10255
rect 24495 -10375 24540 -10255
rect 24660 -10375 24705 -10255
rect 24825 -10375 24870 -10255
rect 24990 -10375 25045 -10255
rect 25165 -10375 25210 -10255
rect 25330 -10375 25375 -10255
rect 25495 -10375 25540 -10255
rect 25660 -10375 25715 -10255
rect 25835 -10375 25880 -10255
rect 26000 -10375 26045 -10255
rect 26165 -10375 26210 -10255
rect 26330 -10375 26385 -10255
rect 26505 -10375 26550 -10255
rect 26670 -10375 26715 -10255
rect 26835 -10375 26880 -10255
rect 27000 -10375 27055 -10255
rect 27175 -10375 27220 -10255
rect 27340 -10375 27385 -10255
rect 27505 -10375 27550 -10255
rect 27670 -10375 27725 -10255
rect 27845 -10375 27890 -10255
rect 28010 -10375 28055 -10255
rect 28175 -10375 28220 -10255
rect 28340 -10375 28395 -10255
rect 28515 -10375 28560 -10255
rect 28680 -10375 28725 -10255
rect 28845 -10375 28890 -10255
rect 29010 -10375 29065 -10255
rect 29185 -10375 29230 -10255
rect 29350 -10375 29395 -10255
rect 29515 -10375 29560 -10255
rect 29680 -10375 29690 -10255
rect 24190 -10420 29690 -10375
rect 24190 -10540 24200 -10420
rect 24320 -10540 24375 -10420
rect 24495 -10540 24540 -10420
rect 24660 -10540 24705 -10420
rect 24825 -10540 24870 -10420
rect 24990 -10540 25045 -10420
rect 25165 -10540 25210 -10420
rect 25330 -10540 25375 -10420
rect 25495 -10540 25540 -10420
rect 25660 -10540 25715 -10420
rect 25835 -10540 25880 -10420
rect 26000 -10540 26045 -10420
rect 26165 -10540 26210 -10420
rect 26330 -10540 26385 -10420
rect 26505 -10540 26550 -10420
rect 26670 -10540 26715 -10420
rect 26835 -10540 26880 -10420
rect 27000 -10540 27055 -10420
rect 27175 -10540 27220 -10420
rect 27340 -10540 27385 -10420
rect 27505 -10540 27550 -10420
rect 27670 -10540 27725 -10420
rect 27845 -10540 27890 -10420
rect 28010 -10540 28055 -10420
rect 28175 -10540 28220 -10420
rect 28340 -10540 28395 -10420
rect 28515 -10540 28560 -10420
rect 28680 -10540 28725 -10420
rect 28845 -10540 28890 -10420
rect 29010 -10540 29065 -10420
rect 29185 -10540 29230 -10420
rect 29350 -10540 29395 -10420
rect 29515 -10540 29560 -10420
rect 29680 -10540 29690 -10420
rect 24190 -10585 29690 -10540
rect 24190 -10705 24200 -10585
rect 24320 -10705 24375 -10585
rect 24495 -10705 24540 -10585
rect 24660 -10705 24705 -10585
rect 24825 -10705 24870 -10585
rect 24990 -10705 25045 -10585
rect 25165 -10705 25210 -10585
rect 25330 -10705 25375 -10585
rect 25495 -10705 25540 -10585
rect 25660 -10705 25715 -10585
rect 25835 -10705 25880 -10585
rect 26000 -10705 26045 -10585
rect 26165 -10705 26210 -10585
rect 26330 -10705 26385 -10585
rect 26505 -10705 26550 -10585
rect 26670 -10705 26715 -10585
rect 26835 -10705 26880 -10585
rect 27000 -10705 27055 -10585
rect 27175 -10705 27220 -10585
rect 27340 -10705 27385 -10585
rect 27505 -10705 27550 -10585
rect 27670 -10705 27725 -10585
rect 27845 -10705 27890 -10585
rect 28010 -10705 28055 -10585
rect 28175 -10705 28220 -10585
rect 28340 -10705 28395 -10585
rect 28515 -10705 28560 -10585
rect 28680 -10705 28725 -10585
rect 28845 -10705 28890 -10585
rect 29010 -10705 29065 -10585
rect 29185 -10705 29230 -10585
rect 29350 -10705 29395 -10585
rect 29515 -10705 29560 -10585
rect 29680 -10705 29690 -10585
rect 24190 -10760 29690 -10705
rect 24190 -10880 24200 -10760
rect 24320 -10880 24375 -10760
rect 24495 -10880 24540 -10760
rect 24660 -10880 24705 -10760
rect 24825 -10880 24870 -10760
rect 24990 -10880 25045 -10760
rect 25165 -10880 25210 -10760
rect 25330 -10880 25375 -10760
rect 25495 -10880 25540 -10760
rect 25660 -10880 25715 -10760
rect 25835 -10880 25880 -10760
rect 26000 -10880 26045 -10760
rect 26165 -10880 26210 -10760
rect 26330 -10880 26385 -10760
rect 26505 -10880 26550 -10760
rect 26670 -10880 26715 -10760
rect 26835 -10880 26880 -10760
rect 27000 -10880 27055 -10760
rect 27175 -10880 27220 -10760
rect 27340 -10880 27385 -10760
rect 27505 -10880 27550 -10760
rect 27670 -10880 27725 -10760
rect 27845 -10880 27890 -10760
rect 28010 -10880 28055 -10760
rect 28175 -10880 28220 -10760
rect 28340 -10880 28395 -10760
rect 28515 -10880 28560 -10760
rect 28680 -10880 28725 -10760
rect 28845 -10880 28890 -10760
rect 29010 -10880 29065 -10760
rect 29185 -10880 29230 -10760
rect 29350 -10880 29395 -10760
rect 29515 -10880 29560 -10760
rect 29680 -10880 29690 -10760
rect 24190 -10925 29690 -10880
rect 24190 -11045 24200 -10925
rect 24320 -11045 24375 -10925
rect 24495 -11045 24540 -10925
rect 24660 -11045 24705 -10925
rect 24825 -11045 24870 -10925
rect 24990 -11045 25045 -10925
rect 25165 -11045 25210 -10925
rect 25330 -11045 25375 -10925
rect 25495 -11045 25540 -10925
rect 25660 -11045 25715 -10925
rect 25835 -11045 25880 -10925
rect 26000 -11045 26045 -10925
rect 26165 -11045 26210 -10925
rect 26330 -11045 26385 -10925
rect 26505 -11045 26550 -10925
rect 26670 -11045 26715 -10925
rect 26835 -11045 26880 -10925
rect 27000 -11045 27055 -10925
rect 27175 -11045 27220 -10925
rect 27340 -11045 27385 -10925
rect 27505 -11045 27550 -10925
rect 27670 -11045 27725 -10925
rect 27845 -11045 27890 -10925
rect 28010 -11045 28055 -10925
rect 28175 -11045 28220 -10925
rect 28340 -11045 28395 -10925
rect 28515 -11045 28560 -10925
rect 28680 -11045 28725 -10925
rect 28845 -11045 28890 -10925
rect 29010 -11045 29065 -10925
rect 29185 -11045 29230 -10925
rect 29350 -11045 29395 -10925
rect 29515 -11045 29560 -10925
rect 29680 -11045 29690 -10925
rect 24190 -11090 29690 -11045
rect 24190 -11210 24200 -11090
rect 24320 -11210 24375 -11090
rect 24495 -11210 24540 -11090
rect 24660 -11210 24705 -11090
rect 24825 -11210 24870 -11090
rect 24990 -11210 25045 -11090
rect 25165 -11210 25210 -11090
rect 25330 -11210 25375 -11090
rect 25495 -11210 25540 -11090
rect 25660 -11210 25715 -11090
rect 25835 -11210 25880 -11090
rect 26000 -11210 26045 -11090
rect 26165 -11210 26210 -11090
rect 26330 -11210 26385 -11090
rect 26505 -11210 26550 -11090
rect 26670 -11210 26715 -11090
rect 26835 -11210 26880 -11090
rect 27000 -11210 27055 -11090
rect 27175 -11210 27220 -11090
rect 27340 -11210 27385 -11090
rect 27505 -11210 27550 -11090
rect 27670 -11210 27725 -11090
rect 27845 -11210 27890 -11090
rect 28010 -11210 28055 -11090
rect 28175 -11210 28220 -11090
rect 28340 -11210 28395 -11090
rect 28515 -11210 28560 -11090
rect 28680 -11210 28725 -11090
rect 28845 -11210 28890 -11090
rect 29010 -11210 29065 -11090
rect 29185 -11210 29230 -11090
rect 29350 -11210 29395 -11090
rect 29515 -11210 29560 -11090
rect 29680 -11210 29690 -11090
rect 24190 -11255 29690 -11210
rect 24190 -11375 24200 -11255
rect 24320 -11375 24375 -11255
rect 24495 -11375 24540 -11255
rect 24660 -11375 24705 -11255
rect 24825 -11375 24870 -11255
rect 24990 -11375 25045 -11255
rect 25165 -11375 25210 -11255
rect 25330 -11375 25375 -11255
rect 25495 -11375 25540 -11255
rect 25660 -11375 25715 -11255
rect 25835 -11375 25880 -11255
rect 26000 -11375 26045 -11255
rect 26165 -11375 26210 -11255
rect 26330 -11375 26385 -11255
rect 26505 -11375 26550 -11255
rect 26670 -11375 26715 -11255
rect 26835 -11375 26880 -11255
rect 27000 -11375 27055 -11255
rect 27175 -11375 27220 -11255
rect 27340 -11375 27385 -11255
rect 27505 -11375 27550 -11255
rect 27670 -11375 27725 -11255
rect 27845 -11375 27890 -11255
rect 28010 -11375 28055 -11255
rect 28175 -11375 28220 -11255
rect 28340 -11375 28395 -11255
rect 28515 -11375 28560 -11255
rect 28680 -11375 28725 -11255
rect 28845 -11375 28890 -11255
rect 29010 -11375 29065 -11255
rect 29185 -11375 29230 -11255
rect 29350 -11375 29395 -11255
rect 29515 -11375 29560 -11255
rect 29680 -11375 29690 -11255
rect 24190 -11430 29690 -11375
rect 24190 -11550 24200 -11430
rect 24320 -11550 24375 -11430
rect 24495 -11550 24540 -11430
rect 24660 -11550 24705 -11430
rect 24825 -11550 24870 -11430
rect 24990 -11550 25045 -11430
rect 25165 -11550 25210 -11430
rect 25330 -11550 25375 -11430
rect 25495 -11550 25540 -11430
rect 25660 -11550 25715 -11430
rect 25835 -11550 25880 -11430
rect 26000 -11550 26045 -11430
rect 26165 -11550 26210 -11430
rect 26330 -11550 26385 -11430
rect 26505 -11550 26550 -11430
rect 26670 -11550 26715 -11430
rect 26835 -11550 26880 -11430
rect 27000 -11550 27055 -11430
rect 27175 -11550 27220 -11430
rect 27340 -11550 27385 -11430
rect 27505 -11550 27550 -11430
rect 27670 -11550 27725 -11430
rect 27845 -11550 27890 -11430
rect 28010 -11550 28055 -11430
rect 28175 -11550 28220 -11430
rect 28340 -11550 28395 -11430
rect 28515 -11550 28560 -11430
rect 28680 -11550 28725 -11430
rect 28845 -11550 28890 -11430
rect 29010 -11550 29065 -11430
rect 29185 -11550 29230 -11430
rect 29350 -11550 29395 -11430
rect 29515 -11550 29560 -11430
rect 29680 -11550 29690 -11430
rect 24190 -11595 29690 -11550
rect 24190 -11715 24200 -11595
rect 24320 -11715 24375 -11595
rect 24495 -11715 24540 -11595
rect 24660 -11715 24705 -11595
rect 24825 -11715 24870 -11595
rect 24990 -11715 25045 -11595
rect 25165 -11715 25210 -11595
rect 25330 -11715 25375 -11595
rect 25495 -11715 25540 -11595
rect 25660 -11715 25715 -11595
rect 25835 -11715 25880 -11595
rect 26000 -11715 26045 -11595
rect 26165 -11715 26210 -11595
rect 26330 -11715 26385 -11595
rect 26505 -11715 26550 -11595
rect 26670 -11715 26715 -11595
rect 26835 -11715 26880 -11595
rect 27000 -11715 27055 -11595
rect 27175 -11715 27220 -11595
rect 27340 -11715 27385 -11595
rect 27505 -11715 27550 -11595
rect 27670 -11715 27725 -11595
rect 27845 -11715 27890 -11595
rect 28010 -11715 28055 -11595
rect 28175 -11715 28220 -11595
rect 28340 -11715 28395 -11595
rect 28515 -11715 28560 -11595
rect 28680 -11715 28725 -11595
rect 28845 -11715 28890 -11595
rect 29010 -11715 29065 -11595
rect 29185 -11715 29230 -11595
rect 29350 -11715 29395 -11595
rect 29515 -11715 29560 -11595
rect 29680 -11715 29690 -11595
rect 24190 -11760 29690 -11715
rect 24190 -11880 24200 -11760
rect 24320 -11880 24375 -11760
rect 24495 -11880 24540 -11760
rect 24660 -11880 24705 -11760
rect 24825 -11880 24870 -11760
rect 24990 -11880 25045 -11760
rect 25165 -11880 25210 -11760
rect 25330 -11880 25375 -11760
rect 25495 -11880 25540 -11760
rect 25660 -11880 25715 -11760
rect 25835 -11880 25880 -11760
rect 26000 -11880 26045 -11760
rect 26165 -11880 26210 -11760
rect 26330 -11880 26385 -11760
rect 26505 -11880 26550 -11760
rect 26670 -11880 26715 -11760
rect 26835 -11880 26880 -11760
rect 27000 -11880 27055 -11760
rect 27175 -11880 27220 -11760
rect 27340 -11880 27385 -11760
rect 27505 -11880 27550 -11760
rect 27670 -11880 27725 -11760
rect 27845 -11880 27890 -11760
rect 28010 -11880 28055 -11760
rect 28175 -11880 28220 -11760
rect 28340 -11880 28395 -11760
rect 28515 -11880 28560 -11760
rect 28680 -11880 28725 -11760
rect 28845 -11880 28890 -11760
rect 29010 -11880 29065 -11760
rect 29185 -11880 29230 -11760
rect 29350 -11880 29395 -11760
rect 29515 -11880 29560 -11760
rect 29680 -11880 29690 -11760
rect 24190 -11925 29690 -11880
rect 24190 -12045 24200 -11925
rect 24320 -12045 24375 -11925
rect 24495 -12045 24540 -11925
rect 24660 -12045 24705 -11925
rect 24825 -12045 24870 -11925
rect 24990 -12045 25045 -11925
rect 25165 -12045 25210 -11925
rect 25330 -12045 25375 -11925
rect 25495 -12045 25540 -11925
rect 25660 -12045 25715 -11925
rect 25835 -12045 25880 -11925
rect 26000 -12045 26045 -11925
rect 26165 -12045 26210 -11925
rect 26330 -12045 26385 -11925
rect 26505 -12045 26550 -11925
rect 26670 -12045 26715 -11925
rect 26835 -12045 26880 -11925
rect 27000 -12045 27055 -11925
rect 27175 -12045 27220 -11925
rect 27340 -12045 27385 -11925
rect 27505 -12045 27550 -11925
rect 27670 -12045 27725 -11925
rect 27845 -12045 27890 -11925
rect 28010 -12045 28055 -11925
rect 28175 -12045 28220 -11925
rect 28340 -12045 28395 -11925
rect 28515 -12045 28560 -11925
rect 28680 -12045 28725 -11925
rect 28845 -12045 28890 -11925
rect 29010 -12045 29065 -11925
rect 29185 -12045 29230 -11925
rect 29350 -12045 29395 -11925
rect 29515 -12045 29560 -11925
rect 29680 -12045 29690 -11925
rect 24190 -12100 29690 -12045
rect 24190 -12220 24200 -12100
rect 24320 -12220 24375 -12100
rect 24495 -12220 24540 -12100
rect 24660 -12220 24705 -12100
rect 24825 -12220 24870 -12100
rect 24990 -12220 25045 -12100
rect 25165 -12220 25210 -12100
rect 25330 -12220 25375 -12100
rect 25495 -12220 25540 -12100
rect 25660 -12220 25715 -12100
rect 25835 -12220 25880 -12100
rect 26000 -12220 26045 -12100
rect 26165 -12220 26210 -12100
rect 26330 -12220 26385 -12100
rect 26505 -12220 26550 -12100
rect 26670 -12220 26715 -12100
rect 26835 -12220 26880 -12100
rect 27000 -12220 27055 -12100
rect 27175 -12220 27220 -12100
rect 27340 -12220 27385 -12100
rect 27505 -12220 27550 -12100
rect 27670 -12220 27725 -12100
rect 27845 -12220 27890 -12100
rect 28010 -12220 28055 -12100
rect 28175 -12220 28220 -12100
rect 28340 -12220 28395 -12100
rect 28515 -12220 28560 -12100
rect 28680 -12220 28725 -12100
rect 28845 -12220 28890 -12100
rect 29010 -12220 29065 -12100
rect 29185 -12220 29230 -12100
rect 29350 -12220 29395 -12100
rect 29515 -12220 29560 -12100
rect 29680 -12220 29690 -12100
rect 24190 -12265 29690 -12220
rect 24190 -12385 24200 -12265
rect 24320 -12385 24375 -12265
rect 24495 -12385 24540 -12265
rect 24660 -12385 24705 -12265
rect 24825 -12385 24870 -12265
rect 24990 -12385 25045 -12265
rect 25165 -12385 25210 -12265
rect 25330 -12385 25375 -12265
rect 25495 -12385 25540 -12265
rect 25660 -12385 25715 -12265
rect 25835 -12385 25880 -12265
rect 26000 -12385 26045 -12265
rect 26165 -12385 26210 -12265
rect 26330 -12385 26385 -12265
rect 26505 -12385 26550 -12265
rect 26670 -12385 26715 -12265
rect 26835 -12385 26880 -12265
rect 27000 -12385 27055 -12265
rect 27175 -12385 27220 -12265
rect 27340 -12385 27385 -12265
rect 27505 -12385 27550 -12265
rect 27670 -12385 27725 -12265
rect 27845 -12385 27890 -12265
rect 28010 -12385 28055 -12265
rect 28175 -12385 28220 -12265
rect 28340 -12385 28395 -12265
rect 28515 -12385 28560 -12265
rect 28680 -12385 28725 -12265
rect 28845 -12385 28890 -12265
rect 29010 -12385 29065 -12265
rect 29185 -12385 29230 -12265
rect 29350 -12385 29395 -12265
rect 29515 -12385 29560 -12265
rect 29680 -12385 29690 -12265
rect 24190 -12430 29690 -12385
rect 24190 -12550 24200 -12430
rect 24320 -12550 24375 -12430
rect 24495 -12550 24540 -12430
rect 24660 -12550 24705 -12430
rect 24825 -12550 24870 -12430
rect 24990 -12550 25045 -12430
rect 25165 -12550 25210 -12430
rect 25330 -12550 25375 -12430
rect 25495 -12550 25540 -12430
rect 25660 -12550 25715 -12430
rect 25835 -12550 25880 -12430
rect 26000 -12550 26045 -12430
rect 26165 -12550 26210 -12430
rect 26330 -12550 26385 -12430
rect 26505 -12550 26550 -12430
rect 26670 -12550 26715 -12430
rect 26835 -12550 26880 -12430
rect 27000 -12550 27055 -12430
rect 27175 -12550 27220 -12430
rect 27340 -12550 27385 -12430
rect 27505 -12550 27550 -12430
rect 27670 -12550 27725 -12430
rect 27845 -12550 27890 -12430
rect 28010 -12550 28055 -12430
rect 28175 -12550 28220 -12430
rect 28340 -12550 28395 -12430
rect 28515 -12550 28560 -12430
rect 28680 -12550 28725 -12430
rect 28845 -12550 28890 -12430
rect 29010 -12550 29065 -12430
rect 29185 -12550 29230 -12430
rect 29350 -12550 29395 -12430
rect 29515 -12550 29560 -12430
rect 29680 -12550 29690 -12430
rect 24190 -12595 29690 -12550
rect 24190 -12715 24200 -12595
rect 24320 -12715 24375 -12595
rect 24495 -12715 24540 -12595
rect 24660 -12715 24705 -12595
rect 24825 -12715 24870 -12595
rect 24990 -12715 25045 -12595
rect 25165 -12715 25210 -12595
rect 25330 -12715 25375 -12595
rect 25495 -12715 25540 -12595
rect 25660 -12715 25715 -12595
rect 25835 -12715 25880 -12595
rect 26000 -12715 26045 -12595
rect 26165 -12715 26210 -12595
rect 26330 -12715 26385 -12595
rect 26505 -12715 26550 -12595
rect 26670 -12715 26715 -12595
rect 26835 -12715 26880 -12595
rect 27000 -12715 27055 -12595
rect 27175 -12715 27220 -12595
rect 27340 -12715 27385 -12595
rect 27505 -12715 27550 -12595
rect 27670 -12715 27725 -12595
rect 27845 -12715 27890 -12595
rect 28010 -12715 28055 -12595
rect 28175 -12715 28220 -12595
rect 28340 -12715 28395 -12595
rect 28515 -12715 28560 -12595
rect 28680 -12715 28725 -12595
rect 28845 -12715 28890 -12595
rect 29010 -12715 29065 -12595
rect 29185 -12715 29230 -12595
rect 29350 -12715 29395 -12595
rect 29515 -12715 29560 -12595
rect 29680 -12715 29690 -12595
rect 24190 -12770 29690 -12715
rect 24190 -12890 24200 -12770
rect 24320 -12890 24375 -12770
rect 24495 -12890 24540 -12770
rect 24660 -12890 24705 -12770
rect 24825 -12890 24870 -12770
rect 24990 -12890 25045 -12770
rect 25165 -12890 25210 -12770
rect 25330 -12890 25375 -12770
rect 25495 -12890 25540 -12770
rect 25660 -12890 25715 -12770
rect 25835 -12890 25880 -12770
rect 26000 -12890 26045 -12770
rect 26165 -12890 26210 -12770
rect 26330 -12890 26385 -12770
rect 26505 -12890 26550 -12770
rect 26670 -12890 26715 -12770
rect 26835 -12890 26880 -12770
rect 27000 -12890 27055 -12770
rect 27175 -12890 27220 -12770
rect 27340 -12890 27385 -12770
rect 27505 -12890 27550 -12770
rect 27670 -12890 27725 -12770
rect 27845 -12890 27890 -12770
rect 28010 -12890 28055 -12770
rect 28175 -12890 28220 -12770
rect 28340 -12890 28395 -12770
rect 28515 -12890 28560 -12770
rect 28680 -12890 28725 -12770
rect 28845 -12890 28890 -12770
rect 29010 -12890 29065 -12770
rect 29185 -12890 29230 -12770
rect 29350 -12890 29395 -12770
rect 29515 -12890 29560 -12770
rect 29680 -12890 29690 -12770
rect 24190 -12935 29690 -12890
rect 24190 -13055 24200 -12935
rect 24320 -13055 24375 -12935
rect 24495 -13055 24540 -12935
rect 24660 -13055 24705 -12935
rect 24825 -13055 24870 -12935
rect 24990 -13055 25045 -12935
rect 25165 -13055 25210 -12935
rect 25330 -13055 25375 -12935
rect 25495 -13055 25540 -12935
rect 25660 -13055 25715 -12935
rect 25835 -13055 25880 -12935
rect 26000 -13055 26045 -12935
rect 26165 -13055 26210 -12935
rect 26330 -13055 26385 -12935
rect 26505 -13055 26550 -12935
rect 26670 -13055 26715 -12935
rect 26835 -13055 26880 -12935
rect 27000 -13055 27055 -12935
rect 27175 -13055 27220 -12935
rect 27340 -13055 27385 -12935
rect 27505 -13055 27550 -12935
rect 27670 -13055 27725 -12935
rect 27845 -13055 27890 -12935
rect 28010 -13055 28055 -12935
rect 28175 -13055 28220 -12935
rect 28340 -13055 28395 -12935
rect 28515 -13055 28560 -12935
rect 28680 -13055 28725 -12935
rect 28845 -13055 28890 -12935
rect 29010 -13055 29065 -12935
rect 29185 -13055 29230 -12935
rect 29350 -13055 29395 -12935
rect 29515 -13055 29560 -12935
rect 29680 -13055 29690 -12935
rect 24190 -13100 29690 -13055
rect 24190 -13220 24200 -13100
rect 24320 -13220 24375 -13100
rect 24495 -13220 24540 -13100
rect 24660 -13220 24705 -13100
rect 24825 -13220 24870 -13100
rect 24990 -13220 25045 -13100
rect 25165 -13220 25210 -13100
rect 25330 -13220 25375 -13100
rect 25495 -13220 25540 -13100
rect 25660 -13220 25715 -13100
rect 25835 -13220 25880 -13100
rect 26000 -13220 26045 -13100
rect 26165 -13220 26210 -13100
rect 26330 -13220 26385 -13100
rect 26505 -13220 26550 -13100
rect 26670 -13220 26715 -13100
rect 26835 -13220 26880 -13100
rect 27000 -13220 27055 -13100
rect 27175 -13220 27220 -13100
rect 27340 -13220 27385 -13100
rect 27505 -13220 27550 -13100
rect 27670 -13220 27725 -13100
rect 27845 -13220 27890 -13100
rect 28010 -13220 28055 -13100
rect 28175 -13220 28220 -13100
rect 28340 -13220 28395 -13100
rect 28515 -13220 28560 -13100
rect 28680 -13220 28725 -13100
rect 28845 -13220 28890 -13100
rect 29010 -13220 29065 -13100
rect 29185 -13220 29230 -13100
rect 29350 -13220 29395 -13100
rect 29515 -13220 29560 -13100
rect 29680 -13220 29690 -13100
rect 24190 -13265 29690 -13220
rect 24190 -13385 24200 -13265
rect 24320 -13385 24375 -13265
rect 24495 -13385 24540 -13265
rect 24660 -13385 24705 -13265
rect 24825 -13385 24870 -13265
rect 24990 -13385 25045 -13265
rect 25165 -13385 25210 -13265
rect 25330 -13385 25375 -13265
rect 25495 -13385 25540 -13265
rect 25660 -13385 25715 -13265
rect 25835 -13385 25880 -13265
rect 26000 -13385 26045 -13265
rect 26165 -13385 26210 -13265
rect 26330 -13385 26385 -13265
rect 26505 -13385 26550 -13265
rect 26670 -13385 26715 -13265
rect 26835 -13385 26880 -13265
rect 27000 -13385 27055 -13265
rect 27175 -13385 27220 -13265
rect 27340 -13385 27385 -13265
rect 27505 -13385 27550 -13265
rect 27670 -13385 27725 -13265
rect 27845 -13385 27890 -13265
rect 28010 -13385 28055 -13265
rect 28175 -13385 28220 -13265
rect 28340 -13385 28395 -13265
rect 28515 -13385 28560 -13265
rect 28680 -13385 28725 -13265
rect 28845 -13385 28890 -13265
rect 29010 -13385 29065 -13265
rect 29185 -13385 29230 -13265
rect 29350 -13385 29395 -13265
rect 29515 -13385 29560 -13265
rect 29680 -13385 29690 -13265
rect 24190 -13440 29690 -13385
rect 24190 -13560 24200 -13440
rect 24320 -13560 24375 -13440
rect 24495 -13560 24540 -13440
rect 24660 -13560 24705 -13440
rect 24825 -13560 24870 -13440
rect 24990 -13560 25045 -13440
rect 25165 -13560 25210 -13440
rect 25330 -13560 25375 -13440
rect 25495 -13560 25540 -13440
rect 25660 -13560 25715 -13440
rect 25835 -13560 25880 -13440
rect 26000 -13560 26045 -13440
rect 26165 -13560 26210 -13440
rect 26330 -13560 26385 -13440
rect 26505 -13560 26550 -13440
rect 26670 -13560 26715 -13440
rect 26835 -13560 26880 -13440
rect 27000 -13560 27055 -13440
rect 27175 -13560 27220 -13440
rect 27340 -13560 27385 -13440
rect 27505 -13560 27550 -13440
rect 27670 -13560 27725 -13440
rect 27845 -13560 27890 -13440
rect 28010 -13560 28055 -13440
rect 28175 -13560 28220 -13440
rect 28340 -13560 28395 -13440
rect 28515 -13560 28560 -13440
rect 28680 -13560 28725 -13440
rect 28845 -13560 28890 -13440
rect 29010 -13560 29065 -13440
rect 29185 -13560 29230 -13440
rect 29350 -13560 29395 -13440
rect 29515 -13560 29560 -13440
rect 29680 -13560 29690 -13440
rect 24190 -13605 29690 -13560
rect 24190 -13725 24200 -13605
rect 24320 -13725 24375 -13605
rect 24495 -13725 24540 -13605
rect 24660 -13725 24705 -13605
rect 24825 -13725 24870 -13605
rect 24990 -13725 25045 -13605
rect 25165 -13725 25210 -13605
rect 25330 -13725 25375 -13605
rect 25495 -13725 25540 -13605
rect 25660 -13725 25715 -13605
rect 25835 -13725 25880 -13605
rect 26000 -13725 26045 -13605
rect 26165 -13725 26210 -13605
rect 26330 -13725 26385 -13605
rect 26505 -13725 26550 -13605
rect 26670 -13725 26715 -13605
rect 26835 -13725 26880 -13605
rect 27000 -13725 27055 -13605
rect 27175 -13725 27220 -13605
rect 27340 -13725 27385 -13605
rect 27505 -13725 27550 -13605
rect 27670 -13725 27725 -13605
rect 27845 -13725 27890 -13605
rect 28010 -13725 28055 -13605
rect 28175 -13725 28220 -13605
rect 28340 -13725 28395 -13605
rect 28515 -13725 28560 -13605
rect 28680 -13725 28725 -13605
rect 28845 -13725 28890 -13605
rect 29010 -13725 29065 -13605
rect 29185 -13725 29230 -13605
rect 29350 -13725 29395 -13605
rect 29515 -13725 29560 -13605
rect 29680 -13725 29690 -13605
rect 24190 -13770 29690 -13725
rect 24190 -13890 24200 -13770
rect 24320 -13890 24375 -13770
rect 24495 -13890 24540 -13770
rect 24660 -13890 24705 -13770
rect 24825 -13890 24870 -13770
rect 24990 -13890 25045 -13770
rect 25165 -13890 25210 -13770
rect 25330 -13890 25375 -13770
rect 25495 -13890 25540 -13770
rect 25660 -13890 25715 -13770
rect 25835 -13890 25880 -13770
rect 26000 -13890 26045 -13770
rect 26165 -13890 26210 -13770
rect 26330 -13890 26385 -13770
rect 26505 -13890 26550 -13770
rect 26670 -13890 26715 -13770
rect 26835 -13890 26880 -13770
rect 27000 -13890 27055 -13770
rect 27175 -13890 27220 -13770
rect 27340 -13890 27385 -13770
rect 27505 -13890 27550 -13770
rect 27670 -13890 27725 -13770
rect 27845 -13890 27890 -13770
rect 28010 -13890 28055 -13770
rect 28175 -13890 28220 -13770
rect 28340 -13890 28395 -13770
rect 28515 -13890 28560 -13770
rect 28680 -13890 28725 -13770
rect 28845 -13890 28890 -13770
rect 29010 -13890 29065 -13770
rect 29185 -13890 29230 -13770
rect 29350 -13890 29395 -13770
rect 29515 -13890 29560 -13770
rect 29680 -13890 29690 -13770
rect 24190 -13935 29690 -13890
rect 24190 -14055 24200 -13935
rect 24320 -14055 24375 -13935
rect 24495 -14055 24540 -13935
rect 24660 -14055 24705 -13935
rect 24825 -14055 24870 -13935
rect 24990 -14055 25045 -13935
rect 25165 -14055 25210 -13935
rect 25330 -14055 25375 -13935
rect 25495 -14055 25540 -13935
rect 25660 -14055 25715 -13935
rect 25835 -14055 25880 -13935
rect 26000 -14055 26045 -13935
rect 26165 -14055 26210 -13935
rect 26330 -14055 26385 -13935
rect 26505 -14055 26550 -13935
rect 26670 -14055 26715 -13935
rect 26835 -14055 26880 -13935
rect 27000 -14055 27055 -13935
rect 27175 -14055 27220 -13935
rect 27340 -14055 27385 -13935
rect 27505 -14055 27550 -13935
rect 27670 -14055 27725 -13935
rect 27845 -14055 27890 -13935
rect 28010 -14055 28055 -13935
rect 28175 -14055 28220 -13935
rect 28340 -14055 28395 -13935
rect 28515 -14055 28560 -13935
rect 28680 -14055 28725 -13935
rect 28845 -14055 28890 -13935
rect 29010 -14055 29065 -13935
rect 29185 -14055 29230 -13935
rect 29350 -14055 29395 -13935
rect 29515 -14055 29560 -13935
rect 29680 -14055 29690 -13935
rect 24190 -14110 29690 -14055
rect 24190 -14230 24200 -14110
rect 24320 -14230 24375 -14110
rect 24495 -14230 24540 -14110
rect 24660 -14230 24705 -14110
rect 24825 -14230 24870 -14110
rect 24990 -14230 25045 -14110
rect 25165 -14230 25210 -14110
rect 25330 -14230 25375 -14110
rect 25495 -14230 25540 -14110
rect 25660 -14230 25715 -14110
rect 25835 -14230 25880 -14110
rect 26000 -14230 26045 -14110
rect 26165 -14230 26210 -14110
rect 26330 -14230 26385 -14110
rect 26505 -14230 26550 -14110
rect 26670 -14230 26715 -14110
rect 26835 -14230 26880 -14110
rect 27000 -14230 27055 -14110
rect 27175 -14230 27220 -14110
rect 27340 -14230 27385 -14110
rect 27505 -14230 27550 -14110
rect 27670 -14230 27725 -14110
rect 27845 -14230 27890 -14110
rect 28010 -14230 28055 -14110
rect 28175 -14230 28220 -14110
rect 28340 -14230 28395 -14110
rect 28515 -14230 28560 -14110
rect 28680 -14230 28725 -14110
rect 28845 -14230 28890 -14110
rect 29010 -14230 29065 -14110
rect 29185 -14230 29230 -14110
rect 29350 -14230 29395 -14110
rect 29515 -14230 29560 -14110
rect 29680 -14230 29690 -14110
rect 24190 -14275 29690 -14230
rect 24190 -14395 24200 -14275
rect 24320 -14395 24375 -14275
rect 24495 -14395 24540 -14275
rect 24660 -14395 24705 -14275
rect 24825 -14395 24870 -14275
rect 24990 -14395 25045 -14275
rect 25165 -14395 25210 -14275
rect 25330 -14395 25375 -14275
rect 25495 -14395 25540 -14275
rect 25660 -14395 25715 -14275
rect 25835 -14395 25880 -14275
rect 26000 -14395 26045 -14275
rect 26165 -14395 26210 -14275
rect 26330 -14395 26385 -14275
rect 26505 -14395 26550 -14275
rect 26670 -14395 26715 -14275
rect 26835 -14395 26880 -14275
rect 27000 -14395 27055 -14275
rect 27175 -14395 27220 -14275
rect 27340 -14395 27385 -14275
rect 27505 -14395 27550 -14275
rect 27670 -14395 27725 -14275
rect 27845 -14395 27890 -14275
rect 28010 -14395 28055 -14275
rect 28175 -14395 28220 -14275
rect 28340 -14395 28395 -14275
rect 28515 -14395 28560 -14275
rect 28680 -14395 28725 -14275
rect 28845 -14395 28890 -14275
rect 29010 -14395 29065 -14275
rect 29185 -14395 29230 -14275
rect 29350 -14395 29395 -14275
rect 29515 -14395 29560 -14275
rect 29680 -14395 29690 -14275
rect 24190 -14440 29690 -14395
rect 24190 -14560 24200 -14440
rect 24320 -14560 24375 -14440
rect 24495 -14560 24540 -14440
rect 24660 -14560 24705 -14440
rect 24825 -14560 24870 -14440
rect 24990 -14560 25045 -14440
rect 25165 -14560 25210 -14440
rect 25330 -14560 25375 -14440
rect 25495 -14560 25540 -14440
rect 25660 -14560 25715 -14440
rect 25835 -14560 25880 -14440
rect 26000 -14560 26045 -14440
rect 26165 -14560 26210 -14440
rect 26330 -14560 26385 -14440
rect 26505 -14560 26550 -14440
rect 26670 -14560 26715 -14440
rect 26835 -14560 26880 -14440
rect 27000 -14560 27055 -14440
rect 27175 -14560 27220 -14440
rect 27340 -14560 27385 -14440
rect 27505 -14560 27550 -14440
rect 27670 -14560 27725 -14440
rect 27845 -14560 27890 -14440
rect 28010 -14560 28055 -14440
rect 28175 -14560 28220 -14440
rect 28340 -14560 28395 -14440
rect 28515 -14560 28560 -14440
rect 28680 -14560 28725 -14440
rect 28845 -14560 28890 -14440
rect 29010 -14560 29065 -14440
rect 29185 -14560 29230 -14440
rect 29350 -14560 29395 -14440
rect 29515 -14560 29560 -14440
rect 29680 -14560 29690 -14440
rect 24190 -14605 29690 -14560
rect 24190 -14725 24200 -14605
rect 24320 -14725 24375 -14605
rect 24495 -14725 24540 -14605
rect 24660 -14725 24705 -14605
rect 24825 -14725 24870 -14605
rect 24990 -14725 25045 -14605
rect 25165 -14725 25210 -14605
rect 25330 -14725 25375 -14605
rect 25495 -14725 25540 -14605
rect 25660 -14725 25715 -14605
rect 25835 -14725 25880 -14605
rect 26000 -14725 26045 -14605
rect 26165 -14725 26210 -14605
rect 26330 -14725 26385 -14605
rect 26505 -14725 26550 -14605
rect 26670 -14725 26715 -14605
rect 26835 -14725 26880 -14605
rect 27000 -14725 27055 -14605
rect 27175 -14725 27220 -14605
rect 27340 -14725 27385 -14605
rect 27505 -14725 27550 -14605
rect 27670 -14725 27725 -14605
rect 27845 -14725 27890 -14605
rect 28010 -14725 28055 -14605
rect 28175 -14725 28220 -14605
rect 28340 -14725 28395 -14605
rect 28515 -14725 28560 -14605
rect 28680 -14725 28725 -14605
rect 28845 -14725 28890 -14605
rect 29010 -14725 29065 -14605
rect 29185 -14725 29230 -14605
rect 29350 -14725 29395 -14605
rect 29515 -14725 29560 -14605
rect 29680 -14725 29690 -14605
rect 24190 -14780 29690 -14725
rect 24190 -14900 24200 -14780
rect 24320 -14900 24375 -14780
rect 24495 -14900 24540 -14780
rect 24660 -14900 24705 -14780
rect 24825 -14900 24870 -14780
rect 24990 -14900 25045 -14780
rect 25165 -14900 25210 -14780
rect 25330 -14900 25375 -14780
rect 25495 -14900 25540 -14780
rect 25660 -14900 25715 -14780
rect 25835 -14900 25880 -14780
rect 26000 -14900 26045 -14780
rect 26165 -14900 26210 -14780
rect 26330 -14900 26385 -14780
rect 26505 -14900 26550 -14780
rect 26670 -14900 26715 -14780
rect 26835 -14900 26880 -14780
rect 27000 -14900 27055 -14780
rect 27175 -14900 27220 -14780
rect 27340 -14900 27385 -14780
rect 27505 -14900 27550 -14780
rect 27670 -14900 27725 -14780
rect 27845 -14900 27890 -14780
rect 28010 -14900 28055 -14780
rect 28175 -14900 28220 -14780
rect 28340 -14900 28395 -14780
rect 28515 -14900 28560 -14780
rect 28680 -14900 28725 -14780
rect 28845 -14900 28890 -14780
rect 29010 -14900 29065 -14780
rect 29185 -14900 29230 -14780
rect 29350 -14900 29395 -14780
rect 29515 -14900 29560 -14780
rect 29680 -14900 29690 -14780
rect 24190 -14945 29690 -14900
rect 24190 -15065 24200 -14945
rect 24320 -15065 24375 -14945
rect 24495 -15065 24540 -14945
rect 24660 -15065 24705 -14945
rect 24825 -15065 24870 -14945
rect 24990 -15065 25045 -14945
rect 25165 -15065 25210 -14945
rect 25330 -15065 25375 -14945
rect 25495 -15065 25540 -14945
rect 25660 -15065 25715 -14945
rect 25835 -15065 25880 -14945
rect 26000 -15065 26045 -14945
rect 26165 -15065 26210 -14945
rect 26330 -15065 26385 -14945
rect 26505 -15065 26550 -14945
rect 26670 -15065 26715 -14945
rect 26835 -15065 26880 -14945
rect 27000 -15065 27055 -14945
rect 27175 -15065 27220 -14945
rect 27340 -15065 27385 -14945
rect 27505 -15065 27550 -14945
rect 27670 -15065 27725 -14945
rect 27845 -15065 27890 -14945
rect 28010 -15065 28055 -14945
rect 28175 -15065 28220 -14945
rect 28340 -15065 28395 -14945
rect 28515 -15065 28560 -14945
rect 28680 -15065 28725 -14945
rect 28845 -15065 28890 -14945
rect 29010 -15065 29065 -14945
rect 29185 -15065 29230 -14945
rect 29350 -15065 29395 -14945
rect 29515 -15065 29560 -14945
rect 29680 -15065 29690 -14945
rect 24190 -15110 29690 -15065
rect 24190 -15230 24200 -15110
rect 24320 -15230 24375 -15110
rect 24495 -15230 24540 -15110
rect 24660 -15230 24705 -15110
rect 24825 -15230 24870 -15110
rect 24990 -15230 25045 -15110
rect 25165 -15230 25210 -15110
rect 25330 -15230 25375 -15110
rect 25495 -15230 25540 -15110
rect 25660 -15230 25715 -15110
rect 25835 -15230 25880 -15110
rect 26000 -15230 26045 -15110
rect 26165 -15230 26210 -15110
rect 26330 -15230 26385 -15110
rect 26505 -15230 26550 -15110
rect 26670 -15230 26715 -15110
rect 26835 -15230 26880 -15110
rect 27000 -15230 27055 -15110
rect 27175 -15230 27220 -15110
rect 27340 -15230 27385 -15110
rect 27505 -15230 27550 -15110
rect 27670 -15230 27725 -15110
rect 27845 -15230 27890 -15110
rect 28010 -15230 28055 -15110
rect 28175 -15230 28220 -15110
rect 28340 -15230 28395 -15110
rect 28515 -15230 28560 -15110
rect 28680 -15230 28725 -15110
rect 28845 -15230 28890 -15110
rect 29010 -15230 29065 -15110
rect 29185 -15230 29230 -15110
rect 29350 -15230 29395 -15110
rect 29515 -15230 29560 -15110
rect 29680 -15230 29690 -15110
rect 24190 -15275 29690 -15230
rect 24190 -15395 24200 -15275
rect 24320 -15395 24375 -15275
rect 24495 -15395 24540 -15275
rect 24660 -15395 24705 -15275
rect 24825 -15395 24870 -15275
rect 24990 -15395 25045 -15275
rect 25165 -15395 25210 -15275
rect 25330 -15395 25375 -15275
rect 25495 -15395 25540 -15275
rect 25660 -15395 25715 -15275
rect 25835 -15395 25880 -15275
rect 26000 -15395 26045 -15275
rect 26165 -15395 26210 -15275
rect 26330 -15395 26385 -15275
rect 26505 -15395 26550 -15275
rect 26670 -15395 26715 -15275
rect 26835 -15395 26880 -15275
rect 27000 -15395 27055 -15275
rect 27175 -15395 27220 -15275
rect 27340 -15395 27385 -15275
rect 27505 -15395 27550 -15275
rect 27670 -15395 27725 -15275
rect 27845 -15395 27890 -15275
rect 28010 -15395 28055 -15275
rect 28175 -15395 28220 -15275
rect 28340 -15395 28395 -15275
rect 28515 -15395 28560 -15275
rect 28680 -15395 28725 -15275
rect 28845 -15395 28890 -15275
rect 29010 -15395 29065 -15275
rect 29185 -15395 29230 -15275
rect 29350 -15395 29395 -15275
rect 29515 -15395 29560 -15275
rect 29680 -15395 29690 -15275
rect 24190 -15450 29690 -15395
rect 24190 -15570 24200 -15450
rect 24320 -15570 24375 -15450
rect 24495 -15570 24540 -15450
rect 24660 -15570 24705 -15450
rect 24825 -15570 24870 -15450
rect 24990 -15570 25045 -15450
rect 25165 -15570 25210 -15450
rect 25330 -15570 25375 -15450
rect 25495 -15570 25540 -15450
rect 25660 -15570 25715 -15450
rect 25835 -15570 25880 -15450
rect 26000 -15570 26045 -15450
rect 26165 -15570 26210 -15450
rect 26330 -15570 26385 -15450
rect 26505 -15570 26550 -15450
rect 26670 -15570 26715 -15450
rect 26835 -15570 26880 -15450
rect 27000 -15570 27055 -15450
rect 27175 -15570 27220 -15450
rect 27340 -15570 27385 -15450
rect 27505 -15570 27550 -15450
rect 27670 -15570 27725 -15450
rect 27845 -15570 27890 -15450
rect 28010 -15570 28055 -15450
rect 28175 -15570 28220 -15450
rect 28340 -15570 28395 -15450
rect 28515 -15570 28560 -15450
rect 28680 -15570 28725 -15450
rect 28845 -15570 28890 -15450
rect 29010 -15570 29065 -15450
rect 29185 -15570 29230 -15450
rect 29350 -15570 29395 -15450
rect 29515 -15570 29560 -15450
rect 29680 -15570 29690 -15450
rect 24190 -15580 29690 -15570
<< mimcapcontact >>
rect 7130 7040 7250 7160
rect 7295 7040 7415 7160
rect 7460 7040 7580 7160
rect 7625 7040 7745 7160
rect 7800 7040 7920 7160
rect 7965 7040 8085 7160
rect 8130 7040 8250 7160
rect 8295 7040 8415 7160
rect 8470 7040 8590 7160
rect 8635 7040 8755 7160
rect 8800 7040 8920 7160
rect 8965 7040 9085 7160
rect 9140 7040 9260 7160
rect 9305 7040 9425 7160
rect 9470 7040 9590 7160
rect 9635 7040 9755 7160
rect 9810 7040 9930 7160
rect 9975 7040 10095 7160
rect 10140 7040 10260 7160
rect 10305 7040 10425 7160
rect 10480 7040 10600 7160
rect 10645 7040 10765 7160
rect 10810 7040 10930 7160
rect 10975 7040 11095 7160
rect 11150 7040 11270 7160
rect 11315 7040 11435 7160
rect 11480 7040 11600 7160
rect 11645 7040 11765 7160
rect 11820 7040 11940 7160
rect 11985 7040 12105 7160
rect 12150 7040 12270 7160
rect 12315 7040 12435 7160
rect 12490 7040 12610 7160
rect 7130 6865 7250 6985
rect 7295 6865 7415 6985
rect 7460 6865 7580 6985
rect 7625 6865 7745 6985
rect 7800 6865 7920 6985
rect 7965 6865 8085 6985
rect 8130 6865 8250 6985
rect 8295 6865 8415 6985
rect 8470 6865 8590 6985
rect 8635 6865 8755 6985
rect 8800 6865 8920 6985
rect 8965 6865 9085 6985
rect 9140 6865 9260 6985
rect 9305 6865 9425 6985
rect 9470 6865 9590 6985
rect 9635 6865 9755 6985
rect 9810 6865 9930 6985
rect 9975 6865 10095 6985
rect 10140 6865 10260 6985
rect 10305 6865 10425 6985
rect 10480 6865 10600 6985
rect 10645 6865 10765 6985
rect 10810 6865 10930 6985
rect 10975 6865 11095 6985
rect 11150 6865 11270 6985
rect 11315 6865 11435 6985
rect 11480 6865 11600 6985
rect 11645 6865 11765 6985
rect 11820 6865 11940 6985
rect 11985 6865 12105 6985
rect 12150 6865 12270 6985
rect 12315 6865 12435 6985
rect 12490 6865 12610 6985
rect 7130 6700 7250 6820
rect 7295 6700 7415 6820
rect 7460 6700 7580 6820
rect 7625 6700 7745 6820
rect 7800 6700 7920 6820
rect 7965 6700 8085 6820
rect 8130 6700 8250 6820
rect 8295 6700 8415 6820
rect 8470 6700 8590 6820
rect 8635 6700 8755 6820
rect 8800 6700 8920 6820
rect 8965 6700 9085 6820
rect 9140 6700 9260 6820
rect 9305 6700 9425 6820
rect 9470 6700 9590 6820
rect 9635 6700 9755 6820
rect 9810 6700 9930 6820
rect 9975 6700 10095 6820
rect 10140 6700 10260 6820
rect 10305 6700 10425 6820
rect 10480 6700 10600 6820
rect 10645 6700 10765 6820
rect 10810 6700 10930 6820
rect 10975 6700 11095 6820
rect 11150 6700 11270 6820
rect 11315 6700 11435 6820
rect 11480 6700 11600 6820
rect 11645 6700 11765 6820
rect 11820 6700 11940 6820
rect 11985 6700 12105 6820
rect 12150 6700 12270 6820
rect 12315 6700 12435 6820
rect 12490 6700 12610 6820
rect 7130 6535 7250 6655
rect 7295 6535 7415 6655
rect 7460 6535 7580 6655
rect 7625 6535 7745 6655
rect 7800 6535 7920 6655
rect 7965 6535 8085 6655
rect 8130 6535 8250 6655
rect 8295 6535 8415 6655
rect 8470 6535 8590 6655
rect 8635 6535 8755 6655
rect 8800 6535 8920 6655
rect 8965 6535 9085 6655
rect 9140 6535 9260 6655
rect 9305 6535 9425 6655
rect 9470 6535 9590 6655
rect 9635 6535 9755 6655
rect 9810 6535 9930 6655
rect 9975 6535 10095 6655
rect 10140 6535 10260 6655
rect 10305 6535 10425 6655
rect 10480 6535 10600 6655
rect 10645 6535 10765 6655
rect 10810 6535 10930 6655
rect 10975 6535 11095 6655
rect 11150 6535 11270 6655
rect 11315 6535 11435 6655
rect 11480 6535 11600 6655
rect 11645 6535 11765 6655
rect 11820 6535 11940 6655
rect 11985 6535 12105 6655
rect 12150 6535 12270 6655
rect 12315 6535 12435 6655
rect 12490 6535 12610 6655
rect 7130 6370 7250 6490
rect 7295 6370 7415 6490
rect 7460 6370 7580 6490
rect 7625 6370 7745 6490
rect 7800 6370 7920 6490
rect 7965 6370 8085 6490
rect 8130 6370 8250 6490
rect 8295 6370 8415 6490
rect 8470 6370 8590 6490
rect 8635 6370 8755 6490
rect 8800 6370 8920 6490
rect 8965 6370 9085 6490
rect 9140 6370 9260 6490
rect 9305 6370 9425 6490
rect 9470 6370 9590 6490
rect 9635 6370 9755 6490
rect 9810 6370 9930 6490
rect 9975 6370 10095 6490
rect 10140 6370 10260 6490
rect 10305 6370 10425 6490
rect 10480 6370 10600 6490
rect 10645 6370 10765 6490
rect 10810 6370 10930 6490
rect 10975 6370 11095 6490
rect 11150 6370 11270 6490
rect 11315 6370 11435 6490
rect 11480 6370 11600 6490
rect 11645 6370 11765 6490
rect 11820 6370 11940 6490
rect 11985 6370 12105 6490
rect 12150 6370 12270 6490
rect 12315 6370 12435 6490
rect 12490 6370 12610 6490
rect 7130 6195 7250 6315
rect 7295 6195 7415 6315
rect 7460 6195 7580 6315
rect 7625 6195 7745 6315
rect 7800 6195 7920 6315
rect 7965 6195 8085 6315
rect 8130 6195 8250 6315
rect 8295 6195 8415 6315
rect 8470 6195 8590 6315
rect 8635 6195 8755 6315
rect 8800 6195 8920 6315
rect 8965 6195 9085 6315
rect 9140 6195 9260 6315
rect 9305 6195 9425 6315
rect 9470 6195 9590 6315
rect 9635 6195 9755 6315
rect 9810 6195 9930 6315
rect 9975 6195 10095 6315
rect 10140 6195 10260 6315
rect 10305 6195 10425 6315
rect 10480 6195 10600 6315
rect 10645 6195 10765 6315
rect 10810 6195 10930 6315
rect 10975 6195 11095 6315
rect 11150 6195 11270 6315
rect 11315 6195 11435 6315
rect 11480 6195 11600 6315
rect 11645 6195 11765 6315
rect 11820 6195 11940 6315
rect 11985 6195 12105 6315
rect 12150 6195 12270 6315
rect 12315 6195 12435 6315
rect 12490 6195 12610 6315
rect 7130 6030 7250 6150
rect 7295 6030 7415 6150
rect 7460 6030 7580 6150
rect 7625 6030 7745 6150
rect 7800 6030 7920 6150
rect 7965 6030 8085 6150
rect 8130 6030 8250 6150
rect 8295 6030 8415 6150
rect 8470 6030 8590 6150
rect 8635 6030 8755 6150
rect 8800 6030 8920 6150
rect 8965 6030 9085 6150
rect 9140 6030 9260 6150
rect 9305 6030 9425 6150
rect 9470 6030 9590 6150
rect 9635 6030 9755 6150
rect 9810 6030 9930 6150
rect 9975 6030 10095 6150
rect 10140 6030 10260 6150
rect 10305 6030 10425 6150
rect 10480 6030 10600 6150
rect 10645 6030 10765 6150
rect 10810 6030 10930 6150
rect 10975 6030 11095 6150
rect 11150 6030 11270 6150
rect 11315 6030 11435 6150
rect 11480 6030 11600 6150
rect 11645 6030 11765 6150
rect 11820 6030 11940 6150
rect 11985 6030 12105 6150
rect 12150 6030 12270 6150
rect 12315 6030 12435 6150
rect 12490 6030 12610 6150
rect 7130 5865 7250 5985
rect 7295 5865 7415 5985
rect 7460 5865 7580 5985
rect 7625 5865 7745 5985
rect 7800 5865 7920 5985
rect 7965 5865 8085 5985
rect 8130 5865 8250 5985
rect 8295 5865 8415 5985
rect 8470 5865 8590 5985
rect 8635 5865 8755 5985
rect 8800 5865 8920 5985
rect 8965 5865 9085 5985
rect 9140 5865 9260 5985
rect 9305 5865 9425 5985
rect 9470 5865 9590 5985
rect 9635 5865 9755 5985
rect 9810 5865 9930 5985
rect 9975 5865 10095 5985
rect 10140 5865 10260 5985
rect 10305 5865 10425 5985
rect 10480 5865 10600 5985
rect 10645 5865 10765 5985
rect 10810 5865 10930 5985
rect 10975 5865 11095 5985
rect 11150 5865 11270 5985
rect 11315 5865 11435 5985
rect 11480 5865 11600 5985
rect 11645 5865 11765 5985
rect 11820 5865 11940 5985
rect 11985 5865 12105 5985
rect 12150 5865 12270 5985
rect 12315 5865 12435 5985
rect 12490 5865 12610 5985
rect 7130 5700 7250 5820
rect 7295 5700 7415 5820
rect 7460 5700 7580 5820
rect 7625 5700 7745 5820
rect 7800 5700 7920 5820
rect 7965 5700 8085 5820
rect 8130 5700 8250 5820
rect 8295 5700 8415 5820
rect 8470 5700 8590 5820
rect 8635 5700 8755 5820
rect 8800 5700 8920 5820
rect 8965 5700 9085 5820
rect 9140 5700 9260 5820
rect 9305 5700 9425 5820
rect 9470 5700 9590 5820
rect 9635 5700 9755 5820
rect 9810 5700 9930 5820
rect 9975 5700 10095 5820
rect 10140 5700 10260 5820
rect 10305 5700 10425 5820
rect 10480 5700 10600 5820
rect 10645 5700 10765 5820
rect 10810 5700 10930 5820
rect 10975 5700 11095 5820
rect 11150 5700 11270 5820
rect 11315 5700 11435 5820
rect 11480 5700 11600 5820
rect 11645 5700 11765 5820
rect 11820 5700 11940 5820
rect 11985 5700 12105 5820
rect 12150 5700 12270 5820
rect 12315 5700 12435 5820
rect 12490 5700 12610 5820
rect 7130 5525 7250 5645
rect 7295 5525 7415 5645
rect 7460 5525 7580 5645
rect 7625 5525 7745 5645
rect 7800 5525 7920 5645
rect 7965 5525 8085 5645
rect 8130 5525 8250 5645
rect 8295 5525 8415 5645
rect 8470 5525 8590 5645
rect 8635 5525 8755 5645
rect 8800 5525 8920 5645
rect 8965 5525 9085 5645
rect 9140 5525 9260 5645
rect 9305 5525 9425 5645
rect 9470 5525 9590 5645
rect 9635 5525 9755 5645
rect 9810 5525 9930 5645
rect 9975 5525 10095 5645
rect 10140 5525 10260 5645
rect 10305 5525 10425 5645
rect 10480 5525 10600 5645
rect 10645 5525 10765 5645
rect 10810 5525 10930 5645
rect 10975 5525 11095 5645
rect 11150 5525 11270 5645
rect 11315 5525 11435 5645
rect 11480 5525 11600 5645
rect 11645 5525 11765 5645
rect 11820 5525 11940 5645
rect 11985 5525 12105 5645
rect 12150 5525 12270 5645
rect 12315 5525 12435 5645
rect 12490 5525 12610 5645
rect 7130 5360 7250 5480
rect 7295 5360 7415 5480
rect 7460 5360 7580 5480
rect 7625 5360 7745 5480
rect 7800 5360 7920 5480
rect 7965 5360 8085 5480
rect 8130 5360 8250 5480
rect 8295 5360 8415 5480
rect 8470 5360 8590 5480
rect 8635 5360 8755 5480
rect 8800 5360 8920 5480
rect 8965 5360 9085 5480
rect 9140 5360 9260 5480
rect 9305 5360 9425 5480
rect 9470 5360 9590 5480
rect 9635 5360 9755 5480
rect 9810 5360 9930 5480
rect 9975 5360 10095 5480
rect 10140 5360 10260 5480
rect 10305 5360 10425 5480
rect 10480 5360 10600 5480
rect 10645 5360 10765 5480
rect 10810 5360 10930 5480
rect 10975 5360 11095 5480
rect 11150 5360 11270 5480
rect 11315 5360 11435 5480
rect 11480 5360 11600 5480
rect 11645 5360 11765 5480
rect 11820 5360 11940 5480
rect 11985 5360 12105 5480
rect 12150 5360 12270 5480
rect 12315 5360 12435 5480
rect 12490 5360 12610 5480
rect 7130 5195 7250 5315
rect 7295 5195 7415 5315
rect 7460 5195 7580 5315
rect 7625 5195 7745 5315
rect 7800 5195 7920 5315
rect 7965 5195 8085 5315
rect 8130 5195 8250 5315
rect 8295 5195 8415 5315
rect 8470 5195 8590 5315
rect 8635 5195 8755 5315
rect 8800 5195 8920 5315
rect 8965 5195 9085 5315
rect 9140 5195 9260 5315
rect 9305 5195 9425 5315
rect 9470 5195 9590 5315
rect 9635 5195 9755 5315
rect 9810 5195 9930 5315
rect 9975 5195 10095 5315
rect 10140 5195 10260 5315
rect 10305 5195 10425 5315
rect 10480 5195 10600 5315
rect 10645 5195 10765 5315
rect 10810 5195 10930 5315
rect 10975 5195 11095 5315
rect 11150 5195 11270 5315
rect 11315 5195 11435 5315
rect 11480 5195 11600 5315
rect 11645 5195 11765 5315
rect 11820 5195 11940 5315
rect 11985 5195 12105 5315
rect 12150 5195 12270 5315
rect 12315 5195 12435 5315
rect 12490 5195 12610 5315
rect 7130 5030 7250 5150
rect 7295 5030 7415 5150
rect 7460 5030 7580 5150
rect 7625 5030 7745 5150
rect 7800 5030 7920 5150
rect 7965 5030 8085 5150
rect 8130 5030 8250 5150
rect 8295 5030 8415 5150
rect 8470 5030 8590 5150
rect 8635 5030 8755 5150
rect 8800 5030 8920 5150
rect 8965 5030 9085 5150
rect 9140 5030 9260 5150
rect 9305 5030 9425 5150
rect 9470 5030 9590 5150
rect 9635 5030 9755 5150
rect 9810 5030 9930 5150
rect 9975 5030 10095 5150
rect 10140 5030 10260 5150
rect 10305 5030 10425 5150
rect 10480 5030 10600 5150
rect 10645 5030 10765 5150
rect 10810 5030 10930 5150
rect 10975 5030 11095 5150
rect 11150 5030 11270 5150
rect 11315 5030 11435 5150
rect 11480 5030 11600 5150
rect 11645 5030 11765 5150
rect 11820 5030 11940 5150
rect 11985 5030 12105 5150
rect 12150 5030 12270 5150
rect 12315 5030 12435 5150
rect 12490 5030 12610 5150
rect 7130 4855 7250 4975
rect 7295 4855 7415 4975
rect 7460 4855 7580 4975
rect 7625 4855 7745 4975
rect 7800 4855 7920 4975
rect 7965 4855 8085 4975
rect 8130 4855 8250 4975
rect 8295 4855 8415 4975
rect 8470 4855 8590 4975
rect 8635 4855 8755 4975
rect 8800 4855 8920 4975
rect 8965 4855 9085 4975
rect 9140 4855 9260 4975
rect 9305 4855 9425 4975
rect 9470 4855 9590 4975
rect 9635 4855 9755 4975
rect 9810 4855 9930 4975
rect 9975 4855 10095 4975
rect 10140 4855 10260 4975
rect 10305 4855 10425 4975
rect 10480 4855 10600 4975
rect 10645 4855 10765 4975
rect 10810 4855 10930 4975
rect 10975 4855 11095 4975
rect 11150 4855 11270 4975
rect 11315 4855 11435 4975
rect 11480 4855 11600 4975
rect 11645 4855 11765 4975
rect 11820 4855 11940 4975
rect 11985 4855 12105 4975
rect 12150 4855 12270 4975
rect 12315 4855 12435 4975
rect 12490 4855 12610 4975
rect 7130 4690 7250 4810
rect 7295 4690 7415 4810
rect 7460 4690 7580 4810
rect 7625 4690 7745 4810
rect 7800 4690 7920 4810
rect 7965 4690 8085 4810
rect 8130 4690 8250 4810
rect 8295 4690 8415 4810
rect 8470 4690 8590 4810
rect 8635 4690 8755 4810
rect 8800 4690 8920 4810
rect 8965 4690 9085 4810
rect 9140 4690 9260 4810
rect 9305 4690 9425 4810
rect 9470 4690 9590 4810
rect 9635 4690 9755 4810
rect 9810 4690 9930 4810
rect 9975 4690 10095 4810
rect 10140 4690 10260 4810
rect 10305 4690 10425 4810
rect 10480 4690 10600 4810
rect 10645 4690 10765 4810
rect 10810 4690 10930 4810
rect 10975 4690 11095 4810
rect 11150 4690 11270 4810
rect 11315 4690 11435 4810
rect 11480 4690 11600 4810
rect 11645 4690 11765 4810
rect 11820 4690 11940 4810
rect 11985 4690 12105 4810
rect 12150 4690 12270 4810
rect 12315 4690 12435 4810
rect 12490 4690 12610 4810
rect 7130 4525 7250 4645
rect 7295 4525 7415 4645
rect 7460 4525 7580 4645
rect 7625 4525 7745 4645
rect 7800 4525 7920 4645
rect 7965 4525 8085 4645
rect 8130 4525 8250 4645
rect 8295 4525 8415 4645
rect 8470 4525 8590 4645
rect 8635 4525 8755 4645
rect 8800 4525 8920 4645
rect 8965 4525 9085 4645
rect 9140 4525 9260 4645
rect 9305 4525 9425 4645
rect 9470 4525 9590 4645
rect 9635 4525 9755 4645
rect 9810 4525 9930 4645
rect 9975 4525 10095 4645
rect 10140 4525 10260 4645
rect 10305 4525 10425 4645
rect 10480 4525 10600 4645
rect 10645 4525 10765 4645
rect 10810 4525 10930 4645
rect 10975 4525 11095 4645
rect 11150 4525 11270 4645
rect 11315 4525 11435 4645
rect 11480 4525 11600 4645
rect 11645 4525 11765 4645
rect 11820 4525 11940 4645
rect 11985 4525 12105 4645
rect 12150 4525 12270 4645
rect 12315 4525 12435 4645
rect 12490 4525 12610 4645
rect 7130 4360 7250 4480
rect 7295 4360 7415 4480
rect 7460 4360 7580 4480
rect 7625 4360 7745 4480
rect 7800 4360 7920 4480
rect 7965 4360 8085 4480
rect 8130 4360 8250 4480
rect 8295 4360 8415 4480
rect 8470 4360 8590 4480
rect 8635 4360 8755 4480
rect 8800 4360 8920 4480
rect 8965 4360 9085 4480
rect 9140 4360 9260 4480
rect 9305 4360 9425 4480
rect 9470 4360 9590 4480
rect 9635 4360 9755 4480
rect 9810 4360 9930 4480
rect 9975 4360 10095 4480
rect 10140 4360 10260 4480
rect 10305 4360 10425 4480
rect 10480 4360 10600 4480
rect 10645 4360 10765 4480
rect 10810 4360 10930 4480
rect 10975 4360 11095 4480
rect 11150 4360 11270 4480
rect 11315 4360 11435 4480
rect 11480 4360 11600 4480
rect 11645 4360 11765 4480
rect 11820 4360 11940 4480
rect 11985 4360 12105 4480
rect 12150 4360 12270 4480
rect 12315 4360 12435 4480
rect 12490 4360 12610 4480
rect 7130 4185 7250 4305
rect 7295 4185 7415 4305
rect 7460 4185 7580 4305
rect 7625 4185 7745 4305
rect 7800 4185 7920 4305
rect 7965 4185 8085 4305
rect 8130 4185 8250 4305
rect 8295 4185 8415 4305
rect 8470 4185 8590 4305
rect 8635 4185 8755 4305
rect 8800 4185 8920 4305
rect 8965 4185 9085 4305
rect 9140 4185 9260 4305
rect 9305 4185 9425 4305
rect 9470 4185 9590 4305
rect 9635 4185 9755 4305
rect 9810 4185 9930 4305
rect 9975 4185 10095 4305
rect 10140 4185 10260 4305
rect 10305 4185 10425 4305
rect 10480 4185 10600 4305
rect 10645 4185 10765 4305
rect 10810 4185 10930 4305
rect 10975 4185 11095 4305
rect 11150 4185 11270 4305
rect 11315 4185 11435 4305
rect 11480 4185 11600 4305
rect 11645 4185 11765 4305
rect 11820 4185 11940 4305
rect 11985 4185 12105 4305
rect 12150 4185 12270 4305
rect 12315 4185 12435 4305
rect 12490 4185 12610 4305
rect 7130 4020 7250 4140
rect 7295 4020 7415 4140
rect 7460 4020 7580 4140
rect 7625 4020 7745 4140
rect 7800 4020 7920 4140
rect 7965 4020 8085 4140
rect 8130 4020 8250 4140
rect 8295 4020 8415 4140
rect 8470 4020 8590 4140
rect 8635 4020 8755 4140
rect 8800 4020 8920 4140
rect 8965 4020 9085 4140
rect 9140 4020 9260 4140
rect 9305 4020 9425 4140
rect 9470 4020 9590 4140
rect 9635 4020 9755 4140
rect 9810 4020 9930 4140
rect 9975 4020 10095 4140
rect 10140 4020 10260 4140
rect 10305 4020 10425 4140
rect 10480 4020 10600 4140
rect 10645 4020 10765 4140
rect 10810 4020 10930 4140
rect 10975 4020 11095 4140
rect 11150 4020 11270 4140
rect 11315 4020 11435 4140
rect 11480 4020 11600 4140
rect 11645 4020 11765 4140
rect 11820 4020 11940 4140
rect 11985 4020 12105 4140
rect 12150 4020 12270 4140
rect 12315 4020 12435 4140
rect 12490 4020 12610 4140
rect 7130 3855 7250 3975
rect 7295 3855 7415 3975
rect 7460 3855 7580 3975
rect 7625 3855 7745 3975
rect 7800 3855 7920 3975
rect 7965 3855 8085 3975
rect 8130 3855 8250 3975
rect 8295 3855 8415 3975
rect 8470 3855 8590 3975
rect 8635 3855 8755 3975
rect 8800 3855 8920 3975
rect 8965 3855 9085 3975
rect 9140 3855 9260 3975
rect 9305 3855 9425 3975
rect 9470 3855 9590 3975
rect 9635 3855 9755 3975
rect 9810 3855 9930 3975
rect 9975 3855 10095 3975
rect 10140 3855 10260 3975
rect 10305 3855 10425 3975
rect 10480 3855 10600 3975
rect 10645 3855 10765 3975
rect 10810 3855 10930 3975
rect 10975 3855 11095 3975
rect 11150 3855 11270 3975
rect 11315 3855 11435 3975
rect 11480 3855 11600 3975
rect 11645 3855 11765 3975
rect 11820 3855 11940 3975
rect 11985 3855 12105 3975
rect 12150 3855 12270 3975
rect 12315 3855 12435 3975
rect 12490 3855 12610 3975
rect 7130 3690 7250 3810
rect 7295 3690 7415 3810
rect 7460 3690 7580 3810
rect 7625 3690 7745 3810
rect 7800 3690 7920 3810
rect 7965 3690 8085 3810
rect 8130 3690 8250 3810
rect 8295 3690 8415 3810
rect 8470 3690 8590 3810
rect 8635 3690 8755 3810
rect 8800 3690 8920 3810
rect 8965 3690 9085 3810
rect 9140 3690 9260 3810
rect 9305 3690 9425 3810
rect 9470 3690 9590 3810
rect 9635 3690 9755 3810
rect 9810 3690 9930 3810
rect 9975 3690 10095 3810
rect 10140 3690 10260 3810
rect 10305 3690 10425 3810
rect 10480 3690 10600 3810
rect 10645 3690 10765 3810
rect 10810 3690 10930 3810
rect 10975 3690 11095 3810
rect 11150 3690 11270 3810
rect 11315 3690 11435 3810
rect 11480 3690 11600 3810
rect 11645 3690 11765 3810
rect 11820 3690 11940 3810
rect 11985 3690 12105 3810
rect 12150 3690 12270 3810
rect 12315 3690 12435 3810
rect 12490 3690 12610 3810
rect 7130 3515 7250 3635
rect 7295 3515 7415 3635
rect 7460 3515 7580 3635
rect 7625 3515 7745 3635
rect 7800 3515 7920 3635
rect 7965 3515 8085 3635
rect 8130 3515 8250 3635
rect 8295 3515 8415 3635
rect 8470 3515 8590 3635
rect 8635 3515 8755 3635
rect 8800 3515 8920 3635
rect 8965 3515 9085 3635
rect 9140 3515 9260 3635
rect 9305 3515 9425 3635
rect 9470 3515 9590 3635
rect 9635 3515 9755 3635
rect 9810 3515 9930 3635
rect 9975 3515 10095 3635
rect 10140 3515 10260 3635
rect 10305 3515 10425 3635
rect 10480 3515 10600 3635
rect 10645 3515 10765 3635
rect 10810 3515 10930 3635
rect 10975 3515 11095 3635
rect 11150 3515 11270 3635
rect 11315 3515 11435 3635
rect 11480 3515 11600 3635
rect 11645 3515 11765 3635
rect 11820 3515 11940 3635
rect 11985 3515 12105 3635
rect 12150 3515 12270 3635
rect 12315 3515 12435 3635
rect 12490 3515 12610 3635
rect 7130 3350 7250 3470
rect 7295 3350 7415 3470
rect 7460 3350 7580 3470
rect 7625 3350 7745 3470
rect 7800 3350 7920 3470
rect 7965 3350 8085 3470
rect 8130 3350 8250 3470
rect 8295 3350 8415 3470
rect 8470 3350 8590 3470
rect 8635 3350 8755 3470
rect 8800 3350 8920 3470
rect 8965 3350 9085 3470
rect 9140 3350 9260 3470
rect 9305 3350 9425 3470
rect 9470 3350 9590 3470
rect 9635 3350 9755 3470
rect 9810 3350 9930 3470
rect 9975 3350 10095 3470
rect 10140 3350 10260 3470
rect 10305 3350 10425 3470
rect 10480 3350 10600 3470
rect 10645 3350 10765 3470
rect 10810 3350 10930 3470
rect 10975 3350 11095 3470
rect 11150 3350 11270 3470
rect 11315 3350 11435 3470
rect 11480 3350 11600 3470
rect 11645 3350 11765 3470
rect 11820 3350 11940 3470
rect 11985 3350 12105 3470
rect 12150 3350 12270 3470
rect 12315 3350 12435 3470
rect 12490 3350 12610 3470
rect 7130 3185 7250 3305
rect 7295 3185 7415 3305
rect 7460 3185 7580 3305
rect 7625 3185 7745 3305
rect 7800 3185 7920 3305
rect 7965 3185 8085 3305
rect 8130 3185 8250 3305
rect 8295 3185 8415 3305
rect 8470 3185 8590 3305
rect 8635 3185 8755 3305
rect 8800 3185 8920 3305
rect 8965 3185 9085 3305
rect 9140 3185 9260 3305
rect 9305 3185 9425 3305
rect 9470 3185 9590 3305
rect 9635 3185 9755 3305
rect 9810 3185 9930 3305
rect 9975 3185 10095 3305
rect 10140 3185 10260 3305
rect 10305 3185 10425 3305
rect 10480 3185 10600 3305
rect 10645 3185 10765 3305
rect 10810 3185 10930 3305
rect 10975 3185 11095 3305
rect 11150 3185 11270 3305
rect 11315 3185 11435 3305
rect 11480 3185 11600 3305
rect 11645 3185 11765 3305
rect 11820 3185 11940 3305
rect 11985 3185 12105 3305
rect 12150 3185 12270 3305
rect 12315 3185 12435 3305
rect 12490 3185 12610 3305
rect 7130 3020 7250 3140
rect 7295 3020 7415 3140
rect 7460 3020 7580 3140
rect 7625 3020 7745 3140
rect 7800 3020 7920 3140
rect 7965 3020 8085 3140
rect 8130 3020 8250 3140
rect 8295 3020 8415 3140
rect 8470 3020 8590 3140
rect 8635 3020 8755 3140
rect 8800 3020 8920 3140
rect 8965 3020 9085 3140
rect 9140 3020 9260 3140
rect 9305 3020 9425 3140
rect 9470 3020 9590 3140
rect 9635 3020 9755 3140
rect 9810 3020 9930 3140
rect 9975 3020 10095 3140
rect 10140 3020 10260 3140
rect 10305 3020 10425 3140
rect 10480 3020 10600 3140
rect 10645 3020 10765 3140
rect 10810 3020 10930 3140
rect 10975 3020 11095 3140
rect 11150 3020 11270 3140
rect 11315 3020 11435 3140
rect 11480 3020 11600 3140
rect 11645 3020 11765 3140
rect 11820 3020 11940 3140
rect 11985 3020 12105 3140
rect 12150 3020 12270 3140
rect 12315 3020 12435 3140
rect 12490 3020 12610 3140
rect 7130 2845 7250 2965
rect 7295 2845 7415 2965
rect 7460 2845 7580 2965
rect 7625 2845 7745 2965
rect 7800 2845 7920 2965
rect 7965 2845 8085 2965
rect 8130 2845 8250 2965
rect 8295 2845 8415 2965
rect 8470 2845 8590 2965
rect 8635 2845 8755 2965
rect 8800 2845 8920 2965
rect 8965 2845 9085 2965
rect 9140 2845 9260 2965
rect 9305 2845 9425 2965
rect 9470 2845 9590 2965
rect 9635 2845 9755 2965
rect 9810 2845 9930 2965
rect 9975 2845 10095 2965
rect 10140 2845 10260 2965
rect 10305 2845 10425 2965
rect 10480 2845 10600 2965
rect 10645 2845 10765 2965
rect 10810 2845 10930 2965
rect 10975 2845 11095 2965
rect 11150 2845 11270 2965
rect 11315 2845 11435 2965
rect 11480 2845 11600 2965
rect 11645 2845 11765 2965
rect 11820 2845 11940 2965
rect 11985 2845 12105 2965
rect 12150 2845 12270 2965
rect 12315 2845 12435 2965
rect 12490 2845 12610 2965
rect 7130 2680 7250 2800
rect 7295 2680 7415 2800
rect 7460 2680 7580 2800
rect 7625 2680 7745 2800
rect 7800 2680 7920 2800
rect 7965 2680 8085 2800
rect 8130 2680 8250 2800
rect 8295 2680 8415 2800
rect 8470 2680 8590 2800
rect 8635 2680 8755 2800
rect 8800 2680 8920 2800
rect 8965 2680 9085 2800
rect 9140 2680 9260 2800
rect 9305 2680 9425 2800
rect 9470 2680 9590 2800
rect 9635 2680 9755 2800
rect 9810 2680 9930 2800
rect 9975 2680 10095 2800
rect 10140 2680 10260 2800
rect 10305 2680 10425 2800
rect 10480 2680 10600 2800
rect 10645 2680 10765 2800
rect 10810 2680 10930 2800
rect 10975 2680 11095 2800
rect 11150 2680 11270 2800
rect 11315 2680 11435 2800
rect 11480 2680 11600 2800
rect 11645 2680 11765 2800
rect 11820 2680 11940 2800
rect 11985 2680 12105 2800
rect 12150 2680 12270 2800
rect 12315 2680 12435 2800
rect 12490 2680 12610 2800
rect 7130 2515 7250 2635
rect 7295 2515 7415 2635
rect 7460 2515 7580 2635
rect 7625 2515 7745 2635
rect 7800 2515 7920 2635
rect 7965 2515 8085 2635
rect 8130 2515 8250 2635
rect 8295 2515 8415 2635
rect 8470 2515 8590 2635
rect 8635 2515 8755 2635
rect 8800 2515 8920 2635
rect 8965 2515 9085 2635
rect 9140 2515 9260 2635
rect 9305 2515 9425 2635
rect 9470 2515 9590 2635
rect 9635 2515 9755 2635
rect 9810 2515 9930 2635
rect 9975 2515 10095 2635
rect 10140 2515 10260 2635
rect 10305 2515 10425 2635
rect 10480 2515 10600 2635
rect 10645 2515 10765 2635
rect 10810 2515 10930 2635
rect 10975 2515 11095 2635
rect 11150 2515 11270 2635
rect 11315 2515 11435 2635
rect 11480 2515 11600 2635
rect 11645 2515 11765 2635
rect 11820 2515 11940 2635
rect 11985 2515 12105 2635
rect 12150 2515 12270 2635
rect 12315 2515 12435 2635
rect 12490 2515 12610 2635
rect 7130 2350 7250 2470
rect 7295 2350 7415 2470
rect 7460 2350 7580 2470
rect 7625 2350 7745 2470
rect 7800 2350 7920 2470
rect 7965 2350 8085 2470
rect 8130 2350 8250 2470
rect 8295 2350 8415 2470
rect 8470 2350 8590 2470
rect 8635 2350 8755 2470
rect 8800 2350 8920 2470
rect 8965 2350 9085 2470
rect 9140 2350 9260 2470
rect 9305 2350 9425 2470
rect 9470 2350 9590 2470
rect 9635 2350 9755 2470
rect 9810 2350 9930 2470
rect 9975 2350 10095 2470
rect 10140 2350 10260 2470
rect 10305 2350 10425 2470
rect 10480 2350 10600 2470
rect 10645 2350 10765 2470
rect 10810 2350 10930 2470
rect 10975 2350 11095 2470
rect 11150 2350 11270 2470
rect 11315 2350 11435 2470
rect 11480 2350 11600 2470
rect 11645 2350 11765 2470
rect 11820 2350 11940 2470
rect 11985 2350 12105 2470
rect 12150 2350 12270 2470
rect 12315 2350 12435 2470
rect 12490 2350 12610 2470
rect 7130 2175 7250 2295
rect 7295 2175 7415 2295
rect 7460 2175 7580 2295
rect 7625 2175 7745 2295
rect 7800 2175 7920 2295
rect 7965 2175 8085 2295
rect 8130 2175 8250 2295
rect 8295 2175 8415 2295
rect 8470 2175 8590 2295
rect 8635 2175 8755 2295
rect 8800 2175 8920 2295
rect 8965 2175 9085 2295
rect 9140 2175 9260 2295
rect 9305 2175 9425 2295
rect 9470 2175 9590 2295
rect 9635 2175 9755 2295
rect 9810 2175 9930 2295
rect 9975 2175 10095 2295
rect 10140 2175 10260 2295
rect 10305 2175 10425 2295
rect 10480 2175 10600 2295
rect 10645 2175 10765 2295
rect 10810 2175 10930 2295
rect 10975 2175 11095 2295
rect 11150 2175 11270 2295
rect 11315 2175 11435 2295
rect 11480 2175 11600 2295
rect 11645 2175 11765 2295
rect 11820 2175 11940 2295
rect 11985 2175 12105 2295
rect 12150 2175 12270 2295
rect 12315 2175 12435 2295
rect 12490 2175 12610 2295
rect 7130 2010 7250 2130
rect 7295 2010 7415 2130
rect 7460 2010 7580 2130
rect 7625 2010 7745 2130
rect 7800 2010 7920 2130
rect 7965 2010 8085 2130
rect 8130 2010 8250 2130
rect 8295 2010 8415 2130
rect 8470 2010 8590 2130
rect 8635 2010 8755 2130
rect 8800 2010 8920 2130
rect 8965 2010 9085 2130
rect 9140 2010 9260 2130
rect 9305 2010 9425 2130
rect 9470 2010 9590 2130
rect 9635 2010 9755 2130
rect 9810 2010 9930 2130
rect 9975 2010 10095 2130
rect 10140 2010 10260 2130
rect 10305 2010 10425 2130
rect 10480 2010 10600 2130
rect 10645 2010 10765 2130
rect 10810 2010 10930 2130
rect 10975 2010 11095 2130
rect 11150 2010 11270 2130
rect 11315 2010 11435 2130
rect 11480 2010 11600 2130
rect 11645 2010 11765 2130
rect 11820 2010 11940 2130
rect 11985 2010 12105 2130
rect 12150 2010 12270 2130
rect 12315 2010 12435 2130
rect 12490 2010 12610 2130
rect 7130 1845 7250 1965
rect 7295 1845 7415 1965
rect 7460 1845 7580 1965
rect 7625 1845 7745 1965
rect 7800 1845 7920 1965
rect 7965 1845 8085 1965
rect 8130 1845 8250 1965
rect 8295 1845 8415 1965
rect 8470 1845 8590 1965
rect 8635 1845 8755 1965
rect 8800 1845 8920 1965
rect 8965 1845 9085 1965
rect 9140 1845 9260 1965
rect 9305 1845 9425 1965
rect 9470 1845 9590 1965
rect 9635 1845 9755 1965
rect 9810 1845 9930 1965
rect 9975 1845 10095 1965
rect 10140 1845 10260 1965
rect 10305 1845 10425 1965
rect 10480 1845 10600 1965
rect 10645 1845 10765 1965
rect 10810 1845 10930 1965
rect 10975 1845 11095 1965
rect 11150 1845 11270 1965
rect 11315 1845 11435 1965
rect 11480 1845 11600 1965
rect 11645 1845 11765 1965
rect 11820 1845 11940 1965
rect 11985 1845 12105 1965
rect 12150 1845 12270 1965
rect 12315 1845 12435 1965
rect 12490 1845 12610 1965
rect 7130 1680 7250 1800
rect 7295 1680 7415 1800
rect 7460 1680 7580 1800
rect 7625 1680 7745 1800
rect 7800 1680 7920 1800
rect 7965 1680 8085 1800
rect 8130 1680 8250 1800
rect 8295 1680 8415 1800
rect 8470 1680 8590 1800
rect 8635 1680 8755 1800
rect 8800 1680 8920 1800
rect 8965 1680 9085 1800
rect 9140 1680 9260 1800
rect 9305 1680 9425 1800
rect 9470 1680 9590 1800
rect 9635 1680 9755 1800
rect 9810 1680 9930 1800
rect 9975 1680 10095 1800
rect 10140 1680 10260 1800
rect 10305 1680 10425 1800
rect 10480 1680 10600 1800
rect 10645 1680 10765 1800
rect 10810 1680 10930 1800
rect 10975 1680 11095 1800
rect 11150 1680 11270 1800
rect 11315 1680 11435 1800
rect 11480 1680 11600 1800
rect 11645 1680 11765 1800
rect 11820 1680 11940 1800
rect 11985 1680 12105 1800
rect 12150 1680 12270 1800
rect 12315 1680 12435 1800
rect 12490 1680 12610 1800
rect 12820 7040 12940 7160
rect 12985 7040 13105 7160
rect 13150 7040 13270 7160
rect 13315 7040 13435 7160
rect 13490 7040 13610 7160
rect 13655 7040 13775 7160
rect 13820 7040 13940 7160
rect 13985 7040 14105 7160
rect 14160 7040 14280 7160
rect 14325 7040 14445 7160
rect 14490 7040 14610 7160
rect 14655 7040 14775 7160
rect 14830 7040 14950 7160
rect 14995 7040 15115 7160
rect 15160 7040 15280 7160
rect 15325 7040 15445 7160
rect 15500 7040 15620 7160
rect 15665 7040 15785 7160
rect 15830 7040 15950 7160
rect 15995 7040 16115 7160
rect 16170 7040 16290 7160
rect 16335 7040 16455 7160
rect 16500 7040 16620 7160
rect 16665 7040 16785 7160
rect 16840 7040 16960 7160
rect 17005 7040 17125 7160
rect 17170 7040 17290 7160
rect 17335 7040 17455 7160
rect 17510 7040 17630 7160
rect 17675 7040 17795 7160
rect 17840 7040 17960 7160
rect 18005 7040 18125 7160
rect 18180 7040 18300 7160
rect 12820 6865 12940 6985
rect 12985 6865 13105 6985
rect 13150 6865 13270 6985
rect 13315 6865 13435 6985
rect 13490 6865 13610 6985
rect 13655 6865 13775 6985
rect 13820 6865 13940 6985
rect 13985 6865 14105 6985
rect 14160 6865 14280 6985
rect 14325 6865 14445 6985
rect 14490 6865 14610 6985
rect 14655 6865 14775 6985
rect 14830 6865 14950 6985
rect 14995 6865 15115 6985
rect 15160 6865 15280 6985
rect 15325 6865 15445 6985
rect 15500 6865 15620 6985
rect 15665 6865 15785 6985
rect 15830 6865 15950 6985
rect 15995 6865 16115 6985
rect 16170 6865 16290 6985
rect 16335 6865 16455 6985
rect 16500 6865 16620 6985
rect 16665 6865 16785 6985
rect 16840 6865 16960 6985
rect 17005 6865 17125 6985
rect 17170 6865 17290 6985
rect 17335 6865 17455 6985
rect 17510 6865 17630 6985
rect 17675 6865 17795 6985
rect 17840 6865 17960 6985
rect 18005 6865 18125 6985
rect 18180 6865 18300 6985
rect 12820 6700 12940 6820
rect 12985 6700 13105 6820
rect 13150 6700 13270 6820
rect 13315 6700 13435 6820
rect 13490 6700 13610 6820
rect 13655 6700 13775 6820
rect 13820 6700 13940 6820
rect 13985 6700 14105 6820
rect 14160 6700 14280 6820
rect 14325 6700 14445 6820
rect 14490 6700 14610 6820
rect 14655 6700 14775 6820
rect 14830 6700 14950 6820
rect 14995 6700 15115 6820
rect 15160 6700 15280 6820
rect 15325 6700 15445 6820
rect 15500 6700 15620 6820
rect 15665 6700 15785 6820
rect 15830 6700 15950 6820
rect 15995 6700 16115 6820
rect 16170 6700 16290 6820
rect 16335 6700 16455 6820
rect 16500 6700 16620 6820
rect 16665 6700 16785 6820
rect 16840 6700 16960 6820
rect 17005 6700 17125 6820
rect 17170 6700 17290 6820
rect 17335 6700 17455 6820
rect 17510 6700 17630 6820
rect 17675 6700 17795 6820
rect 17840 6700 17960 6820
rect 18005 6700 18125 6820
rect 18180 6700 18300 6820
rect 12820 6535 12940 6655
rect 12985 6535 13105 6655
rect 13150 6535 13270 6655
rect 13315 6535 13435 6655
rect 13490 6535 13610 6655
rect 13655 6535 13775 6655
rect 13820 6535 13940 6655
rect 13985 6535 14105 6655
rect 14160 6535 14280 6655
rect 14325 6535 14445 6655
rect 14490 6535 14610 6655
rect 14655 6535 14775 6655
rect 14830 6535 14950 6655
rect 14995 6535 15115 6655
rect 15160 6535 15280 6655
rect 15325 6535 15445 6655
rect 15500 6535 15620 6655
rect 15665 6535 15785 6655
rect 15830 6535 15950 6655
rect 15995 6535 16115 6655
rect 16170 6535 16290 6655
rect 16335 6535 16455 6655
rect 16500 6535 16620 6655
rect 16665 6535 16785 6655
rect 16840 6535 16960 6655
rect 17005 6535 17125 6655
rect 17170 6535 17290 6655
rect 17335 6535 17455 6655
rect 17510 6535 17630 6655
rect 17675 6535 17795 6655
rect 17840 6535 17960 6655
rect 18005 6535 18125 6655
rect 18180 6535 18300 6655
rect 12820 6370 12940 6490
rect 12985 6370 13105 6490
rect 13150 6370 13270 6490
rect 13315 6370 13435 6490
rect 13490 6370 13610 6490
rect 13655 6370 13775 6490
rect 13820 6370 13940 6490
rect 13985 6370 14105 6490
rect 14160 6370 14280 6490
rect 14325 6370 14445 6490
rect 14490 6370 14610 6490
rect 14655 6370 14775 6490
rect 14830 6370 14950 6490
rect 14995 6370 15115 6490
rect 15160 6370 15280 6490
rect 15325 6370 15445 6490
rect 15500 6370 15620 6490
rect 15665 6370 15785 6490
rect 15830 6370 15950 6490
rect 15995 6370 16115 6490
rect 16170 6370 16290 6490
rect 16335 6370 16455 6490
rect 16500 6370 16620 6490
rect 16665 6370 16785 6490
rect 16840 6370 16960 6490
rect 17005 6370 17125 6490
rect 17170 6370 17290 6490
rect 17335 6370 17455 6490
rect 17510 6370 17630 6490
rect 17675 6370 17795 6490
rect 17840 6370 17960 6490
rect 18005 6370 18125 6490
rect 18180 6370 18300 6490
rect 12820 6195 12940 6315
rect 12985 6195 13105 6315
rect 13150 6195 13270 6315
rect 13315 6195 13435 6315
rect 13490 6195 13610 6315
rect 13655 6195 13775 6315
rect 13820 6195 13940 6315
rect 13985 6195 14105 6315
rect 14160 6195 14280 6315
rect 14325 6195 14445 6315
rect 14490 6195 14610 6315
rect 14655 6195 14775 6315
rect 14830 6195 14950 6315
rect 14995 6195 15115 6315
rect 15160 6195 15280 6315
rect 15325 6195 15445 6315
rect 15500 6195 15620 6315
rect 15665 6195 15785 6315
rect 15830 6195 15950 6315
rect 15995 6195 16115 6315
rect 16170 6195 16290 6315
rect 16335 6195 16455 6315
rect 16500 6195 16620 6315
rect 16665 6195 16785 6315
rect 16840 6195 16960 6315
rect 17005 6195 17125 6315
rect 17170 6195 17290 6315
rect 17335 6195 17455 6315
rect 17510 6195 17630 6315
rect 17675 6195 17795 6315
rect 17840 6195 17960 6315
rect 18005 6195 18125 6315
rect 18180 6195 18300 6315
rect 12820 6030 12940 6150
rect 12985 6030 13105 6150
rect 13150 6030 13270 6150
rect 13315 6030 13435 6150
rect 13490 6030 13610 6150
rect 13655 6030 13775 6150
rect 13820 6030 13940 6150
rect 13985 6030 14105 6150
rect 14160 6030 14280 6150
rect 14325 6030 14445 6150
rect 14490 6030 14610 6150
rect 14655 6030 14775 6150
rect 14830 6030 14950 6150
rect 14995 6030 15115 6150
rect 15160 6030 15280 6150
rect 15325 6030 15445 6150
rect 15500 6030 15620 6150
rect 15665 6030 15785 6150
rect 15830 6030 15950 6150
rect 15995 6030 16115 6150
rect 16170 6030 16290 6150
rect 16335 6030 16455 6150
rect 16500 6030 16620 6150
rect 16665 6030 16785 6150
rect 16840 6030 16960 6150
rect 17005 6030 17125 6150
rect 17170 6030 17290 6150
rect 17335 6030 17455 6150
rect 17510 6030 17630 6150
rect 17675 6030 17795 6150
rect 17840 6030 17960 6150
rect 18005 6030 18125 6150
rect 18180 6030 18300 6150
rect 12820 5865 12940 5985
rect 12985 5865 13105 5985
rect 13150 5865 13270 5985
rect 13315 5865 13435 5985
rect 13490 5865 13610 5985
rect 13655 5865 13775 5985
rect 13820 5865 13940 5985
rect 13985 5865 14105 5985
rect 14160 5865 14280 5985
rect 14325 5865 14445 5985
rect 14490 5865 14610 5985
rect 14655 5865 14775 5985
rect 14830 5865 14950 5985
rect 14995 5865 15115 5985
rect 15160 5865 15280 5985
rect 15325 5865 15445 5985
rect 15500 5865 15620 5985
rect 15665 5865 15785 5985
rect 15830 5865 15950 5985
rect 15995 5865 16115 5985
rect 16170 5865 16290 5985
rect 16335 5865 16455 5985
rect 16500 5865 16620 5985
rect 16665 5865 16785 5985
rect 16840 5865 16960 5985
rect 17005 5865 17125 5985
rect 17170 5865 17290 5985
rect 17335 5865 17455 5985
rect 17510 5865 17630 5985
rect 17675 5865 17795 5985
rect 17840 5865 17960 5985
rect 18005 5865 18125 5985
rect 18180 5865 18300 5985
rect 12820 5700 12940 5820
rect 12985 5700 13105 5820
rect 13150 5700 13270 5820
rect 13315 5700 13435 5820
rect 13490 5700 13610 5820
rect 13655 5700 13775 5820
rect 13820 5700 13940 5820
rect 13985 5700 14105 5820
rect 14160 5700 14280 5820
rect 14325 5700 14445 5820
rect 14490 5700 14610 5820
rect 14655 5700 14775 5820
rect 14830 5700 14950 5820
rect 14995 5700 15115 5820
rect 15160 5700 15280 5820
rect 15325 5700 15445 5820
rect 15500 5700 15620 5820
rect 15665 5700 15785 5820
rect 15830 5700 15950 5820
rect 15995 5700 16115 5820
rect 16170 5700 16290 5820
rect 16335 5700 16455 5820
rect 16500 5700 16620 5820
rect 16665 5700 16785 5820
rect 16840 5700 16960 5820
rect 17005 5700 17125 5820
rect 17170 5700 17290 5820
rect 17335 5700 17455 5820
rect 17510 5700 17630 5820
rect 17675 5700 17795 5820
rect 17840 5700 17960 5820
rect 18005 5700 18125 5820
rect 18180 5700 18300 5820
rect 12820 5525 12940 5645
rect 12985 5525 13105 5645
rect 13150 5525 13270 5645
rect 13315 5525 13435 5645
rect 13490 5525 13610 5645
rect 13655 5525 13775 5645
rect 13820 5525 13940 5645
rect 13985 5525 14105 5645
rect 14160 5525 14280 5645
rect 14325 5525 14445 5645
rect 14490 5525 14610 5645
rect 14655 5525 14775 5645
rect 14830 5525 14950 5645
rect 14995 5525 15115 5645
rect 15160 5525 15280 5645
rect 15325 5525 15445 5645
rect 15500 5525 15620 5645
rect 15665 5525 15785 5645
rect 15830 5525 15950 5645
rect 15995 5525 16115 5645
rect 16170 5525 16290 5645
rect 16335 5525 16455 5645
rect 16500 5525 16620 5645
rect 16665 5525 16785 5645
rect 16840 5525 16960 5645
rect 17005 5525 17125 5645
rect 17170 5525 17290 5645
rect 17335 5525 17455 5645
rect 17510 5525 17630 5645
rect 17675 5525 17795 5645
rect 17840 5525 17960 5645
rect 18005 5525 18125 5645
rect 18180 5525 18300 5645
rect 12820 5360 12940 5480
rect 12985 5360 13105 5480
rect 13150 5360 13270 5480
rect 13315 5360 13435 5480
rect 13490 5360 13610 5480
rect 13655 5360 13775 5480
rect 13820 5360 13940 5480
rect 13985 5360 14105 5480
rect 14160 5360 14280 5480
rect 14325 5360 14445 5480
rect 14490 5360 14610 5480
rect 14655 5360 14775 5480
rect 14830 5360 14950 5480
rect 14995 5360 15115 5480
rect 15160 5360 15280 5480
rect 15325 5360 15445 5480
rect 15500 5360 15620 5480
rect 15665 5360 15785 5480
rect 15830 5360 15950 5480
rect 15995 5360 16115 5480
rect 16170 5360 16290 5480
rect 16335 5360 16455 5480
rect 16500 5360 16620 5480
rect 16665 5360 16785 5480
rect 16840 5360 16960 5480
rect 17005 5360 17125 5480
rect 17170 5360 17290 5480
rect 17335 5360 17455 5480
rect 17510 5360 17630 5480
rect 17675 5360 17795 5480
rect 17840 5360 17960 5480
rect 18005 5360 18125 5480
rect 18180 5360 18300 5480
rect 12820 5195 12940 5315
rect 12985 5195 13105 5315
rect 13150 5195 13270 5315
rect 13315 5195 13435 5315
rect 13490 5195 13610 5315
rect 13655 5195 13775 5315
rect 13820 5195 13940 5315
rect 13985 5195 14105 5315
rect 14160 5195 14280 5315
rect 14325 5195 14445 5315
rect 14490 5195 14610 5315
rect 14655 5195 14775 5315
rect 14830 5195 14950 5315
rect 14995 5195 15115 5315
rect 15160 5195 15280 5315
rect 15325 5195 15445 5315
rect 15500 5195 15620 5315
rect 15665 5195 15785 5315
rect 15830 5195 15950 5315
rect 15995 5195 16115 5315
rect 16170 5195 16290 5315
rect 16335 5195 16455 5315
rect 16500 5195 16620 5315
rect 16665 5195 16785 5315
rect 16840 5195 16960 5315
rect 17005 5195 17125 5315
rect 17170 5195 17290 5315
rect 17335 5195 17455 5315
rect 17510 5195 17630 5315
rect 17675 5195 17795 5315
rect 17840 5195 17960 5315
rect 18005 5195 18125 5315
rect 18180 5195 18300 5315
rect 12820 5030 12940 5150
rect 12985 5030 13105 5150
rect 13150 5030 13270 5150
rect 13315 5030 13435 5150
rect 13490 5030 13610 5150
rect 13655 5030 13775 5150
rect 13820 5030 13940 5150
rect 13985 5030 14105 5150
rect 14160 5030 14280 5150
rect 14325 5030 14445 5150
rect 14490 5030 14610 5150
rect 14655 5030 14775 5150
rect 14830 5030 14950 5150
rect 14995 5030 15115 5150
rect 15160 5030 15280 5150
rect 15325 5030 15445 5150
rect 15500 5030 15620 5150
rect 15665 5030 15785 5150
rect 15830 5030 15950 5150
rect 15995 5030 16115 5150
rect 16170 5030 16290 5150
rect 16335 5030 16455 5150
rect 16500 5030 16620 5150
rect 16665 5030 16785 5150
rect 16840 5030 16960 5150
rect 17005 5030 17125 5150
rect 17170 5030 17290 5150
rect 17335 5030 17455 5150
rect 17510 5030 17630 5150
rect 17675 5030 17795 5150
rect 17840 5030 17960 5150
rect 18005 5030 18125 5150
rect 18180 5030 18300 5150
rect 12820 4855 12940 4975
rect 12985 4855 13105 4975
rect 13150 4855 13270 4975
rect 13315 4855 13435 4975
rect 13490 4855 13610 4975
rect 13655 4855 13775 4975
rect 13820 4855 13940 4975
rect 13985 4855 14105 4975
rect 14160 4855 14280 4975
rect 14325 4855 14445 4975
rect 14490 4855 14610 4975
rect 14655 4855 14775 4975
rect 14830 4855 14950 4975
rect 14995 4855 15115 4975
rect 15160 4855 15280 4975
rect 15325 4855 15445 4975
rect 15500 4855 15620 4975
rect 15665 4855 15785 4975
rect 15830 4855 15950 4975
rect 15995 4855 16115 4975
rect 16170 4855 16290 4975
rect 16335 4855 16455 4975
rect 16500 4855 16620 4975
rect 16665 4855 16785 4975
rect 16840 4855 16960 4975
rect 17005 4855 17125 4975
rect 17170 4855 17290 4975
rect 17335 4855 17455 4975
rect 17510 4855 17630 4975
rect 17675 4855 17795 4975
rect 17840 4855 17960 4975
rect 18005 4855 18125 4975
rect 18180 4855 18300 4975
rect 12820 4690 12940 4810
rect 12985 4690 13105 4810
rect 13150 4690 13270 4810
rect 13315 4690 13435 4810
rect 13490 4690 13610 4810
rect 13655 4690 13775 4810
rect 13820 4690 13940 4810
rect 13985 4690 14105 4810
rect 14160 4690 14280 4810
rect 14325 4690 14445 4810
rect 14490 4690 14610 4810
rect 14655 4690 14775 4810
rect 14830 4690 14950 4810
rect 14995 4690 15115 4810
rect 15160 4690 15280 4810
rect 15325 4690 15445 4810
rect 15500 4690 15620 4810
rect 15665 4690 15785 4810
rect 15830 4690 15950 4810
rect 15995 4690 16115 4810
rect 16170 4690 16290 4810
rect 16335 4690 16455 4810
rect 16500 4690 16620 4810
rect 16665 4690 16785 4810
rect 16840 4690 16960 4810
rect 17005 4690 17125 4810
rect 17170 4690 17290 4810
rect 17335 4690 17455 4810
rect 17510 4690 17630 4810
rect 17675 4690 17795 4810
rect 17840 4690 17960 4810
rect 18005 4690 18125 4810
rect 18180 4690 18300 4810
rect 12820 4525 12940 4645
rect 12985 4525 13105 4645
rect 13150 4525 13270 4645
rect 13315 4525 13435 4645
rect 13490 4525 13610 4645
rect 13655 4525 13775 4645
rect 13820 4525 13940 4645
rect 13985 4525 14105 4645
rect 14160 4525 14280 4645
rect 14325 4525 14445 4645
rect 14490 4525 14610 4645
rect 14655 4525 14775 4645
rect 14830 4525 14950 4645
rect 14995 4525 15115 4645
rect 15160 4525 15280 4645
rect 15325 4525 15445 4645
rect 15500 4525 15620 4645
rect 15665 4525 15785 4645
rect 15830 4525 15950 4645
rect 15995 4525 16115 4645
rect 16170 4525 16290 4645
rect 16335 4525 16455 4645
rect 16500 4525 16620 4645
rect 16665 4525 16785 4645
rect 16840 4525 16960 4645
rect 17005 4525 17125 4645
rect 17170 4525 17290 4645
rect 17335 4525 17455 4645
rect 17510 4525 17630 4645
rect 17675 4525 17795 4645
rect 17840 4525 17960 4645
rect 18005 4525 18125 4645
rect 18180 4525 18300 4645
rect 12820 4360 12940 4480
rect 12985 4360 13105 4480
rect 13150 4360 13270 4480
rect 13315 4360 13435 4480
rect 13490 4360 13610 4480
rect 13655 4360 13775 4480
rect 13820 4360 13940 4480
rect 13985 4360 14105 4480
rect 14160 4360 14280 4480
rect 14325 4360 14445 4480
rect 14490 4360 14610 4480
rect 14655 4360 14775 4480
rect 14830 4360 14950 4480
rect 14995 4360 15115 4480
rect 15160 4360 15280 4480
rect 15325 4360 15445 4480
rect 15500 4360 15620 4480
rect 15665 4360 15785 4480
rect 15830 4360 15950 4480
rect 15995 4360 16115 4480
rect 16170 4360 16290 4480
rect 16335 4360 16455 4480
rect 16500 4360 16620 4480
rect 16665 4360 16785 4480
rect 16840 4360 16960 4480
rect 17005 4360 17125 4480
rect 17170 4360 17290 4480
rect 17335 4360 17455 4480
rect 17510 4360 17630 4480
rect 17675 4360 17795 4480
rect 17840 4360 17960 4480
rect 18005 4360 18125 4480
rect 18180 4360 18300 4480
rect 12820 4185 12940 4305
rect 12985 4185 13105 4305
rect 13150 4185 13270 4305
rect 13315 4185 13435 4305
rect 13490 4185 13610 4305
rect 13655 4185 13775 4305
rect 13820 4185 13940 4305
rect 13985 4185 14105 4305
rect 14160 4185 14280 4305
rect 14325 4185 14445 4305
rect 14490 4185 14610 4305
rect 14655 4185 14775 4305
rect 14830 4185 14950 4305
rect 14995 4185 15115 4305
rect 15160 4185 15280 4305
rect 15325 4185 15445 4305
rect 15500 4185 15620 4305
rect 15665 4185 15785 4305
rect 15830 4185 15950 4305
rect 15995 4185 16115 4305
rect 16170 4185 16290 4305
rect 16335 4185 16455 4305
rect 16500 4185 16620 4305
rect 16665 4185 16785 4305
rect 16840 4185 16960 4305
rect 17005 4185 17125 4305
rect 17170 4185 17290 4305
rect 17335 4185 17455 4305
rect 17510 4185 17630 4305
rect 17675 4185 17795 4305
rect 17840 4185 17960 4305
rect 18005 4185 18125 4305
rect 18180 4185 18300 4305
rect 12820 4020 12940 4140
rect 12985 4020 13105 4140
rect 13150 4020 13270 4140
rect 13315 4020 13435 4140
rect 13490 4020 13610 4140
rect 13655 4020 13775 4140
rect 13820 4020 13940 4140
rect 13985 4020 14105 4140
rect 14160 4020 14280 4140
rect 14325 4020 14445 4140
rect 14490 4020 14610 4140
rect 14655 4020 14775 4140
rect 14830 4020 14950 4140
rect 14995 4020 15115 4140
rect 15160 4020 15280 4140
rect 15325 4020 15445 4140
rect 15500 4020 15620 4140
rect 15665 4020 15785 4140
rect 15830 4020 15950 4140
rect 15995 4020 16115 4140
rect 16170 4020 16290 4140
rect 16335 4020 16455 4140
rect 16500 4020 16620 4140
rect 16665 4020 16785 4140
rect 16840 4020 16960 4140
rect 17005 4020 17125 4140
rect 17170 4020 17290 4140
rect 17335 4020 17455 4140
rect 17510 4020 17630 4140
rect 17675 4020 17795 4140
rect 17840 4020 17960 4140
rect 18005 4020 18125 4140
rect 18180 4020 18300 4140
rect 12820 3855 12940 3975
rect 12985 3855 13105 3975
rect 13150 3855 13270 3975
rect 13315 3855 13435 3975
rect 13490 3855 13610 3975
rect 13655 3855 13775 3975
rect 13820 3855 13940 3975
rect 13985 3855 14105 3975
rect 14160 3855 14280 3975
rect 14325 3855 14445 3975
rect 14490 3855 14610 3975
rect 14655 3855 14775 3975
rect 14830 3855 14950 3975
rect 14995 3855 15115 3975
rect 15160 3855 15280 3975
rect 15325 3855 15445 3975
rect 15500 3855 15620 3975
rect 15665 3855 15785 3975
rect 15830 3855 15950 3975
rect 15995 3855 16115 3975
rect 16170 3855 16290 3975
rect 16335 3855 16455 3975
rect 16500 3855 16620 3975
rect 16665 3855 16785 3975
rect 16840 3855 16960 3975
rect 17005 3855 17125 3975
rect 17170 3855 17290 3975
rect 17335 3855 17455 3975
rect 17510 3855 17630 3975
rect 17675 3855 17795 3975
rect 17840 3855 17960 3975
rect 18005 3855 18125 3975
rect 18180 3855 18300 3975
rect 12820 3690 12940 3810
rect 12985 3690 13105 3810
rect 13150 3690 13270 3810
rect 13315 3690 13435 3810
rect 13490 3690 13610 3810
rect 13655 3690 13775 3810
rect 13820 3690 13940 3810
rect 13985 3690 14105 3810
rect 14160 3690 14280 3810
rect 14325 3690 14445 3810
rect 14490 3690 14610 3810
rect 14655 3690 14775 3810
rect 14830 3690 14950 3810
rect 14995 3690 15115 3810
rect 15160 3690 15280 3810
rect 15325 3690 15445 3810
rect 15500 3690 15620 3810
rect 15665 3690 15785 3810
rect 15830 3690 15950 3810
rect 15995 3690 16115 3810
rect 16170 3690 16290 3810
rect 16335 3690 16455 3810
rect 16500 3690 16620 3810
rect 16665 3690 16785 3810
rect 16840 3690 16960 3810
rect 17005 3690 17125 3810
rect 17170 3690 17290 3810
rect 17335 3690 17455 3810
rect 17510 3690 17630 3810
rect 17675 3690 17795 3810
rect 17840 3690 17960 3810
rect 18005 3690 18125 3810
rect 18180 3690 18300 3810
rect 12820 3515 12940 3635
rect 12985 3515 13105 3635
rect 13150 3515 13270 3635
rect 13315 3515 13435 3635
rect 13490 3515 13610 3635
rect 13655 3515 13775 3635
rect 13820 3515 13940 3635
rect 13985 3515 14105 3635
rect 14160 3515 14280 3635
rect 14325 3515 14445 3635
rect 14490 3515 14610 3635
rect 14655 3515 14775 3635
rect 14830 3515 14950 3635
rect 14995 3515 15115 3635
rect 15160 3515 15280 3635
rect 15325 3515 15445 3635
rect 15500 3515 15620 3635
rect 15665 3515 15785 3635
rect 15830 3515 15950 3635
rect 15995 3515 16115 3635
rect 16170 3515 16290 3635
rect 16335 3515 16455 3635
rect 16500 3515 16620 3635
rect 16665 3515 16785 3635
rect 16840 3515 16960 3635
rect 17005 3515 17125 3635
rect 17170 3515 17290 3635
rect 17335 3515 17455 3635
rect 17510 3515 17630 3635
rect 17675 3515 17795 3635
rect 17840 3515 17960 3635
rect 18005 3515 18125 3635
rect 18180 3515 18300 3635
rect 12820 3350 12940 3470
rect 12985 3350 13105 3470
rect 13150 3350 13270 3470
rect 13315 3350 13435 3470
rect 13490 3350 13610 3470
rect 13655 3350 13775 3470
rect 13820 3350 13940 3470
rect 13985 3350 14105 3470
rect 14160 3350 14280 3470
rect 14325 3350 14445 3470
rect 14490 3350 14610 3470
rect 14655 3350 14775 3470
rect 14830 3350 14950 3470
rect 14995 3350 15115 3470
rect 15160 3350 15280 3470
rect 15325 3350 15445 3470
rect 15500 3350 15620 3470
rect 15665 3350 15785 3470
rect 15830 3350 15950 3470
rect 15995 3350 16115 3470
rect 16170 3350 16290 3470
rect 16335 3350 16455 3470
rect 16500 3350 16620 3470
rect 16665 3350 16785 3470
rect 16840 3350 16960 3470
rect 17005 3350 17125 3470
rect 17170 3350 17290 3470
rect 17335 3350 17455 3470
rect 17510 3350 17630 3470
rect 17675 3350 17795 3470
rect 17840 3350 17960 3470
rect 18005 3350 18125 3470
rect 18180 3350 18300 3470
rect 12820 3185 12940 3305
rect 12985 3185 13105 3305
rect 13150 3185 13270 3305
rect 13315 3185 13435 3305
rect 13490 3185 13610 3305
rect 13655 3185 13775 3305
rect 13820 3185 13940 3305
rect 13985 3185 14105 3305
rect 14160 3185 14280 3305
rect 14325 3185 14445 3305
rect 14490 3185 14610 3305
rect 14655 3185 14775 3305
rect 14830 3185 14950 3305
rect 14995 3185 15115 3305
rect 15160 3185 15280 3305
rect 15325 3185 15445 3305
rect 15500 3185 15620 3305
rect 15665 3185 15785 3305
rect 15830 3185 15950 3305
rect 15995 3185 16115 3305
rect 16170 3185 16290 3305
rect 16335 3185 16455 3305
rect 16500 3185 16620 3305
rect 16665 3185 16785 3305
rect 16840 3185 16960 3305
rect 17005 3185 17125 3305
rect 17170 3185 17290 3305
rect 17335 3185 17455 3305
rect 17510 3185 17630 3305
rect 17675 3185 17795 3305
rect 17840 3185 17960 3305
rect 18005 3185 18125 3305
rect 18180 3185 18300 3305
rect 12820 3020 12940 3140
rect 12985 3020 13105 3140
rect 13150 3020 13270 3140
rect 13315 3020 13435 3140
rect 13490 3020 13610 3140
rect 13655 3020 13775 3140
rect 13820 3020 13940 3140
rect 13985 3020 14105 3140
rect 14160 3020 14280 3140
rect 14325 3020 14445 3140
rect 14490 3020 14610 3140
rect 14655 3020 14775 3140
rect 14830 3020 14950 3140
rect 14995 3020 15115 3140
rect 15160 3020 15280 3140
rect 15325 3020 15445 3140
rect 15500 3020 15620 3140
rect 15665 3020 15785 3140
rect 15830 3020 15950 3140
rect 15995 3020 16115 3140
rect 16170 3020 16290 3140
rect 16335 3020 16455 3140
rect 16500 3020 16620 3140
rect 16665 3020 16785 3140
rect 16840 3020 16960 3140
rect 17005 3020 17125 3140
rect 17170 3020 17290 3140
rect 17335 3020 17455 3140
rect 17510 3020 17630 3140
rect 17675 3020 17795 3140
rect 17840 3020 17960 3140
rect 18005 3020 18125 3140
rect 18180 3020 18300 3140
rect 12820 2845 12940 2965
rect 12985 2845 13105 2965
rect 13150 2845 13270 2965
rect 13315 2845 13435 2965
rect 13490 2845 13610 2965
rect 13655 2845 13775 2965
rect 13820 2845 13940 2965
rect 13985 2845 14105 2965
rect 14160 2845 14280 2965
rect 14325 2845 14445 2965
rect 14490 2845 14610 2965
rect 14655 2845 14775 2965
rect 14830 2845 14950 2965
rect 14995 2845 15115 2965
rect 15160 2845 15280 2965
rect 15325 2845 15445 2965
rect 15500 2845 15620 2965
rect 15665 2845 15785 2965
rect 15830 2845 15950 2965
rect 15995 2845 16115 2965
rect 16170 2845 16290 2965
rect 16335 2845 16455 2965
rect 16500 2845 16620 2965
rect 16665 2845 16785 2965
rect 16840 2845 16960 2965
rect 17005 2845 17125 2965
rect 17170 2845 17290 2965
rect 17335 2845 17455 2965
rect 17510 2845 17630 2965
rect 17675 2845 17795 2965
rect 17840 2845 17960 2965
rect 18005 2845 18125 2965
rect 18180 2845 18300 2965
rect 12820 2680 12940 2800
rect 12985 2680 13105 2800
rect 13150 2680 13270 2800
rect 13315 2680 13435 2800
rect 13490 2680 13610 2800
rect 13655 2680 13775 2800
rect 13820 2680 13940 2800
rect 13985 2680 14105 2800
rect 14160 2680 14280 2800
rect 14325 2680 14445 2800
rect 14490 2680 14610 2800
rect 14655 2680 14775 2800
rect 14830 2680 14950 2800
rect 14995 2680 15115 2800
rect 15160 2680 15280 2800
rect 15325 2680 15445 2800
rect 15500 2680 15620 2800
rect 15665 2680 15785 2800
rect 15830 2680 15950 2800
rect 15995 2680 16115 2800
rect 16170 2680 16290 2800
rect 16335 2680 16455 2800
rect 16500 2680 16620 2800
rect 16665 2680 16785 2800
rect 16840 2680 16960 2800
rect 17005 2680 17125 2800
rect 17170 2680 17290 2800
rect 17335 2680 17455 2800
rect 17510 2680 17630 2800
rect 17675 2680 17795 2800
rect 17840 2680 17960 2800
rect 18005 2680 18125 2800
rect 18180 2680 18300 2800
rect 12820 2515 12940 2635
rect 12985 2515 13105 2635
rect 13150 2515 13270 2635
rect 13315 2515 13435 2635
rect 13490 2515 13610 2635
rect 13655 2515 13775 2635
rect 13820 2515 13940 2635
rect 13985 2515 14105 2635
rect 14160 2515 14280 2635
rect 14325 2515 14445 2635
rect 14490 2515 14610 2635
rect 14655 2515 14775 2635
rect 14830 2515 14950 2635
rect 14995 2515 15115 2635
rect 15160 2515 15280 2635
rect 15325 2515 15445 2635
rect 15500 2515 15620 2635
rect 15665 2515 15785 2635
rect 15830 2515 15950 2635
rect 15995 2515 16115 2635
rect 16170 2515 16290 2635
rect 16335 2515 16455 2635
rect 16500 2515 16620 2635
rect 16665 2515 16785 2635
rect 16840 2515 16960 2635
rect 17005 2515 17125 2635
rect 17170 2515 17290 2635
rect 17335 2515 17455 2635
rect 17510 2515 17630 2635
rect 17675 2515 17795 2635
rect 17840 2515 17960 2635
rect 18005 2515 18125 2635
rect 18180 2515 18300 2635
rect 12820 2350 12940 2470
rect 12985 2350 13105 2470
rect 13150 2350 13270 2470
rect 13315 2350 13435 2470
rect 13490 2350 13610 2470
rect 13655 2350 13775 2470
rect 13820 2350 13940 2470
rect 13985 2350 14105 2470
rect 14160 2350 14280 2470
rect 14325 2350 14445 2470
rect 14490 2350 14610 2470
rect 14655 2350 14775 2470
rect 14830 2350 14950 2470
rect 14995 2350 15115 2470
rect 15160 2350 15280 2470
rect 15325 2350 15445 2470
rect 15500 2350 15620 2470
rect 15665 2350 15785 2470
rect 15830 2350 15950 2470
rect 15995 2350 16115 2470
rect 16170 2350 16290 2470
rect 16335 2350 16455 2470
rect 16500 2350 16620 2470
rect 16665 2350 16785 2470
rect 16840 2350 16960 2470
rect 17005 2350 17125 2470
rect 17170 2350 17290 2470
rect 17335 2350 17455 2470
rect 17510 2350 17630 2470
rect 17675 2350 17795 2470
rect 17840 2350 17960 2470
rect 18005 2350 18125 2470
rect 18180 2350 18300 2470
rect 12820 2175 12940 2295
rect 12985 2175 13105 2295
rect 13150 2175 13270 2295
rect 13315 2175 13435 2295
rect 13490 2175 13610 2295
rect 13655 2175 13775 2295
rect 13820 2175 13940 2295
rect 13985 2175 14105 2295
rect 14160 2175 14280 2295
rect 14325 2175 14445 2295
rect 14490 2175 14610 2295
rect 14655 2175 14775 2295
rect 14830 2175 14950 2295
rect 14995 2175 15115 2295
rect 15160 2175 15280 2295
rect 15325 2175 15445 2295
rect 15500 2175 15620 2295
rect 15665 2175 15785 2295
rect 15830 2175 15950 2295
rect 15995 2175 16115 2295
rect 16170 2175 16290 2295
rect 16335 2175 16455 2295
rect 16500 2175 16620 2295
rect 16665 2175 16785 2295
rect 16840 2175 16960 2295
rect 17005 2175 17125 2295
rect 17170 2175 17290 2295
rect 17335 2175 17455 2295
rect 17510 2175 17630 2295
rect 17675 2175 17795 2295
rect 17840 2175 17960 2295
rect 18005 2175 18125 2295
rect 18180 2175 18300 2295
rect 12820 2010 12940 2130
rect 12985 2010 13105 2130
rect 13150 2010 13270 2130
rect 13315 2010 13435 2130
rect 13490 2010 13610 2130
rect 13655 2010 13775 2130
rect 13820 2010 13940 2130
rect 13985 2010 14105 2130
rect 14160 2010 14280 2130
rect 14325 2010 14445 2130
rect 14490 2010 14610 2130
rect 14655 2010 14775 2130
rect 14830 2010 14950 2130
rect 14995 2010 15115 2130
rect 15160 2010 15280 2130
rect 15325 2010 15445 2130
rect 15500 2010 15620 2130
rect 15665 2010 15785 2130
rect 15830 2010 15950 2130
rect 15995 2010 16115 2130
rect 16170 2010 16290 2130
rect 16335 2010 16455 2130
rect 16500 2010 16620 2130
rect 16665 2010 16785 2130
rect 16840 2010 16960 2130
rect 17005 2010 17125 2130
rect 17170 2010 17290 2130
rect 17335 2010 17455 2130
rect 17510 2010 17630 2130
rect 17675 2010 17795 2130
rect 17840 2010 17960 2130
rect 18005 2010 18125 2130
rect 18180 2010 18300 2130
rect 12820 1845 12940 1965
rect 12985 1845 13105 1965
rect 13150 1845 13270 1965
rect 13315 1845 13435 1965
rect 13490 1845 13610 1965
rect 13655 1845 13775 1965
rect 13820 1845 13940 1965
rect 13985 1845 14105 1965
rect 14160 1845 14280 1965
rect 14325 1845 14445 1965
rect 14490 1845 14610 1965
rect 14655 1845 14775 1965
rect 14830 1845 14950 1965
rect 14995 1845 15115 1965
rect 15160 1845 15280 1965
rect 15325 1845 15445 1965
rect 15500 1845 15620 1965
rect 15665 1845 15785 1965
rect 15830 1845 15950 1965
rect 15995 1845 16115 1965
rect 16170 1845 16290 1965
rect 16335 1845 16455 1965
rect 16500 1845 16620 1965
rect 16665 1845 16785 1965
rect 16840 1845 16960 1965
rect 17005 1845 17125 1965
rect 17170 1845 17290 1965
rect 17335 1845 17455 1965
rect 17510 1845 17630 1965
rect 17675 1845 17795 1965
rect 17840 1845 17960 1965
rect 18005 1845 18125 1965
rect 18180 1845 18300 1965
rect 12820 1680 12940 1800
rect 12985 1680 13105 1800
rect 13150 1680 13270 1800
rect 13315 1680 13435 1800
rect 13490 1680 13610 1800
rect 13655 1680 13775 1800
rect 13820 1680 13940 1800
rect 13985 1680 14105 1800
rect 14160 1680 14280 1800
rect 14325 1680 14445 1800
rect 14490 1680 14610 1800
rect 14655 1680 14775 1800
rect 14830 1680 14950 1800
rect 14995 1680 15115 1800
rect 15160 1680 15280 1800
rect 15325 1680 15445 1800
rect 15500 1680 15620 1800
rect 15665 1680 15785 1800
rect 15830 1680 15950 1800
rect 15995 1680 16115 1800
rect 16170 1680 16290 1800
rect 16335 1680 16455 1800
rect 16500 1680 16620 1800
rect 16665 1680 16785 1800
rect 16840 1680 16960 1800
rect 17005 1680 17125 1800
rect 17170 1680 17290 1800
rect 17335 1680 17455 1800
rect 17510 1680 17630 1800
rect 17675 1680 17795 1800
rect 17840 1680 17960 1800
rect 18005 1680 18125 1800
rect 18180 1680 18300 1800
rect 18510 7040 18630 7160
rect 18675 7040 18795 7160
rect 18840 7040 18960 7160
rect 19005 7040 19125 7160
rect 19180 7040 19300 7160
rect 19345 7040 19465 7160
rect 19510 7040 19630 7160
rect 19675 7040 19795 7160
rect 19850 7040 19970 7160
rect 20015 7040 20135 7160
rect 20180 7040 20300 7160
rect 20345 7040 20465 7160
rect 20520 7040 20640 7160
rect 20685 7040 20805 7160
rect 20850 7040 20970 7160
rect 21015 7040 21135 7160
rect 21190 7040 21310 7160
rect 21355 7040 21475 7160
rect 21520 7040 21640 7160
rect 21685 7040 21805 7160
rect 21860 7040 21980 7160
rect 22025 7040 22145 7160
rect 22190 7040 22310 7160
rect 22355 7040 22475 7160
rect 22530 7040 22650 7160
rect 22695 7040 22815 7160
rect 22860 7040 22980 7160
rect 23025 7040 23145 7160
rect 23200 7040 23320 7160
rect 23365 7040 23485 7160
rect 23530 7040 23650 7160
rect 23695 7040 23815 7160
rect 23870 7040 23990 7160
rect 18510 6865 18630 6985
rect 18675 6865 18795 6985
rect 18840 6865 18960 6985
rect 19005 6865 19125 6985
rect 19180 6865 19300 6985
rect 19345 6865 19465 6985
rect 19510 6865 19630 6985
rect 19675 6865 19795 6985
rect 19850 6865 19970 6985
rect 20015 6865 20135 6985
rect 20180 6865 20300 6985
rect 20345 6865 20465 6985
rect 20520 6865 20640 6985
rect 20685 6865 20805 6985
rect 20850 6865 20970 6985
rect 21015 6865 21135 6985
rect 21190 6865 21310 6985
rect 21355 6865 21475 6985
rect 21520 6865 21640 6985
rect 21685 6865 21805 6985
rect 21860 6865 21980 6985
rect 22025 6865 22145 6985
rect 22190 6865 22310 6985
rect 22355 6865 22475 6985
rect 22530 6865 22650 6985
rect 22695 6865 22815 6985
rect 22860 6865 22980 6985
rect 23025 6865 23145 6985
rect 23200 6865 23320 6985
rect 23365 6865 23485 6985
rect 23530 6865 23650 6985
rect 23695 6865 23815 6985
rect 23870 6865 23990 6985
rect 18510 6700 18630 6820
rect 18675 6700 18795 6820
rect 18840 6700 18960 6820
rect 19005 6700 19125 6820
rect 19180 6700 19300 6820
rect 19345 6700 19465 6820
rect 19510 6700 19630 6820
rect 19675 6700 19795 6820
rect 19850 6700 19970 6820
rect 20015 6700 20135 6820
rect 20180 6700 20300 6820
rect 20345 6700 20465 6820
rect 20520 6700 20640 6820
rect 20685 6700 20805 6820
rect 20850 6700 20970 6820
rect 21015 6700 21135 6820
rect 21190 6700 21310 6820
rect 21355 6700 21475 6820
rect 21520 6700 21640 6820
rect 21685 6700 21805 6820
rect 21860 6700 21980 6820
rect 22025 6700 22145 6820
rect 22190 6700 22310 6820
rect 22355 6700 22475 6820
rect 22530 6700 22650 6820
rect 22695 6700 22815 6820
rect 22860 6700 22980 6820
rect 23025 6700 23145 6820
rect 23200 6700 23320 6820
rect 23365 6700 23485 6820
rect 23530 6700 23650 6820
rect 23695 6700 23815 6820
rect 23870 6700 23990 6820
rect 18510 6535 18630 6655
rect 18675 6535 18795 6655
rect 18840 6535 18960 6655
rect 19005 6535 19125 6655
rect 19180 6535 19300 6655
rect 19345 6535 19465 6655
rect 19510 6535 19630 6655
rect 19675 6535 19795 6655
rect 19850 6535 19970 6655
rect 20015 6535 20135 6655
rect 20180 6535 20300 6655
rect 20345 6535 20465 6655
rect 20520 6535 20640 6655
rect 20685 6535 20805 6655
rect 20850 6535 20970 6655
rect 21015 6535 21135 6655
rect 21190 6535 21310 6655
rect 21355 6535 21475 6655
rect 21520 6535 21640 6655
rect 21685 6535 21805 6655
rect 21860 6535 21980 6655
rect 22025 6535 22145 6655
rect 22190 6535 22310 6655
rect 22355 6535 22475 6655
rect 22530 6535 22650 6655
rect 22695 6535 22815 6655
rect 22860 6535 22980 6655
rect 23025 6535 23145 6655
rect 23200 6535 23320 6655
rect 23365 6535 23485 6655
rect 23530 6535 23650 6655
rect 23695 6535 23815 6655
rect 23870 6535 23990 6655
rect 18510 6370 18630 6490
rect 18675 6370 18795 6490
rect 18840 6370 18960 6490
rect 19005 6370 19125 6490
rect 19180 6370 19300 6490
rect 19345 6370 19465 6490
rect 19510 6370 19630 6490
rect 19675 6370 19795 6490
rect 19850 6370 19970 6490
rect 20015 6370 20135 6490
rect 20180 6370 20300 6490
rect 20345 6370 20465 6490
rect 20520 6370 20640 6490
rect 20685 6370 20805 6490
rect 20850 6370 20970 6490
rect 21015 6370 21135 6490
rect 21190 6370 21310 6490
rect 21355 6370 21475 6490
rect 21520 6370 21640 6490
rect 21685 6370 21805 6490
rect 21860 6370 21980 6490
rect 22025 6370 22145 6490
rect 22190 6370 22310 6490
rect 22355 6370 22475 6490
rect 22530 6370 22650 6490
rect 22695 6370 22815 6490
rect 22860 6370 22980 6490
rect 23025 6370 23145 6490
rect 23200 6370 23320 6490
rect 23365 6370 23485 6490
rect 23530 6370 23650 6490
rect 23695 6370 23815 6490
rect 23870 6370 23990 6490
rect 18510 6195 18630 6315
rect 18675 6195 18795 6315
rect 18840 6195 18960 6315
rect 19005 6195 19125 6315
rect 19180 6195 19300 6315
rect 19345 6195 19465 6315
rect 19510 6195 19630 6315
rect 19675 6195 19795 6315
rect 19850 6195 19970 6315
rect 20015 6195 20135 6315
rect 20180 6195 20300 6315
rect 20345 6195 20465 6315
rect 20520 6195 20640 6315
rect 20685 6195 20805 6315
rect 20850 6195 20970 6315
rect 21015 6195 21135 6315
rect 21190 6195 21310 6315
rect 21355 6195 21475 6315
rect 21520 6195 21640 6315
rect 21685 6195 21805 6315
rect 21860 6195 21980 6315
rect 22025 6195 22145 6315
rect 22190 6195 22310 6315
rect 22355 6195 22475 6315
rect 22530 6195 22650 6315
rect 22695 6195 22815 6315
rect 22860 6195 22980 6315
rect 23025 6195 23145 6315
rect 23200 6195 23320 6315
rect 23365 6195 23485 6315
rect 23530 6195 23650 6315
rect 23695 6195 23815 6315
rect 23870 6195 23990 6315
rect 18510 6030 18630 6150
rect 18675 6030 18795 6150
rect 18840 6030 18960 6150
rect 19005 6030 19125 6150
rect 19180 6030 19300 6150
rect 19345 6030 19465 6150
rect 19510 6030 19630 6150
rect 19675 6030 19795 6150
rect 19850 6030 19970 6150
rect 20015 6030 20135 6150
rect 20180 6030 20300 6150
rect 20345 6030 20465 6150
rect 20520 6030 20640 6150
rect 20685 6030 20805 6150
rect 20850 6030 20970 6150
rect 21015 6030 21135 6150
rect 21190 6030 21310 6150
rect 21355 6030 21475 6150
rect 21520 6030 21640 6150
rect 21685 6030 21805 6150
rect 21860 6030 21980 6150
rect 22025 6030 22145 6150
rect 22190 6030 22310 6150
rect 22355 6030 22475 6150
rect 22530 6030 22650 6150
rect 22695 6030 22815 6150
rect 22860 6030 22980 6150
rect 23025 6030 23145 6150
rect 23200 6030 23320 6150
rect 23365 6030 23485 6150
rect 23530 6030 23650 6150
rect 23695 6030 23815 6150
rect 23870 6030 23990 6150
rect 18510 5865 18630 5985
rect 18675 5865 18795 5985
rect 18840 5865 18960 5985
rect 19005 5865 19125 5985
rect 19180 5865 19300 5985
rect 19345 5865 19465 5985
rect 19510 5865 19630 5985
rect 19675 5865 19795 5985
rect 19850 5865 19970 5985
rect 20015 5865 20135 5985
rect 20180 5865 20300 5985
rect 20345 5865 20465 5985
rect 20520 5865 20640 5985
rect 20685 5865 20805 5985
rect 20850 5865 20970 5985
rect 21015 5865 21135 5985
rect 21190 5865 21310 5985
rect 21355 5865 21475 5985
rect 21520 5865 21640 5985
rect 21685 5865 21805 5985
rect 21860 5865 21980 5985
rect 22025 5865 22145 5985
rect 22190 5865 22310 5985
rect 22355 5865 22475 5985
rect 22530 5865 22650 5985
rect 22695 5865 22815 5985
rect 22860 5865 22980 5985
rect 23025 5865 23145 5985
rect 23200 5865 23320 5985
rect 23365 5865 23485 5985
rect 23530 5865 23650 5985
rect 23695 5865 23815 5985
rect 23870 5865 23990 5985
rect 18510 5700 18630 5820
rect 18675 5700 18795 5820
rect 18840 5700 18960 5820
rect 19005 5700 19125 5820
rect 19180 5700 19300 5820
rect 19345 5700 19465 5820
rect 19510 5700 19630 5820
rect 19675 5700 19795 5820
rect 19850 5700 19970 5820
rect 20015 5700 20135 5820
rect 20180 5700 20300 5820
rect 20345 5700 20465 5820
rect 20520 5700 20640 5820
rect 20685 5700 20805 5820
rect 20850 5700 20970 5820
rect 21015 5700 21135 5820
rect 21190 5700 21310 5820
rect 21355 5700 21475 5820
rect 21520 5700 21640 5820
rect 21685 5700 21805 5820
rect 21860 5700 21980 5820
rect 22025 5700 22145 5820
rect 22190 5700 22310 5820
rect 22355 5700 22475 5820
rect 22530 5700 22650 5820
rect 22695 5700 22815 5820
rect 22860 5700 22980 5820
rect 23025 5700 23145 5820
rect 23200 5700 23320 5820
rect 23365 5700 23485 5820
rect 23530 5700 23650 5820
rect 23695 5700 23815 5820
rect 23870 5700 23990 5820
rect 18510 5525 18630 5645
rect 18675 5525 18795 5645
rect 18840 5525 18960 5645
rect 19005 5525 19125 5645
rect 19180 5525 19300 5645
rect 19345 5525 19465 5645
rect 19510 5525 19630 5645
rect 19675 5525 19795 5645
rect 19850 5525 19970 5645
rect 20015 5525 20135 5645
rect 20180 5525 20300 5645
rect 20345 5525 20465 5645
rect 20520 5525 20640 5645
rect 20685 5525 20805 5645
rect 20850 5525 20970 5645
rect 21015 5525 21135 5645
rect 21190 5525 21310 5645
rect 21355 5525 21475 5645
rect 21520 5525 21640 5645
rect 21685 5525 21805 5645
rect 21860 5525 21980 5645
rect 22025 5525 22145 5645
rect 22190 5525 22310 5645
rect 22355 5525 22475 5645
rect 22530 5525 22650 5645
rect 22695 5525 22815 5645
rect 22860 5525 22980 5645
rect 23025 5525 23145 5645
rect 23200 5525 23320 5645
rect 23365 5525 23485 5645
rect 23530 5525 23650 5645
rect 23695 5525 23815 5645
rect 23870 5525 23990 5645
rect 18510 5360 18630 5480
rect 18675 5360 18795 5480
rect 18840 5360 18960 5480
rect 19005 5360 19125 5480
rect 19180 5360 19300 5480
rect 19345 5360 19465 5480
rect 19510 5360 19630 5480
rect 19675 5360 19795 5480
rect 19850 5360 19970 5480
rect 20015 5360 20135 5480
rect 20180 5360 20300 5480
rect 20345 5360 20465 5480
rect 20520 5360 20640 5480
rect 20685 5360 20805 5480
rect 20850 5360 20970 5480
rect 21015 5360 21135 5480
rect 21190 5360 21310 5480
rect 21355 5360 21475 5480
rect 21520 5360 21640 5480
rect 21685 5360 21805 5480
rect 21860 5360 21980 5480
rect 22025 5360 22145 5480
rect 22190 5360 22310 5480
rect 22355 5360 22475 5480
rect 22530 5360 22650 5480
rect 22695 5360 22815 5480
rect 22860 5360 22980 5480
rect 23025 5360 23145 5480
rect 23200 5360 23320 5480
rect 23365 5360 23485 5480
rect 23530 5360 23650 5480
rect 23695 5360 23815 5480
rect 23870 5360 23990 5480
rect 18510 5195 18630 5315
rect 18675 5195 18795 5315
rect 18840 5195 18960 5315
rect 19005 5195 19125 5315
rect 19180 5195 19300 5315
rect 19345 5195 19465 5315
rect 19510 5195 19630 5315
rect 19675 5195 19795 5315
rect 19850 5195 19970 5315
rect 20015 5195 20135 5315
rect 20180 5195 20300 5315
rect 20345 5195 20465 5315
rect 20520 5195 20640 5315
rect 20685 5195 20805 5315
rect 20850 5195 20970 5315
rect 21015 5195 21135 5315
rect 21190 5195 21310 5315
rect 21355 5195 21475 5315
rect 21520 5195 21640 5315
rect 21685 5195 21805 5315
rect 21860 5195 21980 5315
rect 22025 5195 22145 5315
rect 22190 5195 22310 5315
rect 22355 5195 22475 5315
rect 22530 5195 22650 5315
rect 22695 5195 22815 5315
rect 22860 5195 22980 5315
rect 23025 5195 23145 5315
rect 23200 5195 23320 5315
rect 23365 5195 23485 5315
rect 23530 5195 23650 5315
rect 23695 5195 23815 5315
rect 23870 5195 23990 5315
rect 18510 5030 18630 5150
rect 18675 5030 18795 5150
rect 18840 5030 18960 5150
rect 19005 5030 19125 5150
rect 19180 5030 19300 5150
rect 19345 5030 19465 5150
rect 19510 5030 19630 5150
rect 19675 5030 19795 5150
rect 19850 5030 19970 5150
rect 20015 5030 20135 5150
rect 20180 5030 20300 5150
rect 20345 5030 20465 5150
rect 20520 5030 20640 5150
rect 20685 5030 20805 5150
rect 20850 5030 20970 5150
rect 21015 5030 21135 5150
rect 21190 5030 21310 5150
rect 21355 5030 21475 5150
rect 21520 5030 21640 5150
rect 21685 5030 21805 5150
rect 21860 5030 21980 5150
rect 22025 5030 22145 5150
rect 22190 5030 22310 5150
rect 22355 5030 22475 5150
rect 22530 5030 22650 5150
rect 22695 5030 22815 5150
rect 22860 5030 22980 5150
rect 23025 5030 23145 5150
rect 23200 5030 23320 5150
rect 23365 5030 23485 5150
rect 23530 5030 23650 5150
rect 23695 5030 23815 5150
rect 23870 5030 23990 5150
rect 18510 4855 18630 4975
rect 18675 4855 18795 4975
rect 18840 4855 18960 4975
rect 19005 4855 19125 4975
rect 19180 4855 19300 4975
rect 19345 4855 19465 4975
rect 19510 4855 19630 4975
rect 19675 4855 19795 4975
rect 19850 4855 19970 4975
rect 20015 4855 20135 4975
rect 20180 4855 20300 4975
rect 20345 4855 20465 4975
rect 20520 4855 20640 4975
rect 20685 4855 20805 4975
rect 20850 4855 20970 4975
rect 21015 4855 21135 4975
rect 21190 4855 21310 4975
rect 21355 4855 21475 4975
rect 21520 4855 21640 4975
rect 21685 4855 21805 4975
rect 21860 4855 21980 4975
rect 22025 4855 22145 4975
rect 22190 4855 22310 4975
rect 22355 4855 22475 4975
rect 22530 4855 22650 4975
rect 22695 4855 22815 4975
rect 22860 4855 22980 4975
rect 23025 4855 23145 4975
rect 23200 4855 23320 4975
rect 23365 4855 23485 4975
rect 23530 4855 23650 4975
rect 23695 4855 23815 4975
rect 23870 4855 23990 4975
rect 18510 4690 18630 4810
rect 18675 4690 18795 4810
rect 18840 4690 18960 4810
rect 19005 4690 19125 4810
rect 19180 4690 19300 4810
rect 19345 4690 19465 4810
rect 19510 4690 19630 4810
rect 19675 4690 19795 4810
rect 19850 4690 19970 4810
rect 20015 4690 20135 4810
rect 20180 4690 20300 4810
rect 20345 4690 20465 4810
rect 20520 4690 20640 4810
rect 20685 4690 20805 4810
rect 20850 4690 20970 4810
rect 21015 4690 21135 4810
rect 21190 4690 21310 4810
rect 21355 4690 21475 4810
rect 21520 4690 21640 4810
rect 21685 4690 21805 4810
rect 21860 4690 21980 4810
rect 22025 4690 22145 4810
rect 22190 4690 22310 4810
rect 22355 4690 22475 4810
rect 22530 4690 22650 4810
rect 22695 4690 22815 4810
rect 22860 4690 22980 4810
rect 23025 4690 23145 4810
rect 23200 4690 23320 4810
rect 23365 4690 23485 4810
rect 23530 4690 23650 4810
rect 23695 4690 23815 4810
rect 23870 4690 23990 4810
rect 18510 4525 18630 4645
rect 18675 4525 18795 4645
rect 18840 4525 18960 4645
rect 19005 4525 19125 4645
rect 19180 4525 19300 4645
rect 19345 4525 19465 4645
rect 19510 4525 19630 4645
rect 19675 4525 19795 4645
rect 19850 4525 19970 4645
rect 20015 4525 20135 4645
rect 20180 4525 20300 4645
rect 20345 4525 20465 4645
rect 20520 4525 20640 4645
rect 20685 4525 20805 4645
rect 20850 4525 20970 4645
rect 21015 4525 21135 4645
rect 21190 4525 21310 4645
rect 21355 4525 21475 4645
rect 21520 4525 21640 4645
rect 21685 4525 21805 4645
rect 21860 4525 21980 4645
rect 22025 4525 22145 4645
rect 22190 4525 22310 4645
rect 22355 4525 22475 4645
rect 22530 4525 22650 4645
rect 22695 4525 22815 4645
rect 22860 4525 22980 4645
rect 23025 4525 23145 4645
rect 23200 4525 23320 4645
rect 23365 4525 23485 4645
rect 23530 4525 23650 4645
rect 23695 4525 23815 4645
rect 23870 4525 23990 4645
rect 18510 4360 18630 4480
rect 18675 4360 18795 4480
rect 18840 4360 18960 4480
rect 19005 4360 19125 4480
rect 19180 4360 19300 4480
rect 19345 4360 19465 4480
rect 19510 4360 19630 4480
rect 19675 4360 19795 4480
rect 19850 4360 19970 4480
rect 20015 4360 20135 4480
rect 20180 4360 20300 4480
rect 20345 4360 20465 4480
rect 20520 4360 20640 4480
rect 20685 4360 20805 4480
rect 20850 4360 20970 4480
rect 21015 4360 21135 4480
rect 21190 4360 21310 4480
rect 21355 4360 21475 4480
rect 21520 4360 21640 4480
rect 21685 4360 21805 4480
rect 21860 4360 21980 4480
rect 22025 4360 22145 4480
rect 22190 4360 22310 4480
rect 22355 4360 22475 4480
rect 22530 4360 22650 4480
rect 22695 4360 22815 4480
rect 22860 4360 22980 4480
rect 23025 4360 23145 4480
rect 23200 4360 23320 4480
rect 23365 4360 23485 4480
rect 23530 4360 23650 4480
rect 23695 4360 23815 4480
rect 23870 4360 23990 4480
rect 18510 4185 18630 4305
rect 18675 4185 18795 4305
rect 18840 4185 18960 4305
rect 19005 4185 19125 4305
rect 19180 4185 19300 4305
rect 19345 4185 19465 4305
rect 19510 4185 19630 4305
rect 19675 4185 19795 4305
rect 19850 4185 19970 4305
rect 20015 4185 20135 4305
rect 20180 4185 20300 4305
rect 20345 4185 20465 4305
rect 20520 4185 20640 4305
rect 20685 4185 20805 4305
rect 20850 4185 20970 4305
rect 21015 4185 21135 4305
rect 21190 4185 21310 4305
rect 21355 4185 21475 4305
rect 21520 4185 21640 4305
rect 21685 4185 21805 4305
rect 21860 4185 21980 4305
rect 22025 4185 22145 4305
rect 22190 4185 22310 4305
rect 22355 4185 22475 4305
rect 22530 4185 22650 4305
rect 22695 4185 22815 4305
rect 22860 4185 22980 4305
rect 23025 4185 23145 4305
rect 23200 4185 23320 4305
rect 23365 4185 23485 4305
rect 23530 4185 23650 4305
rect 23695 4185 23815 4305
rect 23870 4185 23990 4305
rect 18510 4020 18630 4140
rect 18675 4020 18795 4140
rect 18840 4020 18960 4140
rect 19005 4020 19125 4140
rect 19180 4020 19300 4140
rect 19345 4020 19465 4140
rect 19510 4020 19630 4140
rect 19675 4020 19795 4140
rect 19850 4020 19970 4140
rect 20015 4020 20135 4140
rect 20180 4020 20300 4140
rect 20345 4020 20465 4140
rect 20520 4020 20640 4140
rect 20685 4020 20805 4140
rect 20850 4020 20970 4140
rect 21015 4020 21135 4140
rect 21190 4020 21310 4140
rect 21355 4020 21475 4140
rect 21520 4020 21640 4140
rect 21685 4020 21805 4140
rect 21860 4020 21980 4140
rect 22025 4020 22145 4140
rect 22190 4020 22310 4140
rect 22355 4020 22475 4140
rect 22530 4020 22650 4140
rect 22695 4020 22815 4140
rect 22860 4020 22980 4140
rect 23025 4020 23145 4140
rect 23200 4020 23320 4140
rect 23365 4020 23485 4140
rect 23530 4020 23650 4140
rect 23695 4020 23815 4140
rect 23870 4020 23990 4140
rect 18510 3855 18630 3975
rect 18675 3855 18795 3975
rect 18840 3855 18960 3975
rect 19005 3855 19125 3975
rect 19180 3855 19300 3975
rect 19345 3855 19465 3975
rect 19510 3855 19630 3975
rect 19675 3855 19795 3975
rect 19850 3855 19970 3975
rect 20015 3855 20135 3975
rect 20180 3855 20300 3975
rect 20345 3855 20465 3975
rect 20520 3855 20640 3975
rect 20685 3855 20805 3975
rect 20850 3855 20970 3975
rect 21015 3855 21135 3975
rect 21190 3855 21310 3975
rect 21355 3855 21475 3975
rect 21520 3855 21640 3975
rect 21685 3855 21805 3975
rect 21860 3855 21980 3975
rect 22025 3855 22145 3975
rect 22190 3855 22310 3975
rect 22355 3855 22475 3975
rect 22530 3855 22650 3975
rect 22695 3855 22815 3975
rect 22860 3855 22980 3975
rect 23025 3855 23145 3975
rect 23200 3855 23320 3975
rect 23365 3855 23485 3975
rect 23530 3855 23650 3975
rect 23695 3855 23815 3975
rect 23870 3855 23990 3975
rect 18510 3690 18630 3810
rect 18675 3690 18795 3810
rect 18840 3690 18960 3810
rect 19005 3690 19125 3810
rect 19180 3690 19300 3810
rect 19345 3690 19465 3810
rect 19510 3690 19630 3810
rect 19675 3690 19795 3810
rect 19850 3690 19970 3810
rect 20015 3690 20135 3810
rect 20180 3690 20300 3810
rect 20345 3690 20465 3810
rect 20520 3690 20640 3810
rect 20685 3690 20805 3810
rect 20850 3690 20970 3810
rect 21015 3690 21135 3810
rect 21190 3690 21310 3810
rect 21355 3690 21475 3810
rect 21520 3690 21640 3810
rect 21685 3690 21805 3810
rect 21860 3690 21980 3810
rect 22025 3690 22145 3810
rect 22190 3690 22310 3810
rect 22355 3690 22475 3810
rect 22530 3690 22650 3810
rect 22695 3690 22815 3810
rect 22860 3690 22980 3810
rect 23025 3690 23145 3810
rect 23200 3690 23320 3810
rect 23365 3690 23485 3810
rect 23530 3690 23650 3810
rect 23695 3690 23815 3810
rect 23870 3690 23990 3810
rect 18510 3515 18630 3635
rect 18675 3515 18795 3635
rect 18840 3515 18960 3635
rect 19005 3515 19125 3635
rect 19180 3515 19300 3635
rect 19345 3515 19465 3635
rect 19510 3515 19630 3635
rect 19675 3515 19795 3635
rect 19850 3515 19970 3635
rect 20015 3515 20135 3635
rect 20180 3515 20300 3635
rect 20345 3515 20465 3635
rect 20520 3515 20640 3635
rect 20685 3515 20805 3635
rect 20850 3515 20970 3635
rect 21015 3515 21135 3635
rect 21190 3515 21310 3635
rect 21355 3515 21475 3635
rect 21520 3515 21640 3635
rect 21685 3515 21805 3635
rect 21860 3515 21980 3635
rect 22025 3515 22145 3635
rect 22190 3515 22310 3635
rect 22355 3515 22475 3635
rect 22530 3515 22650 3635
rect 22695 3515 22815 3635
rect 22860 3515 22980 3635
rect 23025 3515 23145 3635
rect 23200 3515 23320 3635
rect 23365 3515 23485 3635
rect 23530 3515 23650 3635
rect 23695 3515 23815 3635
rect 23870 3515 23990 3635
rect 18510 3350 18630 3470
rect 18675 3350 18795 3470
rect 18840 3350 18960 3470
rect 19005 3350 19125 3470
rect 19180 3350 19300 3470
rect 19345 3350 19465 3470
rect 19510 3350 19630 3470
rect 19675 3350 19795 3470
rect 19850 3350 19970 3470
rect 20015 3350 20135 3470
rect 20180 3350 20300 3470
rect 20345 3350 20465 3470
rect 20520 3350 20640 3470
rect 20685 3350 20805 3470
rect 20850 3350 20970 3470
rect 21015 3350 21135 3470
rect 21190 3350 21310 3470
rect 21355 3350 21475 3470
rect 21520 3350 21640 3470
rect 21685 3350 21805 3470
rect 21860 3350 21980 3470
rect 22025 3350 22145 3470
rect 22190 3350 22310 3470
rect 22355 3350 22475 3470
rect 22530 3350 22650 3470
rect 22695 3350 22815 3470
rect 22860 3350 22980 3470
rect 23025 3350 23145 3470
rect 23200 3350 23320 3470
rect 23365 3350 23485 3470
rect 23530 3350 23650 3470
rect 23695 3350 23815 3470
rect 23870 3350 23990 3470
rect 18510 3185 18630 3305
rect 18675 3185 18795 3305
rect 18840 3185 18960 3305
rect 19005 3185 19125 3305
rect 19180 3185 19300 3305
rect 19345 3185 19465 3305
rect 19510 3185 19630 3305
rect 19675 3185 19795 3305
rect 19850 3185 19970 3305
rect 20015 3185 20135 3305
rect 20180 3185 20300 3305
rect 20345 3185 20465 3305
rect 20520 3185 20640 3305
rect 20685 3185 20805 3305
rect 20850 3185 20970 3305
rect 21015 3185 21135 3305
rect 21190 3185 21310 3305
rect 21355 3185 21475 3305
rect 21520 3185 21640 3305
rect 21685 3185 21805 3305
rect 21860 3185 21980 3305
rect 22025 3185 22145 3305
rect 22190 3185 22310 3305
rect 22355 3185 22475 3305
rect 22530 3185 22650 3305
rect 22695 3185 22815 3305
rect 22860 3185 22980 3305
rect 23025 3185 23145 3305
rect 23200 3185 23320 3305
rect 23365 3185 23485 3305
rect 23530 3185 23650 3305
rect 23695 3185 23815 3305
rect 23870 3185 23990 3305
rect 18510 3020 18630 3140
rect 18675 3020 18795 3140
rect 18840 3020 18960 3140
rect 19005 3020 19125 3140
rect 19180 3020 19300 3140
rect 19345 3020 19465 3140
rect 19510 3020 19630 3140
rect 19675 3020 19795 3140
rect 19850 3020 19970 3140
rect 20015 3020 20135 3140
rect 20180 3020 20300 3140
rect 20345 3020 20465 3140
rect 20520 3020 20640 3140
rect 20685 3020 20805 3140
rect 20850 3020 20970 3140
rect 21015 3020 21135 3140
rect 21190 3020 21310 3140
rect 21355 3020 21475 3140
rect 21520 3020 21640 3140
rect 21685 3020 21805 3140
rect 21860 3020 21980 3140
rect 22025 3020 22145 3140
rect 22190 3020 22310 3140
rect 22355 3020 22475 3140
rect 22530 3020 22650 3140
rect 22695 3020 22815 3140
rect 22860 3020 22980 3140
rect 23025 3020 23145 3140
rect 23200 3020 23320 3140
rect 23365 3020 23485 3140
rect 23530 3020 23650 3140
rect 23695 3020 23815 3140
rect 23870 3020 23990 3140
rect 18510 2845 18630 2965
rect 18675 2845 18795 2965
rect 18840 2845 18960 2965
rect 19005 2845 19125 2965
rect 19180 2845 19300 2965
rect 19345 2845 19465 2965
rect 19510 2845 19630 2965
rect 19675 2845 19795 2965
rect 19850 2845 19970 2965
rect 20015 2845 20135 2965
rect 20180 2845 20300 2965
rect 20345 2845 20465 2965
rect 20520 2845 20640 2965
rect 20685 2845 20805 2965
rect 20850 2845 20970 2965
rect 21015 2845 21135 2965
rect 21190 2845 21310 2965
rect 21355 2845 21475 2965
rect 21520 2845 21640 2965
rect 21685 2845 21805 2965
rect 21860 2845 21980 2965
rect 22025 2845 22145 2965
rect 22190 2845 22310 2965
rect 22355 2845 22475 2965
rect 22530 2845 22650 2965
rect 22695 2845 22815 2965
rect 22860 2845 22980 2965
rect 23025 2845 23145 2965
rect 23200 2845 23320 2965
rect 23365 2845 23485 2965
rect 23530 2845 23650 2965
rect 23695 2845 23815 2965
rect 23870 2845 23990 2965
rect 18510 2680 18630 2800
rect 18675 2680 18795 2800
rect 18840 2680 18960 2800
rect 19005 2680 19125 2800
rect 19180 2680 19300 2800
rect 19345 2680 19465 2800
rect 19510 2680 19630 2800
rect 19675 2680 19795 2800
rect 19850 2680 19970 2800
rect 20015 2680 20135 2800
rect 20180 2680 20300 2800
rect 20345 2680 20465 2800
rect 20520 2680 20640 2800
rect 20685 2680 20805 2800
rect 20850 2680 20970 2800
rect 21015 2680 21135 2800
rect 21190 2680 21310 2800
rect 21355 2680 21475 2800
rect 21520 2680 21640 2800
rect 21685 2680 21805 2800
rect 21860 2680 21980 2800
rect 22025 2680 22145 2800
rect 22190 2680 22310 2800
rect 22355 2680 22475 2800
rect 22530 2680 22650 2800
rect 22695 2680 22815 2800
rect 22860 2680 22980 2800
rect 23025 2680 23145 2800
rect 23200 2680 23320 2800
rect 23365 2680 23485 2800
rect 23530 2680 23650 2800
rect 23695 2680 23815 2800
rect 23870 2680 23990 2800
rect 18510 2515 18630 2635
rect 18675 2515 18795 2635
rect 18840 2515 18960 2635
rect 19005 2515 19125 2635
rect 19180 2515 19300 2635
rect 19345 2515 19465 2635
rect 19510 2515 19630 2635
rect 19675 2515 19795 2635
rect 19850 2515 19970 2635
rect 20015 2515 20135 2635
rect 20180 2515 20300 2635
rect 20345 2515 20465 2635
rect 20520 2515 20640 2635
rect 20685 2515 20805 2635
rect 20850 2515 20970 2635
rect 21015 2515 21135 2635
rect 21190 2515 21310 2635
rect 21355 2515 21475 2635
rect 21520 2515 21640 2635
rect 21685 2515 21805 2635
rect 21860 2515 21980 2635
rect 22025 2515 22145 2635
rect 22190 2515 22310 2635
rect 22355 2515 22475 2635
rect 22530 2515 22650 2635
rect 22695 2515 22815 2635
rect 22860 2515 22980 2635
rect 23025 2515 23145 2635
rect 23200 2515 23320 2635
rect 23365 2515 23485 2635
rect 23530 2515 23650 2635
rect 23695 2515 23815 2635
rect 23870 2515 23990 2635
rect 18510 2350 18630 2470
rect 18675 2350 18795 2470
rect 18840 2350 18960 2470
rect 19005 2350 19125 2470
rect 19180 2350 19300 2470
rect 19345 2350 19465 2470
rect 19510 2350 19630 2470
rect 19675 2350 19795 2470
rect 19850 2350 19970 2470
rect 20015 2350 20135 2470
rect 20180 2350 20300 2470
rect 20345 2350 20465 2470
rect 20520 2350 20640 2470
rect 20685 2350 20805 2470
rect 20850 2350 20970 2470
rect 21015 2350 21135 2470
rect 21190 2350 21310 2470
rect 21355 2350 21475 2470
rect 21520 2350 21640 2470
rect 21685 2350 21805 2470
rect 21860 2350 21980 2470
rect 22025 2350 22145 2470
rect 22190 2350 22310 2470
rect 22355 2350 22475 2470
rect 22530 2350 22650 2470
rect 22695 2350 22815 2470
rect 22860 2350 22980 2470
rect 23025 2350 23145 2470
rect 23200 2350 23320 2470
rect 23365 2350 23485 2470
rect 23530 2350 23650 2470
rect 23695 2350 23815 2470
rect 23870 2350 23990 2470
rect 18510 2175 18630 2295
rect 18675 2175 18795 2295
rect 18840 2175 18960 2295
rect 19005 2175 19125 2295
rect 19180 2175 19300 2295
rect 19345 2175 19465 2295
rect 19510 2175 19630 2295
rect 19675 2175 19795 2295
rect 19850 2175 19970 2295
rect 20015 2175 20135 2295
rect 20180 2175 20300 2295
rect 20345 2175 20465 2295
rect 20520 2175 20640 2295
rect 20685 2175 20805 2295
rect 20850 2175 20970 2295
rect 21015 2175 21135 2295
rect 21190 2175 21310 2295
rect 21355 2175 21475 2295
rect 21520 2175 21640 2295
rect 21685 2175 21805 2295
rect 21860 2175 21980 2295
rect 22025 2175 22145 2295
rect 22190 2175 22310 2295
rect 22355 2175 22475 2295
rect 22530 2175 22650 2295
rect 22695 2175 22815 2295
rect 22860 2175 22980 2295
rect 23025 2175 23145 2295
rect 23200 2175 23320 2295
rect 23365 2175 23485 2295
rect 23530 2175 23650 2295
rect 23695 2175 23815 2295
rect 23870 2175 23990 2295
rect 18510 2010 18630 2130
rect 18675 2010 18795 2130
rect 18840 2010 18960 2130
rect 19005 2010 19125 2130
rect 19180 2010 19300 2130
rect 19345 2010 19465 2130
rect 19510 2010 19630 2130
rect 19675 2010 19795 2130
rect 19850 2010 19970 2130
rect 20015 2010 20135 2130
rect 20180 2010 20300 2130
rect 20345 2010 20465 2130
rect 20520 2010 20640 2130
rect 20685 2010 20805 2130
rect 20850 2010 20970 2130
rect 21015 2010 21135 2130
rect 21190 2010 21310 2130
rect 21355 2010 21475 2130
rect 21520 2010 21640 2130
rect 21685 2010 21805 2130
rect 21860 2010 21980 2130
rect 22025 2010 22145 2130
rect 22190 2010 22310 2130
rect 22355 2010 22475 2130
rect 22530 2010 22650 2130
rect 22695 2010 22815 2130
rect 22860 2010 22980 2130
rect 23025 2010 23145 2130
rect 23200 2010 23320 2130
rect 23365 2010 23485 2130
rect 23530 2010 23650 2130
rect 23695 2010 23815 2130
rect 23870 2010 23990 2130
rect 18510 1845 18630 1965
rect 18675 1845 18795 1965
rect 18840 1845 18960 1965
rect 19005 1845 19125 1965
rect 19180 1845 19300 1965
rect 19345 1845 19465 1965
rect 19510 1845 19630 1965
rect 19675 1845 19795 1965
rect 19850 1845 19970 1965
rect 20015 1845 20135 1965
rect 20180 1845 20300 1965
rect 20345 1845 20465 1965
rect 20520 1845 20640 1965
rect 20685 1845 20805 1965
rect 20850 1845 20970 1965
rect 21015 1845 21135 1965
rect 21190 1845 21310 1965
rect 21355 1845 21475 1965
rect 21520 1845 21640 1965
rect 21685 1845 21805 1965
rect 21860 1845 21980 1965
rect 22025 1845 22145 1965
rect 22190 1845 22310 1965
rect 22355 1845 22475 1965
rect 22530 1845 22650 1965
rect 22695 1845 22815 1965
rect 22860 1845 22980 1965
rect 23025 1845 23145 1965
rect 23200 1845 23320 1965
rect 23365 1845 23485 1965
rect 23530 1845 23650 1965
rect 23695 1845 23815 1965
rect 23870 1845 23990 1965
rect 18510 1680 18630 1800
rect 18675 1680 18795 1800
rect 18840 1680 18960 1800
rect 19005 1680 19125 1800
rect 19180 1680 19300 1800
rect 19345 1680 19465 1800
rect 19510 1680 19630 1800
rect 19675 1680 19795 1800
rect 19850 1680 19970 1800
rect 20015 1680 20135 1800
rect 20180 1680 20300 1800
rect 20345 1680 20465 1800
rect 20520 1680 20640 1800
rect 20685 1680 20805 1800
rect 20850 1680 20970 1800
rect 21015 1680 21135 1800
rect 21190 1680 21310 1800
rect 21355 1680 21475 1800
rect 21520 1680 21640 1800
rect 21685 1680 21805 1800
rect 21860 1680 21980 1800
rect 22025 1680 22145 1800
rect 22190 1680 22310 1800
rect 22355 1680 22475 1800
rect 22530 1680 22650 1800
rect 22695 1680 22815 1800
rect 22860 1680 22980 1800
rect 23025 1680 23145 1800
rect 23200 1680 23320 1800
rect 23365 1680 23485 1800
rect 23530 1680 23650 1800
rect 23695 1680 23815 1800
rect 23870 1680 23990 1800
rect 24200 7040 24320 7160
rect 24365 7040 24485 7160
rect 24530 7040 24650 7160
rect 24695 7040 24815 7160
rect 24870 7040 24990 7160
rect 25035 7040 25155 7160
rect 25200 7040 25320 7160
rect 25365 7040 25485 7160
rect 25540 7040 25660 7160
rect 25705 7040 25825 7160
rect 25870 7040 25990 7160
rect 26035 7040 26155 7160
rect 26210 7040 26330 7160
rect 26375 7040 26495 7160
rect 26540 7040 26660 7160
rect 26705 7040 26825 7160
rect 26880 7040 27000 7160
rect 27045 7040 27165 7160
rect 27210 7040 27330 7160
rect 27375 7040 27495 7160
rect 27550 7040 27670 7160
rect 27715 7040 27835 7160
rect 27880 7040 28000 7160
rect 28045 7040 28165 7160
rect 28220 7040 28340 7160
rect 28385 7040 28505 7160
rect 28550 7040 28670 7160
rect 28715 7040 28835 7160
rect 28890 7040 29010 7160
rect 29055 7040 29175 7160
rect 29220 7040 29340 7160
rect 29385 7040 29505 7160
rect 29560 7040 29680 7160
rect 24200 6865 24320 6985
rect 24365 6865 24485 6985
rect 24530 6865 24650 6985
rect 24695 6865 24815 6985
rect 24870 6865 24990 6985
rect 25035 6865 25155 6985
rect 25200 6865 25320 6985
rect 25365 6865 25485 6985
rect 25540 6865 25660 6985
rect 25705 6865 25825 6985
rect 25870 6865 25990 6985
rect 26035 6865 26155 6985
rect 26210 6865 26330 6985
rect 26375 6865 26495 6985
rect 26540 6865 26660 6985
rect 26705 6865 26825 6985
rect 26880 6865 27000 6985
rect 27045 6865 27165 6985
rect 27210 6865 27330 6985
rect 27375 6865 27495 6985
rect 27550 6865 27670 6985
rect 27715 6865 27835 6985
rect 27880 6865 28000 6985
rect 28045 6865 28165 6985
rect 28220 6865 28340 6985
rect 28385 6865 28505 6985
rect 28550 6865 28670 6985
rect 28715 6865 28835 6985
rect 28890 6865 29010 6985
rect 29055 6865 29175 6985
rect 29220 6865 29340 6985
rect 29385 6865 29505 6985
rect 29560 6865 29680 6985
rect 24200 6700 24320 6820
rect 24365 6700 24485 6820
rect 24530 6700 24650 6820
rect 24695 6700 24815 6820
rect 24870 6700 24990 6820
rect 25035 6700 25155 6820
rect 25200 6700 25320 6820
rect 25365 6700 25485 6820
rect 25540 6700 25660 6820
rect 25705 6700 25825 6820
rect 25870 6700 25990 6820
rect 26035 6700 26155 6820
rect 26210 6700 26330 6820
rect 26375 6700 26495 6820
rect 26540 6700 26660 6820
rect 26705 6700 26825 6820
rect 26880 6700 27000 6820
rect 27045 6700 27165 6820
rect 27210 6700 27330 6820
rect 27375 6700 27495 6820
rect 27550 6700 27670 6820
rect 27715 6700 27835 6820
rect 27880 6700 28000 6820
rect 28045 6700 28165 6820
rect 28220 6700 28340 6820
rect 28385 6700 28505 6820
rect 28550 6700 28670 6820
rect 28715 6700 28835 6820
rect 28890 6700 29010 6820
rect 29055 6700 29175 6820
rect 29220 6700 29340 6820
rect 29385 6700 29505 6820
rect 29560 6700 29680 6820
rect 24200 6535 24320 6655
rect 24365 6535 24485 6655
rect 24530 6535 24650 6655
rect 24695 6535 24815 6655
rect 24870 6535 24990 6655
rect 25035 6535 25155 6655
rect 25200 6535 25320 6655
rect 25365 6535 25485 6655
rect 25540 6535 25660 6655
rect 25705 6535 25825 6655
rect 25870 6535 25990 6655
rect 26035 6535 26155 6655
rect 26210 6535 26330 6655
rect 26375 6535 26495 6655
rect 26540 6535 26660 6655
rect 26705 6535 26825 6655
rect 26880 6535 27000 6655
rect 27045 6535 27165 6655
rect 27210 6535 27330 6655
rect 27375 6535 27495 6655
rect 27550 6535 27670 6655
rect 27715 6535 27835 6655
rect 27880 6535 28000 6655
rect 28045 6535 28165 6655
rect 28220 6535 28340 6655
rect 28385 6535 28505 6655
rect 28550 6535 28670 6655
rect 28715 6535 28835 6655
rect 28890 6535 29010 6655
rect 29055 6535 29175 6655
rect 29220 6535 29340 6655
rect 29385 6535 29505 6655
rect 29560 6535 29680 6655
rect 24200 6370 24320 6490
rect 24365 6370 24485 6490
rect 24530 6370 24650 6490
rect 24695 6370 24815 6490
rect 24870 6370 24990 6490
rect 25035 6370 25155 6490
rect 25200 6370 25320 6490
rect 25365 6370 25485 6490
rect 25540 6370 25660 6490
rect 25705 6370 25825 6490
rect 25870 6370 25990 6490
rect 26035 6370 26155 6490
rect 26210 6370 26330 6490
rect 26375 6370 26495 6490
rect 26540 6370 26660 6490
rect 26705 6370 26825 6490
rect 26880 6370 27000 6490
rect 27045 6370 27165 6490
rect 27210 6370 27330 6490
rect 27375 6370 27495 6490
rect 27550 6370 27670 6490
rect 27715 6370 27835 6490
rect 27880 6370 28000 6490
rect 28045 6370 28165 6490
rect 28220 6370 28340 6490
rect 28385 6370 28505 6490
rect 28550 6370 28670 6490
rect 28715 6370 28835 6490
rect 28890 6370 29010 6490
rect 29055 6370 29175 6490
rect 29220 6370 29340 6490
rect 29385 6370 29505 6490
rect 29560 6370 29680 6490
rect 24200 6195 24320 6315
rect 24365 6195 24485 6315
rect 24530 6195 24650 6315
rect 24695 6195 24815 6315
rect 24870 6195 24990 6315
rect 25035 6195 25155 6315
rect 25200 6195 25320 6315
rect 25365 6195 25485 6315
rect 25540 6195 25660 6315
rect 25705 6195 25825 6315
rect 25870 6195 25990 6315
rect 26035 6195 26155 6315
rect 26210 6195 26330 6315
rect 26375 6195 26495 6315
rect 26540 6195 26660 6315
rect 26705 6195 26825 6315
rect 26880 6195 27000 6315
rect 27045 6195 27165 6315
rect 27210 6195 27330 6315
rect 27375 6195 27495 6315
rect 27550 6195 27670 6315
rect 27715 6195 27835 6315
rect 27880 6195 28000 6315
rect 28045 6195 28165 6315
rect 28220 6195 28340 6315
rect 28385 6195 28505 6315
rect 28550 6195 28670 6315
rect 28715 6195 28835 6315
rect 28890 6195 29010 6315
rect 29055 6195 29175 6315
rect 29220 6195 29340 6315
rect 29385 6195 29505 6315
rect 29560 6195 29680 6315
rect 24200 6030 24320 6150
rect 24365 6030 24485 6150
rect 24530 6030 24650 6150
rect 24695 6030 24815 6150
rect 24870 6030 24990 6150
rect 25035 6030 25155 6150
rect 25200 6030 25320 6150
rect 25365 6030 25485 6150
rect 25540 6030 25660 6150
rect 25705 6030 25825 6150
rect 25870 6030 25990 6150
rect 26035 6030 26155 6150
rect 26210 6030 26330 6150
rect 26375 6030 26495 6150
rect 26540 6030 26660 6150
rect 26705 6030 26825 6150
rect 26880 6030 27000 6150
rect 27045 6030 27165 6150
rect 27210 6030 27330 6150
rect 27375 6030 27495 6150
rect 27550 6030 27670 6150
rect 27715 6030 27835 6150
rect 27880 6030 28000 6150
rect 28045 6030 28165 6150
rect 28220 6030 28340 6150
rect 28385 6030 28505 6150
rect 28550 6030 28670 6150
rect 28715 6030 28835 6150
rect 28890 6030 29010 6150
rect 29055 6030 29175 6150
rect 29220 6030 29340 6150
rect 29385 6030 29505 6150
rect 29560 6030 29680 6150
rect 24200 5865 24320 5985
rect 24365 5865 24485 5985
rect 24530 5865 24650 5985
rect 24695 5865 24815 5985
rect 24870 5865 24990 5985
rect 25035 5865 25155 5985
rect 25200 5865 25320 5985
rect 25365 5865 25485 5985
rect 25540 5865 25660 5985
rect 25705 5865 25825 5985
rect 25870 5865 25990 5985
rect 26035 5865 26155 5985
rect 26210 5865 26330 5985
rect 26375 5865 26495 5985
rect 26540 5865 26660 5985
rect 26705 5865 26825 5985
rect 26880 5865 27000 5985
rect 27045 5865 27165 5985
rect 27210 5865 27330 5985
rect 27375 5865 27495 5985
rect 27550 5865 27670 5985
rect 27715 5865 27835 5985
rect 27880 5865 28000 5985
rect 28045 5865 28165 5985
rect 28220 5865 28340 5985
rect 28385 5865 28505 5985
rect 28550 5865 28670 5985
rect 28715 5865 28835 5985
rect 28890 5865 29010 5985
rect 29055 5865 29175 5985
rect 29220 5865 29340 5985
rect 29385 5865 29505 5985
rect 29560 5865 29680 5985
rect 24200 5700 24320 5820
rect 24365 5700 24485 5820
rect 24530 5700 24650 5820
rect 24695 5700 24815 5820
rect 24870 5700 24990 5820
rect 25035 5700 25155 5820
rect 25200 5700 25320 5820
rect 25365 5700 25485 5820
rect 25540 5700 25660 5820
rect 25705 5700 25825 5820
rect 25870 5700 25990 5820
rect 26035 5700 26155 5820
rect 26210 5700 26330 5820
rect 26375 5700 26495 5820
rect 26540 5700 26660 5820
rect 26705 5700 26825 5820
rect 26880 5700 27000 5820
rect 27045 5700 27165 5820
rect 27210 5700 27330 5820
rect 27375 5700 27495 5820
rect 27550 5700 27670 5820
rect 27715 5700 27835 5820
rect 27880 5700 28000 5820
rect 28045 5700 28165 5820
rect 28220 5700 28340 5820
rect 28385 5700 28505 5820
rect 28550 5700 28670 5820
rect 28715 5700 28835 5820
rect 28890 5700 29010 5820
rect 29055 5700 29175 5820
rect 29220 5700 29340 5820
rect 29385 5700 29505 5820
rect 29560 5700 29680 5820
rect 24200 5525 24320 5645
rect 24365 5525 24485 5645
rect 24530 5525 24650 5645
rect 24695 5525 24815 5645
rect 24870 5525 24990 5645
rect 25035 5525 25155 5645
rect 25200 5525 25320 5645
rect 25365 5525 25485 5645
rect 25540 5525 25660 5645
rect 25705 5525 25825 5645
rect 25870 5525 25990 5645
rect 26035 5525 26155 5645
rect 26210 5525 26330 5645
rect 26375 5525 26495 5645
rect 26540 5525 26660 5645
rect 26705 5525 26825 5645
rect 26880 5525 27000 5645
rect 27045 5525 27165 5645
rect 27210 5525 27330 5645
rect 27375 5525 27495 5645
rect 27550 5525 27670 5645
rect 27715 5525 27835 5645
rect 27880 5525 28000 5645
rect 28045 5525 28165 5645
rect 28220 5525 28340 5645
rect 28385 5525 28505 5645
rect 28550 5525 28670 5645
rect 28715 5525 28835 5645
rect 28890 5525 29010 5645
rect 29055 5525 29175 5645
rect 29220 5525 29340 5645
rect 29385 5525 29505 5645
rect 29560 5525 29680 5645
rect 24200 5360 24320 5480
rect 24365 5360 24485 5480
rect 24530 5360 24650 5480
rect 24695 5360 24815 5480
rect 24870 5360 24990 5480
rect 25035 5360 25155 5480
rect 25200 5360 25320 5480
rect 25365 5360 25485 5480
rect 25540 5360 25660 5480
rect 25705 5360 25825 5480
rect 25870 5360 25990 5480
rect 26035 5360 26155 5480
rect 26210 5360 26330 5480
rect 26375 5360 26495 5480
rect 26540 5360 26660 5480
rect 26705 5360 26825 5480
rect 26880 5360 27000 5480
rect 27045 5360 27165 5480
rect 27210 5360 27330 5480
rect 27375 5360 27495 5480
rect 27550 5360 27670 5480
rect 27715 5360 27835 5480
rect 27880 5360 28000 5480
rect 28045 5360 28165 5480
rect 28220 5360 28340 5480
rect 28385 5360 28505 5480
rect 28550 5360 28670 5480
rect 28715 5360 28835 5480
rect 28890 5360 29010 5480
rect 29055 5360 29175 5480
rect 29220 5360 29340 5480
rect 29385 5360 29505 5480
rect 29560 5360 29680 5480
rect 24200 5195 24320 5315
rect 24365 5195 24485 5315
rect 24530 5195 24650 5315
rect 24695 5195 24815 5315
rect 24870 5195 24990 5315
rect 25035 5195 25155 5315
rect 25200 5195 25320 5315
rect 25365 5195 25485 5315
rect 25540 5195 25660 5315
rect 25705 5195 25825 5315
rect 25870 5195 25990 5315
rect 26035 5195 26155 5315
rect 26210 5195 26330 5315
rect 26375 5195 26495 5315
rect 26540 5195 26660 5315
rect 26705 5195 26825 5315
rect 26880 5195 27000 5315
rect 27045 5195 27165 5315
rect 27210 5195 27330 5315
rect 27375 5195 27495 5315
rect 27550 5195 27670 5315
rect 27715 5195 27835 5315
rect 27880 5195 28000 5315
rect 28045 5195 28165 5315
rect 28220 5195 28340 5315
rect 28385 5195 28505 5315
rect 28550 5195 28670 5315
rect 28715 5195 28835 5315
rect 28890 5195 29010 5315
rect 29055 5195 29175 5315
rect 29220 5195 29340 5315
rect 29385 5195 29505 5315
rect 29560 5195 29680 5315
rect 24200 5030 24320 5150
rect 24365 5030 24485 5150
rect 24530 5030 24650 5150
rect 24695 5030 24815 5150
rect 24870 5030 24990 5150
rect 25035 5030 25155 5150
rect 25200 5030 25320 5150
rect 25365 5030 25485 5150
rect 25540 5030 25660 5150
rect 25705 5030 25825 5150
rect 25870 5030 25990 5150
rect 26035 5030 26155 5150
rect 26210 5030 26330 5150
rect 26375 5030 26495 5150
rect 26540 5030 26660 5150
rect 26705 5030 26825 5150
rect 26880 5030 27000 5150
rect 27045 5030 27165 5150
rect 27210 5030 27330 5150
rect 27375 5030 27495 5150
rect 27550 5030 27670 5150
rect 27715 5030 27835 5150
rect 27880 5030 28000 5150
rect 28045 5030 28165 5150
rect 28220 5030 28340 5150
rect 28385 5030 28505 5150
rect 28550 5030 28670 5150
rect 28715 5030 28835 5150
rect 28890 5030 29010 5150
rect 29055 5030 29175 5150
rect 29220 5030 29340 5150
rect 29385 5030 29505 5150
rect 29560 5030 29680 5150
rect 24200 4855 24320 4975
rect 24365 4855 24485 4975
rect 24530 4855 24650 4975
rect 24695 4855 24815 4975
rect 24870 4855 24990 4975
rect 25035 4855 25155 4975
rect 25200 4855 25320 4975
rect 25365 4855 25485 4975
rect 25540 4855 25660 4975
rect 25705 4855 25825 4975
rect 25870 4855 25990 4975
rect 26035 4855 26155 4975
rect 26210 4855 26330 4975
rect 26375 4855 26495 4975
rect 26540 4855 26660 4975
rect 26705 4855 26825 4975
rect 26880 4855 27000 4975
rect 27045 4855 27165 4975
rect 27210 4855 27330 4975
rect 27375 4855 27495 4975
rect 27550 4855 27670 4975
rect 27715 4855 27835 4975
rect 27880 4855 28000 4975
rect 28045 4855 28165 4975
rect 28220 4855 28340 4975
rect 28385 4855 28505 4975
rect 28550 4855 28670 4975
rect 28715 4855 28835 4975
rect 28890 4855 29010 4975
rect 29055 4855 29175 4975
rect 29220 4855 29340 4975
rect 29385 4855 29505 4975
rect 29560 4855 29680 4975
rect 24200 4690 24320 4810
rect 24365 4690 24485 4810
rect 24530 4690 24650 4810
rect 24695 4690 24815 4810
rect 24870 4690 24990 4810
rect 25035 4690 25155 4810
rect 25200 4690 25320 4810
rect 25365 4690 25485 4810
rect 25540 4690 25660 4810
rect 25705 4690 25825 4810
rect 25870 4690 25990 4810
rect 26035 4690 26155 4810
rect 26210 4690 26330 4810
rect 26375 4690 26495 4810
rect 26540 4690 26660 4810
rect 26705 4690 26825 4810
rect 26880 4690 27000 4810
rect 27045 4690 27165 4810
rect 27210 4690 27330 4810
rect 27375 4690 27495 4810
rect 27550 4690 27670 4810
rect 27715 4690 27835 4810
rect 27880 4690 28000 4810
rect 28045 4690 28165 4810
rect 28220 4690 28340 4810
rect 28385 4690 28505 4810
rect 28550 4690 28670 4810
rect 28715 4690 28835 4810
rect 28890 4690 29010 4810
rect 29055 4690 29175 4810
rect 29220 4690 29340 4810
rect 29385 4690 29505 4810
rect 29560 4690 29680 4810
rect 24200 4525 24320 4645
rect 24365 4525 24485 4645
rect 24530 4525 24650 4645
rect 24695 4525 24815 4645
rect 24870 4525 24990 4645
rect 25035 4525 25155 4645
rect 25200 4525 25320 4645
rect 25365 4525 25485 4645
rect 25540 4525 25660 4645
rect 25705 4525 25825 4645
rect 25870 4525 25990 4645
rect 26035 4525 26155 4645
rect 26210 4525 26330 4645
rect 26375 4525 26495 4645
rect 26540 4525 26660 4645
rect 26705 4525 26825 4645
rect 26880 4525 27000 4645
rect 27045 4525 27165 4645
rect 27210 4525 27330 4645
rect 27375 4525 27495 4645
rect 27550 4525 27670 4645
rect 27715 4525 27835 4645
rect 27880 4525 28000 4645
rect 28045 4525 28165 4645
rect 28220 4525 28340 4645
rect 28385 4525 28505 4645
rect 28550 4525 28670 4645
rect 28715 4525 28835 4645
rect 28890 4525 29010 4645
rect 29055 4525 29175 4645
rect 29220 4525 29340 4645
rect 29385 4525 29505 4645
rect 29560 4525 29680 4645
rect 24200 4360 24320 4480
rect 24365 4360 24485 4480
rect 24530 4360 24650 4480
rect 24695 4360 24815 4480
rect 24870 4360 24990 4480
rect 25035 4360 25155 4480
rect 25200 4360 25320 4480
rect 25365 4360 25485 4480
rect 25540 4360 25660 4480
rect 25705 4360 25825 4480
rect 25870 4360 25990 4480
rect 26035 4360 26155 4480
rect 26210 4360 26330 4480
rect 26375 4360 26495 4480
rect 26540 4360 26660 4480
rect 26705 4360 26825 4480
rect 26880 4360 27000 4480
rect 27045 4360 27165 4480
rect 27210 4360 27330 4480
rect 27375 4360 27495 4480
rect 27550 4360 27670 4480
rect 27715 4360 27835 4480
rect 27880 4360 28000 4480
rect 28045 4360 28165 4480
rect 28220 4360 28340 4480
rect 28385 4360 28505 4480
rect 28550 4360 28670 4480
rect 28715 4360 28835 4480
rect 28890 4360 29010 4480
rect 29055 4360 29175 4480
rect 29220 4360 29340 4480
rect 29385 4360 29505 4480
rect 29560 4360 29680 4480
rect 24200 4185 24320 4305
rect 24365 4185 24485 4305
rect 24530 4185 24650 4305
rect 24695 4185 24815 4305
rect 24870 4185 24990 4305
rect 25035 4185 25155 4305
rect 25200 4185 25320 4305
rect 25365 4185 25485 4305
rect 25540 4185 25660 4305
rect 25705 4185 25825 4305
rect 25870 4185 25990 4305
rect 26035 4185 26155 4305
rect 26210 4185 26330 4305
rect 26375 4185 26495 4305
rect 26540 4185 26660 4305
rect 26705 4185 26825 4305
rect 26880 4185 27000 4305
rect 27045 4185 27165 4305
rect 27210 4185 27330 4305
rect 27375 4185 27495 4305
rect 27550 4185 27670 4305
rect 27715 4185 27835 4305
rect 27880 4185 28000 4305
rect 28045 4185 28165 4305
rect 28220 4185 28340 4305
rect 28385 4185 28505 4305
rect 28550 4185 28670 4305
rect 28715 4185 28835 4305
rect 28890 4185 29010 4305
rect 29055 4185 29175 4305
rect 29220 4185 29340 4305
rect 29385 4185 29505 4305
rect 29560 4185 29680 4305
rect 24200 4020 24320 4140
rect 24365 4020 24485 4140
rect 24530 4020 24650 4140
rect 24695 4020 24815 4140
rect 24870 4020 24990 4140
rect 25035 4020 25155 4140
rect 25200 4020 25320 4140
rect 25365 4020 25485 4140
rect 25540 4020 25660 4140
rect 25705 4020 25825 4140
rect 25870 4020 25990 4140
rect 26035 4020 26155 4140
rect 26210 4020 26330 4140
rect 26375 4020 26495 4140
rect 26540 4020 26660 4140
rect 26705 4020 26825 4140
rect 26880 4020 27000 4140
rect 27045 4020 27165 4140
rect 27210 4020 27330 4140
rect 27375 4020 27495 4140
rect 27550 4020 27670 4140
rect 27715 4020 27835 4140
rect 27880 4020 28000 4140
rect 28045 4020 28165 4140
rect 28220 4020 28340 4140
rect 28385 4020 28505 4140
rect 28550 4020 28670 4140
rect 28715 4020 28835 4140
rect 28890 4020 29010 4140
rect 29055 4020 29175 4140
rect 29220 4020 29340 4140
rect 29385 4020 29505 4140
rect 29560 4020 29680 4140
rect 24200 3855 24320 3975
rect 24365 3855 24485 3975
rect 24530 3855 24650 3975
rect 24695 3855 24815 3975
rect 24870 3855 24990 3975
rect 25035 3855 25155 3975
rect 25200 3855 25320 3975
rect 25365 3855 25485 3975
rect 25540 3855 25660 3975
rect 25705 3855 25825 3975
rect 25870 3855 25990 3975
rect 26035 3855 26155 3975
rect 26210 3855 26330 3975
rect 26375 3855 26495 3975
rect 26540 3855 26660 3975
rect 26705 3855 26825 3975
rect 26880 3855 27000 3975
rect 27045 3855 27165 3975
rect 27210 3855 27330 3975
rect 27375 3855 27495 3975
rect 27550 3855 27670 3975
rect 27715 3855 27835 3975
rect 27880 3855 28000 3975
rect 28045 3855 28165 3975
rect 28220 3855 28340 3975
rect 28385 3855 28505 3975
rect 28550 3855 28670 3975
rect 28715 3855 28835 3975
rect 28890 3855 29010 3975
rect 29055 3855 29175 3975
rect 29220 3855 29340 3975
rect 29385 3855 29505 3975
rect 29560 3855 29680 3975
rect 24200 3690 24320 3810
rect 24365 3690 24485 3810
rect 24530 3690 24650 3810
rect 24695 3690 24815 3810
rect 24870 3690 24990 3810
rect 25035 3690 25155 3810
rect 25200 3690 25320 3810
rect 25365 3690 25485 3810
rect 25540 3690 25660 3810
rect 25705 3690 25825 3810
rect 25870 3690 25990 3810
rect 26035 3690 26155 3810
rect 26210 3690 26330 3810
rect 26375 3690 26495 3810
rect 26540 3690 26660 3810
rect 26705 3690 26825 3810
rect 26880 3690 27000 3810
rect 27045 3690 27165 3810
rect 27210 3690 27330 3810
rect 27375 3690 27495 3810
rect 27550 3690 27670 3810
rect 27715 3690 27835 3810
rect 27880 3690 28000 3810
rect 28045 3690 28165 3810
rect 28220 3690 28340 3810
rect 28385 3690 28505 3810
rect 28550 3690 28670 3810
rect 28715 3690 28835 3810
rect 28890 3690 29010 3810
rect 29055 3690 29175 3810
rect 29220 3690 29340 3810
rect 29385 3690 29505 3810
rect 29560 3690 29680 3810
rect 24200 3515 24320 3635
rect 24365 3515 24485 3635
rect 24530 3515 24650 3635
rect 24695 3515 24815 3635
rect 24870 3515 24990 3635
rect 25035 3515 25155 3635
rect 25200 3515 25320 3635
rect 25365 3515 25485 3635
rect 25540 3515 25660 3635
rect 25705 3515 25825 3635
rect 25870 3515 25990 3635
rect 26035 3515 26155 3635
rect 26210 3515 26330 3635
rect 26375 3515 26495 3635
rect 26540 3515 26660 3635
rect 26705 3515 26825 3635
rect 26880 3515 27000 3635
rect 27045 3515 27165 3635
rect 27210 3515 27330 3635
rect 27375 3515 27495 3635
rect 27550 3515 27670 3635
rect 27715 3515 27835 3635
rect 27880 3515 28000 3635
rect 28045 3515 28165 3635
rect 28220 3515 28340 3635
rect 28385 3515 28505 3635
rect 28550 3515 28670 3635
rect 28715 3515 28835 3635
rect 28890 3515 29010 3635
rect 29055 3515 29175 3635
rect 29220 3515 29340 3635
rect 29385 3515 29505 3635
rect 29560 3515 29680 3635
rect 24200 3350 24320 3470
rect 24365 3350 24485 3470
rect 24530 3350 24650 3470
rect 24695 3350 24815 3470
rect 24870 3350 24990 3470
rect 25035 3350 25155 3470
rect 25200 3350 25320 3470
rect 25365 3350 25485 3470
rect 25540 3350 25660 3470
rect 25705 3350 25825 3470
rect 25870 3350 25990 3470
rect 26035 3350 26155 3470
rect 26210 3350 26330 3470
rect 26375 3350 26495 3470
rect 26540 3350 26660 3470
rect 26705 3350 26825 3470
rect 26880 3350 27000 3470
rect 27045 3350 27165 3470
rect 27210 3350 27330 3470
rect 27375 3350 27495 3470
rect 27550 3350 27670 3470
rect 27715 3350 27835 3470
rect 27880 3350 28000 3470
rect 28045 3350 28165 3470
rect 28220 3350 28340 3470
rect 28385 3350 28505 3470
rect 28550 3350 28670 3470
rect 28715 3350 28835 3470
rect 28890 3350 29010 3470
rect 29055 3350 29175 3470
rect 29220 3350 29340 3470
rect 29385 3350 29505 3470
rect 29560 3350 29680 3470
rect 24200 3185 24320 3305
rect 24365 3185 24485 3305
rect 24530 3185 24650 3305
rect 24695 3185 24815 3305
rect 24870 3185 24990 3305
rect 25035 3185 25155 3305
rect 25200 3185 25320 3305
rect 25365 3185 25485 3305
rect 25540 3185 25660 3305
rect 25705 3185 25825 3305
rect 25870 3185 25990 3305
rect 26035 3185 26155 3305
rect 26210 3185 26330 3305
rect 26375 3185 26495 3305
rect 26540 3185 26660 3305
rect 26705 3185 26825 3305
rect 26880 3185 27000 3305
rect 27045 3185 27165 3305
rect 27210 3185 27330 3305
rect 27375 3185 27495 3305
rect 27550 3185 27670 3305
rect 27715 3185 27835 3305
rect 27880 3185 28000 3305
rect 28045 3185 28165 3305
rect 28220 3185 28340 3305
rect 28385 3185 28505 3305
rect 28550 3185 28670 3305
rect 28715 3185 28835 3305
rect 28890 3185 29010 3305
rect 29055 3185 29175 3305
rect 29220 3185 29340 3305
rect 29385 3185 29505 3305
rect 29560 3185 29680 3305
rect 24200 3020 24320 3140
rect 24365 3020 24485 3140
rect 24530 3020 24650 3140
rect 24695 3020 24815 3140
rect 24870 3020 24990 3140
rect 25035 3020 25155 3140
rect 25200 3020 25320 3140
rect 25365 3020 25485 3140
rect 25540 3020 25660 3140
rect 25705 3020 25825 3140
rect 25870 3020 25990 3140
rect 26035 3020 26155 3140
rect 26210 3020 26330 3140
rect 26375 3020 26495 3140
rect 26540 3020 26660 3140
rect 26705 3020 26825 3140
rect 26880 3020 27000 3140
rect 27045 3020 27165 3140
rect 27210 3020 27330 3140
rect 27375 3020 27495 3140
rect 27550 3020 27670 3140
rect 27715 3020 27835 3140
rect 27880 3020 28000 3140
rect 28045 3020 28165 3140
rect 28220 3020 28340 3140
rect 28385 3020 28505 3140
rect 28550 3020 28670 3140
rect 28715 3020 28835 3140
rect 28890 3020 29010 3140
rect 29055 3020 29175 3140
rect 29220 3020 29340 3140
rect 29385 3020 29505 3140
rect 29560 3020 29680 3140
rect 24200 2845 24320 2965
rect 24365 2845 24485 2965
rect 24530 2845 24650 2965
rect 24695 2845 24815 2965
rect 24870 2845 24990 2965
rect 25035 2845 25155 2965
rect 25200 2845 25320 2965
rect 25365 2845 25485 2965
rect 25540 2845 25660 2965
rect 25705 2845 25825 2965
rect 25870 2845 25990 2965
rect 26035 2845 26155 2965
rect 26210 2845 26330 2965
rect 26375 2845 26495 2965
rect 26540 2845 26660 2965
rect 26705 2845 26825 2965
rect 26880 2845 27000 2965
rect 27045 2845 27165 2965
rect 27210 2845 27330 2965
rect 27375 2845 27495 2965
rect 27550 2845 27670 2965
rect 27715 2845 27835 2965
rect 27880 2845 28000 2965
rect 28045 2845 28165 2965
rect 28220 2845 28340 2965
rect 28385 2845 28505 2965
rect 28550 2845 28670 2965
rect 28715 2845 28835 2965
rect 28890 2845 29010 2965
rect 29055 2845 29175 2965
rect 29220 2845 29340 2965
rect 29385 2845 29505 2965
rect 29560 2845 29680 2965
rect 24200 2680 24320 2800
rect 24365 2680 24485 2800
rect 24530 2680 24650 2800
rect 24695 2680 24815 2800
rect 24870 2680 24990 2800
rect 25035 2680 25155 2800
rect 25200 2680 25320 2800
rect 25365 2680 25485 2800
rect 25540 2680 25660 2800
rect 25705 2680 25825 2800
rect 25870 2680 25990 2800
rect 26035 2680 26155 2800
rect 26210 2680 26330 2800
rect 26375 2680 26495 2800
rect 26540 2680 26660 2800
rect 26705 2680 26825 2800
rect 26880 2680 27000 2800
rect 27045 2680 27165 2800
rect 27210 2680 27330 2800
rect 27375 2680 27495 2800
rect 27550 2680 27670 2800
rect 27715 2680 27835 2800
rect 27880 2680 28000 2800
rect 28045 2680 28165 2800
rect 28220 2680 28340 2800
rect 28385 2680 28505 2800
rect 28550 2680 28670 2800
rect 28715 2680 28835 2800
rect 28890 2680 29010 2800
rect 29055 2680 29175 2800
rect 29220 2680 29340 2800
rect 29385 2680 29505 2800
rect 29560 2680 29680 2800
rect 24200 2515 24320 2635
rect 24365 2515 24485 2635
rect 24530 2515 24650 2635
rect 24695 2515 24815 2635
rect 24870 2515 24990 2635
rect 25035 2515 25155 2635
rect 25200 2515 25320 2635
rect 25365 2515 25485 2635
rect 25540 2515 25660 2635
rect 25705 2515 25825 2635
rect 25870 2515 25990 2635
rect 26035 2515 26155 2635
rect 26210 2515 26330 2635
rect 26375 2515 26495 2635
rect 26540 2515 26660 2635
rect 26705 2515 26825 2635
rect 26880 2515 27000 2635
rect 27045 2515 27165 2635
rect 27210 2515 27330 2635
rect 27375 2515 27495 2635
rect 27550 2515 27670 2635
rect 27715 2515 27835 2635
rect 27880 2515 28000 2635
rect 28045 2515 28165 2635
rect 28220 2515 28340 2635
rect 28385 2515 28505 2635
rect 28550 2515 28670 2635
rect 28715 2515 28835 2635
rect 28890 2515 29010 2635
rect 29055 2515 29175 2635
rect 29220 2515 29340 2635
rect 29385 2515 29505 2635
rect 29560 2515 29680 2635
rect 24200 2350 24320 2470
rect 24365 2350 24485 2470
rect 24530 2350 24650 2470
rect 24695 2350 24815 2470
rect 24870 2350 24990 2470
rect 25035 2350 25155 2470
rect 25200 2350 25320 2470
rect 25365 2350 25485 2470
rect 25540 2350 25660 2470
rect 25705 2350 25825 2470
rect 25870 2350 25990 2470
rect 26035 2350 26155 2470
rect 26210 2350 26330 2470
rect 26375 2350 26495 2470
rect 26540 2350 26660 2470
rect 26705 2350 26825 2470
rect 26880 2350 27000 2470
rect 27045 2350 27165 2470
rect 27210 2350 27330 2470
rect 27375 2350 27495 2470
rect 27550 2350 27670 2470
rect 27715 2350 27835 2470
rect 27880 2350 28000 2470
rect 28045 2350 28165 2470
rect 28220 2350 28340 2470
rect 28385 2350 28505 2470
rect 28550 2350 28670 2470
rect 28715 2350 28835 2470
rect 28890 2350 29010 2470
rect 29055 2350 29175 2470
rect 29220 2350 29340 2470
rect 29385 2350 29505 2470
rect 29560 2350 29680 2470
rect 24200 2175 24320 2295
rect 24365 2175 24485 2295
rect 24530 2175 24650 2295
rect 24695 2175 24815 2295
rect 24870 2175 24990 2295
rect 25035 2175 25155 2295
rect 25200 2175 25320 2295
rect 25365 2175 25485 2295
rect 25540 2175 25660 2295
rect 25705 2175 25825 2295
rect 25870 2175 25990 2295
rect 26035 2175 26155 2295
rect 26210 2175 26330 2295
rect 26375 2175 26495 2295
rect 26540 2175 26660 2295
rect 26705 2175 26825 2295
rect 26880 2175 27000 2295
rect 27045 2175 27165 2295
rect 27210 2175 27330 2295
rect 27375 2175 27495 2295
rect 27550 2175 27670 2295
rect 27715 2175 27835 2295
rect 27880 2175 28000 2295
rect 28045 2175 28165 2295
rect 28220 2175 28340 2295
rect 28385 2175 28505 2295
rect 28550 2175 28670 2295
rect 28715 2175 28835 2295
rect 28890 2175 29010 2295
rect 29055 2175 29175 2295
rect 29220 2175 29340 2295
rect 29385 2175 29505 2295
rect 29560 2175 29680 2295
rect 24200 2010 24320 2130
rect 24365 2010 24485 2130
rect 24530 2010 24650 2130
rect 24695 2010 24815 2130
rect 24870 2010 24990 2130
rect 25035 2010 25155 2130
rect 25200 2010 25320 2130
rect 25365 2010 25485 2130
rect 25540 2010 25660 2130
rect 25705 2010 25825 2130
rect 25870 2010 25990 2130
rect 26035 2010 26155 2130
rect 26210 2010 26330 2130
rect 26375 2010 26495 2130
rect 26540 2010 26660 2130
rect 26705 2010 26825 2130
rect 26880 2010 27000 2130
rect 27045 2010 27165 2130
rect 27210 2010 27330 2130
rect 27375 2010 27495 2130
rect 27550 2010 27670 2130
rect 27715 2010 27835 2130
rect 27880 2010 28000 2130
rect 28045 2010 28165 2130
rect 28220 2010 28340 2130
rect 28385 2010 28505 2130
rect 28550 2010 28670 2130
rect 28715 2010 28835 2130
rect 28890 2010 29010 2130
rect 29055 2010 29175 2130
rect 29220 2010 29340 2130
rect 29385 2010 29505 2130
rect 29560 2010 29680 2130
rect 24200 1845 24320 1965
rect 24365 1845 24485 1965
rect 24530 1845 24650 1965
rect 24695 1845 24815 1965
rect 24870 1845 24990 1965
rect 25035 1845 25155 1965
rect 25200 1845 25320 1965
rect 25365 1845 25485 1965
rect 25540 1845 25660 1965
rect 25705 1845 25825 1965
rect 25870 1845 25990 1965
rect 26035 1845 26155 1965
rect 26210 1845 26330 1965
rect 26375 1845 26495 1965
rect 26540 1845 26660 1965
rect 26705 1845 26825 1965
rect 26880 1845 27000 1965
rect 27045 1845 27165 1965
rect 27210 1845 27330 1965
rect 27375 1845 27495 1965
rect 27550 1845 27670 1965
rect 27715 1845 27835 1965
rect 27880 1845 28000 1965
rect 28045 1845 28165 1965
rect 28220 1845 28340 1965
rect 28385 1845 28505 1965
rect 28550 1845 28670 1965
rect 28715 1845 28835 1965
rect 28890 1845 29010 1965
rect 29055 1845 29175 1965
rect 29220 1845 29340 1965
rect 29385 1845 29505 1965
rect 29560 1845 29680 1965
rect 24200 1680 24320 1800
rect 24365 1680 24485 1800
rect 24530 1680 24650 1800
rect 24695 1680 24815 1800
rect 24870 1680 24990 1800
rect 25035 1680 25155 1800
rect 25200 1680 25320 1800
rect 25365 1680 25485 1800
rect 25540 1680 25660 1800
rect 25705 1680 25825 1800
rect 25870 1680 25990 1800
rect 26035 1680 26155 1800
rect 26210 1680 26330 1800
rect 26375 1680 26495 1800
rect 26540 1680 26660 1800
rect 26705 1680 26825 1800
rect 26880 1680 27000 1800
rect 27045 1680 27165 1800
rect 27210 1680 27330 1800
rect 27375 1680 27495 1800
rect 27550 1680 27670 1800
rect 27715 1680 27835 1800
rect 27880 1680 28000 1800
rect 28045 1680 28165 1800
rect 28220 1680 28340 1800
rect 28385 1680 28505 1800
rect 28550 1680 28670 1800
rect 28715 1680 28835 1800
rect 28890 1680 29010 1800
rect 29055 1680 29175 1800
rect 29220 1680 29340 1800
rect 29385 1680 29505 1800
rect 29560 1680 29680 1800
rect 7130 1260 7250 1380
rect 7305 1260 7425 1380
rect 7470 1260 7590 1380
rect 7635 1260 7755 1380
rect 7800 1260 7920 1380
rect 7975 1260 8095 1380
rect 8140 1260 8260 1380
rect 8305 1260 8425 1380
rect 8470 1260 8590 1380
rect 8645 1260 8765 1380
rect 8810 1260 8930 1380
rect 8975 1260 9095 1380
rect 9140 1260 9260 1380
rect 9315 1260 9435 1380
rect 9480 1260 9600 1380
rect 9645 1260 9765 1380
rect 9810 1260 9930 1380
rect 9985 1260 10105 1380
rect 10150 1260 10270 1380
rect 10315 1260 10435 1380
rect 10480 1260 10600 1380
rect 10655 1260 10775 1380
rect 10820 1260 10940 1380
rect 10985 1260 11105 1380
rect 11150 1260 11270 1380
rect 11325 1260 11445 1380
rect 11490 1260 11610 1380
rect 11655 1260 11775 1380
rect 11820 1260 11940 1380
rect 11995 1260 12115 1380
rect 12160 1260 12280 1380
rect 12325 1260 12445 1380
rect 12490 1260 12610 1380
rect 7130 1095 7250 1215
rect 7305 1095 7425 1215
rect 7470 1095 7590 1215
rect 7635 1095 7755 1215
rect 7800 1095 7920 1215
rect 7975 1095 8095 1215
rect 8140 1095 8260 1215
rect 8305 1095 8425 1215
rect 8470 1095 8590 1215
rect 8645 1095 8765 1215
rect 8810 1095 8930 1215
rect 8975 1095 9095 1215
rect 9140 1095 9260 1215
rect 9315 1095 9435 1215
rect 9480 1095 9600 1215
rect 9645 1095 9765 1215
rect 9810 1095 9930 1215
rect 9985 1095 10105 1215
rect 10150 1095 10270 1215
rect 10315 1095 10435 1215
rect 10480 1095 10600 1215
rect 10655 1095 10775 1215
rect 10820 1095 10940 1215
rect 10985 1095 11105 1215
rect 11150 1095 11270 1215
rect 11325 1095 11445 1215
rect 11490 1095 11610 1215
rect 11655 1095 11775 1215
rect 11820 1095 11940 1215
rect 11995 1095 12115 1215
rect 12160 1095 12280 1215
rect 12325 1095 12445 1215
rect 12490 1095 12610 1215
rect 7130 930 7250 1050
rect 7305 930 7425 1050
rect 7470 930 7590 1050
rect 7635 930 7755 1050
rect 7800 930 7920 1050
rect 7975 930 8095 1050
rect 8140 930 8260 1050
rect 8305 930 8425 1050
rect 8470 930 8590 1050
rect 8645 930 8765 1050
rect 8810 930 8930 1050
rect 8975 930 9095 1050
rect 9140 930 9260 1050
rect 9315 930 9435 1050
rect 9480 930 9600 1050
rect 9645 930 9765 1050
rect 9810 930 9930 1050
rect 9985 930 10105 1050
rect 10150 930 10270 1050
rect 10315 930 10435 1050
rect 10480 930 10600 1050
rect 10655 930 10775 1050
rect 10820 930 10940 1050
rect 10985 930 11105 1050
rect 11150 930 11270 1050
rect 11325 930 11445 1050
rect 11490 930 11610 1050
rect 11655 930 11775 1050
rect 11820 930 11940 1050
rect 11995 930 12115 1050
rect 12160 930 12280 1050
rect 12325 930 12445 1050
rect 12490 930 12610 1050
rect 7130 765 7250 885
rect 7305 765 7425 885
rect 7470 765 7590 885
rect 7635 765 7755 885
rect 7800 765 7920 885
rect 7975 765 8095 885
rect 8140 765 8260 885
rect 8305 765 8425 885
rect 8470 765 8590 885
rect 8645 765 8765 885
rect 8810 765 8930 885
rect 8975 765 9095 885
rect 9140 765 9260 885
rect 9315 765 9435 885
rect 9480 765 9600 885
rect 9645 765 9765 885
rect 9810 765 9930 885
rect 9985 765 10105 885
rect 10150 765 10270 885
rect 10315 765 10435 885
rect 10480 765 10600 885
rect 10655 765 10775 885
rect 10820 765 10940 885
rect 10985 765 11105 885
rect 11150 765 11270 885
rect 11325 765 11445 885
rect 11490 765 11610 885
rect 11655 765 11775 885
rect 11820 765 11940 885
rect 11995 765 12115 885
rect 12160 765 12280 885
rect 12325 765 12445 885
rect 12490 765 12610 885
rect 7130 590 7250 710
rect 7305 590 7425 710
rect 7470 590 7590 710
rect 7635 590 7755 710
rect 7800 590 7920 710
rect 7975 590 8095 710
rect 8140 590 8260 710
rect 8305 590 8425 710
rect 8470 590 8590 710
rect 8645 590 8765 710
rect 8810 590 8930 710
rect 8975 590 9095 710
rect 9140 590 9260 710
rect 9315 590 9435 710
rect 9480 590 9600 710
rect 9645 590 9765 710
rect 9810 590 9930 710
rect 9985 590 10105 710
rect 10150 590 10270 710
rect 10315 590 10435 710
rect 10480 590 10600 710
rect 10655 590 10775 710
rect 10820 590 10940 710
rect 10985 590 11105 710
rect 11150 590 11270 710
rect 11325 590 11445 710
rect 11490 590 11610 710
rect 11655 590 11775 710
rect 11820 590 11940 710
rect 11995 590 12115 710
rect 12160 590 12280 710
rect 12325 590 12445 710
rect 12490 590 12610 710
rect 7130 425 7250 545
rect 7305 425 7425 545
rect 7470 425 7590 545
rect 7635 425 7755 545
rect 7800 425 7920 545
rect 7975 425 8095 545
rect 8140 425 8260 545
rect 8305 425 8425 545
rect 8470 425 8590 545
rect 8645 425 8765 545
rect 8810 425 8930 545
rect 8975 425 9095 545
rect 9140 425 9260 545
rect 9315 425 9435 545
rect 9480 425 9600 545
rect 9645 425 9765 545
rect 9810 425 9930 545
rect 9985 425 10105 545
rect 10150 425 10270 545
rect 10315 425 10435 545
rect 10480 425 10600 545
rect 10655 425 10775 545
rect 10820 425 10940 545
rect 10985 425 11105 545
rect 11150 425 11270 545
rect 11325 425 11445 545
rect 11490 425 11610 545
rect 11655 425 11775 545
rect 11820 425 11940 545
rect 11995 425 12115 545
rect 12160 425 12280 545
rect 12325 425 12445 545
rect 12490 425 12610 545
rect 7130 260 7250 380
rect 7305 260 7425 380
rect 7470 260 7590 380
rect 7635 260 7755 380
rect 7800 260 7920 380
rect 7975 260 8095 380
rect 8140 260 8260 380
rect 8305 260 8425 380
rect 8470 260 8590 380
rect 8645 260 8765 380
rect 8810 260 8930 380
rect 8975 260 9095 380
rect 9140 260 9260 380
rect 9315 260 9435 380
rect 9480 260 9600 380
rect 9645 260 9765 380
rect 9810 260 9930 380
rect 9985 260 10105 380
rect 10150 260 10270 380
rect 10315 260 10435 380
rect 10480 260 10600 380
rect 10655 260 10775 380
rect 10820 260 10940 380
rect 10985 260 11105 380
rect 11150 260 11270 380
rect 11325 260 11445 380
rect 11490 260 11610 380
rect 11655 260 11775 380
rect 11820 260 11940 380
rect 11995 260 12115 380
rect 12160 260 12280 380
rect 12325 260 12445 380
rect 12490 260 12610 380
rect 7130 95 7250 215
rect 7305 95 7425 215
rect 7470 95 7590 215
rect 7635 95 7755 215
rect 7800 95 7920 215
rect 7975 95 8095 215
rect 8140 95 8260 215
rect 8305 95 8425 215
rect 8470 95 8590 215
rect 8645 95 8765 215
rect 8810 95 8930 215
rect 8975 95 9095 215
rect 9140 95 9260 215
rect 9315 95 9435 215
rect 9480 95 9600 215
rect 9645 95 9765 215
rect 9810 95 9930 215
rect 9985 95 10105 215
rect 10150 95 10270 215
rect 10315 95 10435 215
rect 10480 95 10600 215
rect 10655 95 10775 215
rect 10820 95 10940 215
rect 10985 95 11105 215
rect 11150 95 11270 215
rect 11325 95 11445 215
rect 11490 95 11610 215
rect 11655 95 11775 215
rect 11820 95 11940 215
rect 11995 95 12115 215
rect 12160 95 12280 215
rect 12325 95 12445 215
rect 12490 95 12610 215
rect 7130 -80 7250 40
rect 7305 -80 7425 40
rect 7470 -80 7590 40
rect 7635 -80 7755 40
rect 7800 -80 7920 40
rect 7975 -80 8095 40
rect 8140 -80 8260 40
rect 8305 -80 8425 40
rect 8470 -80 8590 40
rect 8645 -80 8765 40
rect 8810 -80 8930 40
rect 8975 -80 9095 40
rect 9140 -80 9260 40
rect 9315 -80 9435 40
rect 9480 -80 9600 40
rect 9645 -80 9765 40
rect 9810 -80 9930 40
rect 9985 -80 10105 40
rect 10150 -80 10270 40
rect 10315 -80 10435 40
rect 10480 -80 10600 40
rect 10655 -80 10775 40
rect 10820 -80 10940 40
rect 10985 -80 11105 40
rect 11150 -80 11270 40
rect 11325 -80 11445 40
rect 11490 -80 11610 40
rect 11655 -80 11775 40
rect 11820 -80 11940 40
rect 11995 -80 12115 40
rect 12160 -80 12280 40
rect 12325 -80 12445 40
rect 12490 -80 12610 40
rect 7130 -245 7250 -125
rect 7305 -245 7425 -125
rect 7470 -245 7590 -125
rect 7635 -245 7755 -125
rect 7800 -245 7920 -125
rect 7975 -245 8095 -125
rect 8140 -245 8260 -125
rect 8305 -245 8425 -125
rect 8470 -245 8590 -125
rect 8645 -245 8765 -125
rect 8810 -245 8930 -125
rect 8975 -245 9095 -125
rect 9140 -245 9260 -125
rect 9315 -245 9435 -125
rect 9480 -245 9600 -125
rect 9645 -245 9765 -125
rect 9810 -245 9930 -125
rect 9985 -245 10105 -125
rect 10150 -245 10270 -125
rect 10315 -245 10435 -125
rect 10480 -245 10600 -125
rect 10655 -245 10775 -125
rect 10820 -245 10940 -125
rect 10985 -245 11105 -125
rect 11150 -245 11270 -125
rect 11325 -245 11445 -125
rect 11490 -245 11610 -125
rect 11655 -245 11775 -125
rect 11820 -245 11940 -125
rect 11995 -245 12115 -125
rect 12160 -245 12280 -125
rect 12325 -245 12445 -125
rect 12490 -245 12610 -125
rect 7130 -410 7250 -290
rect 7305 -410 7425 -290
rect 7470 -410 7590 -290
rect 7635 -410 7755 -290
rect 7800 -410 7920 -290
rect 7975 -410 8095 -290
rect 8140 -410 8260 -290
rect 8305 -410 8425 -290
rect 8470 -410 8590 -290
rect 8645 -410 8765 -290
rect 8810 -410 8930 -290
rect 8975 -410 9095 -290
rect 9140 -410 9260 -290
rect 9315 -410 9435 -290
rect 9480 -410 9600 -290
rect 9645 -410 9765 -290
rect 9810 -410 9930 -290
rect 9985 -410 10105 -290
rect 10150 -410 10270 -290
rect 10315 -410 10435 -290
rect 10480 -410 10600 -290
rect 10655 -410 10775 -290
rect 10820 -410 10940 -290
rect 10985 -410 11105 -290
rect 11150 -410 11270 -290
rect 11325 -410 11445 -290
rect 11490 -410 11610 -290
rect 11655 -410 11775 -290
rect 11820 -410 11940 -290
rect 11995 -410 12115 -290
rect 12160 -410 12280 -290
rect 12325 -410 12445 -290
rect 12490 -410 12610 -290
rect 7130 -575 7250 -455
rect 7305 -575 7425 -455
rect 7470 -575 7590 -455
rect 7635 -575 7755 -455
rect 7800 -575 7920 -455
rect 7975 -575 8095 -455
rect 8140 -575 8260 -455
rect 8305 -575 8425 -455
rect 8470 -575 8590 -455
rect 8645 -575 8765 -455
rect 8810 -575 8930 -455
rect 8975 -575 9095 -455
rect 9140 -575 9260 -455
rect 9315 -575 9435 -455
rect 9480 -575 9600 -455
rect 9645 -575 9765 -455
rect 9810 -575 9930 -455
rect 9985 -575 10105 -455
rect 10150 -575 10270 -455
rect 10315 -575 10435 -455
rect 10480 -575 10600 -455
rect 10655 -575 10775 -455
rect 10820 -575 10940 -455
rect 10985 -575 11105 -455
rect 11150 -575 11270 -455
rect 11325 -575 11445 -455
rect 11490 -575 11610 -455
rect 11655 -575 11775 -455
rect 11820 -575 11940 -455
rect 11995 -575 12115 -455
rect 12160 -575 12280 -455
rect 12325 -575 12445 -455
rect 12490 -575 12610 -455
rect 7130 -750 7250 -630
rect 7305 -750 7425 -630
rect 7470 -750 7590 -630
rect 7635 -750 7755 -630
rect 7800 -750 7920 -630
rect 7975 -750 8095 -630
rect 8140 -750 8260 -630
rect 8305 -750 8425 -630
rect 8470 -750 8590 -630
rect 8645 -750 8765 -630
rect 8810 -750 8930 -630
rect 8975 -750 9095 -630
rect 9140 -750 9260 -630
rect 9315 -750 9435 -630
rect 9480 -750 9600 -630
rect 9645 -750 9765 -630
rect 9810 -750 9930 -630
rect 9985 -750 10105 -630
rect 10150 -750 10270 -630
rect 10315 -750 10435 -630
rect 10480 -750 10600 -630
rect 10655 -750 10775 -630
rect 10820 -750 10940 -630
rect 10985 -750 11105 -630
rect 11150 -750 11270 -630
rect 11325 -750 11445 -630
rect 11490 -750 11610 -630
rect 11655 -750 11775 -630
rect 11820 -750 11940 -630
rect 11995 -750 12115 -630
rect 12160 -750 12280 -630
rect 12325 -750 12445 -630
rect 12490 -750 12610 -630
rect 7130 -915 7250 -795
rect 7305 -915 7425 -795
rect 7470 -915 7590 -795
rect 7635 -915 7755 -795
rect 7800 -915 7920 -795
rect 7975 -915 8095 -795
rect 8140 -915 8260 -795
rect 8305 -915 8425 -795
rect 8470 -915 8590 -795
rect 8645 -915 8765 -795
rect 8810 -915 8930 -795
rect 8975 -915 9095 -795
rect 9140 -915 9260 -795
rect 9315 -915 9435 -795
rect 9480 -915 9600 -795
rect 9645 -915 9765 -795
rect 9810 -915 9930 -795
rect 9985 -915 10105 -795
rect 10150 -915 10270 -795
rect 10315 -915 10435 -795
rect 10480 -915 10600 -795
rect 10655 -915 10775 -795
rect 10820 -915 10940 -795
rect 10985 -915 11105 -795
rect 11150 -915 11270 -795
rect 11325 -915 11445 -795
rect 11490 -915 11610 -795
rect 11655 -915 11775 -795
rect 11820 -915 11940 -795
rect 11995 -915 12115 -795
rect 12160 -915 12280 -795
rect 12325 -915 12445 -795
rect 12490 -915 12610 -795
rect 7130 -1080 7250 -960
rect 7305 -1080 7425 -960
rect 7470 -1080 7590 -960
rect 7635 -1080 7755 -960
rect 7800 -1080 7920 -960
rect 7975 -1080 8095 -960
rect 8140 -1080 8260 -960
rect 8305 -1080 8425 -960
rect 8470 -1080 8590 -960
rect 8645 -1080 8765 -960
rect 8810 -1080 8930 -960
rect 8975 -1080 9095 -960
rect 9140 -1080 9260 -960
rect 9315 -1080 9435 -960
rect 9480 -1080 9600 -960
rect 9645 -1080 9765 -960
rect 9810 -1080 9930 -960
rect 9985 -1080 10105 -960
rect 10150 -1080 10270 -960
rect 10315 -1080 10435 -960
rect 10480 -1080 10600 -960
rect 10655 -1080 10775 -960
rect 10820 -1080 10940 -960
rect 10985 -1080 11105 -960
rect 11150 -1080 11270 -960
rect 11325 -1080 11445 -960
rect 11490 -1080 11610 -960
rect 11655 -1080 11775 -960
rect 11820 -1080 11940 -960
rect 11995 -1080 12115 -960
rect 12160 -1080 12280 -960
rect 12325 -1080 12445 -960
rect 12490 -1080 12610 -960
rect 7130 -1245 7250 -1125
rect 7305 -1245 7425 -1125
rect 7470 -1245 7590 -1125
rect 7635 -1245 7755 -1125
rect 7800 -1245 7920 -1125
rect 7975 -1245 8095 -1125
rect 8140 -1245 8260 -1125
rect 8305 -1245 8425 -1125
rect 8470 -1245 8590 -1125
rect 8645 -1245 8765 -1125
rect 8810 -1245 8930 -1125
rect 8975 -1245 9095 -1125
rect 9140 -1245 9260 -1125
rect 9315 -1245 9435 -1125
rect 9480 -1245 9600 -1125
rect 9645 -1245 9765 -1125
rect 9810 -1245 9930 -1125
rect 9985 -1245 10105 -1125
rect 10150 -1245 10270 -1125
rect 10315 -1245 10435 -1125
rect 10480 -1245 10600 -1125
rect 10655 -1245 10775 -1125
rect 10820 -1245 10940 -1125
rect 10985 -1245 11105 -1125
rect 11150 -1245 11270 -1125
rect 11325 -1245 11445 -1125
rect 11490 -1245 11610 -1125
rect 11655 -1245 11775 -1125
rect 11820 -1245 11940 -1125
rect 11995 -1245 12115 -1125
rect 12160 -1245 12280 -1125
rect 12325 -1245 12445 -1125
rect 12490 -1245 12610 -1125
rect 7130 -1420 7250 -1300
rect 7305 -1420 7425 -1300
rect 7470 -1420 7590 -1300
rect 7635 -1420 7755 -1300
rect 7800 -1420 7920 -1300
rect 7975 -1420 8095 -1300
rect 8140 -1420 8260 -1300
rect 8305 -1420 8425 -1300
rect 8470 -1420 8590 -1300
rect 8645 -1420 8765 -1300
rect 8810 -1420 8930 -1300
rect 8975 -1420 9095 -1300
rect 9140 -1420 9260 -1300
rect 9315 -1420 9435 -1300
rect 9480 -1420 9600 -1300
rect 9645 -1420 9765 -1300
rect 9810 -1420 9930 -1300
rect 9985 -1420 10105 -1300
rect 10150 -1420 10270 -1300
rect 10315 -1420 10435 -1300
rect 10480 -1420 10600 -1300
rect 10655 -1420 10775 -1300
rect 10820 -1420 10940 -1300
rect 10985 -1420 11105 -1300
rect 11150 -1420 11270 -1300
rect 11325 -1420 11445 -1300
rect 11490 -1420 11610 -1300
rect 11655 -1420 11775 -1300
rect 11820 -1420 11940 -1300
rect 11995 -1420 12115 -1300
rect 12160 -1420 12280 -1300
rect 12325 -1420 12445 -1300
rect 12490 -1420 12610 -1300
rect 7130 -1585 7250 -1465
rect 7305 -1585 7425 -1465
rect 7470 -1585 7590 -1465
rect 7635 -1585 7755 -1465
rect 7800 -1585 7920 -1465
rect 7975 -1585 8095 -1465
rect 8140 -1585 8260 -1465
rect 8305 -1585 8425 -1465
rect 8470 -1585 8590 -1465
rect 8645 -1585 8765 -1465
rect 8810 -1585 8930 -1465
rect 8975 -1585 9095 -1465
rect 9140 -1585 9260 -1465
rect 9315 -1585 9435 -1465
rect 9480 -1585 9600 -1465
rect 9645 -1585 9765 -1465
rect 9810 -1585 9930 -1465
rect 9985 -1585 10105 -1465
rect 10150 -1585 10270 -1465
rect 10315 -1585 10435 -1465
rect 10480 -1585 10600 -1465
rect 10655 -1585 10775 -1465
rect 10820 -1585 10940 -1465
rect 10985 -1585 11105 -1465
rect 11150 -1585 11270 -1465
rect 11325 -1585 11445 -1465
rect 11490 -1585 11610 -1465
rect 11655 -1585 11775 -1465
rect 11820 -1585 11940 -1465
rect 11995 -1585 12115 -1465
rect 12160 -1585 12280 -1465
rect 12325 -1585 12445 -1465
rect 12490 -1585 12610 -1465
rect 7130 -1750 7250 -1630
rect 7305 -1750 7425 -1630
rect 7470 -1750 7590 -1630
rect 7635 -1750 7755 -1630
rect 7800 -1750 7920 -1630
rect 7975 -1750 8095 -1630
rect 8140 -1750 8260 -1630
rect 8305 -1750 8425 -1630
rect 8470 -1750 8590 -1630
rect 8645 -1750 8765 -1630
rect 8810 -1750 8930 -1630
rect 8975 -1750 9095 -1630
rect 9140 -1750 9260 -1630
rect 9315 -1750 9435 -1630
rect 9480 -1750 9600 -1630
rect 9645 -1750 9765 -1630
rect 9810 -1750 9930 -1630
rect 9985 -1750 10105 -1630
rect 10150 -1750 10270 -1630
rect 10315 -1750 10435 -1630
rect 10480 -1750 10600 -1630
rect 10655 -1750 10775 -1630
rect 10820 -1750 10940 -1630
rect 10985 -1750 11105 -1630
rect 11150 -1750 11270 -1630
rect 11325 -1750 11445 -1630
rect 11490 -1750 11610 -1630
rect 11655 -1750 11775 -1630
rect 11820 -1750 11940 -1630
rect 11995 -1750 12115 -1630
rect 12160 -1750 12280 -1630
rect 12325 -1750 12445 -1630
rect 12490 -1750 12610 -1630
rect 7130 -1915 7250 -1795
rect 7305 -1915 7425 -1795
rect 7470 -1915 7590 -1795
rect 7635 -1915 7755 -1795
rect 7800 -1915 7920 -1795
rect 7975 -1915 8095 -1795
rect 8140 -1915 8260 -1795
rect 8305 -1915 8425 -1795
rect 8470 -1915 8590 -1795
rect 8645 -1915 8765 -1795
rect 8810 -1915 8930 -1795
rect 8975 -1915 9095 -1795
rect 9140 -1915 9260 -1795
rect 9315 -1915 9435 -1795
rect 9480 -1915 9600 -1795
rect 9645 -1915 9765 -1795
rect 9810 -1915 9930 -1795
rect 9985 -1915 10105 -1795
rect 10150 -1915 10270 -1795
rect 10315 -1915 10435 -1795
rect 10480 -1915 10600 -1795
rect 10655 -1915 10775 -1795
rect 10820 -1915 10940 -1795
rect 10985 -1915 11105 -1795
rect 11150 -1915 11270 -1795
rect 11325 -1915 11445 -1795
rect 11490 -1915 11610 -1795
rect 11655 -1915 11775 -1795
rect 11820 -1915 11940 -1795
rect 11995 -1915 12115 -1795
rect 12160 -1915 12280 -1795
rect 12325 -1915 12445 -1795
rect 12490 -1915 12610 -1795
rect 7130 -2090 7250 -1970
rect 7305 -2090 7425 -1970
rect 7470 -2090 7590 -1970
rect 7635 -2090 7755 -1970
rect 7800 -2090 7920 -1970
rect 7975 -2090 8095 -1970
rect 8140 -2090 8260 -1970
rect 8305 -2090 8425 -1970
rect 8470 -2090 8590 -1970
rect 8645 -2090 8765 -1970
rect 8810 -2090 8930 -1970
rect 8975 -2090 9095 -1970
rect 9140 -2090 9260 -1970
rect 9315 -2090 9435 -1970
rect 9480 -2090 9600 -1970
rect 9645 -2090 9765 -1970
rect 9810 -2090 9930 -1970
rect 9985 -2090 10105 -1970
rect 10150 -2090 10270 -1970
rect 10315 -2090 10435 -1970
rect 10480 -2090 10600 -1970
rect 10655 -2090 10775 -1970
rect 10820 -2090 10940 -1970
rect 10985 -2090 11105 -1970
rect 11150 -2090 11270 -1970
rect 11325 -2090 11445 -1970
rect 11490 -2090 11610 -1970
rect 11655 -2090 11775 -1970
rect 11820 -2090 11940 -1970
rect 11995 -2090 12115 -1970
rect 12160 -2090 12280 -1970
rect 12325 -2090 12445 -1970
rect 12490 -2090 12610 -1970
rect 7130 -2255 7250 -2135
rect 7305 -2255 7425 -2135
rect 7470 -2255 7590 -2135
rect 7635 -2255 7755 -2135
rect 7800 -2255 7920 -2135
rect 7975 -2255 8095 -2135
rect 8140 -2255 8260 -2135
rect 8305 -2255 8425 -2135
rect 8470 -2255 8590 -2135
rect 8645 -2255 8765 -2135
rect 8810 -2255 8930 -2135
rect 8975 -2255 9095 -2135
rect 9140 -2255 9260 -2135
rect 9315 -2255 9435 -2135
rect 9480 -2255 9600 -2135
rect 9645 -2255 9765 -2135
rect 9810 -2255 9930 -2135
rect 9985 -2255 10105 -2135
rect 10150 -2255 10270 -2135
rect 10315 -2255 10435 -2135
rect 10480 -2255 10600 -2135
rect 10655 -2255 10775 -2135
rect 10820 -2255 10940 -2135
rect 10985 -2255 11105 -2135
rect 11150 -2255 11270 -2135
rect 11325 -2255 11445 -2135
rect 11490 -2255 11610 -2135
rect 11655 -2255 11775 -2135
rect 11820 -2255 11940 -2135
rect 11995 -2255 12115 -2135
rect 12160 -2255 12280 -2135
rect 12325 -2255 12445 -2135
rect 12490 -2255 12610 -2135
rect 7130 -2420 7250 -2300
rect 7305 -2420 7425 -2300
rect 7470 -2420 7590 -2300
rect 7635 -2420 7755 -2300
rect 7800 -2420 7920 -2300
rect 7975 -2420 8095 -2300
rect 8140 -2420 8260 -2300
rect 8305 -2420 8425 -2300
rect 8470 -2420 8590 -2300
rect 8645 -2420 8765 -2300
rect 8810 -2420 8930 -2300
rect 8975 -2420 9095 -2300
rect 9140 -2420 9260 -2300
rect 9315 -2420 9435 -2300
rect 9480 -2420 9600 -2300
rect 9645 -2420 9765 -2300
rect 9810 -2420 9930 -2300
rect 9985 -2420 10105 -2300
rect 10150 -2420 10270 -2300
rect 10315 -2420 10435 -2300
rect 10480 -2420 10600 -2300
rect 10655 -2420 10775 -2300
rect 10820 -2420 10940 -2300
rect 10985 -2420 11105 -2300
rect 11150 -2420 11270 -2300
rect 11325 -2420 11445 -2300
rect 11490 -2420 11610 -2300
rect 11655 -2420 11775 -2300
rect 11820 -2420 11940 -2300
rect 11995 -2420 12115 -2300
rect 12160 -2420 12280 -2300
rect 12325 -2420 12445 -2300
rect 12490 -2420 12610 -2300
rect 7130 -2585 7250 -2465
rect 7305 -2585 7425 -2465
rect 7470 -2585 7590 -2465
rect 7635 -2585 7755 -2465
rect 7800 -2585 7920 -2465
rect 7975 -2585 8095 -2465
rect 8140 -2585 8260 -2465
rect 8305 -2585 8425 -2465
rect 8470 -2585 8590 -2465
rect 8645 -2585 8765 -2465
rect 8810 -2585 8930 -2465
rect 8975 -2585 9095 -2465
rect 9140 -2585 9260 -2465
rect 9315 -2585 9435 -2465
rect 9480 -2585 9600 -2465
rect 9645 -2585 9765 -2465
rect 9810 -2585 9930 -2465
rect 9985 -2585 10105 -2465
rect 10150 -2585 10270 -2465
rect 10315 -2585 10435 -2465
rect 10480 -2585 10600 -2465
rect 10655 -2585 10775 -2465
rect 10820 -2585 10940 -2465
rect 10985 -2585 11105 -2465
rect 11150 -2585 11270 -2465
rect 11325 -2585 11445 -2465
rect 11490 -2585 11610 -2465
rect 11655 -2585 11775 -2465
rect 11820 -2585 11940 -2465
rect 11995 -2585 12115 -2465
rect 12160 -2585 12280 -2465
rect 12325 -2585 12445 -2465
rect 12490 -2585 12610 -2465
rect 7130 -2760 7250 -2640
rect 7305 -2760 7425 -2640
rect 7470 -2760 7590 -2640
rect 7635 -2760 7755 -2640
rect 7800 -2760 7920 -2640
rect 7975 -2760 8095 -2640
rect 8140 -2760 8260 -2640
rect 8305 -2760 8425 -2640
rect 8470 -2760 8590 -2640
rect 8645 -2760 8765 -2640
rect 8810 -2760 8930 -2640
rect 8975 -2760 9095 -2640
rect 9140 -2760 9260 -2640
rect 9315 -2760 9435 -2640
rect 9480 -2760 9600 -2640
rect 9645 -2760 9765 -2640
rect 9810 -2760 9930 -2640
rect 9985 -2760 10105 -2640
rect 10150 -2760 10270 -2640
rect 10315 -2760 10435 -2640
rect 10480 -2760 10600 -2640
rect 10655 -2760 10775 -2640
rect 10820 -2760 10940 -2640
rect 10985 -2760 11105 -2640
rect 11150 -2760 11270 -2640
rect 11325 -2760 11445 -2640
rect 11490 -2760 11610 -2640
rect 11655 -2760 11775 -2640
rect 11820 -2760 11940 -2640
rect 11995 -2760 12115 -2640
rect 12160 -2760 12280 -2640
rect 12325 -2760 12445 -2640
rect 12490 -2760 12610 -2640
rect 7130 -2925 7250 -2805
rect 7305 -2925 7425 -2805
rect 7470 -2925 7590 -2805
rect 7635 -2925 7755 -2805
rect 7800 -2925 7920 -2805
rect 7975 -2925 8095 -2805
rect 8140 -2925 8260 -2805
rect 8305 -2925 8425 -2805
rect 8470 -2925 8590 -2805
rect 8645 -2925 8765 -2805
rect 8810 -2925 8930 -2805
rect 8975 -2925 9095 -2805
rect 9140 -2925 9260 -2805
rect 9315 -2925 9435 -2805
rect 9480 -2925 9600 -2805
rect 9645 -2925 9765 -2805
rect 9810 -2925 9930 -2805
rect 9985 -2925 10105 -2805
rect 10150 -2925 10270 -2805
rect 10315 -2925 10435 -2805
rect 10480 -2925 10600 -2805
rect 10655 -2925 10775 -2805
rect 10820 -2925 10940 -2805
rect 10985 -2925 11105 -2805
rect 11150 -2925 11270 -2805
rect 11325 -2925 11445 -2805
rect 11490 -2925 11610 -2805
rect 11655 -2925 11775 -2805
rect 11820 -2925 11940 -2805
rect 11995 -2925 12115 -2805
rect 12160 -2925 12280 -2805
rect 12325 -2925 12445 -2805
rect 12490 -2925 12610 -2805
rect 7130 -3090 7250 -2970
rect 7305 -3090 7425 -2970
rect 7470 -3090 7590 -2970
rect 7635 -3090 7755 -2970
rect 7800 -3090 7920 -2970
rect 7975 -3090 8095 -2970
rect 8140 -3090 8260 -2970
rect 8305 -3090 8425 -2970
rect 8470 -3090 8590 -2970
rect 8645 -3090 8765 -2970
rect 8810 -3090 8930 -2970
rect 8975 -3090 9095 -2970
rect 9140 -3090 9260 -2970
rect 9315 -3090 9435 -2970
rect 9480 -3090 9600 -2970
rect 9645 -3090 9765 -2970
rect 9810 -3090 9930 -2970
rect 9985 -3090 10105 -2970
rect 10150 -3090 10270 -2970
rect 10315 -3090 10435 -2970
rect 10480 -3090 10600 -2970
rect 10655 -3090 10775 -2970
rect 10820 -3090 10940 -2970
rect 10985 -3090 11105 -2970
rect 11150 -3090 11270 -2970
rect 11325 -3090 11445 -2970
rect 11490 -3090 11610 -2970
rect 11655 -3090 11775 -2970
rect 11820 -3090 11940 -2970
rect 11995 -3090 12115 -2970
rect 12160 -3090 12280 -2970
rect 12325 -3090 12445 -2970
rect 12490 -3090 12610 -2970
rect 7130 -3255 7250 -3135
rect 7305 -3255 7425 -3135
rect 7470 -3255 7590 -3135
rect 7635 -3255 7755 -3135
rect 7800 -3255 7920 -3135
rect 7975 -3255 8095 -3135
rect 8140 -3255 8260 -3135
rect 8305 -3255 8425 -3135
rect 8470 -3255 8590 -3135
rect 8645 -3255 8765 -3135
rect 8810 -3255 8930 -3135
rect 8975 -3255 9095 -3135
rect 9140 -3255 9260 -3135
rect 9315 -3255 9435 -3135
rect 9480 -3255 9600 -3135
rect 9645 -3255 9765 -3135
rect 9810 -3255 9930 -3135
rect 9985 -3255 10105 -3135
rect 10150 -3255 10270 -3135
rect 10315 -3255 10435 -3135
rect 10480 -3255 10600 -3135
rect 10655 -3255 10775 -3135
rect 10820 -3255 10940 -3135
rect 10985 -3255 11105 -3135
rect 11150 -3255 11270 -3135
rect 11325 -3255 11445 -3135
rect 11490 -3255 11610 -3135
rect 11655 -3255 11775 -3135
rect 11820 -3255 11940 -3135
rect 11995 -3255 12115 -3135
rect 12160 -3255 12280 -3135
rect 12325 -3255 12445 -3135
rect 12490 -3255 12610 -3135
rect 7130 -3430 7250 -3310
rect 7305 -3430 7425 -3310
rect 7470 -3430 7590 -3310
rect 7635 -3430 7755 -3310
rect 7800 -3430 7920 -3310
rect 7975 -3430 8095 -3310
rect 8140 -3430 8260 -3310
rect 8305 -3430 8425 -3310
rect 8470 -3430 8590 -3310
rect 8645 -3430 8765 -3310
rect 8810 -3430 8930 -3310
rect 8975 -3430 9095 -3310
rect 9140 -3430 9260 -3310
rect 9315 -3430 9435 -3310
rect 9480 -3430 9600 -3310
rect 9645 -3430 9765 -3310
rect 9810 -3430 9930 -3310
rect 9985 -3430 10105 -3310
rect 10150 -3430 10270 -3310
rect 10315 -3430 10435 -3310
rect 10480 -3430 10600 -3310
rect 10655 -3430 10775 -3310
rect 10820 -3430 10940 -3310
rect 10985 -3430 11105 -3310
rect 11150 -3430 11270 -3310
rect 11325 -3430 11445 -3310
rect 11490 -3430 11610 -3310
rect 11655 -3430 11775 -3310
rect 11820 -3430 11940 -3310
rect 11995 -3430 12115 -3310
rect 12160 -3430 12280 -3310
rect 12325 -3430 12445 -3310
rect 12490 -3430 12610 -3310
rect 7130 -3595 7250 -3475
rect 7305 -3595 7425 -3475
rect 7470 -3595 7590 -3475
rect 7635 -3595 7755 -3475
rect 7800 -3595 7920 -3475
rect 7975 -3595 8095 -3475
rect 8140 -3595 8260 -3475
rect 8305 -3595 8425 -3475
rect 8470 -3595 8590 -3475
rect 8645 -3595 8765 -3475
rect 8810 -3595 8930 -3475
rect 8975 -3595 9095 -3475
rect 9140 -3595 9260 -3475
rect 9315 -3595 9435 -3475
rect 9480 -3595 9600 -3475
rect 9645 -3595 9765 -3475
rect 9810 -3595 9930 -3475
rect 9985 -3595 10105 -3475
rect 10150 -3595 10270 -3475
rect 10315 -3595 10435 -3475
rect 10480 -3595 10600 -3475
rect 10655 -3595 10775 -3475
rect 10820 -3595 10940 -3475
rect 10985 -3595 11105 -3475
rect 11150 -3595 11270 -3475
rect 11325 -3595 11445 -3475
rect 11490 -3595 11610 -3475
rect 11655 -3595 11775 -3475
rect 11820 -3595 11940 -3475
rect 11995 -3595 12115 -3475
rect 12160 -3595 12280 -3475
rect 12325 -3595 12445 -3475
rect 12490 -3595 12610 -3475
rect 7130 -3760 7250 -3640
rect 7305 -3760 7425 -3640
rect 7470 -3760 7590 -3640
rect 7635 -3760 7755 -3640
rect 7800 -3760 7920 -3640
rect 7975 -3760 8095 -3640
rect 8140 -3760 8260 -3640
rect 8305 -3760 8425 -3640
rect 8470 -3760 8590 -3640
rect 8645 -3760 8765 -3640
rect 8810 -3760 8930 -3640
rect 8975 -3760 9095 -3640
rect 9140 -3760 9260 -3640
rect 9315 -3760 9435 -3640
rect 9480 -3760 9600 -3640
rect 9645 -3760 9765 -3640
rect 9810 -3760 9930 -3640
rect 9985 -3760 10105 -3640
rect 10150 -3760 10270 -3640
rect 10315 -3760 10435 -3640
rect 10480 -3760 10600 -3640
rect 10655 -3760 10775 -3640
rect 10820 -3760 10940 -3640
rect 10985 -3760 11105 -3640
rect 11150 -3760 11270 -3640
rect 11325 -3760 11445 -3640
rect 11490 -3760 11610 -3640
rect 11655 -3760 11775 -3640
rect 11820 -3760 11940 -3640
rect 11995 -3760 12115 -3640
rect 12160 -3760 12280 -3640
rect 12325 -3760 12445 -3640
rect 12490 -3760 12610 -3640
rect 7130 -3925 7250 -3805
rect 7305 -3925 7425 -3805
rect 7470 -3925 7590 -3805
rect 7635 -3925 7755 -3805
rect 7800 -3925 7920 -3805
rect 7975 -3925 8095 -3805
rect 8140 -3925 8260 -3805
rect 8305 -3925 8425 -3805
rect 8470 -3925 8590 -3805
rect 8645 -3925 8765 -3805
rect 8810 -3925 8930 -3805
rect 8975 -3925 9095 -3805
rect 9140 -3925 9260 -3805
rect 9315 -3925 9435 -3805
rect 9480 -3925 9600 -3805
rect 9645 -3925 9765 -3805
rect 9810 -3925 9930 -3805
rect 9985 -3925 10105 -3805
rect 10150 -3925 10270 -3805
rect 10315 -3925 10435 -3805
rect 10480 -3925 10600 -3805
rect 10655 -3925 10775 -3805
rect 10820 -3925 10940 -3805
rect 10985 -3925 11105 -3805
rect 11150 -3925 11270 -3805
rect 11325 -3925 11445 -3805
rect 11490 -3925 11610 -3805
rect 11655 -3925 11775 -3805
rect 11820 -3925 11940 -3805
rect 11995 -3925 12115 -3805
rect 12160 -3925 12280 -3805
rect 12325 -3925 12445 -3805
rect 12490 -3925 12610 -3805
rect 7130 -4100 7250 -3980
rect 7305 -4100 7425 -3980
rect 7470 -4100 7590 -3980
rect 7635 -4100 7755 -3980
rect 7800 -4100 7920 -3980
rect 7975 -4100 8095 -3980
rect 8140 -4100 8260 -3980
rect 8305 -4100 8425 -3980
rect 8470 -4100 8590 -3980
rect 8645 -4100 8765 -3980
rect 8810 -4100 8930 -3980
rect 8975 -4100 9095 -3980
rect 9140 -4100 9260 -3980
rect 9315 -4100 9435 -3980
rect 9480 -4100 9600 -3980
rect 9645 -4100 9765 -3980
rect 9810 -4100 9930 -3980
rect 9985 -4100 10105 -3980
rect 10150 -4100 10270 -3980
rect 10315 -4100 10435 -3980
rect 10480 -4100 10600 -3980
rect 10655 -4100 10775 -3980
rect 10820 -4100 10940 -3980
rect 10985 -4100 11105 -3980
rect 11150 -4100 11270 -3980
rect 11325 -4100 11445 -3980
rect 11490 -4100 11610 -3980
rect 11655 -4100 11775 -3980
rect 11820 -4100 11940 -3980
rect 11995 -4100 12115 -3980
rect 12160 -4100 12280 -3980
rect 12325 -4100 12445 -3980
rect 12490 -4100 12610 -3980
rect 12820 1260 12940 1380
rect 12995 1260 13115 1380
rect 13160 1260 13280 1380
rect 13325 1260 13445 1380
rect 13490 1260 13610 1380
rect 13665 1260 13785 1380
rect 13830 1260 13950 1380
rect 13995 1260 14115 1380
rect 14160 1260 14280 1380
rect 14335 1260 14455 1380
rect 14500 1260 14620 1380
rect 14665 1260 14785 1380
rect 14830 1260 14950 1380
rect 15005 1260 15125 1380
rect 15170 1260 15290 1380
rect 15335 1260 15455 1380
rect 15500 1260 15620 1380
rect 15675 1260 15795 1380
rect 15840 1260 15960 1380
rect 16005 1260 16125 1380
rect 16170 1260 16290 1380
rect 16345 1260 16465 1380
rect 16510 1260 16630 1380
rect 16675 1260 16795 1380
rect 16840 1260 16960 1380
rect 17015 1260 17135 1380
rect 17180 1260 17300 1380
rect 17345 1260 17465 1380
rect 17510 1260 17630 1380
rect 17685 1260 17805 1380
rect 17850 1260 17970 1380
rect 18015 1260 18135 1380
rect 18180 1260 18300 1380
rect 12820 1095 12940 1215
rect 12995 1095 13115 1215
rect 13160 1095 13280 1215
rect 13325 1095 13445 1215
rect 13490 1095 13610 1215
rect 13665 1095 13785 1215
rect 13830 1095 13950 1215
rect 13995 1095 14115 1215
rect 14160 1095 14280 1215
rect 14335 1095 14455 1215
rect 14500 1095 14620 1215
rect 14665 1095 14785 1215
rect 14830 1095 14950 1215
rect 15005 1095 15125 1215
rect 15170 1095 15290 1215
rect 15335 1095 15455 1215
rect 15500 1095 15620 1215
rect 15675 1095 15795 1215
rect 15840 1095 15960 1215
rect 16005 1095 16125 1215
rect 16170 1095 16290 1215
rect 16345 1095 16465 1215
rect 16510 1095 16630 1215
rect 16675 1095 16795 1215
rect 16840 1095 16960 1215
rect 17015 1095 17135 1215
rect 17180 1095 17300 1215
rect 17345 1095 17465 1215
rect 17510 1095 17630 1215
rect 17685 1095 17805 1215
rect 17850 1095 17970 1215
rect 18015 1095 18135 1215
rect 18180 1095 18300 1215
rect 12820 930 12940 1050
rect 12995 930 13115 1050
rect 13160 930 13280 1050
rect 13325 930 13445 1050
rect 13490 930 13610 1050
rect 13665 930 13785 1050
rect 13830 930 13950 1050
rect 13995 930 14115 1050
rect 14160 930 14280 1050
rect 14335 930 14455 1050
rect 14500 930 14620 1050
rect 14665 930 14785 1050
rect 14830 930 14950 1050
rect 15005 930 15125 1050
rect 15170 930 15290 1050
rect 15335 930 15455 1050
rect 15500 930 15620 1050
rect 15675 930 15795 1050
rect 15840 930 15960 1050
rect 16005 930 16125 1050
rect 16170 930 16290 1050
rect 16345 930 16465 1050
rect 16510 930 16630 1050
rect 16675 930 16795 1050
rect 16840 930 16960 1050
rect 17015 930 17135 1050
rect 17180 930 17300 1050
rect 17345 930 17465 1050
rect 17510 930 17630 1050
rect 17685 930 17805 1050
rect 17850 930 17970 1050
rect 18015 930 18135 1050
rect 18180 930 18300 1050
rect 12820 765 12940 885
rect 12995 765 13115 885
rect 13160 765 13280 885
rect 13325 765 13445 885
rect 13490 765 13610 885
rect 13665 765 13785 885
rect 13830 765 13950 885
rect 13995 765 14115 885
rect 14160 765 14280 885
rect 14335 765 14455 885
rect 14500 765 14620 885
rect 14665 765 14785 885
rect 14830 765 14950 885
rect 15005 765 15125 885
rect 15170 765 15290 885
rect 15335 765 15455 885
rect 15500 765 15620 885
rect 15675 765 15795 885
rect 15840 765 15960 885
rect 16005 765 16125 885
rect 16170 765 16290 885
rect 16345 765 16465 885
rect 16510 765 16630 885
rect 16675 765 16795 885
rect 16840 765 16960 885
rect 17015 765 17135 885
rect 17180 765 17300 885
rect 17345 765 17465 885
rect 17510 765 17630 885
rect 17685 765 17805 885
rect 17850 765 17970 885
rect 18015 765 18135 885
rect 18180 765 18300 885
rect 12820 590 12940 710
rect 12995 590 13115 710
rect 13160 590 13280 710
rect 13325 590 13445 710
rect 13490 590 13610 710
rect 13665 590 13785 710
rect 13830 590 13950 710
rect 13995 590 14115 710
rect 14160 590 14280 710
rect 14335 590 14455 710
rect 14500 590 14620 710
rect 14665 590 14785 710
rect 14830 590 14950 710
rect 15005 590 15125 710
rect 15170 590 15290 710
rect 15335 590 15455 710
rect 15500 590 15620 710
rect 15675 590 15795 710
rect 15840 590 15960 710
rect 16005 590 16125 710
rect 16170 590 16290 710
rect 16345 590 16465 710
rect 16510 590 16630 710
rect 16675 590 16795 710
rect 16840 590 16960 710
rect 17015 590 17135 710
rect 17180 590 17300 710
rect 17345 590 17465 710
rect 17510 590 17630 710
rect 17685 590 17805 710
rect 17850 590 17970 710
rect 18015 590 18135 710
rect 18180 590 18300 710
rect 12820 425 12940 545
rect 12995 425 13115 545
rect 13160 425 13280 545
rect 13325 425 13445 545
rect 13490 425 13610 545
rect 13665 425 13785 545
rect 13830 425 13950 545
rect 13995 425 14115 545
rect 14160 425 14280 545
rect 14335 425 14455 545
rect 14500 425 14620 545
rect 14665 425 14785 545
rect 14830 425 14950 545
rect 15005 425 15125 545
rect 15170 425 15290 545
rect 15335 425 15455 545
rect 15500 425 15620 545
rect 15675 425 15795 545
rect 15840 425 15960 545
rect 16005 425 16125 545
rect 16170 425 16290 545
rect 16345 425 16465 545
rect 16510 425 16630 545
rect 16675 425 16795 545
rect 16840 425 16960 545
rect 17015 425 17135 545
rect 17180 425 17300 545
rect 17345 425 17465 545
rect 17510 425 17630 545
rect 17685 425 17805 545
rect 17850 425 17970 545
rect 18015 425 18135 545
rect 18180 425 18300 545
rect 12820 260 12940 380
rect 12995 260 13115 380
rect 13160 260 13280 380
rect 13325 260 13445 380
rect 13490 260 13610 380
rect 13665 260 13785 380
rect 13830 260 13950 380
rect 13995 260 14115 380
rect 14160 260 14280 380
rect 14335 260 14455 380
rect 14500 260 14620 380
rect 14665 260 14785 380
rect 14830 260 14950 380
rect 15005 260 15125 380
rect 15170 260 15290 380
rect 15335 260 15455 380
rect 15500 260 15620 380
rect 15675 260 15795 380
rect 15840 260 15960 380
rect 16005 260 16125 380
rect 16170 260 16290 380
rect 16345 260 16465 380
rect 16510 260 16630 380
rect 16675 260 16795 380
rect 16840 260 16960 380
rect 17015 260 17135 380
rect 17180 260 17300 380
rect 17345 260 17465 380
rect 17510 260 17630 380
rect 17685 260 17805 380
rect 17850 260 17970 380
rect 18015 260 18135 380
rect 18180 260 18300 380
rect 12820 95 12940 215
rect 12995 95 13115 215
rect 13160 95 13280 215
rect 13325 95 13445 215
rect 13490 95 13610 215
rect 13665 95 13785 215
rect 13830 95 13950 215
rect 13995 95 14115 215
rect 14160 95 14280 215
rect 14335 95 14455 215
rect 14500 95 14620 215
rect 14665 95 14785 215
rect 14830 95 14950 215
rect 15005 95 15125 215
rect 15170 95 15290 215
rect 15335 95 15455 215
rect 15500 95 15620 215
rect 15675 95 15795 215
rect 15840 95 15960 215
rect 16005 95 16125 215
rect 16170 95 16290 215
rect 16345 95 16465 215
rect 16510 95 16630 215
rect 16675 95 16795 215
rect 16840 95 16960 215
rect 17015 95 17135 215
rect 17180 95 17300 215
rect 17345 95 17465 215
rect 17510 95 17630 215
rect 17685 95 17805 215
rect 17850 95 17970 215
rect 18015 95 18135 215
rect 18180 95 18300 215
rect 12820 -80 12940 40
rect 12995 -80 13115 40
rect 13160 -80 13280 40
rect 13325 -80 13445 40
rect 13490 -80 13610 40
rect 13665 -80 13785 40
rect 13830 -80 13950 40
rect 13995 -80 14115 40
rect 14160 -80 14280 40
rect 14335 -80 14455 40
rect 14500 -80 14620 40
rect 14665 -80 14785 40
rect 14830 -80 14950 40
rect 15005 -80 15125 40
rect 15170 -80 15290 40
rect 15335 -80 15455 40
rect 15500 -80 15620 40
rect 15675 -80 15795 40
rect 15840 -80 15960 40
rect 16005 -80 16125 40
rect 16170 -80 16290 40
rect 16345 -80 16465 40
rect 16510 -80 16630 40
rect 16675 -80 16795 40
rect 16840 -80 16960 40
rect 17015 -80 17135 40
rect 17180 -80 17300 40
rect 17345 -80 17465 40
rect 17510 -80 17630 40
rect 17685 -80 17805 40
rect 17850 -80 17970 40
rect 18015 -80 18135 40
rect 18180 -80 18300 40
rect 12820 -245 12940 -125
rect 12995 -245 13115 -125
rect 13160 -245 13280 -125
rect 13325 -245 13445 -125
rect 13490 -245 13610 -125
rect 13665 -245 13785 -125
rect 13830 -245 13950 -125
rect 13995 -245 14115 -125
rect 14160 -245 14280 -125
rect 14335 -245 14455 -125
rect 14500 -245 14620 -125
rect 14665 -245 14785 -125
rect 14830 -245 14950 -125
rect 15005 -245 15125 -125
rect 15170 -245 15290 -125
rect 15335 -245 15455 -125
rect 15500 -245 15620 -125
rect 15675 -245 15795 -125
rect 15840 -245 15960 -125
rect 16005 -245 16125 -125
rect 16170 -245 16290 -125
rect 16345 -245 16465 -125
rect 16510 -245 16630 -125
rect 16675 -245 16795 -125
rect 16840 -245 16960 -125
rect 17015 -245 17135 -125
rect 17180 -245 17300 -125
rect 17345 -245 17465 -125
rect 17510 -245 17630 -125
rect 17685 -245 17805 -125
rect 17850 -245 17970 -125
rect 18015 -245 18135 -125
rect 18180 -245 18300 -125
rect 12820 -410 12940 -290
rect 12995 -410 13115 -290
rect 13160 -410 13280 -290
rect 13325 -410 13445 -290
rect 13490 -410 13610 -290
rect 13665 -410 13785 -290
rect 13830 -410 13950 -290
rect 13995 -410 14115 -290
rect 14160 -410 14280 -290
rect 14335 -410 14455 -290
rect 14500 -410 14620 -290
rect 14665 -410 14785 -290
rect 14830 -410 14950 -290
rect 15005 -410 15125 -290
rect 15170 -410 15290 -290
rect 15335 -410 15455 -290
rect 15500 -410 15620 -290
rect 15675 -410 15795 -290
rect 15840 -410 15960 -290
rect 16005 -410 16125 -290
rect 16170 -410 16290 -290
rect 16345 -410 16465 -290
rect 16510 -410 16630 -290
rect 16675 -410 16795 -290
rect 16840 -410 16960 -290
rect 17015 -410 17135 -290
rect 17180 -410 17300 -290
rect 17345 -410 17465 -290
rect 17510 -410 17630 -290
rect 17685 -410 17805 -290
rect 17850 -410 17970 -290
rect 18015 -410 18135 -290
rect 18180 -410 18300 -290
rect 12820 -575 12940 -455
rect 12995 -575 13115 -455
rect 13160 -575 13280 -455
rect 13325 -575 13445 -455
rect 13490 -575 13610 -455
rect 13665 -575 13785 -455
rect 13830 -575 13950 -455
rect 13995 -575 14115 -455
rect 14160 -575 14280 -455
rect 14335 -575 14455 -455
rect 14500 -575 14620 -455
rect 14665 -575 14785 -455
rect 14830 -575 14950 -455
rect 15005 -575 15125 -455
rect 15170 -575 15290 -455
rect 15335 -575 15455 -455
rect 15500 -575 15620 -455
rect 15675 -575 15795 -455
rect 15840 -575 15960 -455
rect 16005 -575 16125 -455
rect 16170 -575 16290 -455
rect 16345 -575 16465 -455
rect 16510 -575 16630 -455
rect 16675 -575 16795 -455
rect 16840 -575 16960 -455
rect 17015 -575 17135 -455
rect 17180 -575 17300 -455
rect 17345 -575 17465 -455
rect 17510 -575 17630 -455
rect 17685 -575 17805 -455
rect 17850 -575 17970 -455
rect 18015 -575 18135 -455
rect 18180 -575 18300 -455
rect 12820 -750 12940 -630
rect 12995 -750 13115 -630
rect 13160 -750 13280 -630
rect 13325 -750 13445 -630
rect 13490 -750 13610 -630
rect 13665 -750 13785 -630
rect 13830 -750 13950 -630
rect 13995 -750 14115 -630
rect 14160 -750 14280 -630
rect 14335 -750 14455 -630
rect 14500 -750 14620 -630
rect 14665 -750 14785 -630
rect 14830 -750 14950 -630
rect 15005 -750 15125 -630
rect 15170 -750 15290 -630
rect 15335 -750 15455 -630
rect 15500 -750 15620 -630
rect 15675 -750 15795 -630
rect 15840 -750 15960 -630
rect 16005 -750 16125 -630
rect 16170 -750 16290 -630
rect 16345 -750 16465 -630
rect 16510 -750 16630 -630
rect 16675 -750 16795 -630
rect 16840 -750 16960 -630
rect 17015 -750 17135 -630
rect 17180 -750 17300 -630
rect 17345 -750 17465 -630
rect 17510 -750 17630 -630
rect 17685 -750 17805 -630
rect 17850 -750 17970 -630
rect 18015 -750 18135 -630
rect 18180 -750 18300 -630
rect 12820 -915 12940 -795
rect 12995 -915 13115 -795
rect 13160 -915 13280 -795
rect 13325 -915 13445 -795
rect 13490 -915 13610 -795
rect 13665 -915 13785 -795
rect 13830 -915 13950 -795
rect 13995 -915 14115 -795
rect 14160 -915 14280 -795
rect 14335 -915 14455 -795
rect 14500 -915 14620 -795
rect 14665 -915 14785 -795
rect 14830 -915 14950 -795
rect 15005 -915 15125 -795
rect 15170 -915 15290 -795
rect 15335 -915 15455 -795
rect 15500 -915 15620 -795
rect 15675 -915 15795 -795
rect 15840 -915 15960 -795
rect 16005 -915 16125 -795
rect 16170 -915 16290 -795
rect 16345 -915 16465 -795
rect 16510 -915 16630 -795
rect 16675 -915 16795 -795
rect 16840 -915 16960 -795
rect 17015 -915 17135 -795
rect 17180 -915 17300 -795
rect 17345 -915 17465 -795
rect 17510 -915 17630 -795
rect 17685 -915 17805 -795
rect 17850 -915 17970 -795
rect 18015 -915 18135 -795
rect 18180 -915 18300 -795
rect 12820 -1080 12940 -960
rect 12995 -1080 13115 -960
rect 13160 -1080 13280 -960
rect 13325 -1080 13445 -960
rect 13490 -1080 13610 -960
rect 13665 -1080 13785 -960
rect 13830 -1080 13950 -960
rect 13995 -1080 14115 -960
rect 14160 -1080 14280 -960
rect 14335 -1080 14455 -960
rect 14500 -1080 14620 -960
rect 14665 -1080 14785 -960
rect 14830 -1080 14950 -960
rect 15005 -1080 15125 -960
rect 15170 -1080 15290 -960
rect 15335 -1080 15455 -960
rect 15500 -1080 15620 -960
rect 15675 -1080 15795 -960
rect 15840 -1080 15960 -960
rect 16005 -1080 16125 -960
rect 16170 -1080 16290 -960
rect 16345 -1080 16465 -960
rect 16510 -1080 16630 -960
rect 16675 -1080 16795 -960
rect 16840 -1080 16960 -960
rect 17015 -1080 17135 -960
rect 17180 -1080 17300 -960
rect 17345 -1080 17465 -960
rect 17510 -1080 17630 -960
rect 17685 -1080 17805 -960
rect 17850 -1080 17970 -960
rect 18015 -1080 18135 -960
rect 18180 -1080 18300 -960
rect 12820 -1245 12940 -1125
rect 12995 -1245 13115 -1125
rect 13160 -1245 13280 -1125
rect 13325 -1245 13445 -1125
rect 13490 -1245 13610 -1125
rect 13665 -1245 13785 -1125
rect 13830 -1245 13950 -1125
rect 13995 -1245 14115 -1125
rect 14160 -1245 14280 -1125
rect 14335 -1245 14455 -1125
rect 14500 -1245 14620 -1125
rect 14665 -1245 14785 -1125
rect 14830 -1245 14950 -1125
rect 15005 -1245 15125 -1125
rect 15170 -1245 15290 -1125
rect 15335 -1245 15455 -1125
rect 15500 -1245 15620 -1125
rect 15675 -1245 15795 -1125
rect 15840 -1245 15960 -1125
rect 16005 -1245 16125 -1125
rect 16170 -1245 16290 -1125
rect 16345 -1245 16465 -1125
rect 16510 -1245 16630 -1125
rect 16675 -1245 16795 -1125
rect 16840 -1245 16960 -1125
rect 17015 -1245 17135 -1125
rect 17180 -1245 17300 -1125
rect 17345 -1245 17465 -1125
rect 17510 -1245 17630 -1125
rect 17685 -1245 17805 -1125
rect 17850 -1245 17970 -1125
rect 18015 -1245 18135 -1125
rect 18180 -1245 18300 -1125
rect 12820 -1420 12940 -1300
rect 12995 -1420 13115 -1300
rect 13160 -1420 13280 -1300
rect 13325 -1420 13445 -1300
rect 13490 -1420 13610 -1300
rect 13665 -1420 13785 -1300
rect 13830 -1420 13950 -1300
rect 13995 -1420 14115 -1300
rect 14160 -1420 14280 -1300
rect 14335 -1420 14455 -1300
rect 14500 -1420 14620 -1300
rect 14665 -1420 14785 -1300
rect 14830 -1420 14950 -1300
rect 15005 -1420 15125 -1300
rect 15170 -1420 15290 -1300
rect 15335 -1420 15455 -1300
rect 15500 -1420 15620 -1300
rect 15675 -1420 15795 -1300
rect 15840 -1420 15960 -1300
rect 16005 -1420 16125 -1300
rect 16170 -1420 16290 -1300
rect 16345 -1420 16465 -1300
rect 16510 -1420 16630 -1300
rect 16675 -1420 16795 -1300
rect 16840 -1420 16960 -1300
rect 17015 -1420 17135 -1300
rect 17180 -1420 17300 -1300
rect 17345 -1420 17465 -1300
rect 17510 -1420 17630 -1300
rect 17685 -1420 17805 -1300
rect 17850 -1420 17970 -1300
rect 18015 -1420 18135 -1300
rect 18180 -1420 18300 -1300
rect 12820 -1585 12940 -1465
rect 12995 -1585 13115 -1465
rect 13160 -1585 13280 -1465
rect 13325 -1585 13445 -1465
rect 13490 -1585 13610 -1465
rect 13665 -1585 13785 -1465
rect 13830 -1585 13950 -1465
rect 13995 -1585 14115 -1465
rect 14160 -1585 14280 -1465
rect 14335 -1585 14455 -1465
rect 14500 -1585 14620 -1465
rect 14665 -1585 14785 -1465
rect 14830 -1585 14950 -1465
rect 15005 -1585 15125 -1465
rect 15170 -1585 15290 -1465
rect 15335 -1585 15455 -1465
rect 15500 -1585 15620 -1465
rect 15675 -1585 15795 -1465
rect 15840 -1585 15960 -1465
rect 16005 -1585 16125 -1465
rect 16170 -1585 16290 -1465
rect 16345 -1585 16465 -1465
rect 16510 -1585 16630 -1465
rect 16675 -1585 16795 -1465
rect 16840 -1585 16960 -1465
rect 17015 -1585 17135 -1465
rect 17180 -1585 17300 -1465
rect 17345 -1585 17465 -1465
rect 17510 -1585 17630 -1465
rect 17685 -1585 17805 -1465
rect 17850 -1585 17970 -1465
rect 18015 -1585 18135 -1465
rect 18180 -1585 18300 -1465
rect 12820 -1750 12940 -1630
rect 12995 -1750 13115 -1630
rect 13160 -1750 13280 -1630
rect 13325 -1750 13445 -1630
rect 13490 -1750 13610 -1630
rect 13665 -1750 13785 -1630
rect 13830 -1750 13950 -1630
rect 13995 -1750 14115 -1630
rect 14160 -1750 14280 -1630
rect 14335 -1750 14455 -1630
rect 14500 -1750 14620 -1630
rect 14665 -1750 14785 -1630
rect 14830 -1750 14950 -1630
rect 15005 -1750 15125 -1630
rect 15170 -1750 15290 -1630
rect 15335 -1750 15455 -1630
rect 15500 -1750 15620 -1630
rect 15675 -1750 15795 -1630
rect 15840 -1750 15960 -1630
rect 16005 -1750 16125 -1630
rect 16170 -1750 16290 -1630
rect 16345 -1750 16465 -1630
rect 16510 -1750 16630 -1630
rect 16675 -1750 16795 -1630
rect 16840 -1750 16960 -1630
rect 17015 -1750 17135 -1630
rect 17180 -1750 17300 -1630
rect 17345 -1750 17465 -1630
rect 17510 -1750 17630 -1630
rect 17685 -1750 17805 -1630
rect 17850 -1750 17970 -1630
rect 18015 -1750 18135 -1630
rect 18180 -1750 18300 -1630
rect 12820 -1915 12940 -1795
rect 12995 -1915 13115 -1795
rect 13160 -1915 13280 -1795
rect 13325 -1915 13445 -1795
rect 13490 -1915 13610 -1795
rect 13665 -1915 13785 -1795
rect 13830 -1915 13950 -1795
rect 13995 -1915 14115 -1795
rect 14160 -1915 14280 -1795
rect 14335 -1915 14455 -1795
rect 14500 -1915 14620 -1795
rect 14665 -1915 14785 -1795
rect 14830 -1915 14950 -1795
rect 15005 -1915 15125 -1795
rect 15170 -1915 15290 -1795
rect 15335 -1915 15455 -1795
rect 15500 -1915 15620 -1795
rect 15675 -1915 15795 -1795
rect 15840 -1915 15960 -1795
rect 16005 -1915 16125 -1795
rect 16170 -1915 16290 -1795
rect 16345 -1915 16465 -1795
rect 16510 -1915 16630 -1795
rect 16675 -1915 16795 -1795
rect 16840 -1915 16960 -1795
rect 17015 -1915 17135 -1795
rect 17180 -1915 17300 -1795
rect 17345 -1915 17465 -1795
rect 17510 -1915 17630 -1795
rect 17685 -1915 17805 -1795
rect 17850 -1915 17970 -1795
rect 18015 -1915 18135 -1795
rect 18180 -1915 18300 -1795
rect 12820 -2090 12940 -1970
rect 12995 -2090 13115 -1970
rect 13160 -2090 13280 -1970
rect 13325 -2090 13445 -1970
rect 13490 -2090 13610 -1970
rect 13665 -2090 13785 -1970
rect 13830 -2090 13950 -1970
rect 13995 -2090 14115 -1970
rect 14160 -2090 14280 -1970
rect 14335 -2090 14455 -1970
rect 14500 -2090 14620 -1970
rect 14665 -2090 14785 -1970
rect 14830 -2090 14950 -1970
rect 15005 -2090 15125 -1970
rect 15170 -2090 15290 -1970
rect 15335 -2090 15455 -1970
rect 15500 -2090 15620 -1970
rect 15675 -2090 15795 -1970
rect 15840 -2090 15960 -1970
rect 16005 -2090 16125 -1970
rect 16170 -2090 16290 -1970
rect 16345 -2090 16465 -1970
rect 16510 -2090 16630 -1970
rect 16675 -2090 16795 -1970
rect 16840 -2090 16960 -1970
rect 17015 -2090 17135 -1970
rect 17180 -2090 17300 -1970
rect 17345 -2090 17465 -1970
rect 17510 -2090 17630 -1970
rect 17685 -2090 17805 -1970
rect 17850 -2090 17970 -1970
rect 18015 -2090 18135 -1970
rect 18180 -2090 18300 -1970
rect 12820 -2255 12940 -2135
rect 12995 -2255 13115 -2135
rect 13160 -2255 13280 -2135
rect 13325 -2255 13445 -2135
rect 13490 -2255 13610 -2135
rect 13665 -2255 13785 -2135
rect 13830 -2255 13950 -2135
rect 13995 -2255 14115 -2135
rect 14160 -2255 14280 -2135
rect 14335 -2255 14455 -2135
rect 14500 -2255 14620 -2135
rect 14665 -2255 14785 -2135
rect 14830 -2255 14950 -2135
rect 15005 -2255 15125 -2135
rect 15170 -2255 15290 -2135
rect 15335 -2255 15455 -2135
rect 15500 -2255 15620 -2135
rect 15675 -2255 15795 -2135
rect 15840 -2255 15960 -2135
rect 16005 -2255 16125 -2135
rect 16170 -2255 16290 -2135
rect 16345 -2255 16465 -2135
rect 16510 -2255 16630 -2135
rect 16675 -2255 16795 -2135
rect 16840 -2255 16960 -2135
rect 17015 -2255 17135 -2135
rect 17180 -2255 17300 -2135
rect 17345 -2255 17465 -2135
rect 17510 -2255 17630 -2135
rect 17685 -2255 17805 -2135
rect 17850 -2255 17970 -2135
rect 18015 -2255 18135 -2135
rect 18180 -2255 18300 -2135
rect 12820 -2420 12940 -2300
rect 12995 -2420 13115 -2300
rect 13160 -2420 13280 -2300
rect 13325 -2420 13445 -2300
rect 13490 -2420 13610 -2300
rect 13665 -2420 13785 -2300
rect 13830 -2420 13950 -2300
rect 13995 -2420 14115 -2300
rect 14160 -2420 14280 -2300
rect 14335 -2420 14455 -2300
rect 14500 -2420 14620 -2300
rect 14665 -2420 14785 -2300
rect 14830 -2420 14950 -2300
rect 15005 -2420 15125 -2300
rect 15170 -2420 15290 -2300
rect 15335 -2420 15455 -2300
rect 15500 -2420 15620 -2300
rect 15675 -2420 15795 -2300
rect 15840 -2420 15960 -2300
rect 16005 -2420 16125 -2300
rect 16170 -2420 16290 -2300
rect 16345 -2420 16465 -2300
rect 16510 -2420 16630 -2300
rect 16675 -2420 16795 -2300
rect 16840 -2420 16960 -2300
rect 17015 -2420 17135 -2300
rect 17180 -2420 17300 -2300
rect 17345 -2420 17465 -2300
rect 17510 -2420 17630 -2300
rect 17685 -2420 17805 -2300
rect 17850 -2420 17970 -2300
rect 18015 -2420 18135 -2300
rect 18180 -2420 18300 -2300
rect 12820 -2585 12940 -2465
rect 12995 -2585 13115 -2465
rect 13160 -2585 13280 -2465
rect 13325 -2585 13445 -2465
rect 13490 -2585 13610 -2465
rect 13665 -2585 13785 -2465
rect 13830 -2585 13950 -2465
rect 13995 -2585 14115 -2465
rect 14160 -2585 14280 -2465
rect 14335 -2585 14455 -2465
rect 14500 -2585 14620 -2465
rect 14665 -2585 14785 -2465
rect 14830 -2585 14950 -2465
rect 15005 -2585 15125 -2465
rect 15170 -2585 15290 -2465
rect 15335 -2585 15455 -2465
rect 15500 -2585 15620 -2465
rect 15675 -2585 15795 -2465
rect 15840 -2585 15960 -2465
rect 16005 -2585 16125 -2465
rect 16170 -2585 16290 -2465
rect 16345 -2585 16465 -2465
rect 16510 -2585 16630 -2465
rect 16675 -2585 16795 -2465
rect 16840 -2585 16960 -2465
rect 17015 -2585 17135 -2465
rect 17180 -2585 17300 -2465
rect 17345 -2585 17465 -2465
rect 17510 -2585 17630 -2465
rect 17685 -2585 17805 -2465
rect 17850 -2585 17970 -2465
rect 18015 -2585 18135 -2465
rect 18180 -2585 18300 -2465
rect 12820 -2760 12940 -2640
rect 12995 -2760 13115 -2640
rect 13160 -2760 13280 -2640
rect 13325 -2760 13445 -2640
rect 13490 -2760 13610 -2640
rect 13665 -2760 13785 -2640
rect 13830 -2760 13950 -2640
rect 13995 -2760 14115 -2640
rect 14160 -2760 14280 -2640
rect 14335 -2760 14455 -2640
rect 14500 -2760 14620 -2640
rect 14665 -2760 14785 -2640
rect 14830 -2760 14950 -2640
rect 15005 -2760 15125 -2640
rect 15170 -2760 15290 -2640
rect 15335 -2760 15455 -2640
rect 15500 -2760 15620 -2640
rect 15675 -2760 15795 -2640
rect 15840 -2760 15960 -2640
rect 16005 -2760 16125 -2640
rect 16170 -2760 16290 -2640
rect 16345 -2760 16465 -2640
rect 16510 -2760 16630 -2640
rect 16675 -2760 16795 -2640
rect 16840 -2760 16960 -2640
rect 17015 -2760 17135 -2640
rect 17180 -2760 17300 -2640
rect 17345 -2760 17465 -2640
rect 17510 -2760 17630 -2640
rect 17685 -2760 17805 -2640
rect 17850 -2760 17970 -2640
rect 18015 -2760 18135 -2640
rect 18180 -2760 18300 -2640
rect 12820 -2925 12940 -2805
rect 12995 -2925 13115 -2805
rect 13160 -2925 13280 -2805
rect 13325 -2925 13445 -2805
rect 13490 -2925 13610 -2805
rect 13665 -2925 13785 -2805
rect 13830 -2925 13950 -2805
rect 13995 -2925 14115 -2805
rect 14160 -2925 14280 -2805
rect 14335 -2925 14455 -2805
rect 14500 -2925 14620 -2805
rect 14665 -2925 14785 -2805
rect 14830 -2925 14950 -2805
rect 15005 -2925 15125 -2805
rect 15170 -2925 15290 -2805
rect 15335 -2925 15455 -2805
rect 15500 -2925 15620 -2805
rect 15675 -2925 15795 -2805
rect 15840 -2925 15960 -2805
rect 16005 -2925 16125 -2805
rect 16170 -2925 16290 -2805
rect 16345 -2925 16465 -2805
rect 16510 -2925 16630 -2805
rect 16675 -2925 16795 -2805
rect 16840 -2925 16960 -2805
rect 17015 -2925 17135 -2805
rect 17180 -2925 17300 -2805
rect 17345 -2925 17465 -2805
rect 17510 -2925 17630 -2805
rect 17685 -2925 17805 -2805
rect 17850 -2925 17970 -2805
rect 18015 -2925 18135 -2805
rect 18180 -2925 18300 -2805
rect 12820 -3090 12940 -2970
rect 12995 -3090 13115 -2970
rect 13160 -3090 13280 -2970
rect 13325 -3090 13445 -2970
rect 13490 -3090 13610 -2970
rect 13665 -3090 13785 -2970
rect 13830 -3090 13950 -2970
rect 13995 -3090 14115 -2970
rect 14160 -3090 14280 -2970
rect 14335 -3090 14455 -2970
rect 14500 -3090 14620 -2970
rect 14665 -3090 14785 -2970
rect 14830 -3090 14950 -2970
rect 15005 -3090 15125 -2970
rect 15170 -3090 15290 -2970
rect 15335 -3090 15455 -2970
rect 15500 -3090 15620 -2970
rect 15675 -3090 15795 -2970
rect 15840 -3090 15960 -2970
rect 16005 -3090 16125 -2970
rect 16170 -3090 16290 -2970
rect 16345 -3090 16465 -2970
rect 16510 -3090 16630 -2970
rect 16675 -3090 16795 -2970
rect 16840 -3090 16960 -2970
rect 17015 -3090 17135 -2970
rect 17180 -3090 17300 -2970
rect 17345 -3090 17465 -2970
rect 17510 -3090 17630 -2970
rect 17685 -3090 17805 -2970
rect 17850 -3090 17970 -2970
rect 18015 -3090 18135 -2970
rect 18180 -3090 18300 -2970
rect 12820 -3255 12940 -3135
rect 12995 -3255 13115 -3135
rect 13160 -3255 13280 -3135
rect 13325 -3255 13445 -3135
rect 13490 -3255 13610 -3135
rect 13665 -3255 13785 -3135
rect 13830 -3255 13950 -3135
rect 13995 -3255 14115 -3135
rect 14160 -3255 14280 -3135
rect 14335 -3255 14455 -3135
rect 14500 -3255 14620 -3135
rect 14665 -3255 14785 -3135
rect 14830 -3255 14950 -3135
rect 15005 -3255 15125 -3135
rect 15170 -3255 15290 -3135
rect 15335 -3255 15455 -3135
rect 15500 -3255 15620 -3135
rect 15675 -3255 15795 -3135
rect 15840 -3255 15960 -3135
rect 16005 -3255 16125 -3135
rect 16170 -3255 16290 -3135
rect 16345 -3255 16465 -3135
rect 16510 -3255 16630 -3135
rect 16675 -3255 16795 -3135
rect 16840 -3255 16960 -3135
rect 17015 -3255 17135 -3135
rect 17180 -3255 17300 -3135
rect 17345 -3255 17465 -3135
rect 17510 -3255 17630 -3135
rect 17685 -3255 17805 -3135
rect 17850 -3255 17970 -3135
rect 18015 -3255 18135 -3135
rect 18180 -3255 18300 -3135
rect 12820 -3430 12940 -3310
rect 12995 -3430 13115 -3310
rect 13160 -3430 13280 -3310
rect 13325 -3430 13445 -3310
rect 13490 -3430 13610 -3310
rect 13665 -3430 13785 -3310
rect 13830 -3430 13950 -3310
rect 13995 -3430 14115 -3310
rect 14160 -3430 14280 -3310
rect 14335 -3430 14455 -3310
rect 14500 -3430 14620 -3310
rect 14665 -3430 14785 -3310
rect 14830 -3430 14950 -3310
rect 15005 -3430 15125 -3310
rect 15170 -3430 15290 -3310
rect 15335 -3430 15455 -3310
rect 15500 -3430 15620 -3310
rect 15675 -3430 15795 -3310
rect 15840 -3430 15960 -3310
rect 16005 -3430 16125 -3310
rect 16170 -3430 16290 -3310
rect 16345 -3430 16465 -3310
rect 16510 -3430 16630 -3310
rect 16675 -3430 16795 -3310
rect 16840 -3430 16960 -3310
rect 17015 -3430 17135 -3310
rect 17180 -3430 17300 -3310
rect 17345 -3430 17465 -3310
rect 17510 -3430 17630 -3310
rect 17685 -3430 17805 -3310
rect 17850 -3430 17970 -3310
rect 18015 -3430 18135 -3310
rect 18180 -3430 18300 -3310
rect 12820 -3595 12940 -3475
rect 12995 -3595 13115 -3475
rect 13160 -3595 13280 -3475
rect 13325 -3595 13445 -3475
rect 13490 -3595 13610 -3475
rect 13665 -3595 13785 -3475
rect 13830 -3595 13950 -3475
rect 13995 -3595 14115 -3475
rect 14160 -3595 14280 -3475
rect 14335 -3595 14455 -3475
rect 14500 -3595 14620 -3475
rect 14665 -3595 14785 -3475
rect 14830 -3595 14950 -3475
rect 15005 -3595 15125 -3475
rect 15170 -3595 15290 -3475
rect 15335 -3595 15455 -3475
rect 15500 -3595 15620 -3475
rect 15675 -3595 15795 -3475
rect 15840 -3595 15960 -3475
rect 16005 -3595 16125 -3475
rect 16170 -3595 16290 -3475
rect 16345 -3595 16465 -3475
rect 16510 -3595 16630 -3475
rect 16675 -3595 16795 -3475
rect 16840 -3595 16960 -3475
rect 17015 -3595 17135 -3475
rect 17180 -3595 17300 -3475
rect 17345 -3595 17465 -3475
rect 17510 -3595 17630 -3475
rect 17685 -3595 17805 -3475
rect 17850 -3595 17970 -3475
rect 18015 -3595 18135 -3475
rect 18180 -3595 18300 -3475
rect 12820 -3760 12940 -3640
rect 12995 -3760 13115 -3640
rect 13160 -3760 13280 -3640
rect 13325 -3760 13445 -3640
rect 13490 -3760 13610 -3640
rect 13665 -3760 13785 -3640
rect 13830 -3760 13950 -3640
rect 13995 -3760 14115 -3640
rect 14160 -3760 14280 -3640
rect 14335 -3760 14455 -3640
rect 14500 -3760 14620 -3640
rect 14665 -3760 14785 -3640
rect 14830 -3760 14950 -3640
rect 15005 -3760 15125 -3640
rect 15170 -3760 15290 -3640
rect 15335 -3760 15455 -3640
rect 15500 -3760 15620 -3640
rect 15675 -3760 15795 -3640
rect 15840 -3760 15960 -3640
rect 16005 -3760 16125 -3640
rect 16170 -3760 16290 -3640
rect 16345 -3760 16465 -3640
rect 16510 -3760 16630 -3640
rect 16675 -3760 16795 -3640
rect 16840 -3760 16960 -3640
rect 17015 -3760 17135 -3640
rect 17180 -3760 17300 -3640
rect 17345 -3760 17465 -3640
rect 17510 -3760 17630 -3640
rect 17685 -3760 17805 -3640
rect 17850 -3760 17970 -3640
rect 18015 -3760 18135 -3640
rect 18180 -3760 18300 -3640
rect 12820 -3925 12940 -3805
rect 12995 -3925 13115 -3805
rect 13160 -3925 13280 -3805
rect 13325 -3925 13445 -3805
rect 13490 -3925 13610 -3805
rect 13665 -3925 13785 -3805
rect 13830 -3925 13950 -3805
rect 13995 -3925 14115 -3805
rect 14160 -3925 14280 -3805
rect 14335 -3925 14455 -3805
rect 14500 -3925 14620 -3805
rect 14665 -3925 14785 -3805
rect 14830 -3925 14950 -3805
rect 15005 -3925 15125 -3805
rect 15170 -3925 15290 -3805
rect 15335 -3925 15455 -3805
rect 15500 -3925 15620 -3805
rect 15675 -3925 15795 -3805
rect 15840 -3925 15960 -3805
rect 16005 -3925 16125 -3805
rect 16170 -3925 16290 -3805
rect 16345 -3925 16465 -3805
rect 16510 -3925 16630 -3805
rect 16675 -3925 16795 -3805
rect 16840 -3925 16960 -3805
rect 17015 -3925 17135 -3805
rect 17180 -3925 17300 -3805
rect 17345 -3925 17465 -3805
rect 17510 -3925 17630 -3805
rect 17685 -3925 17805 -3805
rect 17850 -3925 17970 -3805
rect 18015 -3925 18135 -3805
rect 18180 -3925 18300 -3805
rect 12820 -4100 12940 -3980
rect 12995 -4100 13115 -3980
rect 13160 -4100 13280 -3980
rect 13325 -4100 13445 -3980
rect 13490 -4100 13610 -3980
rect 13665 -4100 13785 -3980
rect 13830 -4100 13950 -3980
rect 13995 -4100 14115 -3980
rect 14160 -4100 14280 -3980
rect 14335 -4100 14455 -3980
rect 14500 -4100 14620 -3980
rect 14665 -4100 14785 -3980
rect 14830 -4100 14950 -3980
rect 15005 -4100 15125 -3980
rect 15170 -4100 15290 -3980
rect 15335 -4100 15455 -3980
rect 15500 -4100 15620 -3980
rect 15675 -4100 15795 -3980
rect 15840 -4100 15960 -3980
rect 16005 -4100 16125 -3980
rect 16170 -4100 16290 -3980
rect 16345 -4100 16465 -3980
rect 16510 -4100 16630 -3980
rect 16675 -4100 16795 -3980
rect 16840 -4100 16960 -3980
rect 17015 -4100 17135 -3980
rect 17180 -4100 17300 -3980
rect 17345 -4100 17465 -3980
rect 17510 -4100 17630 -3980
rect 17685 -4100 17805 -3980
rect 17850 -4100 17970 -3980
rect 18015 -4100 18135 -3980
rect 18180 -4100 18300 -3980
rect 18510 1260 18630 1380
rect 18685 1260 18805 1380
rect 18850 1260 18970 1380
rect 19015 1260 19135 1380
rect 19180 1260 19300 1380
rect 19355 1260 19475 1380
rect 19520 1260 19640 1380
rect 19685 1260 19805 1380
rect 19850 1260 19970 1380
rect 20025 1260 20145 1380
rect 20190 1260 20310 1380
rect 20355 1260 20475 1380
rect 20520 1260 20640 1380
rect 20695 1260 20815 1380
rect 20860 1260 20980 1380
rect 21025 1260 21145 1380
rect 21190 1260 21310 1380
rect 21365 1260 21485 1380
rect 21530 1260 21650 1380
rect 21695 1260 21815 1380
rect 21860 1260 21980 1380
rect 22035 1260 22155 1380
rect 22200 1260 22320 1380
rect 22365 1260 22485 1380
rect 22530 1260 22650 1380
rect 22705 1260 22825 1380
rect 22870 1260 22990 1380
rect 23035 1260 23155 1380
rect 23200 1260 23320 1380
rect 23375 1260 23495 1380
rect 23540 1260 23660 1380
rect 23705 1260 23825 1380
rect 23870 1260 23990 1380
rect 18510 1095 18630 1215
rect 18685 1095 18805 1215
rect 18850 1095 18970 1215
rect 19015 1095 19135 1215
rect 19180 1095 19300 1215
rect 19355 1095 19475 1215
rect 19520 1095 19640 1215
rect 19685 1095 19805 1215
rect 19850 1095 19970 1215
rect 20025 1095 20145 1215
rect 20190 1095 20310 1215
rect 20355 1095 20475 1215
rect 20520 1095 20640 1215
rect 20695 1095 20815 1215
rect 20860 1095 20980 1215
rect 21025 1095 21145 1215
rect 21190 1095 21310 1215
rect 21365 1095 21485 1215
rect 21530 1095 21650 1215
rect 21695 1095 21815 1215
rect 21860 1095 21980 1215
rect 22035 1095 22155 1215
rect 22200 1095 22320 1215
rect 22365 1095 22485 1215
rect 22530 1095 22650 1215
rect 22705 1095 22825 1215
rect 22870 1095 22990 1215
rect 23035 1095 23155 1215
rect 23200 1095 23320 1215
rect 23375 1095 23495 1215
rect 23540 1095 23660 1215
rect 23705 1095 23825 1215
rect 23870 1095 23990 1215
rect 18510 930 18630 1050
rect 18685 930 18805 1050
rect 18850 930 18970 1050
rect 19015 930 19135 1050
rect 19180 930 19300 1050
rect 19355 930 19475 1050
rect 19520 930 19640 1050
rect 19685 930 19805 1050
rect 19850 930 19970 1050
rect 20025 930 20145 1050
rect 20190 930 20310 1050
rect 20355 930 20475 1050
rect 20520 930 20640 1050
rect 20695 930 20815 1050
rect 20860 930 20980 1050
rect 21025 930 21145 1050
rect 21190 930 21310 1050
rect 21365 930 21485 1050
rect 21530 930 21650 1050
rect 21695 930 21815 1050
rect 21860 930 21980 1050
rect 22035 930 22155 1050
rect 22200 930 22320 1050
rect 22365 930 22485 1050
rect 22530 930 22650 1050
rect 22705 930 22825 1050
rect 22870 930 22990 1050
rect 23035 930 23155 1050
rect 23200 930 23320 1050
rect 23375 930 23495 1050
rect 23540 930 23660 1050
rect 23705 930 23825 1050
rect 23870 930 23990 1050
rect 18510 765 18630 885
rect 18685 765 18805 885
rect 18850 765 18970 885
rect 19015 765 19135 885
rect 19180 765 19300 885
rect 19355 765 19475 885
rect 19520 765 19640 885
rect 19685 765 19805 885
rect 19850 765 19970 885
rect 20025 765 20145 885
rect 20190 765 20310 885
rect 20355 765 20475 885
rect 20520 765 20640 885
rect 20695 765 20815 885
rect 20860 765 20980 885
rect 21025 765 21145 885
rect 21190 765 21310 885
rect 21365 765 21485 885
rect 21530 765 21650 885
rect 21695 765 21815 885
rect 21860 765 21980 885
rect 22035 765 22155 885
rect 22200 765 22320 885
rect 22365 765 22485 885
rect 22530 765 22650 885
rect 22705 765 22825 885
rect 22870 765 22990 885
rect 23035 765 23155 885
rect 23200 765 23320 885
rect 23375 765 23495 885
rect 23540 765 23660 885
rect 23705 765 23825 885
rect 23870 765 23990 885
rect 18510 590 18630 710
rect 18685 590 18805 710
rect 18850 590 18970 710
rect 19015 590 19135 710
rect 19180 590 19300 710
rect 19355 590 19475 710
rect 19520 590 19640 710
rect 19685 590 19805 710
rect 19850 590 19970 710
rect 20025 590 20145 710
rect 20190 590 20310 710
rect 20355 590 20475 710
rect 20520 590 20640 710
rect 20695 590 20815 710
rect 20860 590 20980 710
rect 21025 590 21145 710
rect 21190 590 21310 710
rect 21365 590 21485 710
rect 21530 590 21650 710
rect 21695 590 21815 710
rect 21860 590 21980 710
rect 22035 590 22155 710
rect 22200 590 22320 710
rect 22365 590 22485 710
rect 22530 590 22650 710
rect 22705 590 22825 710
rect 22870 590 22990 710
rect 23035 590 23155 710
rect 23200 590 23320 710
rect 23375 590 23495 710
rect 23540 590 23660 710
rect 23705 590 23825 710
rect 23870 590 23990 710
rect 18510 425 18630 545
rect 18685 425 18805 545
rect 18850 425 18970 545
rect 19015 425 19135 545
rect 19180 425 19300 545
rect 19355 425 19475 545
rect 19520 425 19640 545
rect 19685 425 19805 545
rect 19850 425 19970 545
rect 20025 425 20145 545
rect 20190 425 20310 545
rect 20355 425 20475 545
rect 20520 425 20640 545
rect 20695 425 20815 545
rect 20860 425 20980 545
rect 21025 425 21145 545
rect 21190 425 21310 545
rect 21365 425 21485 545
rect 21530 425 21650 545
rect 21695 425 21815 545
rect 21860 425 21980 545
rect 22035 425 22155 545
rect 22200 425 22320 545
rect 22365 425 22485 545
rect 22530 425 22650 545
rect 22705 425 22825 545
rect 22870 425 22990 545
rect 23035 425 23155 545
rect 23200 425 23320 545
rect 23375 425 23495 545
rect 23540 425 23660 545
rect 23705 425 23825 545
rect 23870 425 23990 545
rect 18510 260 18630 380
rect 18685 260 18805 380
rect 18850 260 18970 380
rect 19015 260 19135 380
rect 19180 260 19300 380
rect 19355 260 19475 380
rect 19520 260 19640 380
rect 19685 260 19805 380
rect 19850 260 19970 380
rect 20025 260 20145 380
rect 20190 260 20310 380
rect 20355 260 20475 380
rect 20520 260 20640 380
rect 20695 260 20815 380
rect 20860 260 20980 380
rect 21025 260 21145 380
rect 21190 260 21310 380
rect 21365 260 21485 380
rect 21530 260 21650 380
rect 21695 260 21815 380
rect 21860 260 21980 380
rect 22035 260 22155 380
rect 22200 260 22320 380
rect 22365 260 22485 380
rect 22530 260 22650 380
rect 22705 260 22825 380
rect 22870 260 22990 380
rect 23035 260 23155 380
rect 23200 260 23320 380
rect 23375 260 23495 380
rect 23540 260 23660 380
rect 23705 260 23825 380
rect 23870 260 23990 380
rect 18510 95 18630 215
rect 18685 95 18805 215
rect 18850 95 18970 215
rect 19015 95 19135 215
rect 19180 95 19300 215
rect 19355 95 19475 215
rect 19520 95 19640 215
rect 19685 95 19805 215
rect 19850 95 19970 215
rect 20025 95 20145 215
rect 20190 95 20310 215
rect 20355 95 20475 215
rect 20520 95 20640 215
rect 20695 95 20815 215
rect 20860 95 20980 215
rect 21025 95 21145 215
rect 21190 95 21310 215
rect 21365 95 21485 215
rect 21530 95 21650 215
rect 21695 95 21815 215
rect 21860 95 21980 215
rect 22035 95 22155 215
rect 22200 95 22320 215
rect 22365 95 22485 215
rect 22530 95 22650 215
rect 22705 95 22825 215
rect 22870 95 22990 215
rect 23035 95 23155 215
rect 23200 95 23320 215
rect 23375 95 23495 215
rect 23540 95 23660 215
rect 23705 95 23825 215
rect 23870 95 23990 215
rect 18510 -80 18630 40
rect 18685 -80 18805 40
rect 18850 -80 18970 40
rect 19015 -80 19135 40
rect 19180 -80 19300 40
rect 19355 -80 19475 40
rect 19520 -80 19640 40
rect 19685 -80 19805 40
rect 19850 -80 19970 40
rect 20025 -80 20145 40
rect 20190 -80 20310 40
rect 20355 -80 20475 40
rect 20520 -80 20640 40
rect 20695 -80 20815 40
rect 20860 -80 20980 40
rect 21025 -80 21145 40
rect 21190 -80 21310 40
rect 21365 -80 21485 40
rect 21530 -80 21650 40
rect 21695 -80 21815 40
rect 21860 -80 21980 40
rect 22035 -80 22155 40
rect 22200 -80 22320 40
rect 22365 -80 22485 40
rect 22530 -80 22650 40
rect 22705 -80 22825 40
rect 22870 -80 22990 40
rect 23035 -80 23155 40
rect 23200 -80 23320 40
rect 23375 -80 23495 40
rect 23540 -80 23660 40
rect 23705 -80 23825 40
rect 23870 -80 23990 40
rect 18510 -245 18630 -125
rect 18685 -245 18805 -125
rect 18850 -245 18970 -125
rect 19015 -245 19135 -125
rect 19180 -245 19300 -125
rect 19355 -245 19475 -125
rect 19520 -245 19640 -125
rect 19685 -245 19805 -125
rect 19850 -245 19970 -125
rect 20025 -245 20145 -125
rect 20190 -245 20310 -125
rect 20355 -245 20475 -125
rect 20520 -245 20640 -125
rect 20695 -245 20815 -125
rect 20860 -245 20980 -125
rect 21025 -245 21145 -125
rect 21190 -245 21310 -125
rect 21365 -245 21485 -125
rect 21530 -245 21650 -125
rect 21695 -245 21815 -125
rect 21860 -245 21980 -125
rect 22035 -245 22155 -125
rect 22200 -245 22320 -125
rect 22365 -245 22485 -125
rect 22530 -245 22650 -125
rect 22705 -245 22825 -125
rect 22870 -245 22990 -125
rect 23035 -245 23155 -125
rect 23200 -245 23320 -125
rect 23375 -245 23495 -125
rect 23540 -245 23660 -125
rect 23705 -245 23825 -125
rect 23870 -245 23990 -125
rect 18510 -410 18630 -290
rect 18685 -410 18805 -290
rect 18850 -410 18970 -290
rect 19015 -410 19135 -290
rect 19180 -410 19300 -290
rect 19355 -410 19475 -290
rect 19520 -410 19640 -290
rect 19685 -410 19805 -290
rect 19850 -410 19970 -290
rect 20025 -410 20145 -290
rect 20190 -410 20310 -290
rect 20355 -410 20475 -290
rect 20520 -410 20640 -290
rect 20695 -410 20815 -290
rect 20860 -410 20980 -290
rect 21025 -410 21145 -290
rect 21190 -410 21310 -290
rect 21365 -410 21485 -290
rect 21530 -410 21650 -290
rect 21695 -410 21815 -290
rect 21860 -410 21980 -290
rect 22035 -410 22155 -290
rect 22200 -410 22320 -290
rect 22365 -410 22485 -290
rect 22530 -410 22650 -290
rect 22705 -410 22825 -290
rect 22870 -410 22990 -290
rect 23035 -410 23155 -290
rect 23200 -410 23320 -290
rect 23375 -410 23495 -290
rect 23540 -410 23660 -290
rect 23705 -410 23825 -290
rect 23870 -410 23990 -290
rect 18510 -575 18630 -455
rect 18685 -575 18805 -455
rect 18850 -575 18970 -455
rect 19015 -575 19135 -455
rect 19180 -575 19300 -455
rect 19355 -575 19475 -455
rect 19520 -575 19640 -455
rect 19685 -575 19805 -455
rect 19850 -575 19970 -455
rect 20025 -575 20145 -455
rect 20190 -575 20310 -455
rect 20355 -575 20475 -455
rect 20520 -575 20640 -455
rect 20695 -575 20815 -455
rect 20860 -575 20980 -455
rect 21025 -575 21145 -455
rect 21190 -575 21310 -455
rect 21365 -575 21485 -455
rect 21530 -575 21650 -455
rect 21695 -575 21815 -455
rect 21860 -575 21980 -455
rect 22035 -575 22155 -455
rect 22200 -575 22320 -455
rect 22365 -575 22485 -455
rect 22530 -575 22650 -455
rect 22705 -575 22825 -455
rect 22870 -575 22990 -455
rect 23035 -575 23155 -455
rect 23200 -575 23320 -455
rect 23375 -575 23495 -455
rect 23540 -575 23660 -455
rect 23705 -575 23825 -455
rect 23870 -575 23990 -455
rect 18510 -750 18630 -630
rect 18685 -750 18805 -630
rect 18850 -750 18970 -630
rect 19015 -750 19135 -630
rect 19180 -750 19300 -630
rect 19355 -750 19475 -630
rect 19520 -750 19640 -630
rect 19685 -750 19805 -630
rect 19850 -750 19970 -630
rect 20025 -750 20145 -630
rect 20190 -750 20310 -630
rect 20355 -750 20475 -630
rect 20520 -750 20640 -630
rect 20695 -750 20815 -630
rect 20860 -750 20980 -630
rect 21025 -750 21145 -630
rect 21190 -750 21310 -630
rect 21365 -750 21485 -630
rect 21530 -750 21650 -630
rect 21695 -750 21815 -630
rect 21860 -750 21980 -630
rect 22035 -750 22155 -630
rect 22200 -750 22320 -630
rect 22365 -750 22485 -630
rect 22530 -750 22650 -630
rect 22705 -750 22825 -630
rect 22870 -750 22990 -630
rect 23035 -750 23155 -630
rect 23200 -750 23320 -630
rect 23375 -750 23495 -630
rect 23540 -750 23660 -630
rect 23705 -750 23825 -630
rect 23870 -750 23990 -630
rect 18510 -915 18630 -795
rect 18685 -915 18805 -795
rect 18850 -915 18970 -795
rect 19015 -915 19135 -795
rect 19180 -915 19300 -795
rect 19355 -915 19475 -795
rect 19520 -915 19640 -795
rect 19685 -915 19805 -795
rect 19850 -915 19970 -795
rect 20025 -915 20145 -795
rect 20190 -915 20310 -795
rect 20355 -915 20475 -795
rect 20520 -915 20640 -795
rect 20695 -915 20815 -795
rect 20860 -915 20980 -795
rect 21025 -915 21145 -795
rect 21190 -915 21310 -795
rect 21365 -915 21485 -795
rect 21530 -915 21650 -795
rect 21695 -915 21815 -795
rect 21860 -915 21980 -795
rect 22035 -915 22155 -795
rect 22200 -915 22320 -795
rect 22365 -915 22485 -795
rect 22530 -915 22650 -795
rect 22705 -915 22825 -795
rect 22870 -915 22990 -795
rect 23035 -915 23155 -795
rect 23200 -915 23320 -795
rect 23375 -915 23495 -795
rect 23540 -915 23660 -795
rect 23705 -915 23825 -795
rect 23870 -915 23990 -795
rect 18510 -1080 18630 -960
rect 18685 -1080 18805 -960
rect 18850 -1080 18970 -960
rect 19015 -1080 19135 -960
rect 19180 -1080 19300 -960
rect 19355 -1080 19475 -960
rect 19520 -1080 19640 -960
rect 19685 -1080 19805 -960
rect 19850 -1080 19970 -960
rect 20025 -1080 20145 -960
rect 20190 -1080 20310 -960
rect 20355 -1080 20475 -960
rect 20520 -1080 20640 -960
rect 20695 -1080 20815 -960
rect 20860 -1080 20980 -960
rect 21025 -1080 21145 -960
rect 21190 -1080 21310 -960
rect 21365 -1080 21485 -960
rect 21530 -1080 21650 -960
rect 21695 -1080 21815 -960
rect 21860 -1080 21980 -960
rect 22035 -1080 22155 -960
rect 22200 -1080 22320 -960
rect 22365 -1080 22485 -960
rect 22530 -1080 22650 -960
rect 22705 -1080 22825 -960
rect 22870 -1080 22990 -960
rect 23035 -1080 23155 -960
rect 23200 -1080 23320 -960
rect 23375 -1080 23495 -960
rect 23540 -1080 23660 -960
rect 23705 -1080 23825 -960
rect 23870 -1080 23990 -960
rect 18510 -1245 18630 -1125
rect 18685 -1245 18805 -1125
rect 18850 -1245 18970 -1125
rect 19015 -1245 19135 -1125
rect 19180 -1245 19300 -1125
rect 19355 -1245 19475 -1125
rect 19520 -1245 19640 -1125
rect 19685 -1245 19805 -1125
rect 19850 -1245 19970 -1125
rect 20025 -1245 20145 -1125
rect 20190 -1245 20310 -1125
rect 20355 -1245 20475 -1125
rect 20520 -1245 20640 -1125
rect 20695 -1245 20815 -1125
rect 20860 -1245 20980 -1125
rect 21025 -1245 21145 -1125
rect 21190 -1245 21310 -1125
rect 21365 -1245 21485 -1125
rect 21530 -1245 21650 -1125
rect 21695 -1245 21815 -1125
rect 21860 -1245 21980 -1125
rect 22035 -1245 22155 -1125
rect 22200 -1245 22320 -1125
rect 22365 -1245 22485 -1125
rect 22530 -1245 22650 -1125
rect 22705 -1245 22825 -1125
rect 22870 -1245 22990 -1125
rect 23035 -1245 23155 -1125
rect 23200 -1245 23320 -1125
rect 23375 -1245 23495 -1125
rect 23540 -1245 23660 -1125
rect 23705 -1245 23825 -1125
rect 23870 -1245 23990 -1125
rect 18510 -1420 18630 -1300
rect 18685 -1420 18805 -1300
rect 18850 -1420 18970 -1300
rect 19015 -1420 19135 -1300
rect 19180 -1420 19300 -1300
rect 19355 -1420 19475 -1300
rect 19520 -1420 19640 -1300
rect 19685 -1420 19805 -1300
rect 19850 -1420 19970 -1300
rect 20025 -1420 20145 -1300
rect 20190 -1420 20310 -1300
rect 20355 -1420 20475 -1300
rect 20520 -1420 20640 -1300
rect 20695 -1420 20815 -1300
rect 20860 -1420 20980 -1300
rect 21025 -1420 21145 -1300
rect 21190 -1420 21310 -1300
rect 21365 -1420 21485 -1300
rect 21530 -1420 21650 -1300
rect 21695 -1420 21815 -1300
rect 21860 -1420 21980 -1300
rect 22035 -1420 22155 -1300
rect 22200 -1420 22320 -1300
rect 22365 -1420 22485 -1300
rect 22530 -1420 22650 -1300
rect 22705 -1420 22825 -1300
rect 22870 -1420 22990 -1300
rect 23035 -1420 23155 -1300
rect 23200 -1420 23320 -1300
rect 23375 -1420 23495 -1300
rect 23540 -1420 23660 -1300
rect 23705 -1420 23825 -1300
rect 23870 -1420 23990 -1300
rect 18510 -1585 18630 -1465
rect 18685 -1585 18805 -1465
rect 18850 -1585 18970 -1465
rect 19015 -1585 19135 -1465
rect 19180 -1585 19300 -1465
rect 19355 -1585 19475 -1465
rect 19520 -1585 19640 -1465
rect 19685 -1585 19805 -1465
rect 19850 -1585 19970 -1465
rect 20025 -1585 20145 -1465
rect 20190 -1585 20310 -1465
rect 20355 -1585 20475 -1465
rect 20520 -1585 20640 -1465
rect 20695 -1585 20815 -1465
rect 20860 -1585 20980 -1465
rect 21025 -1585 21145 -1465
rect 21190 -1585 21310 -1465
rect 21365 -1585 21485 -1465
rect 21530 -1585 21650 -1465
rect 21695 -1585 21815 -1465
rect 21860 -1585 21980 -1465
rect 22035 -1585 22155 -1465
rect 22200 -1585 22320 -1465
rect 22365 -1585 22485 -1465
rect 22530 -1585 22650 -1465
rect 22705 -1585 22825 -1465
rect 22870 -1585 22990 -1465
rect 23035 -1585 23155 -1465
rect 23200 -1585 23320 -1465
rect 23375 -1585 23495 -1465
rect 23540 -1585 23660 -1465
rect 23705 -1585 23825 -1465
rect 23870 -1585 23990 -1465
rect 18510 -1750 18630 -1630
rect 18685 -1750 18805 -1630
rect 18850 -1750 18970 -1630
rect 19015 -1750 19135 -1630
rect 19180 -1750 19300 -1630
rect 19355 -1750 19475 -1630
rect 19520 -1750 19640 -1630
rect 19685 -1750 19805 -1630
rect 19850 -1750 19970 -1630
rect 20025 -1750 20145 -1630
rect 20190 -1750 20310 -1630
rect 20355 -1750 20475 -1630
rect 20520 -1750 20640 -1630
rect 20695 -1750 20815 -1630
rect 20860 -1750 20980 -1630
rect 21025 -1750 21145 -1630
rect 21190 -1750 21310 -1630
rect 21365 -1750 21485 -1630
rect 21530 -1750 21650 -1630
rect 21695 -1750 21815 -1630
rect 21860 -1750 21980 -1630
rect 22035 -1750 22155 -1630
rect 22200 -1750 22320 -1630
rect 22365 -1750 22485 -1630
rect 22530 -1750 22650 -1630
rect 22705 -1750 22825 -1630
rect 22870 -1750 22990 -1630
rect 23035 -1750 23155 -1630
rect 23200 -1750 23320 -1630
rect 23375 -1750 23495 -1630
rect 23540 -1750 23660 -1630
rect 23705 -1750 23825 -1630
rect 23870 -1750 23990 -1630
rect 18510 -1915 18630 -1795
rect 18685 -1915 18805 -1795
rect 18850 -1915 18970 -1795
rect 19015 -1915 19135 -1795
rect 19180 -1915 19300 -1795
rect 19355 -1915 19475 -1795
rect 19520 -1915 19640 -1795
rect 19685 -1915 19805 -1795
rect 19850 -1915 19970 -1795
rect 20025 -1915 20145 -1795
rect 20190 -1915 20310 -1795
rect 20355 -1915 20475 -1795
rect 20520 -1915 20640 -1795
rect 20695 -1915 20815 -1795
rect 20860 -1915 20980 -1795
rect 21025 -1915 21145 -1795
rect 21190 -1915 21310 -1795
rect 21365 -1915 21485 -1795
rect 21530 -1915 21650 -1795
rect 21695 -1915 21815 -1795
rect 21860 -1915 21980 -1795
rect 22035 -1915 22155 -1795
rect 22200 -1915 22320 -1795
rect 22365 -1915 22485 -1795
rect 22530 -1915 22650 -1795
rect 22705 -1915 22825 -1795
rect 22870 -1915 22990 -1795
rect 23035 -1915 23155 -1795
rect 23200 -1915 23320 -1795
rect 23375 -1915 23495 -1795
rect 23540 -1915 23660 -1795
rect 23705 -1915 23825 -1795
rect 23870 -1915 23990 -1795
rect 18510 -2090 18630 -1970
rect 18685 -2090 18805 -1970
rect 18850 -2090 18970 -1970
rect 19015 -2090 19135 -1970
rect 19180 -2090 19300 -1970
rect 19355 -2090 19475 -1970
rect 19520 -2090 19640 -1970
rect 19685 -2090 19805 -1970
rect 19850 -2090 19970 -1970
rect 20025 -2090 20145 -1970
rect 20190 -2090 20310 -1970
rect 20355 -2090 20475 -1970
rect 20520 -2090 20640 -1970
rect 20695 -2090 20815 -1970
rect 20860 -2090 20980 -1970
rect 21025 -2090 21145 -1970
rect 21190 -2090 21310 -1970
rect 21365 -2090 21485 -1970
rect 21530 -2090 21650 -1970
rect 21695 -2090 21815 -1970
rect 21860 -2090 21980 -1970
rect 22035 -2090 22155 -1970
rect 22200 -2090 22320 -1970
rect 22365 -2090 22485 -1970
rect 22530 -2090 22650 -1970
rect 22705 -2090 22825 -1970
rect 22870 -2090 22990 -1970
rect 23035 -2090 23155 -1970
rect 23200 -2090 23320 -1970
rect 23375 -2090 23495 -1970
rect 23540 -2090 23660 -1970
rect 23705 -2090 23825 -1970
rect 23870 -2090 23990 -1970
rect 18510 -2255 18630 -2135
rect 18685 -2255 18805 -2135
rect 18850 -2255 18970 -2135
rect 19015 -2255 19135 -2135
rect 19180 -2255 19300 -2135
rect 19355 -2255 19475 -2135
rect 19520 -2255 19640 -2135
rect 19685 -2255 19805 -2135
rect 19850 -2255 19970 -2135
rect 20025 -2255 20145 -2135
rect 20190 -2255 20310 -2135
rect 20355 -2255 20475 -2135
rect 20520 -2255 20640 -2135
rect 20695 -2255 20815 -2135
rect 20860 -2255 20980 -2135
rect 21025 -2255 21145 -2135
rect 21190 -2255 21310 -2135
rect 21365 -2255 21485 -2135
rect 21530 -2255 21650 -2135
rect 21695 -2255 21815 -2135
rect 21860 -2255 21980 -2135
rect 22035 -2255 22155 -2135
rect 22200 -2255 22320 -2135
rect 22365 -2255 22485 -2135
rect 22530 -2255 22650 -2135
rect 22705 -2255 22825 -2135
rect 22870 -2255 22990 -2135
rect 23035 -2255 23155 -2135
rect 23200 -2255 23320 -2135
rect 23375 -2255 23495 -2135
rect 23540 -2255 23660 -2135
rect 23705 -2255 23825 -2135
rect 23870 -2255 23990 -2135
rect 18510 -2420 18630 -2300
rect 18685 -2420 18805 -2300
rect 18850 -2420 18970 -2300
rect 19015 -2420 19135 -2300
rect 19180 -2420 19300 -2300
rect 19355 -2420 19475 -2300
rect 19520 -2420 19640 -2300
rect 19685 -2420 19805 -2300
rect 19850 -2420 19970 -2300
rect 20025 -2420 20145 -2300
rect 20190 -2420 20310 -2300
rect 20355 -2420 20475 -2300
rect 20520 -2420 20640 -2300
rect 20695 -2420 20815 -2300
rect 20860 -2420 20980 -2300
rect 21025 -2420 21145 -2300
rect 21190 -2420 21310 -2300
rect 21365 -2420 21485 -2300
rect 21530 -2420 21650 -2300
rect 21695 -2420 21815 -2300
rect 21860 -2420 21980 -2300
rect 22035 -2420 22155 -2300
rect 22200 -2420 22320 -2300
rect 22365 -2420 22485 -2300
rect 22530 -2420 22650 -2300
rect 22705 -2420 22825 -2300
rect 22870 -2420 22990 -2300
rect 23035 -2420 23155 -2300
rect 23200 -2420 23320 -2300
rect 23375 -2420 23495 -2300
rect 23540 -2420 23660 -2300
rect 23705 -2420 23825 -2300
rect 23870 -2420 23990 -2300
rect 18510 -2585 18630 -2465
rect 18685 -2585 18805 -2465
rect 18850 -2585 18970 -2465
rect 19015 -2585 19135 -2465
rect 19180 -2585 19300 -2465
rect 19355 -2585 19475 -2465
rect 19520 -2585 19640 -2465
rect 19685 -2585 19805 -2465
rect 19850 -2585 19970 -2465
rect 20025 -2585 20145 -2465
rect 20190 -2585 20310 -2465
rect 20355 -2585 20475 -2465
rect 20520 -2585 20640 -2465
rect 20695 -2585 20815 -2465
rect 20860 -2585 20980 -2465
rect 21025 -2585 21145 -2465
rect 21190 -2585 21310 -2465
rect 21365 -2585 21485 -2465
rect 21530 -2585 21650 -2465
rect 21695 -2585 21815 -2465
rect 21860 -2585 21980 -2465
rect 22035 -2585 22155 -2465
rect 22200 -2585 22320 -2465
rect 22365 -2585 22485 -2465
rect 22530 -2585 22650 -2465
rect 22705 -2585 22825 -2465
rect 22870 -2585 22990 -2465
rect 23035 -2585 23155 -2465
rect 23200 -2585 23320 -2465
rect 23375 -2585 23495 -2465
rect 23540 -2585 23660 -2465
rect 23705 -2585 23825 -2465
rect 23870 -2585 23990 -2465
rect 18510 -2760 18630 -2640
rect 18685 -2760 18805 -2640
rect 18850 -2760 18970 -2640
rect 19015 -2760 19135 -2640
rect 19180 -2760 19300 -2640
rect 19355 -2760 19475 -2640
rect 19520 -2760 19640 -2640
rect 19685 -2760 19805 -2640
rect 19850 -2760 19970 -2640
rect 20025 -2760 20145 -2640
rect 20190 -2760 20310 -2640
rect 20355 -2760 20475 -2640
rect 20520 -2760 20640 -2640
rect 20695 -2760 20815 -2640
rect 20860 -2760 20980 -2640
rect 21025 -2760 21145 -2640
rect 21190 -2760 21310 -2640
rect 21365 -2760 21485 -2640
rect 21530 -2760 21650 -2640
rect 21695 -2760 21815 -2640
rect 21860 -2760 21980 -2640
rect 22035 -2760 22155 -2640
rect 22200 -2760 22320 -2640
rect 22365 -2760 22485 -2640
rect 22530 -2760 22650 -2640
rect 22705 -2760 22825 -2640
rect 22870 -2760 22990 -2640
rect 23035 -2760 23155 -2640
rect 23200 -2760 23320 -2640
rect 23375 -2760 23495 -2640
rect 23540 -2760 23660 -2640
rect 23705 -2760 23825 -2640
rect 23870 -2760 23990 -2640
rect 18510 -2925 18630 -2805
rect 18685 -2925 18805 -2805
rect 18850 -2925 18970 -2805
rect 19015 -2925 19135 -2805
rect 19180 -2925 19300 -2805
rect 19355 -2925 19475 -2805
rect 19520 -2925 19640 -2805
rect 19685 -2925 19805 -2805
rect 19850 -2925 19970 -2805
rect 20025 -2925 20145 -2805
rect 20190 -2925 20310 -2805
rect 20355 -2925 20475 -2805
rect 20520 -2925 20640 -2805
rect 20695 -2925 20815 -2805
rect 20860 -2925 20980 -2805
rect 21025 -2925 21145 -2805
rect 21190 -2925 21310 -2805
rect 21365 -2925 21485 -2805
rect 21530 -2925 21650 -2805
rect 21695 -2925 21815 -2805
rect 21860 -2925 21980 -2805
rect 22035 -2925 22155 -2805
rect 22200 -2925 22320 -2805
rect 22365 -2925 22485 -2805
rect 22530 -2925 22650 -2805
rect 22705 -2925 22825 -2805
rect 22870 -2925 22990 -2805
rect 23035 -2925 23155 -2805
rect 23200 -2925 23320 -2805
rect 23375 -2925 23495 -2805
rect 23540 -2925 23660 -2805
rect 23705 -2925 23825 -2805
rect 23870 -2925 23990 -2805
rect 18510 -3090 18630 -2970
rect 18685 -3090 18805 -2970
rect 18850 -3090 18970 -2970
rect 19015 -3090 19135 -2970
rect 19180 -3090 19300 -2970
rect 19355 -3090 19475 -2970
rect 19520 -3090 19640 -2970
rect 19685 -3090 19805 -2970
rect 19850 -3090 19970 -2970
rect 20025 -3090 20145 -2970
rect 20190 -3090 20310 -2970
rect 20355 -3090 20475 -2970
rect 20520 -3090 20640 -2970
rect 20695 -3090 20815 -2970
rect 20860 -3090 20980 -2970
rect 21025 -3090 21145 -2970
rect 21190 -3090 21310 -2970
rect 21365 -3090 21485 -2970
rect 21530 -3090 21650 -2970
rect 21695 -3090 21815 -2970
rect 21860 -3090 21980 -2970
rect 22035 -3090 22155 -2970
rect 22200 -3090 22320 -2970
rect 22365 -3090 22485 -2970
rect 22530 -3090 22650 -2970
rect 22705 -3090 22825 -2970
rect 22870 -3090 22990 -2970
rect 23035 -3090 23155 -2970
rect 23200 -3090 23320 -2970
rect 23375 -3090 23495 -2970
rect 23540 -3090 23660 -2970
rect 23705 -3090 23825 -2970
rect 23870 -3090 23990 -2970
rect 18510 -3255 18630 -3135
rect 18685 -3255 18805 -3135
rect 18850 -3255 18970 -3135
rect 19015 -3255 19135 -3135
rect 19180 -3255 19300 -3135
rect 19355 -3255 19475 -3135
rect 19520 -3255 19640 -3135
rect 19685 -3255 19805 -3135
rect 19850 -3255 19970 -3135
rect 20025 -3255 20145 -3135
rect 20190 -3255 20310 -3135
rect 20355 -3255 20475 -3135
rect 20520 -3255 20640 -3135
rect 20695 -3255 20815 -3135
rect 20860 -3255 20980 -3135
rect 21025 -3255 21145 -3135
rect 21190 -3255 21310 -3135
rect 21365 -3255 21485 -3135
rect 21530 -3255 21650 -3135
rect 21695 -3255 21815 -3135
rect 21860 -3255 21980 -3135
rect 22035 -3255 22155 -3135
rect 22200 -3255 22320 -3135
rect 22365 -3255 22485 -3135
rect 22530 -3255 22650 -3135
rect 22705 -3255 22825 -3135
rect 22870 -3255 22990 -3135
rect 23035 -3255 23155 -3135
rect 23200 -3255 23320 -3135
rect 23375 -3255 23495 -3135
rect 23540 -3255 23660 -3135
rect 23705 -3255 23825 -3135
rect 23870 -3255 23990 -3135
rect 18510 -3430 18630 -3310
rect 18685 -3430 18805 -3310
rect 18850 -3430 18970 -3310
rect 19015 -3430 19135 -3310
rect 19180 -3430 19300 -3310
rect 19355 -3430 19475 -3310
rect 19520 -3430 19640 -3310
rect 19685 -3430 19805 -3310
rect 19850 -3430 19970 -3310
rect 20025 -3430 20145 -3310
rect 20190 -3430 20310 -3310
rect 20355 -3430 20475 -3310
rect 20520 -3430 20640 -3310
rect 20695 -3430 20815 -3310
rect 20860 -3430 20980 -3310
rect 21025 -3430 21145 -3310
rect 21190 -3430 21310 -3310
rect 21365 -3430 21485 -3310
rect 21530 -3430 21650 -3310
rect 21695 -3430 21815 -3310
rect 21860 -3430 21980 -3310
rect 22035 -3430 22155 -3310
rect 22200 -3430 22320 -3310
rect 22365 -3430 22485 -3310
rect 22530 -3430 22650 -3310
rect 22705 -3430 22825 -3310
rect 22870 -3430 22990 -3310
rect 23035 -3430 23155 -3310
rect 23200 -3430 23320 -3310
rect 23375 -3430 23495 -3310
rect 23540 -3430 23660 -3310
rect 23705 -3430 23825 -3310
rect 23870 -3430 23990 -3310
rect 18510 -3595 18630 -3475
rect 18685 -3595 18805 -3475
rect 18850 -3595 18970 -3475
rect 19015 -3595 19135 -3475
rect 19180 -3595 19300 -3475
rect 19355 -3595 19475 -3475
rect 19520 -3595 19640 -3475
rect 19685 -3595 19805 -3475
rect 19850 -3595 19970 -3475
rect 20025 -3595 20145 -3475
rect 20190 -3595 20310 -3475
rect 20355 -3595 20475 -3475
rect 20520 -3595 20640 -3475
rect 20695 -3595 20815 -3475
rect 20860 -3595 20980 -3475
rect 21025 -3595 21145 -3475
rect 21190 -3595 21310 -3475
rect 21365 -3595 21485 -3475
rect 21530 -3595 21650 -3475
rect 21695 -3595 21815 -3475
rect 21860 -3595 21980 -3475
rect 22035 -3595 22155 -3475
rect 22200 -3595 22320 -3475
rect 22365 -3595 22485 -3475
rect 22530 -3595 22650 -3475
rect 22705 -3595 22825 -3475
rect 22870 -3595 22990 -3475
rect 23035 -3595 23155 -3475
rect 23200 -3595 23320 -3475
rect 23375 -3595 23495 -3475
rect 23540 -3595 23660 -3475
rect 23705 -3595 23825 -3475
rect 23870 -3595 23990 -3475
rect 18510 -3760 18630 -3640
rect 18685 -3760 18805 -3640
rect 18850 -3760 18970 -3640
rect 19015 -3760 19135 -3640
rect 19180 -3760 19300 -3640
rect 19355 -3760 19475 -3640
rect 19520 -3760 19640 -3640
rect 19685 -3760 19805 -3640
rect 19850 -3760 19970 -3640
rect 20025 -3760 20145 -3640
rect 20190 -3760 20310 -3640
rect 20355 -3760 20475 -3640
rect 20520 -3760 20640 -3640
rect 20695 -3760 20815 -3640
rect 20860 -3760 20980 -3640
rect 21025 -3760 21145 -3640
rect 21190 -3760 21310 -3640
rect 21365 -3760 21485 -3640
rect 21530 -3760 21650 -3640
rect 21695 -3760 21815 -3640
rect 21860 -3760 21980 -3640
rect 22035 -3760 22155 -3640
rect 22200 -3760 22320 -3640
rect 22365 -3760 22485 -3640
rect 22530 -3760 22650 -3640
rect 22705 -3760 22825 -3640
rect 22870 -3760 22990 -3640
rect 23035 -3760 23155 -3640
rect 23200 -3760 23320 -3640
rect 23375 -3760 23495 -3640
rect 23540 -3760 23660 -3640
rect 23705 -3760 23825 -3640
rect 23870 -3760 23990 -3640
rect 18510 -3925 18630 -3805
rect 18685 -3925 18805 -3805
rect 18850 -3925 18970 -3805
rect 19015 -3925 19135 -3805
rect 19180 -3925 19300 -3805
rect 19355 -3925 19475 -3805
rect 19520 -3925 19640 -3805
rect 19685 -3925 19805 -3805
rect 19850 -3925 19970 -3805
rect 20025 -3925 20145 -3805
rect 20190 -3925 20310 -3805
rect 20355 -3925 20475 -3805
rect 20520 -3925 20640 -3805
rect 20695 -3925 20815 -3805
rect 20860 -3925 20980 -3805
rect 21025 -3925 21145 -3805
rect 21190 -3925 21310 -3805
rect 21365 -3925 21485 -3805
rect 21530 -3925 21650 -3805
rect 21695 -3925 21815 -3805
rect 21860 -3925 21980 -3805
rect 22035 -3925 22155 -3805
rect 22200 -3925 22320 -3805
rect 22365 -3925 22485 -3805
rect 22530 -3925 22650 -3805
rect 22705 -3925 22825 -3805
rect 22870 -3925 22990 -3805
rect 23035 -3925 23155 -3805
rect 23200 -3925 23320 -3805
rect 23375 -3925 23495 -3805
rect 23540 -3925 23660 -3805
rect 23705 -3925 23825 -3805
rect 23870 -3925 23990 -3805
rect 18510 -4100 18630 -3980
rect 18685 -4100 18805 -3980
rect 18850 -4100 18970 -3980
rect 19015 -4100 19135 -3980
rect 19180 -4100 19300 -3980
rect 19355 -4100 19475 -3980
rect 19520 -4100 19640 -3980
rect 19685 -4100 19805 -3980
rect 19850 -4100 19970 -3980
rect 20025 -4100 20145 -3980
rect 20190 -4100 20310 -3980
rect 20355 -4100 20475 -3980
rect 20520 -4100 20640 -3980
rect 20695 -4100 20815 -3980
rect 20860 -4100 20980 -3980
rect 21025 -4100 21145 -3980
rect 21190 -4100 21310 -3980
rect 21365 -4100 21485 -3980
rect 21530 -4100 21650 -3980
rect 21695 -4100 21815 -3980
rect 21860 -4100 21980 -3980
rect 22035 -4100 22155 -3980
rect 22200 -4100 22320 -3980
rect 22365 -4100 22485 -3980
rect 22530 -4100 22650 -3980
rect 22705 -4100 22825 -3980
rect 22870 -4100 22990 -3980
rect 23035 -4100 23155 -3980
rect 23200 -4100 23320 -3980
rect 23375 -4100 23495 -3980
rect 23540 -4100 23660 -3980
rect 23705 -4100 23825 -3980
rect 23870 -4100 23990 -3980
rect 24200 1260 24320 1380
rect 24375 1260 24495 1380
rect 24540 1260 24660 1380
rect 24705 1260 24825 1380
rect 24870 1260 24990 1380
rect 25045 1260 25165 1380
rect 25210 1260 25330 1380
rect 25375 1260 25495 1380
rect 25540 1260 25660 1380
rect 25715 1260 25835 1380
rect 25880 1260 26000 1380
rect 26045 1260 26165 1380
rect 26210 1260 26330 1380
rect 26385 1260 26505 1380
rect 26550 1260 26670 1380
rect 26715 1260 26835 1380
rect 26880 1260 27000 1380
rect 27055 1260 27175 1380
rect 27220 1260 27340 1380
rect 27385 1260 27505 1380
rect 27550 1260 27670 1380
rect 27725 1260 27845 1380
rect 27890 1260 28010 1380
rect 28055 1260 28175 1380
rect 28220 1260 28340 1380
rect 28395 1260 28515 1380
rect 28560 1260 28680 1380
rect 28725 1260 28845 1380
rect 28890 1260 29010 1380
rect 29065 1260 29185 1380
rect 29230 1260 29350 1380
rect 29395 1260 29515 1380
rect 29560 1260 29680 1380
rect 24200 1095 24320 1215
rect 24375 1095 24495 1215
rect 24540 1095 24660 1215
rect 24705 1095 24825 1215
rect 24870 1095 24990 1215
rect 25045 1095 25165 1215
rect 25210 1095 25330 1215
rect 25375 1095 25495 1215
rect 25540 1095 25660 1215
rect 25715 1095 25835 1215
rect 25880 1095 26000 1215
rect 26045 1095 26165 1215
rect 26210 1095 26330 1215
rect 26385 1095 26505 1215
rect 26550 1095 26670 1215
rect 26715 1095 26835 1215
rect 26880 1095 27000 1215
rect 27055 1095 27175 1215
rect 27220 1095 27340 1215
rect 27385 1095 27505 1215
rect 27550 1095 27670 1215
rect 27725 1095 27845 1215
rect 27890 1095 28010 1215
rect 28055 1095 28175 1215
rect 28220 1095 28340 1215
rect 28395 1095 28515 1215
rect 28560 1095 28680 1215
rect 28725 1095 28845 1215
rect 28890 1095 29010 1215
rect 29065 1095 29185 1215
rect 29230 1095 29350 1215
rect 29395 1095 29515 1215
rect 29560 1095 29680 1215
rect 24200 930 24320 1050
rect 24375 930 24495 1050
rect 24540 930 24660 1050
rect 24705 930 24825 1050
rect 24870 930 24990 1050
rect 25045 930 25165 1050
rect 25210 930 25330 1050
rect 25375 930 25495 1050
rect 25540 930 25660 1050
rect 25715 930 25835 1050
rect 25880 930 26000 1050
rect 26045 930 26165 1050
rect 26210 930 26330 1050
rect 26385 930 26505 1050
rect 26550 930 26670 1050
rect 26715 930 26835 1050
rect 26880 930 27000 1050
rect 27055 930 27175 1050
rect 27220 930 27340 1050
rect 27385 930 27505 1050
rect 27550 930 27670 1050
rect 27725 930 27845 1050
rect 27890 930 28010 1050
rect 28055 930 28175 1050
rect 28220 930 28340 1050
rect 28395 930 28515 1050
rect 28560 930 28680 1050
rect 28725 930 28845 1050
rect 28890 930 29010 1050
rect 29065 930 29185 1050
rect 29230 930 29350 1050
rect 29395 930 29515 1050
rect 29560 930 29680 1050
rect 24200 765 24320 885
rect 24375 765 24495 885
rect 24540 765 24660 885
rect 24705 765 24825 885
rect 24870 765 24990 885
rect 25045 765 25165 885
rect 25210 765 25330 885
rect 25375 765 25495 885
rect 25540 765 25660 885
rect 25715 765 25835 885
rect 25880 765 26000 885
rect 26045 765 26165 885
rect 26210 765 26330 885
rect 26385 765 26505 885
rect 26550 765 26670 885
rect 26715 765 26835 885
rect 26880 765 27000 885
rect 27055 765 27175 885
rect 27220 765 27340 885
rect 27385 765 27505 885
rect 27550 765 27670 885
rect 27725 765 27845 885
rect 27890 765 28010 885
rect 28055 765 28175 885
rect 28220 765 28340 885
rect 28395 765 28515 885
rect 28560 765 28680 885
rect 28725 765 28845 885
rect 28890 765 29010 885
rect 29065 765 29185 885
rect 29230 765 29350 885
rect 29395 765 29515 885
rect 29560 765 29680 885
rect 24200 590 24320 710
rect 24375 590 24495 710
rect 24540 590 24660 710
rect 24705 590 24825 710
rect 24870 590 24990 710
rect 25045 590 25165 710
rect 25210 590 25330 710
rect 25375 590 25495 710
rect 25540 590 25660 710
rect 25715 590 25835 710
rect 25880 590 26000 710
rect 26045 590 26165 710
rect 26210 590 26330 710
rect 26385 590 26505 710
rect 26550 590 26670 710
rect 26715 590 26835 710
rect 26880 590 27000 710
rect 27055 590 27175 710
rect 27220 590 27340 710
rect 27385 590 27505 710
rect 27550 590 27670 710
rect 27725 590 27845 710
rect 27890 590 28010 710
rect 28055 590 28175 710
rect 28220 590 28340 710
rect 28395 590 28515 710
rect 28560 590 28680 710
rect 28725 590 28845 710
rect 28890 590 29010 710
rect 29065 590 29185 710
rect 29230 590 29350 710
rect 29395 590 29515 710
rect 29560 590 29680 710
rect 24200 425 24320 545
rect 24375 425 24495 545
rect 24540 425 24660 545
rect 24705 425 24825 545
rect 24870 425 24990 545
rect 25045 425 25165 545
rect 25210 425 25330 545
rect 25375 425 25495 545
rect 25540 425 25660 545
rect 25715 425 25835 545
rect 25880 425 26000 545
rect 26045 425 26165 545
rect 26210 425 26330 545
rect 26385 425 26505 545
rect 26550 425 26670 545
rect 26715 425 26835 545
rect 26880 425 27000 545
rect 27055 425 27175 545
rect 27220 425 27340 545
rect 27385 425 27505 545
rect 27550 425 27670 545
rect 27725 425 27845 545
rect 27890 425 28010 545
rect 28055 425 28175 545
rect 28220 425 28340 545
rect 28395 425 28515 545
rect 28560 425 28680 545
rect 28725 425 28845 545
rect 28890 425 29010 545
rect 29065 425 29185 545
rect 29230 425 29350 545
rect 29395 425 29515 545
rect 29560 425 29680 545
rect 24200 260 24320 380
rect 24375 260 24495 380
rect 24540 260 24660 380
rect 24705 260 24825 380
rect 24870 260 24990 380
rect 25045 260 25165 380
rect 25210 260 25330 380
rect 25375 260 25495 380
rect 25540 260 25660 380
rect 25715 260 25835 380
rect 25880 260 26000 380
rect 26045 260 26165 380
rect 26210 260 26330 380
rect 26385 260 26505 380
rect 26550 260 26670 380
rect 26715 260 26835 380
rect 26880 260 27000 380
rect 27055 260 27175 380
rect 27220 260 27340 380
rect 27385 260 27505 380
rect 27550 260 27670 380
rect 27725 260 27845 380
rect 27890 260 28010 380
rect 28055 260 28175 380
rect 28220 260 28340 380
rect 28395 260 28515 380
rect 28560 260 28680 380
rect 28725 260 28845 380
rect 28890 260 29010 380
rect 29065 260 29185 380
rect 29230 260 29350 380
rect 29395 260 29515 380
rect 29560 260 29680 380
rect 24200 95 24320 215
rect 24375 95 24495 215
rect 24540 95 24660 215
rect 24705 95 24825 215
rect 24870 95 24990 215
rect 25045 95 25165 215
rect 25210 95 25330 215
rect 25375 95 25495 215
rect 25540 95 25660 215
rect 25715 95 25835 215
rect 25880 95 26000 215
rect 26045 95 26165 215
rect 26210 95 26330 215
rect 26385 95 26505 215
rect 26550 95 26670 215
rect 26715 95 26835 215
rect 26880 95 27000 215
rect 27055 95 27175 215
rect 27220 95 27340 215
rect 27385 95 27505 215
rect 27550 95 27670 215
rect 27725 95 27845 215
rect 27890 95 28010 215
rect 28055 95 28175 215
rect 28220 95 28340 215
rect 28395 95 28515 215
rect 28560 95 28680 215
rect 28725 95 28845 215
rect 28890 95 29010 215
rect 29065 95 29185 215
rect 29230 95 29350 215
rect 29395 95 29515 215
rect 29560 95 29680 215
rect 24200 -80 24320 40
rect 24375 -80 24495 40
rect 24540 -80 24660 40
rect 24705 -80 24825 40
rect 24870 -80 24990 40
rect 25045 -80 25165 40
rect 25210 -80 25330 40
rect 25375 -80 25495 40
rect 25540 -80 25660 40
rect 25715 -80 25835 40
rect 25880 -80 26000 40
rect 26045 -80 26165 40
rect 26210 -80 26330 40
rect 26385 -80 26505 40
rect 26550 -80 26670 40
rect 26715 -80 26835 40
rect 26880 -80 27000 40
rect 27055 -80 27175 40
rect 27220 -80 27340 40
rect 27385 -80 27505 40
rect 27550 -80 27670 40
rect 27725 -80 27845 40
rect 27890 -80 28010 40
rect 28055 -80 28175 40
rect 28220 -80 28340 40
rect 28395 -80 28515 40
rect 28560 -80 28680 40
rect 28725 -80 28845 40
rect 28890 -80 29010 40
rect 29065 -80 29185 40
rect 29230 -80 29350 40
rect 29395 -80 29515 40
rect 29560 -80 29680 40
rect 24200 -245 24320 -125
rect 24375 -245 24495 -125
rect 24540 -245 24660 -125
rect 24705 -245 24825 -125
rect 24870 -245 24990 -125
rect 25045 -245 25165 -125
rect 25210 -245 25330 -125
rect 25375 -245 25495 -125
rect 25540 -245 25660 -125
rect 25715 -245 25835 -125
rect 25880 -245 26000 -125
rect 26045 -245 26165 -125
rect 26210 -245 26330 -125
rect 26385 -245 26505 -125
rect 26550 -245 26670 -125
rect 26715 -245 26835 -125
rect 26880 -245 27000 -125
rect 27055 -245 27175 -125
rect 27220 -245 27340 -125
rect 27385 -245 27505 -125
rect 27550 -245 27670 -125
rect 27725 -245 27845 -125
rect 27890 -245 28010 -125
rect 28055 -245 28175 -125
rect 28220 -245 28340 -125
rect 28395 -245 28515 -125
rect 28560 -245 28680 -125
rect 28725 -245 28845 -125
rect 28890 -245 29010 -125
rect 29065 -245 29185 -125
rect 29230 -245 29350 -125
rect 29395 -245 29515 -125
rect 29560 -245 29680 -125
rect 24200 -410 24320 -290
rect 24375 -410 24495 -290
rect 24540 -410 24660 -290
rect 24705 -410 24825 -290
rect 24870 -410 24990 -290
rect 25045 -410 25165 -290
rect 25210 -410 25330 -290
rect 25375 -410 25495 -290
rect 25540 -410 25660 -290
rect 25715 -410 25835 -290
rect 25880 -410 26000 -290
rect 26045 -410 26165 -290
rect 26210 -410 26330 -290
rect 26385 -410 26505 -290
rect 26550 -410 26670 -290
rect 26715 -410 26835 -290
rect 26880 -410 27000 -290
rect 27055 -410 27175 -290
rect 27220 -410 27340 -290
rect 27385 -410 27505 -290
rect 27550 -410 27670 -290
rect 27725 -410 27845 -290
rect 27890 -410 28010 -290
rect 28055 -410 28175 -290
rect 28220 -410 28340 -290
rect 28395 -410 28515 -290
rect 28560 -410 28680 -290
rect 28725 -410 28845 -290
rect 28890 -410 29010 -290
rect 29065 -410 29185 -290
rect 29230 -410 29350 -290
rect 29395 -410 29515 -290
rect 29560 -410 29680 -290
rect 24200 -575 24320 -455
rect 24375 -575 24495 -455
rect 24540 -575 24660 -455
rect 24705 -575 24825 -455
rect 24870 -575 24990 -455
rect 25045 -575 25165 -455
rect 25210 -575 25330 -455
rect 25375 -575 25495 -455
rect 25540 -575 25660 -455
rect 25715 -575 25835 -455
rect 25880 -575 26000 -455
rect 26045 -575 26165 -455
rect 26210 -575 26330 -455
rect 26385 -575 26505 -455
rect 26550 -575 26670 -455
rect 26715 -575 26835 -455
rect 26880 -575 27000 -455
rect 27055 -575 27175 -455
rect 27220 -575 27340 -455
rect 27385 -575 27505 -455
rect 27550 -575 27670 -455
rect 27725 -575 27845 -455
rect 27890 -575 28010 -455
rect 28055 -575 28175 -455
rect 28220 -575 28340 -455
rect 28395 -575 28515 -455
rect 28560 -575 28680 -455
rect 28725 -575 28845 -455
rect 28890 -575 29010 -455
rect 29065 -575 29185 -455
rect 29230 -575 29350 -455
rect 29395 -575 29515 -455
rect 29560 -575 29680 -455
rect 24200 -750 24320 -630
rect 24375 -750 24495 -630
rect 24540 -750 24660 -630
rect 24705 -750 24825 -630
rect 24870 -750 24990 -630
rect 25045 -750 25165 -630
rect 25210 -750 25330 -630
rect 25375 -750 25495 -630
rect 25540 -750 25660 -630
rect 25715 -750 25835 -630
rect 25880 -750 26000 -630
rect 26045 -750 26165 -630
rect 26210 -750 26330 -630
rect 26385 -750 26505 -630
rect 26550 -750 26670 -630
rect 26715 -750 26835 -630
rect 26880 -750 27000 -630
rect 27055 -750 27175 -630
rect 27220 -750 27340 -630
rect 27385 -750 27505 -630
rect 27550 -750 27670 -630
rect 27725 -750 27845 -630
rect 27890 -750 28010 -630
rect 28055 -750 28175 -630
rect 28220 -750 28340 -630
rect 28395 -750 28515 -630
rect 28560 -750 28680 -630
rect 28725 -750 28845 -630
rect 28890 -750 29010 -630
rect 29065 -750 29185 -630
rect 29230 -750 29350 -630
rect 29395 -750 29515 -630
rect 29560 -750 29680 -630
rect 24200 -915 24320 -795
rect 24375 -915 24495 -795
rect 24540 -915 24660 -795
rect 24705 -915 24825 -795
rect 24870 -915 24990 -795
rect 25045 -915 25165 -795
rect 25210 -915 25330 -795
rect 25375 -915 25495 -795
rect 25540 -915 25660 -795
rect 25715 -915 25835 -795
rect 25880 -915 26000 -795
rect 26045 -915 26165 -795
rect 26210 -915 26330 -795
rect 26385 -915 26505 -795
rect 26550 -915 26670 -795
rect 26715 -915 26835 -795
rect 26880 -915 27000 -795
rect 27055 -915 27175 -795
rect 27220 -915 27340 -795
rect 27385 -915 27505 -795
rect 27550 -915 27670 -795
rect 27725 -915 27845 -795
rect 27890 -915 28010 -795
rect 28055 -915 28175 -795
rect 28220 -915 28340 -795
rect 28395 -915 28515 -795
rect 28560 -915 28680 -795
rect 28725 -915 28845 -795
rect 28890 -915 29010 -795
rect 29065 -915 29185 -795
rect 29230 -915 29350 -795
rect 29395 -915 29515 -795
rect 29560 -915 29680 -795
rect 24200 -1080 24320 -960
rect 24375 -1080 24495 -960
rect 24540 -1080 24660 -960
rect 24705 -1080 24825 -960
rect 24870 -1080 24990 -960
rect 25045 -1080 25165 -960
rect 25210 -1080 25330 -960
rect 25375 -1080 25495 -960
rect 25540 -1080 25660 -960
rect 25715 -1080 25835 -960
rect 25880 -1080 26000 -960
rect 26045 -1080 26165 -960
rect 26210 -1080 26330 -960
rect 26385 -1080 26505 -960
rect 26550 -1080 26670 -960
rect 26715 -1080 26835 -960
rect 26880 -1080 27000 -960
rect 27055 -1080 27175 -960
rect 27220 -1080 27340 -960
rect 27385 -1080 27505 -960
rect 27550 -1080 27670 -960
rect 27725 -1080 27845 -960
rect 27890 -1080 28010 -960
rect 28055 -1080 28175 -960
rect 28220 -1080 28340 -960
rect 28395 -1080 28515 -960
rect 28560 -1080 28680 -960
rect 28725 -1080 28845 -960
rect 28890 -1080 29010 -960
rect 29065 -1080 29185 -960
rect 29230 -1080 29350 -960
rect 29395 -1080 29515 -960
rect 29560 -1080 29680 -960
rect 24200 -1245 24320 -1125
rect 24375 -1245 24495 -1125
rect 24540 -1245 24660 -1125
rect 24705 -1245 24825 -1125
rect 24870 -1245 24990 -1125
rect 25045 -1245 25165 -1125
rect 25210 -1245 25330 -1125
rect 25375 -1245 25495 -1125
rect 25540 -1245 25660 -1125
rect 25715 -1245 25835 -1125
rect 25880 -1245 26000 -1125
rect 26045 -1245 26165 -1125
rect 26210 -1245 26330 -1125
rect 26385 -1245 26505 -1125
rect 26550 -1245 26670 -1125
rect 26715 -1245 26835 -1125
rect 26880 -1245 27000 -1125
rect 27055 -1245 27175 -1125
rect 27220 -1245 27340 -1125
rect 27385 -1245 27505 -1125
rect 27550 -1245 27670 -1125
rect 27725 -1245 27845 -1125
rect 27890 -1245 28010 -1125
rect 28055 -1245 28175 -1125
rect 28220 -1245 28340 -1125
rect 28395 -1245 28515 -1125
rect 28560 -1245 28680 -1125
rect 28725 -1245 28845 -1125
rect 28890 -1245 29010 -1125
rect 29065 -1245 29185 -1125
rect 29230 -1245 29350 -1125
rect 29395 -1245 29515 -1125
rect 29560 -1245 29680 -1125
rect 24200 -1420 24320 -1300
rect 24375 -1420 24495 -1300
rect 24540 -1420 24660 -1300
rect 24705 -1420 24825 -1300
rect 24870 -1420 24990 -1300
rect 25045 -1420 25165 -1300
rect 25210 -1420 25330 -1300
rect 25375 -1420 25495 -1300
rect 25540 -1420 25660 -1300
rect 25715 -1420 25835 -1300
rect 25880 -1420 26000 -1300
rect 26045 -1420 26165 -1300
rect 26210 -1420 26330 -1300
rect 26385 -1420 26505 -1300
rect 26550 -1420 26670 -1300
rect 26715 -1420 26835 -1300
rect 26880 -1420 27000 -1300
rect 27055 -1420 27175 -1300
rect 27220 -1420 27340 -1300
rect 27385 -1420 27505 -1300
rect 27550 -1420 27670 -1300
rect 27725 -1420 27845 -1300
rect 27890 -1420 28010 -1300
rect 28055 -1420 28175 -1300
rect 28220 -1420 28340 -1300
rect 28395 -1420 28515 -1300
rect 28560 -1420 28680 -1300
rect 28725 -1420 28845 -1300
rect 28890 -1420 29010 -1300
rect 29065 -1420 29185 -1300
rect 29230 -1420 29350 -1300
rect 29395 -1420 29515 -1300
rect 29560 -1420 29680 -1300
rect 24200 -1585 24320 -1465
rect 24375 -1585 24495 -1465
rect 24540 -1585 24660 -1465
rect 24705 -1585 24825 -1465
rect 24870 -1585 24990 -1465
rect 25045 -1585 25165 -1465
rect 25210 -1585 25330 -1465
rect 25375 -1585 25495 -1465
rect 25540 -1585 25660 -1465
rect 25715 -1585 25835 -1465
rect 25880 -1585 26000 -1465
rect 26045 -1585 26165 -1465
rect 26210 -1585 26330 -1465
rect 26385 -1585 26505 -1465
rect 26550 -1585 26670 -1465
rect 26715 -1585 26835 -1465
rect 26880 -1585 27000 -1465
rect 27055 -1585 27175 -1465
rect 27220 -1585 27340 -1465
rect 27385 -1585 27505 -1465
rect 27550 -1585 27670 -1465
rect 27725 -1585 27845 -1465
rect 27890 -1585 28010 -1465
rect 28055 -1585 28175 -1465
rect 28220 -1585 28340 -1465
rect 28395 -1585 28515 -1465
rect 28560 -1585 28680 -1465
rect 28725 -1585 28845 -1465
rect 28890 -1585 29010 -1465
rect 29065 -1585 29185 -1465
rect 29230 -1585 29350 -1465
rect 29395 -1585 29515 -1465
rect 29560 -1585 29680 -1465
rect 24200 -1750 24320 -1630
rect 24375 -1750 24495 -1630
rect 24540 -1750 24660 -1630
rect 24705 -1750 24825 -1630
rect 24870 -1750 24990 -1630
rect 25045 -1750 25165 -1630
rect 25210 -1750 25330 -1630
rect 25375 -1750 25495 -1630
rect 25540 -1750 25660 -1630
rect 25715 -1750 25835 -1630
rect 25880 -1750 26000 -1630
rect 26045 -1750 26165 -1630
rect 26210 -1750 26330 -1630
rect 26385 -1750 26505 -1630
rect 26550 -1750 26670 -1630
rect 26715 -1750 26835 -1630
rect 26880 -1750 27000 -1630
rect 27055 -1750 27175 -1630
rect 27220 -1750 27340 -1630
rect 27385 -1750 27505 -1630
rect 27550 -1750 27670 -1630
rect 27725 -1750 27845 -1630
rect 27890 -1750 28010 -1630
rect 28055 -1750 28175 -1630
rect 28220 -1750 28340 -1630
rect 28395 -1750 28515 -1630
rect 28560 -1750 28680 -1630
rect 28725 -1750 28845 -1630
rect 28890 -1750 29010 -1630
rect 29065 -1750 29185 -1630
rect 29230 -1750 29350 -1630
rect 29395 -1750 29515 -1630
rect 29560 -1750 29680 -1630
rect 24200 -1915 24320 -1795
rect 24375 -1915 24495 -1795
rect 24540 -1915 24660 -1795
rect 24705 -1915 24825 -1795
rect 24870 -1915 24990 -1795
rect 25045 -1915 25165 -1795
rect 25210 -1915 25330 -1795
rect 25375 -1915 25495 -1795
rect 25540 -1915 25660 -1795
rect 25715 -1915 25835 -1795
rect 25880 -1915 26000 -1795
rect 26045 -1915 26165 -1795
rect 26210 -1915 26330 -1795
rect 26385 -1915 26505 -1795
rect 26550 -1915 26670 -1795
rect 26715 -1915 26835 -1795
rect 26880 -1915 27000 -1795
rect 27055 -1915 27175 -1795
rect 27220 -1915 27340 -1795
rect 27385 -1915 27505 -1795
rect 27550 -1915 27670 -1795
rect 27725 -1915 27845 -1795
rect 27890 -1915 28010 -1795
rect 28055 -1915 28175 -1795
rect 28220 -1915 28340 -1795
rect 28395 -1915 28515 -1795
rect 28560 -1915 28680 -1795
rect 28725 -1915 28845 -1795
rect 28890 -1915 29010 -1795
rect 29065 -1915 29185 -1795
rect 29230 -1915 29350 -1795
rect 29395 -1915 29515 -1795
rect 29560 -1915 29680 -1795
rect 24200 -2090 24320 -1970
rect 24375 -2090 24495 -1970
rect 24540 -2090 24660 -1970
rect 24705 -2090 24825 -1970
rect 24870 -2090 24990 -1970
rect 25045 -2090 25165 -1970
rect 25210 -2090 25330 -1970
rect 25375 -2090 25495 -1970
rect 25540 -2090 25660 -1970
rect 25715 -2090 25835 -1970
rect 25880 -2090 26000 -1970
rect 26045 -2090 26165 -1970
rect 26210 -2090 26330 -1970
rect 26385 -2090 26505 -1970
rect 26550 -2090 26670 -1970
rect 26715 -2090 26835 -1970
rect 26880 -2090 27000 -1970
rect 27055 -2090 27175 -1970
rect 27220 -2090 27340 -1970
rect 27385 -2090 27505 -1970
rect 27550 -2090 27670 -1970
rect 27725 -2090 27845 -1970
rect 27890 -2090 28010 -1970
rect 28055 -2090 28175 -1970
rect 28220 -2090 28340 -1970
rect 28395 -2090 28515 -1970
rect 28560 -2090 28680 -1970
rect 28725 -2090 28845 -1970
rect 28890 -2090 29010 -1970
rect 29065 -2090 29185 -1970
rect 29230 -2090 29350 -1970
rect 29395 -2090 29515 -1970
rect 29560 -2090 29680 -1970
rect 24200 -2255 24320 -2135
rect 24375 -2255 24495 -2135
rect 24540 -2255 24660 -2135
rect 24705 -2255 24825 -2135
rect 24870 -2255 24990 -2135
rect 25045 -2255 25165 -2135
rect 25210 -2255 25330 -2135
rect 25375 -2255 25495 -2135
rect 25540 -2255 25660 -2135
rect 25715 -2255 25835 -2135
rect 25880 -2255 26000 -2135
rect 26045 -2255 26165 -2135
rect 26210 -2255 26330 -2135
rect 26385 -2255 26505 -2135
rect 26550 -2255 26670 -2135
rect 26715 -2255 26835 -2135
rect 26880 -2255 27000 -2135
rect 27055 -2255 27175 -2135
rect 27220 -2255 27340 -2135
rect 27385 -2255 27505 -2135
rect 27550 -2255 27670 -2135
rect 27725 -2255 27845 -2135
rect 27890 -2255 28010 -2135
rect 28055 -2255 28175 -2135
rect 28220 -2255 28340 -2135
rect 28395 -2255 28515 -2135
rect 28560 -2255 28680 -2135
rect 28725 -2255 28845 -2135
rect 28890 -2255 29010 -2135
rect 29065 -2255 29185 -2135
rect 29230 -2255 29350 -2135
rect 29395 -2255 29515 -2135
rect 29560 -2255 29680 -2135
rect 24200 -2420 24320 -2300
rect 24375 -2420 24495 -2300
rect 24540 -2420 24660 -2300
rect 24705 -2420 24825 -2300
rect 24870 -2420 24990 -2300
rect 25045 -2420 25165 -2300
rect 25210 -2420 25330 -2300
rect 25375 -2420 25495 -2300
rect 25540 -2420 25660 -2300
rect 25715 -2420 25835 -2300
rect 25880 -2420 26000 -2300
rect 26045 -2420 26165 -2300
rect 26210 -2420 26330 -2300
rect 26385 -2420 26505 -2300
rect 26550 -2420 26670 -2300
rect 26715 -2420 26835 -2300
rect 26880 -2420 27000 -2300
rect 27055 -2420 27175 -2300
rect 27220 -2420 27340 -2300
rect 27385 -2420 27505 -2300
rect 27550 -2420 27670 -2300
rect 27725 -2420 27845 -2300
rect 27890 -2420 28010 -2300
rect 28055 -2420 28175 -2300
rect 28220 -2420 28340 -2300
rect 28395 -2420 28515 -2300
rect 28560 -2420 28680 -2300
rect 28725 -2420 28845 -2300
rect 28890 -2420 29010 -2300
rect 29065 -2420 29185 -2300
rect 29230 -2420 29350 -2300
rect 29395 -2420 29515 -2300
rect 29560 -2420 29680 -2300
rect 24200 -2585 24320 -2465
rect 24375 -2585 24495 -2465
rect 24540 -2585 24660 -2465
rect 24705 -2585 24825 -2465
rect 24870 -2585 24990 -2465
rect 25045 -2585 25165 -2465
rect 25210 -2585 25330 -2465
rect 25375 -2585 25495 -2465
rect 25540 -2585 25660 -2465
rect 25715 -2585 25835 -2465
rect 25880 -2585 26000 -2465
rect 26045 -2585 26165 -2465
rect 26210 -2585 26330 -2465
rect 26385 -2585 26505 -2465
rect 26550 -2585 26670 -2465
rect 26715 -2585 26835 -2465
rect 26880 -2585 27000 -2465
rect 27055 -2585 27175 -2465
rect 27220 -2585 27340 -2465
rect 27385 -2585 27505 -2465
rect 27550 -2585 27670 -2465
rect 27725 -2585 27845 -2465
rect 27890 -2585 28010 -2465
rect 28055 -2585 28175 -2465
rect 28220 -2585 28340 -2465
rect 28395 -2585 28515 -2465
rect 28560 -2585 28680 -2465
rect 28725 -2585 28845 -2465
rect 28890 -2585 29010 -2465
rect 29065 -2585 29185 -2465
rect 29230 -2585 29350 -2465
rect 29395 -2585 29515 -2465
rect 29560 -2585 29680 -2465
rect 24200 -2760 24320 -2640
rect 24375 -2760 24495 -2640
rect 24540 -2760 24660 -2640
rect 24705 -2760 24825 -2640
rect 24870 -2760 24990 -2640
rect 25045 -2760 25165 -2640
rect 25210 -2760 25330 -2640
rect 25375 -2760 25495 -2640
rect 25540 -2760 25660 -2640
rect 25715 -2760 25835 -2640
rect 25880 -2760 26000 -2640
rect 26045 -2760 26165 -2640
rect 26210 -2760 26330 -2640
rect 26385 -2760 26505 -2640
rect 26550 -2760 26670 -2640
rect 26715 -2760 26835 -2640
rect 26880 -2760 27000 -2640
rect 27055 -2760 27175 -2640
rect 27220 -2760 27340 -2640
rect 27385 -2760 27505 -2640
rect 27550 -2760 27670 -2640
rect 27725 -2760 27845 -2640
rect 27890 -2760 28010 -2640
rect 28055 -2760 28175 -2640
rect 28220 -2760 28340 -2640
rect 28395 -2760 28515 -2640
rect 28560 -2760 28680 -2640
rect 28725 -2760 28845 -2640
rect 28890 -2760 29010 -2640
rect 29065 -2760 29185 -2640
rect 29230 -2760 29350 -2640
rect 29395 -2760 29515 -2640
rect 29560 -2760 29680 -2640
rect 24200 -2925 24320 -2805
rect 24375 -2925 24495 -2805
rect 24540 -2925 24660 -2805
rect 24705 -2925 24825 -2805
rect 24870 -2925 24990 -2805
rect 25045 -2925 25165 -2805
rect 25210 -2925 25330 -2805
rect 25375 -2925 25495 -2805
rect 25540 -2925 25660 -2805
rect 25715 -2925 25835 -2805
rect 25880 -2925 26000 -2805
rect 26045 -2925 26165 -2805
rect 26210 -2925 26330 -2805
rect 26385 -2925 26505 -2805
rect 26550 -2925 26670 -2805
rect 26715 -2925 26835 -2805
rect 26880 -2925 27000 -2805
rect 27055 -2925 27175 -2805
rect 27220 -2925 27340 -2805
rect 27385 -2925 27505 -2805
rect 27550 -2925 27670 -2805
rect 27725 -2925 27845 -2805
rect 27890 -2925 28010 -2805
rect 28055 -2925 28175 -2805
rect 28220 -2925 28340 -2805
rect 28395 -2925 28515 -2805
rect 28560 -2925 28680 -2805
rect 28725 -2925 28845 -2805
rect 28890 -2925 29010 -2805
rect 29065 -2925 29185 -2805
rect 29230 -2925 29350 -2805
rect 29395 -2925 29515 -2805
rect 29560 -2925 29680 -2805
rect 24200 -3090 24320 -2970
rect 24375 -3090 24495 -2970
rect 24540 -3090 24660 -2970
rect 24705 -3090 24825 -2970
rect 24870 -3090 24990 -2970
rect 25045 -3090 25165 -2970
rect 25210 -3090 25330 -2970
rect 25375 -3090 25495 -2970
rect 25540 -3090 25660 -2970
rect 25715 -3090 25835 -2970
rect 25880 -3090 26000 -2970
rect 26045 -3090 26165 -2970
rect 26210 -3090 26330 -2970
rect 26385 -3090 26505 -2970
rect 26550 -3090 26670 -2970
rect 26715 -3090 26835 -2970
rect 26880 -3090 27000 -2970
rect 27055 -3090 27175 -2970
rect 27220 -3090 27340 -2970
rect 27385 -3090 27505 -2970
rect 27550 -3090 27670 -2970
rect 27725 -3090 27845 -2970
rect 27890 -3090 28010 -2970
rect 28055 -3090 28175 -2970
rect 28220 -3090 28340 -2970
rect 28395 -3090 28515 -2970
rect 28560 -3090 28680 -2970
rect 28725 -3090 28845 -2970
rect 28890 -3090 29010 -2970
rect 29065 -3090 29185 -2970
rect 29230 -3090 29350 -2970
rect 29395 -3090 29515 -2970
rect 29560 -3090 29680 -2970
rect 24200 -3255 24320 -3135
rect 24375 -3255 24495 -3135
rect 24540 -3255 24660 -3135
rect 24705 -3255 24825 -3135
rect 24870 -3255 24990 -3135
rect 25045 -3255 25165 -3135
rect 25210 -3255 25330 -3135
rect 25375 -3255 25495 -3135
rect 25540 -3255 25660 -3135
rect 25715 -3255 25835 -3135
rect 25880 -3255 26000 -3135
rect 26045 -3255 26165 -3135
rect 26210 -3255 26330 -3135
rect 26385 -3255 26505 -3135
rect 26550 -3255 26670 -3135
rect 26715 -3255 26835 -3135
rect 26880 -3255 27000 -3135
rect 27055 -3255 27175 -3135
rect 27220 -3255 27340 -3135
rect 27385 -3255 27505 -3135
rect 27550 -3255 27670 -3135
rect 27725 -3255 27845 -3135
rect 27890 -3255 28010 -3135
rect 28055 -3255 28175 -3135
rect 28220 -3255 28340 -3135
rect 28395 -3255 28515 -3135
rect 28560 -3255 28680 -3135
rect 28725 -3255 28845 -3135
rect 28890 -3255 29010 -3135
rect 29065 -3255 29185 -3135
rect 29230 -3255 29350 -3135
rect 29395 -3255 29515 -3135
rect 29560 -3255 29680 -3135
rect 24200 -3430 24320 -3310
rect 24375 -3430 24495 -3310
rect 24540 -3430 24660 -3310
rect 24705 -3430 24825 -3310
rect 24870 -3430 24990 -3310
rect 25045 -3430 25165 -3310
rect 25210 -3430 25330 -3310
rect 25375 -3430 25495 -3310
rect 25540 -3430 25660 -3310
rect 25715 -3430 25835 -3310
rect 25880 -3430 26000 -3310
rect 26045 -3430 26165 -3310
rect 26210 -3430 26330 -3310
rect 26385 -3430 26505 -3310
rect 26550 -3430 26670 -3310
rect 26715 -3430 26835 -3310
rect 26880 -3430 27000 -3310
rect 27055 -3430 27175 -3310
rect 27220 -3430 27340 -3310
rect 27385 -3430 27505 -3310
rect 27550 -3430 27670 -3310
rect 27725 -3430 27845 -3310
rect 27890 -3430 28010 -3310
rect 28055 -3430 28175 -3310
rect 28220 -3430 28340 -3310
rect 28395 -3430 28515 -3310
rect 28560 -3430 28680 -3310
rect 28725 -3430 28845 -3310
rect 28890 -3430 29010 -3310
rect 29065 -3430 29185 -3310
rect 29230 -3430 29350 -3310
rect 29395 -3430 29515 -3310
rect 29560 -3430 29680 -3310
rect 24200 -3595 24320 -3475
rect 24375 -3595 24495 -3475
rect 24540 -3595 24660 -3475
rect 24705 -3595 24825 -3475
rect 24870 -3595 24990 -3475
rect 25045 -3595 25165 -3475
rect 25210 -3595 25330 -3475
rect 25375 -3595 25495 -3475
rect 25540 -3595 25660 -3475
rect 25715 -3595 25835 -3475
rect 25880 -3595 26000 -3475
rect 26045 -3595 26165 -3475
rect 26210 -3595 26330 -3475
rect 26385 -3595 26505 -3475
rect 26550 -3595 26670 -3475
rect 26715 -3595 26835 -3475
rect 26880 -3595 27000 -3475
rect 27055 -3595 27175 -3475
rect 27220 -3595 27340 -3475
rect 27385 -3595 27505 -3475
rect 27550 -3595 27670 -3475
rect 27725 -3595 27845 -3475
rect 27890 -3595 28010 -3475
rect 28055 -3595 28175 -3475
rect 28220 -3595 28340 -3475
rect 28395 -3595 28515 -3475
rect 28560 -3595 28680 -3475
rect 28725 -3595 28845 -3475
rect 28890 -3595 29010 -3475
rect 29065 -3595 29185 -3475
rect 29230 -3595 29350 -3475
rect 29395 -3595 29515 -3475
rect 29560 -3595 29680 -3475
rect 24200 -3760 24320 -3640
rect 24375 -3760 24495 -3640
rect 24540 -3760 24660 -3640
rect 24705 -3760 24825 -3640
rect 24870 -3760 24990 -3640
rect 25045 -3760 25165 -3640
rect 25210 -3760 25330 -3640
rect 25375 -3760 25495 -3640
rect 25540 -3760 25660 -3640
rect 25715 -3760 25835 -3640
rect 25880 -3760 26000 -3640
rect 26045 -3760 26165 -3640
rect 26210 -3760 26330 -3640
rect 26385 -3760 26505 -3640
rect 26550 -3760 26670 -3640
rect 26715 -3760 26835 -3640
rect 26880 -3760 27000 -3640
rect 27055 -3760 27175 -3640
rect 27220 -3760 27340 -3640
rect 27385 -3760 27505 -3640
rect 27550 -3760 27670 -3640
rect 27725 -3760 27845 -3640
rect 27890 -3760 28010 -3640
rect 28055 -3760 28175 -3640
rect 28220 -3760 28340 -3640
rect 28395 -3760 28515 -3640
rect 28560 -3760 28680 -3640
rect 28725 -3760 28845 -3640
rect 28890 -3760 29010 -3640
rect 29065 -3760 29185 -3640
rect 29230 -3760 29350 -3640
rect 29395 -3760 29515 -3640
rect 29560 -3760 29680 -3640
rect 24200 -3925 24320 -3805
rect 24375 -3925 24495 -3805
rect 24540 -3925 24660 -3805
rect 24705 -3925 24825 -3805
rect 24870 -3925 24990 -3805
rect 25045 -3925 25165 -3805
rect 25210 -3925 25330 -3805
rect 25375 -3925 25495 -3805
rect 25540 -3925 25660 -3805
rect 25715 -3925 25835 -3805
rect 25880 -3925 26000 -3805
rect 26045 -3925 26165 -3805
rect 26210 -3925 26330 -3805
rect 26385 -3925 26505 -3805
rect 26550 -3925 26670 -3805
rect 26715 -3925 26835 -3805
rect 26880 -3925 27000 -3805
rect 27055 -3925 27175 -3805
rect 27220 -3925 27340 -3805
rect 27385 -3925 27505 -3805
rect 27550 -3925 27670 -3805
rect 27725 -3925 27845 -3805
rect 27890 -3925 28010 -3805
rect 28055 -3925 28175 -3805
rect 28220 -3925 28340 -3805
rect 28395 -3925 28515 -3805
rect 28560 -3925 28680 -3805
rect 28725 -3925 28845 -3805
rect 28890 -3925 29010 -3805
rect 29065 -3925 29185 -3805
rect 29230 -3925 29350 -3805
rect 29395 -3925 29515 -3805
rect 29560 -3925 29680 -3805
rect 24200 -4100 24320 -3980
rect 24375 -4100 24495 -3980
rect 24540 -4100 24660 -3980
rect 24705 -4100 24825 -3980
rect 24870 -4100 24990 -3980
rect 25045 -4100 25165 -3980
rect 25210 -4100 25330 -3980
rect 25375 -4100 25495 -3980
rect 25540 -4100 25660 -3980
rect 25715 -4100 25835 -3980
rect 25880 -4100 26000 -3980
rect 26045 -4100 26165 -3980
rect 26210 -4100 26330 -3980
rect 26385 -4100 26505 -3980
rect 26550 -4100 26670 -3980
rect 26715 -4100 26835 -3980
rect 26880 -4100 27000 -3980
rect 27055 -4100 27175 -3980
rect 27220 -4100 27340 -3980
rect 27385 -4100 27505 -3980
rect 27550 -4100 27670 -3980
rect 27725 -4100 27845 -3980
rect 27890 -4100 28010 -3980
rect 28055 -4100 28175 -3980
rect 28220 -4100 28340 -3980
rect 28395 -4100 28515 -3980
rect 28560 -4100 28680 -3980
rect 28725 -4100 28845 -3980
rect 28890 -4100 29010 -3980
rect 29065 -4100 29185 -3980
rect 29230 -4100 29350 -3980
rect 29395 -4100 29515 -3980
rect 29560 -4100 29680 -3980
rect 7130 -4430 7250 -4310
rect 7295 -4430 7415 -4310
rect 7460 -4430 7580 -4310
rect 7625 -4430 7745 -4310
rect 7800 -4430 7920 -4310
rect 7965 -4430 8085 -4310
rect 8130 -4430 8250 -4310
rect 8295 -4430 8415 -4310
rect 8470 -4430 8590 -4310
rect 8635 -4430 8755 -4310
rect 8800 -4430 8920 -4310
rect 8965 -4430 9085 -4310
rect 9140 -4430 9260 -4310
rect 9305 -4430 9425 -4310
rect 9470 -4430 9590 -4310
rect 9635 -4430 9755 -4310
rect 9810 -4430 9930 -4310
rect 9975 -4430 10095 -4310
rect 10140 -4430 10260 -4310
rect 10305 -4430 10425 -4310
rect 10480 -4430 10600 -4310
rect 10645 -4430 10765 -4310
rect 10810 -4430 10930 -4310
rect 10975 -4430 11095 -4310
rect 11150 -4430 11270 -4310
rect 11315 -4430 11435 -4310
rect 11480 -4430 11600 -4310
rect 11645 -4430 11765 -4310
rect 11820 -4430 11940 -4310
rect 11985 -4430 12105 -4310
rect 12150 -4430 12270 -4310
rect 12315 -4430 12435 -4310
rect 12490 -4430 12610 -4310
rect 7130 -4605 7250 -4485
rect 7295 -4605 7415 -4485
rect 7460 -4605 7580 -4485
rect 7625 -4605 7745 -4485
rect 7800 -4605 7920 -4485
rect 7965 -4605 8085 -4485
rect 8130 -4605 8250 -4485
rect 8295 -4605 8415 -4485
rect 8470 -4605 8590 -4485
rect 8635 -4605 8755 -4485
rect 8800 -4605 8920 -4485
rect 8965 -4605 9085 -4485
rect 9140 -4605 9260 -4485
rect 9305 -4605 9425 -4485
rect 9470 -4605 9590 -4485
rect 9635 -4605 9755 -4485
rect 9810 -4605 9930 -4485
rect 9975 -4605 10095 -4485
rect 10140 -4605 10260 -4485
rect 10305 -4605 10425 -4485
rect 10480 -4605 10600 -4485
rect 10645 -4605 10765 -4485
rect 10810 -4605 10930 -4485
rect 10975 -4605 11095 -4485
rect 11150 -4605 11270 -4485
rect 11315 -4605 11435 -4485
rect 11480 -4605 11600 -4485
rect 11645 -4605 11765 -4485
rect 11820 -4605 11940 -4485
rect 11985 -4605 12105 -4485
rect 12150 -4605 12270 -4485
rect 12315 -4605 12435 -4485
rect 12490 -4605 12610 -4485
rect 7130 -4770 7250 -4650
rect 7295 -4770 7415 -4650
rect 7460 -4770 7580 -4650
rect 7625 -4770 7745 -4650
rect 7800 -4770 7920 -4650
rect 7965 -4770 8085 -4650
rect 8130 -4770 8250 -4650
rect 8295 -4770 8415 -4650
rect 8470 -4770 8590 -4650
rect 8635 -4770 8755 -4650
rect 8800 -4770 8920 -4650
rect 8965 -4770 9085 -4650
rect 9140 -4770 9260 -4650
rect 9305 -4770 9425 -4650
rect 9470 -4770 9590 -4650
rect 9635 -4770 9755 -4650
rect 9810 -4770 9930 -4650
rect 9975 -4770 10095 -4650
rect 10140 -4770 10260 -4650
rect 10305 -4770 10425 -4650
rect 10480 -4770 10600 -4650
rect 10645 -4770 10765 -4650
rect 10810 -4770 10930 -4650
rect 10975 -4770 11095 -4650
rect 11150 -4770 11270 -4650
rect 11315 -4770 11435 -4650
rect 11480 -4770 11600 -4650
rect 11645 -4770 11765 -4650
rect 11820 -4770 11940 -4650
rect 11985 -4770 12105 -4650
rect 12150 -4770 12270 -4650
rect 12315 -4770 12435 -4650
rect 12490 -4770 12610 -4650
rect 7130 -4935 7250 -4815
rect 7295 -4935 7415 -4815
rect 7460 -4935 7580 -4815
rect 7625 -4935 7745 -4815
rect 7800 -4935 7920 -4815
rect 7965 -4935 8085 -4815
rect 8130 -4935 8250 -4815
rect 8295 -4935 8415 -4815
rect 8470 -4935 8590 -4815
rect 8635 -4935 8755 -4815
rect 8800 -4935 8920 -4815
rect 8965 -4935 9085 -4815
rect 9140 -4935 9260 -4815
rect 9305 -4935 9425 -4815
rect 9470 -4935 9590 -4815
rect 9635 -4935 9755 -4815
rect 9810 -4935 9930 -4815
rect 9975 -4935 10095 -4815
rect 10140 -4935 10260 -4815
rect 10305 -4935 10425 -4815
rect 10480 -4935 10600 -4815
rect 10645 -4935 10765 -4815
rect 10810 -4935 10930 -4815
rect 10975 -4935 11095 -4815
rect 11150 -4935 11270 -4815
rect 11315 -4935 11435 -4815
rect 11480 -4935 11600 -4815
rect 11645 -4935 11765 -4815
rect 11820 -4935 11940 -4815
rect 11985 -4935 12105 -4815
rect 12150 -4935 12270 -4815
rect 12315 -4935 12435 -4815
rect 12490 -4935 12610 -4815
rect 7130 -5100 7250 -4980
rect 7295 -5100 7415 -4980
rect 7460 -5100 7580 -4980
rect 7625 -5100 7745 -4980
rect 7800 -5100 7920 -4980
rect 7965 -5100 8085 -4980
rect 8130 -5100 8250 -4980
rect 8295 -5100 8415 -4980
rect 8470 -5100 8590 -4980
rect 8635 -5100 8755 -4980
rect 8800 -5100 8920 -4980
rect 8965 -5100 9085 -4980
rect 9140 -5100 9260 -4980
rect 9305 -5100 9425 -4980
rect 9470 -5100 9590 -4980
rect 9635 -5100 9755 -4980
rect 9810 -5100 9930 -4980
rect 9975 -5100 10095 -4980
rect 10140 -5100 10260 -4980
rect 10305 -5100 10425 -4980
rect 10480 -5100 10600 -4980
rect 10645 -5100 10765 -4980
rect 10810 -5100 10930 -4980
rect 10975 -5100 11095 -4980
rect 11150 -5100 11270 -4980
rect 11315 -5100 11435 -4980
rect 11480 -5100 11600 -4980
rect 11645 -5100 11765 -4980
rect 11820 -5100 11940 -4980
rect 11985 -5100 12105 -4980
rect 12150 -5100 12270 -4980
rect 12315 -5100 12435 -4980
rect 12490 -5100 12610 -4980
rect 7130 -5275 7250 -5155
rect 7295 -5275 7415 -5155
rect 7460 -5275 7580 -5155
rect 7625 -5275 7745 -5155
rect 7800 -5275 7920 -5155
rect 7965 -5275 8085 -5155
rect 8130 -5275 8250 -5155
rect 8295 -5275 8415 -5155
rect 8470 -5275 8590 -5155
rect 8635 -5275 8755 -5155
rect 8800 -5275 8920 -5155
rect 8965 -5275 9085 -5155
rect 9140 -5275 9260 -5155
rect 9305 -5275 9425 -5155
rect 9470 -5275 9590 -5155
rect 9635 -5275 9755 -5155
rect 9810 -5275 9930 -5155
rect 9975 -5275 10095 -5155
rect 10140 -5275 10260 -5155
rect 10305 -5275 10425 -5155
rect 10480 -5275 10600 -5155
rect 10645 -5275 10765 -5155
rect 10810 -5275 10930 -5155
rect 10975 -5275 11095 -5155
rect 11150 -5275 11270 -5155
rect 11315 -5275 11435 -5155
rect 11480 -5275 11600 -5155
rect 11645 -5275 11765 -5155
rect 11820 -5275 11940 -5155
rect 11985 -5275 12105 -5155
rect 12150 -5275 12270 -5155
rect 12315 -5275 12435 -5155
rect 12490 -5275 12610 -5155
rect 7130 -5440 7250 -5320
rect 7295 -5440 7415 -5320
rect 7460 -5440 7580 -5320
rect 7625 -5440 7745 -5320
rect 7800 -5440 7920 -5320
rect 7965 -5440 8085 -5320
rect 8130 -5440 8250 -5320
rect 8295 -5440 8415 -5320
rect 8470 -5440 8590 -5320
rect 8635 -5440 8755 -5320
rect 8800 -5440 8920 -5320
rect 8965 -5440 9085 -5320
rect 9140 -5440 9260 -5320
rect 9305 -5440 9425 -5320
rect 9470 -5440 9590 -5320
rect 9635 -5440 9755 -5320
rect 9810 -5440 9930 -5320
rect 9975 -5440 10095 -5320
rect 10140 -5440 10260 -5320
rect 10305 -5440 10425 -5320
rect 10480 -5440 10600 -5320
rect 10645 -5440 10765 -5320
rect 10810 -5440 10930 -5320
rect 10975 -5440 11095 -5320
rect 11150 -5440 11270 -5320
rect 11315 -5440 11435 -5320
rect 11480 -5440 11600 -5320
rect 11645 -5440 11765 -5320
rect 11820 -5440 11940 -5320
rect 11985 -5440 12105 -5320
rect 12150 -5440 12270 -5320
rect 12315 -5440 12435 -5320
rect 12490 -5440 12610 -5320
rect 7130 -5605 7250 -5485
rect 7295 -5605 7415 -5485
rect 7460 -5605 7580 -5485
rect 7625 -5605 7745 -5485
rect 7800 -5605 7920 -5485
rect 7965 -5605 8085 -5485
rect 8130 -5605 8250 -5485
rect 8295 -5605 8415 -5485
rect 8470 -5605 8590 -5485
rect 8635 -5605 8755 -5485
rect 8800 -5605 8920 -5485
rect 8965 -5605 9085 -5485
rect 9140 -5605 9260 -5485
rect 9305 -5605 9425 -5485
rect 9470 -5605 9590 -5485
rect 9635 -5605 9755 -5485
rect 9810 -5605 9930 -5485
rect 9975 -5605 10095 -5485
rect 10140 -5605 10260 -5485
rect 10305 -5605 10425 -5485
rect 10480 -5605 10600 -5485
rect 10645 -5605 10765 -5485
rect 10810 -5605 10930 -5485
rect 10975 -5605 11095 -5485
rect 11150 -5605 11270 -5485
rect 11315 -5605 11435 -5485
rect 11480 -5605 11600 -5485
rect 11645 -5605 11765 -5485
rect 11820 -5605 11940 -5485
rect 11985 -5605 12105 -5485
rect 12150 -5605 12270 -5485
rect 12315 -5605 12435 -5485
rect 12490 -5605 12610 -5485
rect 7130 -5770 7250 -5650
rect 7295 -5770 7415 -5650
rect 7460 -5770 7580 -5650
rect 7625 -5770 7745 -5650
rect 7800 -5770 7920 -5650
rect 7965 -5770 8085 -5650
rect 8130 -5770 8250 -5650
rect 8295 -5770 8415 -5650
rect 8470 -5770 8590 -5650
rect 8635 -5770 8755 -5650
rect 8800 -5770 8920 -5650
rect 8965 -5770 9085 -5650
rect 9140 -5770 9260 -5650
rect 9305 -5770 9425 -5650
rect 9470 -5770 9590 -5650
rect 9635 -5770 9755 -5650
rect 9810 -5770 9930 -5650
rect 9975 -5770 10095 -5650
rect 10140 -5770 10260 -5650
rect 10305 -5770 10425 -5650
rect 10480 -5770 10600 -5650
rect 10645 -5770 10765 -5650
rect 10810 -5770 10930 -5650
rect 10975 -5770 11095 -5650
rect 11150 -5770 11270 -5650
rect 11315 -5770 11435 -5650
rect 11480 -5770 11600 -5650
rect 11645 -5770 11765 -5650
rect 11820 -5770 11940 -5650
rect 11985 -5770 12105 -5650
rect 12150 -5770 12270 -5650
rect 12315 -5770 12435 -5650
rect 12490 -5770 12610 -5650
rect 7130 -5945 7250 -5825
rect 7295 -5945 7415 -5825
rect 7460 -5945 7580 -5825
rect 7625 -5945 7745 -5825
rect 7800 -5945 7920 -5825
rect 7965 -5945 8085 -5825
rect 8130 -5945 8250 -5825
rect 8295 -5945 8415 -5825
rect 8470 -5945 8590 -5825
rect 8635 -5945 8755 -5825
rect 8800 -5945 8920 -5825
rect 8965 -5945 9085 -5825
rect 9140 -5945 9260 -5825
rect 9305 -5945 9425 -5825
rect 9470 -5945 9590 -5825
rect 9635 -5945 9755 -5825
rect 9810 -5945 9930 -5825
rect 9975 -5945 10095 -5825
rect 10140 -5945 10260 -5825
rect 10305 -5945 10425 -5825
rect 10480 -5945 10600 -5825
rect 10645 -5945 10765 -5825
rect 10810 -5945 10930 -5825
rect 10975 -5945 11095 -5825
rect 11150 -5945 11270 -5825
rect 11315 -5945 11435 -5825
rect 11480 -5945 11600 -5825
rect 11645 -5945 11765 -5825
rect 11820 -5945 11940 -5825
rect 11985 -5945 12105 -5825
rect 12150 -5945 12270 -5825
rect 12315 -5945 12435 -5825
rect 12490 -5945 12610 -5825
rect 7130 -6110 7250 -5990
rect 7295 -6110 7415 -5990
rect 7460 -6110 7580 -5990
rect 7625 -6110 7745 -5990
rect 7800 -6110 7920 -5990
rect 7965 -6110 8085 -5990
rect 8130 -6110 8250 -5990
rect 8295 -6110 8415 -5990
rect 8470 -6110 8590 -5990
rect 8635 -6110 8755 -5990
rect 8800 -6110 8920 -5990
rect 8965 -6110 9085 -5990
rect 9140 -6110 9260 -5990
rect 9305 -6110 9425 -5990
rect 9470 -6110 9590 -5990
rect 9635 -6110 9755 -5990
rect 9810 -6110 9930 -5990
rect 9975 -6110 10095 -5990
rect 10140 -6110 10260 -5990
rect 10305 -6110 10425 -5990
rect 10480 -6110 10600 -5990
rect 10645 -6110 10765 -5990
rect 10810 -6110 10930 -5990
rect 10975 -6110 11095 -5990
rect 11150 -6110 11270 -5990
rect 11315 -6110 11435 -5990
rect 11480 -6110 11600 -5990
rect 11645 -6110 11765 -5990
rect 11820 -6110 11940 -5990
rect 11985 -6110 12105 -5990
rect 12150 -6110 12270 -5990
rect 12315 -6110 12435 -5990
rect 12490 -6110 12610 -5990
rect 7130 -6275 7250 -6155
rect 7295 -6275 7415 -6155
rect 7460 -6275 7580 -6155
rect 7625 -6275 7745 -6155
rect 7800 -6275 7920 -6155
rect 7965 -6275 8085 -6155
rect 8130 -6275 8250 -6155
rect 8295 -6275 8415 -6155
rect 8470 -6275 8590 -6155
rect 8635 -6275 8755 -6155
rect 8800 -6275 8920 -6155
rect 8965 -6275 9085 -6155
rect 9140 -6275 9260 -6155
rect 9305 -6275 9425 -6155
rect 9470 -6275 9590 -6155
rect 9635 -6275 9755 -6155
rect 9810 -6275 9930 -6155
rect 9975 -6275 10095 -6155
rect 10140 -6275 10260 -6155
rect 10305 -6275 10425 -6155
rect 10480 -6275 10600 -6155
rect 10645 -6275 10765 -6155
rect 10810 -6275 10930 -6155
rect 10975 -6275 11095 -6155
rect 11150 -6275 11270 -6155
rect 11315 -6275 11435 -6155
rect 11480 -6275 11600 -6155
rect 11645 -6275 11765 -6155
rect 11820 -6275 11940 -6155
rect 11985 -6275 12105 -6155
rect 12150 -6275 12270 -6155
rect 12315 -6275 12435 -6155
rect 12490 -6275 12610 -6155
rect 7130 -6440 7250 -6320
rect 7295 -6440 7415 -6320
rect 7460 -6440 7580 -6320
rect 7625 -6440 7745 -6320
rect 7800 -6440 7920 -6320
rect 7965 -6440 8085 -6320
rect 8130 -6440 8250 -6320
rect 8295 -6440 8415 -6320
rect 8470 -6440 8590 -6320
rect 8635 -6440 8755 -6320
rect 8800 -6440 8920 -6320
rect 8965 -6440 9085 -6320
rect 9140 -6440 9260 -6320
rect 9305 -6440 9425 -6320
rect 9470 -6440 9590 -6320
rect 9635 -6440 9755 -6320
rect 9810 -6440 9930 -6320
rect 9975 -6440 10095 -6320
rect 10140 -6440 10260 -6320
rect 10305 -6440 10425 -6320
rect 10480 -6440 10600 -6320
rect 10645 -6440 10765 -6320
rect 10810 -6440 10930 -6320
rect 10975 -6440 11095 -6320
rect 11150 -6440 11270 -6320
rect 11315 -6440 11435 -6320
rect 11480 -6440 11600 -6320
rect 11645 -6440 11765 -6320
rect 11820 -6440 11940 -6320
rect 11985 -6440 12105 -6320
rect 12150 -6440 12270 -6320
rect 12315 -6440 12435 -6320
rect 12490 -6440 12610 -6320
rect 7130 -6615 7250 -6495
rect 7295 -6615 7415 -6495
rect 7460 -6615 7580 -6495
rect 7625 -6615 7745 -6495
rect 7800 -6615 7920 -6495
rect 7965 -6615 8085 -6495
rect 8130 -6615 8250 -6495
rect 8295 -6615 8415 -6495
rect 8470 -6615 8590 -6495
rect 8635 -6615 8755 -6495
rect 8800 -6615 8920 -6495
rect 8965 -6615 9085 -6495
rect 9140 -6615 9260 -6495
rect 9305 -6615 9425 -6495
rect 9470 -6615 9590 -6495
rect 9635 -6615 9755 -6495
rect 9810 -6615 9930 -6495
rect 9975 -6615 10095 -6495
rect 10140 -6615 10260 -6495
rect 10305 -6615 10425 -6495
rect 10480 -6615 10600 -6495
rect 10645 -6615 10765 -6495
rect 10810 -6615 10930 -6495
rect 10975 -6615 11095 -6495
rect 11150 -6615 11270 -6495
rect 11315 -6615 11435 -6495
rect 11480 -6615 11600 -6495
rect 11645 -6615 11765 -6495
rect 11820 -6615 11940 -6495
rect 11985 -6615 12105 -6495
rect 12150 -6615 12270 -6495
rect 12315 -6615 12435 -6495
rect 12490 -6615 12610 -6495
rect 7130 -6780 7250 -6660
rect 7295 -6780 7415 -6660
rect 7460 -6780 7580 -6660
rect 7625 -6780 7745 -6660
rect 7800 -6780 7920 -6660
rect 7965 -6780 8085 -6660
rect 8130 -6780 8250 -6660
rect 8295 -6780 8415 -6660
rect 8470 -6780 8590 -6660
rect 8635 -6780 8755 -6660
rect 8800 -6780 8920 -6660
rect 8965 -6780 9085 -6660
rect 9140 -6780 9260 -6660
rect 9305 -6780 9425 -6660
rect 9470 -6780 9590 -6660
rect 9635 -6780 9755 -6660
rect 9810 -6780 9930 -6660
rect 9975 -6780 10095 -6660
rect 10140 -6780 10260 -6660
rect 10305 -6780 10425 -6660
rect 10480 -6780 10600 -6660
rect 10645 -6780 10765 -6660
rect 10810 -6780 10930 -6660
rect 10975 -6780 11095 -6660
rect 11150 -6780 11270 -6660
rect 11315 -6780 11435 -6660
rect 11480 -6780 11600 -6660
rect 11645 -6780 11765 -6660
rect 11820 -6780 11940 -6660
rect 11985 -6780 12105 -6660
rect 12150 -6780 12270 -6660
rect 12315 -6780 12435 -6660
rect 12490 -6780 12610 -6660
rect 7130 -6945 7250 -6825
rect 7295 -6945 7415 -6825
rect 7460 -6945 7580 -6825
rect 7625 -6945 7745 -6825
rect 7800 -6945 7920 -6825
rect 7965 -6945 8085 -6825
rect 8130 -6945 8250 -6825
rect 8295 -6945 8415 -6825
rect 8470 -6945 8590 -6825
rect 8635 -6945 8755 -6825
rect 8800 -6945 8920 -6825
rect 8965 -6945 9085 -6825
rect 9140 -6945 9260 -6825
rect 9305 -6945 9425 -6825
rect 9470 -6945 9590 -6825
rect 9635 -6945 9755 -6825
rect 9810 -6945 9930 -6825
rect 9975 -6945 10095 -6825
rect 10140 -6945 10260 -6825
rect 10305 -6945 10425 -6825
rect 10480 -6945 10600 -6825
rect 10645 -6945 10765 -6825
rect 10810 -6945 10930 -6825
rect 10975 -6945 11095 -6825
rect 11150 -6945 11270 -6825
rect 11315 -6945 11435 -6825
rect 11480 -6945 11600 -6825
rect 11645 -6945 11765 -6825
rect 11820 -6945 11940 -6825
rect 11985 -6945 12105 -6825
rect 12150 -6945 12270 -6825
rect 12315 -6945 12435 -6825
rect 12490 -6945 12610 -6825
rect 7130 -7110 7250 -6990
rect 7295 -7110 7415 -6990
rect 7460 -7110 7580 -6990
rect 7625 -7110 7745 -6990
rect 7800 -7110 7920 -6990
rect 7965 -7110 8085 -6990
rect 8130 -7110 8250 -6990
rect 8295 -7110 8415 -6990
rect 8470 -7110 8590 -6990
rect 8635 -7110 8755 -6990
rect 8800 -7110 8920 -6990
rect 8965 -7110 9085 -6990
rect 9140 -7110 9260 -6990
rect 9305 -7110 9425 -6990
rect 9470 -7110 9590 -6990
rect 9635 -7110 9755 -6990
rect 9810 -7110 9930 -6990
rect 9975 -7110 10095 -6990
rect 10140 -7110 10260 -6990
rect 10305 -7110 10425 -6990
rect 10480 -7110 10600 -6990
rect 10645 -7110 10765 -6990
rect 10810 -7110 10930 -6990
rect 10975 -7110 11095 -6990
rect 11150 -7110 11270 -6990
rect 11315 -7110 11435 -6990
rect 11480 -7110 11600 -6990
rect 11645 -7110 11765 -6990
rect 11820 -7110 11940 -6990
rect 11985 -7110 12105 -6990
rect 12150 -7110 12270 -6990
rect 12315 -7110 12435 -6990
rect 12490 -7110 12610 -6990
rect 7130 -7285 7250 -7165
rect 7295 -7285 7415 -7165
rect 7460 -7285 7580 -7165
rect 7625 -7285 7745 -7165
rect 7800 -7285 7920 -7165
rect 7965 -7285 8085 -7165
rect 8130 -7285 8250 -7165
rect 8295 -7285 8415 -7165
rect 8470 -7285 8590 -7165
rect 8635 -7285 8755 -7165
rect 8800 -7285 8920 -7165
rect 8965 -7285 9085 -7165
rect 9140 -7285 9260 -7165
rect 9305 -7285 9425 -7165
rect 9470 -7285 9590 -7165
rect 9635 -7285 9755 -7165
rect 9810 -7285 9930 -7165
rect 9975 -7285 10095 -7165
rect 10140 -7285 10260 -7165
rect 10305 -7285 10425 -7165
rect 10480 -7285 10600 -7165
rect 10645 -7285 10765 -7165
rect 10810 -7285 10930 -7165
rect 10975 -7285 11095 -7165
rect 11150 -7285 11270 -7165
rect 11315 -7285 11435 -7165
rect 11480 -7285 11600 -7165
rect 11645 -7285 11765 -7165
rect 11820 -7285 11940 -7165
rect 11985 -7285 12105 -7165
rect 12150 -7285 12270 -7165
rect 12315 -7285 12435 -7165
rect 12490 -7285 12610 -7165
rect 7130 -7450 7250 -7330
rect 7295 -7450 7415 -7330
rect 7460 -7450 7580 -7330
rect 7625 -7450 7745 -7330
rect 7800 -7450 7920 -7330
rect 7965 -7450 8085 -7330
rect 8130 -7450 8250 -7330
rect 8295 -7450 8415 -7330
rect 8470 -7450 8590 -7330
rect 8635 -7450 8755 -7330
rect 8800 -7450 8920 -7330
rect 8965 -7450 9085 -7330
rect 9140 -7450 9260 -7330
rect 9305 -7450 9425 -7330
rect 9470 -7450 9590 -7330
rect 9635 -7450 9755 -7330
rect 9810 -7450 9930 -7330
rect 9975 -7450 10095 -7330
rect 10140 -7450 10260 -7330
rect 10305 -7450 10425 -7330
rect 10480 -7450 10600 -7330
rect 10645 -7450 10765 -7330
rect 10810 -7450 10930 -7330
rect 10975 -7450 11095 -7330
rect 11150 -7450 11270 -7330
rect 11315 -7450 11435 -7330
rect 11480 -7450 11600 -7330
rect 11645 -7450 11765 -7330
rect 11820 -7450 11940 -7330
rect 11985 -7450 12105 -7330
rect 12150 -7450 12270 -7330
rect 12315 -7450 12435 -7330
rect 12490 -7450 12610 -7330
rect 7130 -7615 7250 -7495
rect 7295 -7615 7415 -7495
rect 7460 -7615 7580 -7495
rect 7625 -7615 7745 -7495
rect 7800 -7615 7920 -7495
rect 7965 -7615 8085 -7495
rect 8130 -7615 8250 -7495
rect 8295 -7615 8415 -7495
rect 8470 -7615 8590 -7495
rect 8635 -7615 8755 -7495
rect 8800 -7615 8920 -7495
rect 8965 -7615 9085 -7495
rect 9140 -7615 9260 -7495
rect 9305 -7615 9425 -7495
rect 9470 -7615 9590 -7495
rect 9635 -7615 9755 -7495
rect 9810 -7615 9930 -7495
rect 9975 -7615 10095 -7495
rect 10140 -7615 10260 -7495
rect 10305 -7615 10425 -7495
rect 10480 -7615 10600 -7495
rect 10645 -7615 10765 -7495
rect 10810 -7615 10930 -7495
rect 10975 -7615 11095 -7495
rect 11150 -7615 11270 -7495
rect 11315 -7615 11435 -7495
rect 11480 -7615 11600 -7495
rect 11645 -7615 11765 -7495
rect 11820 -7615 11940 -7495
rect 11985 -7615 12105 -7495
rect 12150 -7615 12270 -7495
rect 12315 -7615 12435 -7495
rect 12490 -7615 12610 -7495
rect 7130 -7780 7250 -7660
rect 7295 -7780 7415 -7660
rect 7460 -7780 7580 -7660
rect 7625 -7780 7745 -7660
rect 7800 -7780 7920 -7660
rect 7965 -7780 8085 -7660
rect 8130 -7780 8250 -7660
rect 8295 -7780 8415 -7660
rect 8470 -7780 8590 -7660
rect 8635 -7780 8755 -7660
rect 8800 -7780 8920 -7660
rect 8965 -7780 9085 -7660
rect 9140 -7780 9260 -7660
rect 9305 -7780 9425 -7660
rect 9470 -7780 9590 -7660
rect 9635 -7780 9755 -7660
rect 9810 -7780 9930 -7660
rect 9975 -7780 10095 -7660
rect 10140 -7780 10260 -7660
rect 10305 -7780 10425 -7660
rect 10480 -7780 10600 -7660
rect 10645 -7780 10765 -7660
rect 10810 -7780 10930 -7660
rect 10975 -7780 11095 -7660
rect 11150 -7780 11270 -7660
rect 11315 -7780 11435 -7660
rect 11480 -7780 11600 -7660
rect 11645 -7780 11765 -7660
rect 11820 -7780 11940 -7660
rect 11985 -7780 12105 -7660
rect 12150 -7780 12270 -7660
rect 12315 -7780 12435 -7660
rect 12490 -7780 12610 -7660
rect 7130 -7955 7250 -7835
rect 7295 -7955 7415 -7835
rect 7460 -7955 7580 -7835
rect 7625 -7955 7745 -7835
rect 7800 -7955 7920 -7835
rect 7965 -7955 8085 -7835
rect 8130 -7955 8250 -7835
rect 8295 -7955 8415 -7835
rect 8470 -7955 8590 -7835
rect 8635 -7955 8755 -7835
rect 8800 -7955 8920 -7835
rect 8965 -7955 9085 -7835
rect 9140 -7955 9260 -7835
rect 9305 -7955 9425 -7835
rect 9470 -7955 9590 -7835
rect 9635 -7955 9755 -7835
rect 9810 -7955 9930 -7835
rect 9975 -7955 10095 -7835
rect 10140 -7955 10260 -7835
rect 10305 -7955 10425 -7835
rect 10480 -7955 10600 -7835
rect 10645 -7955 10765 -7835
rect 10810 -7955 10930 -7835
rect 10975 -7955 11095 -7835
rect 11150 -7955 11270 -7835
rect 11315 -7955 11435 -7835
rect 11480 -7955 11600 -7835
rect 11645 -7955 11765 -7835
rect 11820 -7955 11940 -7835
rect 11985 -7955 12105 -7835
rect 12150 -7955 12270 -7835
rect 12315 -7955 12435 -7835
rect 12490 -7955 12610 -7835
rect 7130 -8120 7250 -8000
rect 7295 -8120 7415 -8000
rect 7460 -8120 7580 -8000
rect 7625 -8120 7745 -8000
rect 7800 -8120 7920 -8000
rect 7965 -8120 8085 -8000
rect 8130 -8120 8250 -8000
rect 8295 -8120 8415 -8000
rect 8470 -8120 8590 -8000
rect 8635 -8120 8755 -8000
rect 8800 -8120 8920 -8000
rect 8965 -8120 9085 -8000
rect 9140 -8120 9260 -8000
rect 9305 -8120 9425 -8000
rect 9470 -8120 9590 -8000
rect 9635 -8120 9755 -8000
rect 9810 -8120 9930 -8000
rect 9975 -8120 10095 -8000
rect 10140 -8120 10260 -8000
rect 10305 -8120 10425 -8000
rect 10480 -8120 10600 -8000
rect 10645 -8120 10765 -8000
rect 10810 -8120 10930 -8000
rect 10975 -8120 11095 -8000
rect 11150 -8120 11270 -8000
rect 11315 -8120 11435 -8000
rect 11480 -8120 11600 -8000
rect 11645 -8120 11765 -8000
rect 11820 -8120 11940 -8000
rect 11985 -8120 12105 -8000
rect 12150 -8120 12270 -8000
rect 12315 -8120 12435 -8000
rect 12490 -8120 12610 -8000
rect 7130 -8285 7250 -8165
rect 7295 -8285 7415 -8165
rect 7460 -8285 7580 -8165
rect 7625 -8285 7745 -8165
rect 7800 -8285 7920 -8165
rect 7965 -8285 8085 -8165
rect 8130 -8285 8250 -8165
rect 8295 -8285 8415 -8165
rect 8470 -8285 8590 -8165
rect 8635 -8285 8755 -8165
rect 8800 -8285 8920 -8165
rect 8965 -8285 9085 -8165
rect 9140 -8285 9260 -8165
rect 9305 -8285 9425 -8165
rect 9470 -8285 9590 -8165
rect 9635 -8285 9755 -8165
rect 9810 -8285 9930 -8165
rect 9975 -8285 10095 -8165
rect 10140 -8285 10260 -8165
rect 10305 -8285 10425 -8165
rect 10480 -8285 10600 -8165
rect 10645 -8285 10765 -8165
rect 10810 -8285 10930 -8165
rect 10975 -8285 11095 -8165
rect 11150 -8285 11270 -8165
rect 11315 -8285 11435 -8165
rect 11480 -8285 11600 -8165
rect 11645 -8285 11765 -8165
rect 11820 -8285 11940 -8165
rect 11985 -8285 12105 -8165
rect 12150 -8285 12270 -8165
rect 12315 -8285 12435 -8165
rect 12490 -8285 12610 -8165
rect 7130 -8450 7250 -8330
rect 7295 -8450 7415 -8330
rect 7460 -8450 7580 -8330
rect 7625 -8450 7745 -8330
rect 7800 -8450 7920 -8330
rect 7965 -8450 8085 -8330
rect 8130 -8450 8250 -8330
rect 8295 -8450 8415 -8330
rect 8470 -8450 8590 -8330
rect 8635 -8450 8755 -8330
rect 8800 -8450 8920 -8330
rect 8965 -8450 9085 -8330
rect 9140 -8450 9260 -8330
rect 9305 -8450 9425 -8330
rect 9470 -8450 9590 -8330
rect 9635 -8450 9755 -8330
rect 9810 -8450 9930 -8330
rect 9975 -8450 10095 -8330
rect 10140 -8450 10260 -8330
rect 10305 -8450 10425 -8330
rect 10480 -8450 10600 -8330
rect 10645 -8450 10765 -8330
rect 10810 -8450 10930 -8330
rect 10975 -8450 11095 -8330
rect 11150 -8450 11270 -8330
rect 11315 -8450 11435 -8330
rect 11480 -8450 11600 -8330
rect 11645 -8450 11765 -8330
rect 11820 -8450 11940 -8330
rect 11985 -8450 12105 -8330
rect 12150 -8450 12270 -8330
rect 12315 -8450 12435 -8330
rect 12490 -8450 12610 -8330
rect 7130 -8625 7250 -8505
rect 7295 -8625 7415 -8505
rect 7460 -8625 7580 -8505
rect 7625 -8625 7745 -8505
rect 7800 -8625 7920 -8505
rect 7965 -8625 8085 -8505
rect 8130 -8625 8250 -8505
rect 8295 -8625 8415 -8505
rect 8470 -8625 8590 -8505
rect 8635 -8625 8755 -8505
rect 8800 -8625 8920 -8505
rect 8965 -8625 9085 -8505
rect 9140 -8625 9260 -8505
rect 9305 -8625 9425 -8505
rect 9470 -8625 9590 -8505
rect 9635 -8625 9755 -8505
rect 9810 -8625 9930 -8505
rect 9975 -8625 10095 -8505
rect 10140 -8625 10260 -8505
rect 10305 -8625 10425 -8505
rect 10480 -8625 10600 -8505
rect 10645 -8625 10765 -8505
rect 10810 -8625 10930 -8505
rect 10975 -8625 11095 -8505
rect 11150 -8625 11270 -8505
rect 11315 -8625 11435 -8505
rect 11480 -8625 11600 -8505
rect 11645 -8625 11765 -8505
rect 11820 -8625 11940 -8505
rect 11985 -8625 12105 -8505
rect 12150 -8625 12270 -8505
rect 12315 -8625 12435 -8505
rect 12490 -8625 12610 -8505
rect 7130 -8790 7250 -8670
rect 7295 -8790 7415 -8670
rect 7460 -8790 7580 -8670
rect 7625 -8790 7745 -8670
rect 7800 -8790 7920 -8670
rect 7965 -8790 8085 -8670
rect 8130 -8790 8250 -8670
rect 8295 -8790 8415 -8670
rect 8470 -8790 8590 -8670
rect 8635 -8790 8755 -8670
rect 8800 -8790 8920 -8670
rect 8965 -8790 9085 -8670
rect 9140 -8790 9260 -8670
rect 9305 -8790 9425 -8670
rect 9470 -8790 9590 -8670
rect 9635 -8790 9755 -8670
rect 9810 -8790 9930 -8670
rect 9975 -8790 10095 -8670
rect 10140 -8790 10260 -8670
rect 10305 -8790 10425 -8670
rect 10480 -8790 10600 -8670
rect 10645 -8790 10765 -8670
rect 10810 -8790 10930 -8670
rect 10975 -8790 11095 -8670
rect 11150 -8790 11270 -8670
rect 11315 -8790 11435 -8670
rect 11480 -8790 11600 -8670
rect 11645 -8790 11765 -8670
rect 11820 -8790 11940 -8670
rect 11985 -8790 12105 -8670
rect 12150 -8790 12270 -8670
rect 12315 -8790 12435 -8670
rect 12490 -8790 12610 -8670
rect 7130 -8955 7250 -8835
rect 7295 -8955 7415 -8835
rect 7460 -8955 7580 -8835
rect 7625 -8955 7745 -8835
rect 7800 -8955 7920 -8835
rect 7965 -8955 8085 -8835
rect 8130 -8955 8250 -8835
rect 8295 -8955 8415 -8835
rect 8470 -8955 8590 -8835
rect 8635 -8955 8755 -8835
rect 8800 -8955 8920 -8835
rect 8965 -8955 9085 -8835
rect 9140 -8955 9260 -8835
rect 9305 -8955 9425 -8835
rect 9470 -8955 9590 -8835
rect 9635 -8955 9755 -8835
rect 9810 -8955 9930 -8835
rect 9975 -8955 10095 -8835
rect 10140 -8955 10260 -8835
rect 10305 -8955 10425 -8835
rect 10480 -8955 10600 -8835
rect 10645 -8955 10765 -8835
rect 10810 -8955 10930 -8835
rect 10975 -8955 11095 -8835
rect 11150 -8955 11270 -8835
rect 11315 -8955 11435 -8835
rect 11480 -8955 11600 -8835
rect 11645 -8955 11765 -8835
rect 11820 -8955 11940 -8835
rect 11985 -8955 12105 -8835
rect 12150 -8955 12270 -8835
rect 12315 -8955 12435 -8835
rect 12490 -8955 12610 -8835
rect 7130 -9120 7250 -9000
rect 7295 -9120 7415 -9000
rect 7460 -9120 7580 -9000
rect 7625 -9120 7745 -9000
rect 7800 -9120 7920 -9000
rect 7965 -9120 8085 -9000
rect 8130 -9120 8250 -9000
rect 8295 -9120 8415 -9000
rect 8470 -9120 8590 -9000
rect 8635 -9120 8755 -9000
rect 8800 -9120 8920 -9000
rect 8965 -9120 9085 -9000
rect 9140 -9120 9260 -9000
rect 9305 -9120 9425 -9000
rect 9470 -9120 9590 -9000
rect 9635 -9120 9755 -9000
rect 9810 -9120 9930 -9000
rect 9975 -9120 10095 -9000
rect 10140 -9120 10260 -9000
rect 10305 -9120 10425 -9000
rect 10480 -9120 10600 -9000
rect 10645 -9120 10765 -9000
rect 10810 -9120 10930 -9000
rect 10975 -9120 11095 -9000
rect 11150 -9120 11270 -9000
rect 11315 -9120 11435 -9000
rect 11480 -9120 11600 -9000
rect 11645 -9120 11765 -9000
rect 11820 -9120 11940 -9000
rect 11985 -9120 12105 -9000
rect 12150 -9120 12270 -9000
rect 12315 -9120 12435 -9000
rect 12490 -9120 12610 -9000
rect 7130 -9295 7250 -9175
rect 7295 -9295 7415 -9175
rect 7460 -9295 7580 -9175
rect 7625 -9295 7745 -9175
rect 7800 -9295 7920 -9175
rect 7965 -9295 8085 -9175
rect 8130 -9295 8250 -9175
rect 8295 -9295 8415 -9175
rect 8470 -9295 8590 -9175
rect 8635 -9295 8755 -9175
rect 8800 -9295 8920 -9175
rect 8965 -9295 9085 -9175
rect 9140 -9295 9260 -9175
rect 9305 -9295 9425 -9175
rect 9470 -9295 9590 -9175
rect 9635 -9295 9755 -9175
rect 9810 -9295 9930 -9175
rect 9975 -9295 10095 -9175
rect 10140 -9295 10260 -9175
rect 10305 -9295 10425 -9175
rect 10480 -9295 10600 -9175
rect 10645 -9295 10765 -9175
rect 10810 -9295 10930 -9175
rect 10975 -9295 11095 -9175
rect 11150 -9295 11270 -9175
rect 11315 -9295 11435 -9175
rect 11480 -9295 11600 -9175
rect 11645 -9295 11765 -9175
rect 11820 -9295 11940 -9175
rect 11985 -9295 12105 -9175
rect 12150 -9295 12270 -9175
rect 12315 -9295 12435 -9175
rect 12490 -9295 12610 -9175
rect 7130 -9460 7250 -9340
rect 7295 -9460 7415 -9340
rect 7460 -9460 7580 -9340
rect 7625 -9460 7745 -9340
rect 7800 -9460 7920 -9340
rect 7965 -9460 8085 -9340
rect 8130 -9460 8250 -9340
rect 8295 -9460 8415 -9340
rect 8470 -9460 8590 -9340
rect 8635 -9460 8755 -9340
rect 8800 -9460 8920 -9340
rect 8965 -9460 9085 -9340
rect 9140 -9460 9260 -9340
rect 9305 -9460 9425 -9340
rect 9470 -9460 9590 -9340
rect 9635 -9460 9755 -9340
rect 9810 -9460 9930 -9340
rect 9975 -9460 10095 -9340
rect 10140 -9460 10260 -9340
rect 10305 -9460 10425 -9340
rect 10480 -9460 10600 -9340
rect 10645 -9460 10765 -9340
rect 10810 -9460 10930 -9340
rect 10975 -9460 11095 -9340
rect 11150 -9460 11270 -9340
rect 11315 -9460 11435 -9340
rect 11480 -9460 11600 -9340
rect 11645 -9460 11765 -9340
rect 11820 -9460 11940 -9340
rect 11985 -9460 12105 -9340
rect 12150 -9460 12270 -9340
rect 12315 -9460 12435 -9340
rect 12490 -9460 12610 -9340
rect 7130 -9625 7250 -9505
rect 7295 -9625 7415 -9505
rect 7460 -9625 7580 -9505
rect 7625 -9625 7745 -9505
rect 7800 -9625 7920 -9505
rect 7965 -9625 8085 -9505
rect 8130 -9625 8250 -9505
rect 8295 -9625 8415 -9505
rect 8470 -9625 8590 -9505
rect 8635 -9625 8755 -9505
rect 8800 -9625 8920 -9505
rect 8965 -9625 9085 -9505
rect 9140 -9625 9260 -9505
rect 9305 -9625 9425 -9505
rect 9470 -9625 9590 -9505
rect 9635 -9625 9755 -9505
rect 9810 -9625 9930 -9505
rect 9975 -9625 10095 -9505
rect 10140 -9625 10260 -9505
rect 10305 -9625 10425 -9505
rect 10480 -9625 10600 -9505
rect 10645 -9625 10765 -9505
rect 10810 -9625 10930 -9505
rect 10975 -9625 11095 -9505
rect 11150 -9625 11270 -9505
rect 11315 -9625 11435 -9505
rect 11480 -9625 11600 -9505
rect 11645 -9625 11765 -9505
rect 11820 -9625 11940 -9505
rect 11985 -9625 12105 -9505
rect 12150 -9625 12270 -9505
rect 12315 -9625 12435 -9505
rect 12490 -9625 12610 -9505
rect 7130 -9790 7250 -9670
rect 7295 -9790 7415 -9670
rect 7460 -9790 7580 -9670
rect 7625 -9790 7745 -9670
rect 7800 -9790 7920 -9670
rect 7965 -9790 8085 -9670
rect 8130 -9790 8250 -9670
rect 8295 -9790 8415 -9670
rect 8470 -9790 8590 -9670
rect 8635 -9790 8755 -9670
rect 8800 -9790 8920 -9670
rect 8965 -9790 9085 -9670
rect 9140 -9790 9260 -9670
rect 9305 -9790 9425 -9670
rect 9470 -9790 9590 -9670
rect 9635 -9790 9755 -9670
rect 9810 -9790 9930 -9670
rect 9975 -9790 10095 -9670
rect 10140 -9790 10260 -9670
rect 10305 -9790 10425 -9670
rect 10480 -9790 10600 -9670
rect 10645 -9790 10765 -9670
rect 10810 -9790 10930 -9670
rect 10975 -9790 11095 -9670
rect 11150 -9790 11270 -9670
rect 11315 -9790 11435 -9670
rect 11480 -9790 11600 -9670
rect 11645 -9790 11765 -9670
rect 11820 -9790 11940 -9670
rect 11985 -9790 12105 -9670
rect 12150 -9790 12270 -9670
rect 12315 -9790 12435 -9670
rect 12490 -9790 12610 -9670
rect 12820 -4430 12940 -4310
rect 12985 -4430 13105 -4310
rect 13150 -4430 13270 -4310
rect 13315 -4430 13435 -4310
rect 13490 -4430 13610 -4310
rect 13655 -4430 13775 -4310
rect 13820 -4430 13940 -4310
rect 13985 -4430 14105 -4310
rect 14160 -4430 14280 -4310
rect 14325 -4430 14445 -4310
rect 14490 -4430 14610 -4310
rect 14655 -4430 14775 -4310
rect 14830 -4430 14950 -4310
rect 14995 -4430 15115 -4310
rect 15160 -4430 15280 -4310
rect 15325 -4430 15445 -4310
rect 15500 -4430 15620 -4310
rect 15665 -4430 15785 -4310
rect 15830 -4430 15950 -4310
rect 15995 -4430 16115 -4310
rect 16170 -4430 16290 -4310
rect 16335 -4430 16455 -4310
rect 16500 -4430 16620 -4310
rect 16665 -4430 16785 -4310
rect 16840 -4430 16960 -4310
rect 17005 -4430 17125 -4310
rect 17170 -4430 17290 -4310
rect 17335 -4430 17455 -4310
rect 17510 -4430 17630 -4310
rect 17675 -4430 17795 -4310
rect 17840 -4430 17960 -4310
rect 18005 -4430 18125 -4310
rect 18180 -4430 18300 -4310
rect 12820 -4605 12940 -4485
rect 12985 -4605 13105 -4485
rect 13150 -4605 13270 -4485
rect 13315 -4605 13435 -4485
rect 13490 -4605 13610 -4485
rect 13655 -4605 13775 -4485
rect 13820 -4605 13940 -4485
rect 13985 -4605 14105 -4485
rect 14160 -4605 14280 -4485
rect 14325 -4605 14445 -4485
rect 14490 -4605 14610 -4485
rect 14655 -4605 14775 -4485
rect 14830 -4605 14950 -4485
rect 14995 -4605 15115 -4485
rect 15160 -4605 15280 -4485
rect 15325 -4605 15445 -4485
rect 15500 -4605 15620 -4485
rect 15665 -4605 15785 -4485
rect 15830 -4605 15950 -4485
rect 15995 -4605 16115 -4485
rect 16170 -4605 16290 -4485
rect 16335 -4605 16455 -4485
rect 16500 -4605 16620 -4485
rect 16665 -4605 16785 -4485
rect 16840 -4605 16960 -4485
rect 17005 -4605 17125 -4485
rect 17170 -4605 17290 -4485
rect 17335 -4605 17455 -4485
rect 17510 -4605 17630 -4485
rect 17675 -4605 17795 -4485
rect 17840 -4605 17960 -4485
rect 18005 -4605 18125 -4485
rect 18180 -4605 18300 -4485
rect 12820 -4770 12940 -4650
rect 12985 -4770 13105 -4650
rect 13150 -4770 13270 -4650
rect 13315 -4770 13435 -4650
rect 13490 -4770 13610 -4650
rect 13655 -4770 13775 -4650
rect 13820 -4770 13940 -4650
rect 13985 -4770 14105 -4650
rect 14160 -4770 14280 -4650
rect 14325 -4770 14445 -4650
rect 14490 -4770 14610 -4650
rect 14655 -4770 14775 -4650
rect 14830 -4770 14950 -4650
rect 14995 -4770 15115 -4650
rect 15160 -4770 15280 -4650
rect 15325 -4770 15445 -4650
rect 15500 -4770 15620 -4650
rect 15665 -4770 15785 -4650
rect 15830 -4770 15950 -4650
rect 15995 -4770 16115 -4650
rect 16170 -4770 16290 -4650
rect 16335 -4770 16455 -4650
rect 16500 -4770 16620 -4650
rect 16665 -4770 16785 -4650
rect 16840 -4770 16960 -4650
rect 17005 -4770 17125 -4650
rect 17170 -4770 17290 -4650
rect 17335 -4770 17455 -4650
rect 17510 -4770 17630 -4650
rect 17675 -4770 17795 -4650
rect 17840 -4770 17960 -4650
rect 18005 -4770 18125 -4650
rect 18180 -4770 18300 -4650
rect 12820 -4935 12940 -4815
rect 12985 -4935 13105 -4815
rect 13150 -4935 13270 -4815
rect 13315 -4935 13435 -4815
rect 13490 -4935 13610 -4815
rect 13655 -4935 13775 -4815
rect 13820 -4935 13940 -4815
rect 13985 -4935 14105 -4815
rect 14160 -4935 14280 -4815
rect 14325 -4935 14445 -4815
rect 14490 -4935 14610 -4815
rect 14655 -4935 14775 -4815
rect 14830 -4935 14950 -4815
rect 14995 -4935 15115 -4815
rect 15160 -4935 15280 -4815
rect 15325 -4935 15445 -4815
rect 15500 -4935 15620 -4815
rect 15665 -4935 15785 -4815
rect 15830 -4935 15950 -4815
rect 15995 -4935 16115 -4815
rect 16170 -4935 16290 -4815
rect 16335 -4935 16455 -4815
rect 16500 -4935 16620 -4815
rect 16665 -4935 16785 -4815
rect 16840 -4935 16960 -4815
rect 17005 -4935 17125 -4815
rect 17170 -4935 17290 -4815
rect 17335 -4935 17455 -4815
rect 17510 -4935 17630 -4815
rect 17675 -4935 17795 -4815
rect 17840 -4935 17960 -4815
rect 18005 -4935 18125 -4815
rect 18180 -4935 18300 -4815
rect 12820 -5100 12940 -4980
rect 12985 -5100 13105 -4980
rect 13150 -5100 13270 -4980
rect 13315 -5100 13435 -4980
rect 13490 -5100 13610 -4980
rect 13655 -5100 13775 -4980
rect 13820 -5100 13940 -4980
rect 13985 -5100 14105 -4980
rect 14160 -5100 14280 -4980
rect 14325 -5100 14445 -4980
rect 14490 -5100 14610 -4980
rect 14655 -5100 14775 -4980
rect 14830 -5100 14950 -4980
rect 14995 -5100 15115 -4980
rect 15160 -5100 15280 -4980
rect 15325 -5100 15445 -4980
rect 15500 -5100 15620 -4980
rect 15665 -5100 15785 -4980
rect 15830 -5100 15950 -4980
rect 15995 -5100 16115 -4980
rect 16170 -5100 16290 -4980
rect 16335 -5100 16455 -4980
rect 16500 -5100 16620 -4980
rect 16665 -5100 16785 -4980
rect 16840 -5100 16960 -4980
rect 17005 -5100 17125 -4980
rect 17170 -5100 17290 -4980
rect 17335 -5100 17455 -4980
rect 17510 -5100 17630 -4980
rect 17675 -5100 17795 -4980
rect 17840 -5100 17960 -4980
rect 18005 -5100 18125 -4980
rect 18180 -5100 18300 -4980
rect 12820 -5275 12940 -5155
rect 12985 -5275 13105 -5155
rect 13150 -5275 13270 -5155
rect 13315 -5275 13435 -5155
rect 13490 -5275 13610 -5155
rect 13655 -5275 13775 -5155
rect 13820 -5275 13940 -5155
rect 13985 -5275 14105 -5155
rect 14160 -5275 14280 -5155
rect 14325 -5275 14445 -5155
rect 14490 -5275 14610 -5155
rect 14655 -5275 14775 -5155
rect 14830 -5275 14950 -5155
rect 14995 -5275 15115 -5155
rect 15160 -5275 15280 -5155
rect 15325 -5275 15445 -5155
rect 15500 -5275 15620 -5155
rect 15665 -5275 15785 -5155
rect 15830 -5275 15950 -5155
rect 15995 -5275 16115 -5155
rect 16170 -5275 16290 -5155
rect 16335 -5275 16455 -5155
rect 16500 -5275 16620 -5155
rect 16665 -5275 16785 -5155
rect 16840 -5275 16960 -5155
rect 17005 -5275 17125 -5155
rect 17170 -5275 17290 -5155
rect 17335 -5275 17455 -5155
rect 17510 -5275 17630 -5155
rect 17675 -5275 17795 -5155
rect 17840 -5275 17960 -5155
rect 18005 -5275 18125 -5155
rect 18180 -5275 18300 -5155
rect 12820 -5440 12940 -5320
rect 12985 -5440 13105 -5320
rect 13150 -5440 13270 -5320
rect 13315 -5440 13435 -5320
rect 13490 -5440 13610 -5320
rect 13655 -5440 13775 -5320
rect 13820 -5440 13940 -5320
rect 13985 -5440 14105 -5320
rect 14160 -5440 14280 -5320
rect 14325 -5440 14445 -5320
rect 14490 -5440 14610 -5320
rect 14655 -5440 14775 -5320
rect 14830 -5440 14950 -5320
rect 14995 -5440 15115 -5320
rect 15160 -5440 15280 -5320
rect 15325 -5440 15445 -5320
rect 15500 -5440 15620 -5320
rect 15665 -5440 15785 -5320
rect 15830 -5440 15950 -5320
rect 15995 -5440 16115 -5320
rect 16170 -5440 16290 -5320
rect 16335 -5440 16455 -5320
rect 16500 -5440 16620 -5320
rect 16665 -5440 16785 -5320
rect 16840 -5440 16960 -5320
rect 17005 -5440 17125 -5320
rect 17170 -5440 17290 -5320
rect 17335 -5440 17455 -5320
rect 17510 -5440 17630 -5320
rect 17675 -5440 17795 -5320
rect 17840 -5440 17960 -5320
rect 18005 -5440 18125 -5320
rect 18180 -5440 18300 -5320
rect 12820 -5605 12940 -5485
rect 12985 -5605 13105 -5485
rect 13150 -5605 13270 -5485
rect 13315 -5605 13435 -5485
rect 13490 -5605 13610 -5485
rect 13655 -5605 13775 -5485
rect 13820 -5605 13940 -5485
rect 13985 -5605 14105 -5485
rect 14160 -5605 14280 -5485
rect 14325 -5605 14445 -5485
rect 14490 -5605 14610 -5485
rect 14655 -5605 14775 -5485
rect 14830 -5605 14950 -5485
rect 14995 -5605 15115 -5485
rect 15160 -5605 15280 -5485
rect 15325 -5605 15445 -5485
rect 15500 -5605 15620 -5485
rect 15665 -5605 15785 -5485
rect 15830 -5605 15950 -5485
rect 15995 -5605 16115 -5485
rect 16170 -5605 16290 -5485
rect 16335 -5605 16455 -5485
rect 16500 -5605 16620 -5485
rect 16665 -5605 16785 -5485
rect 16840 -5605 16960 -5485
rect 17005 -5605 17125 -5485
rect 17170 -5605 17290 -5485
rect 17335 -5605 17455 -5485
rect 17510 -5605 17630 -5485
rect 17675 -5605 17795 -5485
rect 17840 -5605 17960 -5485
rect 18005 -5605 18125 -5485
rect 18180 -5605 18300 -5485
rect 12820 -5770 12940 -5650
rect 12985 -5770 13105 -5650
rect 13150 -5770 13270 -5650
rect 13315 -5770 13435 -5650
rect 13490 -5770 13610 -5650
rect 13655 -5770 13775 -5650
rect 13820 -5770 13940 -5650
rect 13985 -5770 14105 -5650
rect 14160 -5770 14280 -5650
rect 14325 -5770 14445 -5650
rect 14490 -5770 14610 -5650
rect 14655 -5770 14775 -5650
rect 14830 -5770 14950 -5650
rect 14995 -5770 15115 -5650
rect 15160 -5770 15280 -5650
rect 15325 -5770 15445 -5650
rect 15500 -5770 15620 -5650
rect 15665 -5770 15785 -5650
rect 15830 -5770 15950 -5650
rect 15995 -5770 16115 -5650
rect 16170 -5770 16290 -5650
rect 16335 -5770 16455 -5650
rect 16500 -5770 16620 -5650
rect 16665 -5770 16785 -5650
rect 16840 -5770 16960 -5650
rect 17005 -5770 17125 -5650
rect 17170 -5770 17290 -5650
rect 17335 -5770 17455 -5650
rect 17510 -5770 17630 -5650
rect 17675 -5770 17795 -5650
rect 17840 -5770 17960 -5650
rect 18005 -5770 18125 -5650
rect 18180 -5770 18300 -5650
rect 12820 -5945 12940 -5825
rect 12985 -5945 13105 -5825
rect 13150 -5945 13270 -5825
rect 13315 -5945 13435 -5825
rect 13490 -5945 13610 -5825
rect 13655 -5945 13775 -5825
rect 13820 -5945 13940 -5825
rect 13985 -5945 14105 -5825
rect 14160 -5945 14280 -5825
rect 14325 -5945 14445 -5825
rect 14490 -5945 14610 -5825
rect 14655 -5945 14775 -5825
rect 14830 -5945 14950 -5825
rect 14995 -5945 15115 -5825
rect 15160 -5945 15280 -5825
rect 15325 -5945 15445 -5825
rect 15500 -5945 15620 -5825
rect 15665 -5945 15785 -5825
rect 15830 -5945 15950 -5825
rect 15995 -5945 16115 -5825
rect 16170 -5945 16290 -5825
rect 16335 -5945 16455 -5825
rect 16500 -5945 16620 -5825
rect 16665 -5945 16785 -5825
rect 16840 -5945 16960 -5825
rect 17005 -5945 17125 -5825
rect 17170 -5945 17290 -5825
rect 17335 -5945 17455 -5825
rect 17510 -5945 17630 -5825
rect 17675 -5945 17795 -5825
rect 17840 -5945 17960 -5825
rect 18005 -5945 18125 -5825
rect 18180 -5945 18300 -5825
rect 12820 -6110 12940 -5990
rect 12985 -6110 13105 -5990
rect 13150 -6110 13270 -5990
rect 13315 -6110 13435 -5990
rect 13490 -6110 13610 -5990
rect 13655 -6110 13775 -5990
rect 13820 -6110 13940 -5990
rect 13985 -6110 14105 -5990
rect 14160 -6110 14280 -5990
rect 14325 -6110 14445 -5990
rect 14490 -6110 14610 -5990
rect 14655 -6110 14775 -5990
rect 14830 -6110 14950 -5990
rect 14995 -6110 15115 -5990
rect 15160 -6110 15280 -5990
rect 15325 -6110 15445 -5990
rect 15500 -6110 15620 -5990
rect 15665 -6110 15785 -5990
rect 15830 -6110 15950 -5990
rect 15995 -6110 16115 -5990
rect 16170 -6110 16290 -5990
rect 16335 -6110 16455 -5990
rect 16500 -6110 16620 -5990
rect 16665 -6110 16785 -5990
rect 16840 -6110 16960 -5990
rect 17005 -6110 17125 -5990
rect 17170 -6110 17290 -5990
rect 17335 -6110 17455 -5990
rect 17510 -6110 17630 -5990
rect 17675 -6110 17795 -5990
rect 17840 -6110 17960 -5990
rect 18005 -6110 18125 -5990
rect 18180 -6110 18300 -5990
rect 12820 -6275 12940 -6155
rect 12985 -6275 13105 -6155
rect 13150 -6275 13270 -6155
rect 13315 -6275 13435 -6155
rect 13490 -6275 13610 -6155
rect 13655 -6275 13775 -6155
rect 13820 -6275 13940 -6155
rect 13985 -6275 14105 -6155
rect 14160 -6275 14280 -6155
rect 14325 -6275 14445 -6155
rect 14490 -6275 14610 -6155
rect 14655 -6275 14775 -6155
rect 14830 -6275 14950 -6155
rect 14995 -6275 15115 -6155
rect 15160 -6275 15280 -6155
rect 15325 -6275 15445 -6155
rect 15500 -6275 15620 -6155
rect 15665 -6275 15785 -6155
rect 15830 -6275 15950 -6155
rect 15995 -6275 16115 -6155
rect 16170 -6275 16290 -6155
rect 16335 -6275 16455 -6155
rect 16500 -6275 16620 -6155
rect 16665 -6275 16785 -6155
rect 16840 -6275 16960 -6155
rect 17005 -6275 17125 -6155
rect 17170 -6275 17290 -6155
rect 17335 -6275 17455 -6155
rect 17510 -6275 17630 -6155
rect 17675 -6275 17795 -6155
rect 17840 -6275 17960 -6155
rect 18005 -6275 18125 -6155
rect 18180 -6275 18300 -6155
rect 12820 -6440 12940 -6320
rect 12985 -6440 13105 -6320
rect 13150 -6440 13270 -6320
rect 13315 -6440 13435 -6320
rect 13490 -6440 13610 -6320
rect 13655 -6440 13775 -6320
rect 13820 -6440 13940 -6320
rect 13985 -6440 14105 -6320
rect 14160 -6440 14280 -6320
rect 14325 -6440 14445 -6320
rect 14490 -6440 14610 -6320
rect 14655 -6440 14775 -6320
rect 14830 -6440 14950 -6320
rect 14995 -6440 15115 -6320
rect 15160 -6440 15280 -6320
rect 15325 -6440 15445 -6320
rect 15500 -6440 15620 -6320
rect 15665 -6440 15785 -6320
rect 15830 -6440 15950 -6320
rect 15995 -6440 16115 -6320
rect 16170 -6440 16290 -6320
rect 16335 -6440 16455 -6320
rect 16500 -6440 16620 -6320
rect 16665 -6440 16785 -6320
rect 16840 -6440 16960 -6320
rect 17005 -6440 17125 -6320
rect 17170 -6440 17290 -6320
rect 17335 -6440 17455 -6320
rect 17510 -6440 17630 -6320
rect 17675 -6440 17795 -6320
rect 17840 -6440 17960 -6320
rect 18005 -6440 18125 -6320
rect 18180 -6440 18300 -6320
rect 12820 -6615 12940 -6495
rect 12985 -6615 13105 -6495
rect 13150 -6615 13270 -6495
rect 13315 -6615 13435 -6495
rect 13490 -6615 13610 -6495
rect 13655 -6615 13775 -6495
rect 13820 -6615 13940 -6495
rect 13985 -6615 14105 -6495
rect 14160 -6615 14280 -6495
rect 14325 -6615 14445 -6495
rect 14490 -6615 14610 -6495
rect 14655 -6615 14775 -6495
rect 14830 -6615 14950 -6495
rect 14995 -6615 15115 -6495
rect 15160 -6615 15280 -6495
rect 15325 -6615 15445 -6495
rect 15500 -6615 15620 -6495
rect 15665 -6615 15785 -6495
rect 15830 -6615 15950 -6495
rect 15995 -6615 16115 -6495
rect 16170 -6615 16290 -6495
rect 16335 -6615 16455 -6495
rect 16500 -6615 16620 -6495
rect 16665 -6615 16785 -6495
rect 16840 -6615 16960 -6495
rect 17005 -6615 17125 -6495
rect 17170 -6615 17290 -6495
rect 17335 -6615 17455 -6495
rect 17510 -6615 17630 -6495
rect 17675 -6615 17795 -6495
rect 17840 -6615 17960 -6495
rect 18005 -6615 18125 -6495
rect 18180 -6615 18300 -6495
rect 12820 -6780 12940 -6660
rect 12985 -6780 13105 -6660
rect 13150 -6780 13270 -6660
rect 13315 -6780 13435 -6660
rect 13490 -6780 13610 -6660
rect 13655 -6780 13775 -6660
rect 13820 -6780 13940 -6660
rect 13985 -6780 14105 -6660
rect 14160 -6780 14280 -6660
rect 14325 -6780 14445 -6660
rect 14490 -6780 14610 -6660
rect 14655 -6780 14775 -6660
rect 14830 -6780 14950 -6660
rect 14995 -6780 15115 -6660
rect 15160 -6780 15280 -6660
rect 15325 -6780 15445 -6660
rect 15500 -6780 15620 -6660
rect 15665 -6780 15785 -6660
rect 15830 -6780 15950 -6660
rect 15995 -6780 16115 -6660
rect 16170 -6780 16290 -6660
rect 16335 -6780 16455 -6660
rect 16500 -6780 16620 -6660
rect 16665 -6780 16785 -6660
rect 16840 -6780 16960 -6660
rect 17005 -6780 17125 -6660
rect 17170 -6780 17290 -6660
rect 17335 -6780 17455 -6660
rect 17510 -6780 17630 -6660
rect 17675 -6780 17795 -6660
rect 17840 -6780 17960 -6660
rect 18005 -6780 18125 -6660
rect 18180 -6780 18300 -6660
rect 12820 -6945 12940 -6825
rect 12985 -6945 13105 -6825
rect 13150 -6945 13270 -6825
rect 13315 -6945 13435 -6825
rect 13490 -6945 13610 -6825
rect 13655 -6945 13775 -6825
rect 13820 -6945 13940 -6825
rect 13985 -6945 14105 -6825
rect 14160 -6945 14280 -6825
rect 14325 -6945 14445 -6825
rect 14490 -6945 14610 -6825
rect 14655 -6945 14775 -6825
rect 14830 -6945 14950 -6825
rect 14995 -6945 15115 -6825
rect 15160 -6945 15280 -6825
rect 15325 -6945 15445 -6825
rect 15500 -6945 15620 -6825
rect 15665 -6945 15785 -6825
rect 15830 -6945 15950 -6825
rect 15995 -6945 16115 -6825
rect 16170 -6945 16290 -6825
rect 16335 -6945 16455 -6825
rect 16500 -6945 16620 -6825
rect 16665 -6945 16785 -6825
rect 16840 -6945 16960 -6825
rect 17005 -6945 17125 -6825
rect 17170 -6945 17290 -6825
rect 17335 -6945 17455 -6825
rect 17510 -6945 17630 -6825
rect 17675 -6945 17795 -6825
rect 17840 -6945 17960 -6825
rect 18005 -6945 18125 -6825
rect 18180 -6945 18300 -6825
rect 12820 -7110 12940 -6990
rect 12985 -7110 13105 -6990
rect 13150 -7110 13270 -6990
rect 13315 -7110 13435 -6990
rect 13490 -7110 13610 -6990
rect 13655 -7110 13775 -6990
rect 13820 -7110 13940 -6990
rect 13985 -7110 14105 -6990
rect 14160 -7110 14280 -6990
rect 14325 -7110 14445 -6990
rect 14490 -7110 14610 -6990
rect 14655 -7110 14775 -6990
rect 14830 -7110 14950 -6990
rect 14995 -7110 15115 -6990
rect 15160 -7110 15280 -6990
rect 15325 -7110 15445 -6990
rect 15500 -7110 15620 -6990
rect 15665 -7110 15785 -6990
rect 15830 -7110 15950 -6990
rect 15995 -7110 16115 -6990
rect 16170 -7110 16290 -6990
rect 16335 -7110 16455 -6990
rect 16500 -7110 16620 -6990
rect 16665 -7110 16785 -6990
rect 16840 -7110 16960 -6990
rect 17005 -7110 17125 -6990
rect 17170 -7110 17290 -6990
rect 17335 -7110 17455 -6990
rect 17510 -7110 17630 -6990
rect 17675 -7110 17795 -6990
rect 17840 -7110 17960 -6990
rect 18005 -7110 18125 -6990
rect 18180 -7110 18300 -6990
rect 12820 -7285 12940 -7165
rect 12985 -7285 13105 -7165
rect 13150 -7285 13270 -7165
rect 13315 -7285 13435 -7165
rect 13490 -7285 13610 -7165
rect 13655 -7285 13775 -7165
rect 13820 -7285 13940 -7165
rect 13985 -7285 14105 -7165
rect 14160 -7285 14280 -7165
rect 14325 -7285 14445 -7165
rect 14490 -7285 14610 -7165
rect 14655 -7285 14775 -7165
rect 14830 -7285 14950 -7165
rect 14995 -7285 15115 -7165
rect 15160 -7285 15280 -7165
rect 15325 -7285 15445 -7165
rect 15500 -7285 15620 -7165
rect 15665 -7285 15785 -7165
rect 15830 -7285 15950 -7165
rect 15995 -7285 16115 -7165
rect 16170 -7285 16290 -7165
rect 16335 -7285 16455 -7165
rect 16500 -7285 16620 -7165
rect 16665 -7285 16785 -7165
rect 16840 -7285 16960 -7165
rect 17005 -7285 17125 -7165
rect 17170 -7285 17290 -7165
rect 17335 -7285 17455 -7165
rect 17510 -7285 17630 -7165
rect 17675 -7285 17795 -7165
rect 17840 -7285 17960 -7165
rect 18005 -7285 18125 -7165
rect 18180 -7285 18300 -7165
rect 12820 -7450 12940 -7330
rect 12985 -7450 13105 -7330
rect 13150 -7450 13270 -7330
rect 13315 -7450 13435 -7330
rect 13490 -7450 13610 -7330
rect 13655 -7450 13775 -7330
rect 13820 -7450 13940 -7330
rect 13985 -7450 14105 -7330
rect 14160 -7450 14280 -7330
rect 14325 -7450 14445 -7330
rect 14490 -7450 14610 -7330
rect 14655 -7450 14775 -7330
rect 14830 -7450 14950 -7330
rect 14995 -7450 15115 -7330
rect 15160 -7450 15280 -7330
rect 15325 -7450 15445 -7330
rect 15500 -7450 15620 -7330
rect 15665 -7450 15785 -7330
rect 15830 -7450 15950 -7330
rect 15995 -7450 16115 -7330
rect 16170 -7450 16290 -7330
rect 16335 -7450 16455 -7330
rect 16500 -7450 16620 -7330
rect 16665 -7450 16785 -7330
rect 16840 -7450 16960 -7330
rect 17005 -7450 17125 -7330
rect 17170 -7450 17290 -7330
rect 17335 -7450 17455 -7330
rect 17510 -7450 17630 -7330
rect 17675 -7450 17795 -7330
rect 17840 -7450 17960 -7330
rect 18005 -7450 18125 -7330
rect 18180 -7450 18300 -7330
rect 12820 -7615 12940 -7495
rect 12985 -7615 13105 -7495
rect 13150 -7615 13270 -7495
rect 13315 -7615 13435 -7495
rect 13490 -7615 13610 -7495
rect 13655 -7615 13775 -7495
rect 13820 -7615 13940 -7495
rect 13985 -7615 14105 -7495
rect 14160 -7615 14280 -7495
rect 14325 -7615 14445 -7495
rect 14490 -7615 14610 -7495
rect 14655 -7615 14775 -7495
rect 14830 -7615 14950 -7495
rect 14995 -7615 15115 -7495
rect 15160 -7615 15280 -7495
rect 15325 -7615 15445 -7495
rect 15500 -7615 15620 -7495
rect 15665 -7615 15785 -7495
rect 15830 -7615 15950 -7495
rect 15995 -7615 16115 -7495
rect 16170 -7615 16290 -7495
rect 16335 -7615 16455 -7495
rect 16500 -7615 16620 -7495
rect 16665 -7615 16785 -7495
rect 16840 -7615 16960 -7495
rect 17005 -7615 17125 -7495
rect 17170 -7615 17290 -7495
rect 17335 -7615 17455 -7495
rect 17510 -7615 17630 -7495
rect 17675 -7615 17795 -7495
rect 17840 -7615 17960 -7495
rect 18005 -7615 18125 -7495
rect 18180 -7615 18300 -7495
rect 12820 -7780 12940 -7660
rect 12985 -7780 13105 -7660
rect 13150 -7780 13270 -7660
rect 13315 -7780 13435 -7660
rect 13490 -7780 13610 -7660
rect 13655 -7780 13775 -7660
rect 13820 -7780 13940 -7660
rect 13985 -7780 14105 -7660
rect 14160 -7780 14280 -7660
rect 14325 -7780 14445 -7660
rect 14490 -7780 14610 -7660
rect 14655 -7780 14775 -7660
rect 14830 -7780 14950 -7660
rect 14995 -7780 15115 -7660
rect 15160 -7780 15280 -7660
rect 15325 -7780 15445 -7660
rect 15500 -7780 15620 -7660
rect 15665 -7780 15785 -7660
rect 15830 -7780 15950 -7660
rect 15995 -7780 16115 -7660
rect 16170 -7780 16290 -7660
rect 16335 -7780 16455 -7660
rect 16500 -7780 16620 -7660
rect 16665 -7780 16785 -7660
rect 16840 -7780 16960 -7660
rect 17005 -7780 17125 -7660
rect 17170 -7780 17290 -7660
rect 17335 -7780 17455 -7660
rect 17510 -7780 17630 -7660
rect 17675 -7780 17795 -7660
rect 17840 -7780 17960 -7660
rect 18005 -7780 18125 -7660
rect 18180 -7780 18300 -7660
rect 12820 -7955 12940 -7835
rect 12985 -7955 13105 -7835
rect 13150 -7955 13270 -7835
rect 13315 -7955 13435 -7835
rect 13490 -7955 13610 -7835
rect 13655 -7955 13775 -7835
rect 13820 -7955 13940 -7835
rect 13985 -7955 14105 -7835
rect 14160 -7955 14280 -7835
rect 14325 -7955 14445 -7835
rect 14490 -7955 14610 -7835
rect 14655 -7955 14775 -7835
rect 14830 -7955 14950 -7835
rect 14995 -7955 15115 -7835
rect 15160 -7955 15280 -7835
rect 15325 -7955 15445 -7835
rect 15500 -7955 15620 -7835
rect 15665 -7955 15785 -7835
rect 15830 -7955 15950 -7835
rect 15995 -7955 16115 -7835
rect 16170 -7955 16290 -7835
rect 16335 -7955 16455 -7835
rect 16500 -7955 16620 -7835
rect 16665 -7955 16785 -7835
rect 16840 -7955 16960 -7835
rect 17005 -7955 17125 -7835
rect 17170 -7955 17290 -7835
rect 17335 -7955 17455 -7835
rect 17510 -7955 17630 -7835
rect 17675 -7955 17795 -7835
rect 17840 -7955 17960 -7835
rect 18005 -7955 18125 -7835
rect 18180 -7955 18300 -7835
rect 12820 -8120 12940 -8000
rect 12985 -8120 13105 -8000
rect 13150 -8120 13270 -8000
rect 13315 -8120 13435 -8000
rect 13490 -8120 13610 -8000
rect 13655 -8120 13775 -8000
rect 13820 -8120 13940 -8000
rect 13985 -8120 14105 -8000
rect 14160 -8120 14280 -8000
rect 14325 -8120 14445 -8000
rect 14490 -8120 14610 -8000
rect 14655 -8120 14775 -8000
rect 14830 -8120 14950 -8000
rect 14995 -8120 15115 -8000
rect 15160 -8120 15280 -8000
rect 15325 -8120 15445 -8000
rect 15500 -8120 15620 -8000
rect 15665 -8120 15785 -8000
rect 15830 -8120 15950 -8000
rect 15995 -8120 16115 -8000
rect 16170 -8120 16290 -8000
rect 16335 -8120 16455 -8000
rect 16500 -8120 16620 -8000
rect 16665 -8120 16785 -8000
rect 16840 -8120 16960 -8000
rect 17005 -8120 17125 -8000
rect 17170 -8120 17290 -8000
rect 17335 -8120 17455 -8000
rect 17510 -8120 17630 -8000
rect 17675 -8120 17795 -8000
rect 17840 -8120 17960 -8000
rect 18005 -8120 18125 -8000
rect 18180 -8120 18300 -8000
rect 12820 -8285 12940 -8165
rect 12985 -8285 13105 -8165
rect 13150 -8285 13270 -8165
rect 13315 -8285 13435 -8165
rect 13490 -8285 13610 -8165
rect 13655 -8285 13775 -8165
rect 13820 -8285 13940 -8165
rect 13985 -8285 14105 -8165
rect 14160 -8285 14280 -8165
rect 14325 -8285 14445 -8165
rect 14490 -8285 14610 -8165
rect 14655 -8285 14775 -8165
rect 14830 -8285 14950 -8165
rect 14995 -8285 15115 -8165
rect 15160 -8285 15280 -8165
rect 15325 -8285 15445 -8165
rect 15500 -8285 15620 -8165
rect 15665 -8285 15785 -8165
rect 15830 -8285 15950 -8165
rect 15995 -8285 16115 -8165
rect 16170 -8285 16290 -8165
rect 16335 -8285 16455 -8165
rect 16500 -8285 16620 -8165
rect 16665 -8285 16785 -8165
rect 16840 -8285 16960 -8165
rect 17005 -8285 17125 -8165
rect 17170 -8285 17290 -8165
rect 17335 -8285 17455 -8165
rect 17510 -8285 17630 -8165
rect 17675 -8285 17795 -8165
rect 17840 -8285 17960 -8165
rect 18005 -8285 18125 -8165
rect 18180 -8285 18300 -8165
rect 12820 -8450 12940 -8330
rect 12985 -8450 13105 -8330
rect 13150 -8450 13270 -8330
rect 13315 -8450 13435 -8330
rect 13490 -8450 13610 -8330
rect 13655 -8450 13775 -8330
rect 13820 -8450 13940 -8330
rect 13985 -8450 14105 -8330
rect 14160 -8450 14280 -8330
rect 14325 -8450 14445 -8330
rect 14490 -8450 14610 -8330
rect 14655 -8450 14775 -8330
rect 14830 -8450 14950 -8330
rect 14995 -8450 15115 -8330
rect 15160 -8450 15280 -8330
rect 15325 -8450 15445 -8330
rect 15500 -8450 15620 -8330
rect 15665 -8450 15785 -8330
rect 15830 -8450 15950 -8330
rect 15995 -8450 16115 -8330
rect 16170 -8450 16290 -8330
rect 16335 -8450 16455 -8330
rect 16500 -8450 16620 -8330
rect 16665 -8450 16785 -8330
rect 16840 -8450 16960 -8330
rect 17005 -8450 17125 -8330
rect 17170 -8450 17290 -8330
rect 17335 -8450 17455 -8330
rect 17510 -8450 17630 -8330
rect 17675 -8450 17795 -8330
rect 17840 -8450 17960 -8330
rect 18005 -8450 18125 -8330
rect 18180 -8450 18300 -8330
rect 12820 -8625 12940 -8505
rect 12985 -8625 13105 -8505
rect 13150 -8625 13270 -8505
rect 13315 -8625 13435 -8505
rect 13490 -8625 13610 -8505
rect 13655 -8625 13775 -8505
rect 13820 -8625 13940 -8505
rect 13985 -8625 14105 -8505
rect 14160 -8625 14280 -8505
rect 14325 -8625 14445 -8505
rect 14490 -8625 14610 -8505
rect 14655 -8625 14775 -8505
rect 14830 -8625 14950 -8505
rect 14995 -8625 15115 -8505
rect 15160 -8625 15280 -8505
rect 15325 -8625 15445 -8505
rect 15500 -8625 15620 -8505
rect 15665 -8625 15785 -8505
rect 15830 -8625 15950 -8505
rect 15995 -8625 16115 -8505
rect 16170 -8625 16290 -8505
rect 16335 -8625 16455 -8505
rect 16500 -8625 16620 -8505
rect 16665 -8625 16785 -8505
rect 16840 -8625 16960 -8505
rect 17005 -8625 17125 -8505
rect 17170 -8625 17290 -8505
rect 17335 -8625 17455 -8505
rect 17510 -8625 17630 -8505
rect 17675 -8625 17795 -8505
rect 17840 -8625 17960 -8505
rect 18005 -8625 18125 -8505
rect 18180 -8625 18300 -8505
rect 12820 -8790 12940 -8670
rect 12985 -8790 13105 -8670
rect 13150 -8790 13270 -8670
rect 13315 -8790 13435 -8670
rect 13490 -8790 13610 -8670
rect 13655 -8790 13775 -8670
rect 13820 -8790 13940 -8670
rect 13985 -8790 14105 -8670
rect 14160 -8790 14280 -8670
rect 14325 -8790 14445 -8670
rect 14490 -8790 14610 -8670
rect 14655 -8790 14775 -8670
rect 14830 -8790 14950 -8670
rect 14995 -8790 15115 -8670
rect 15160 -8790 15280 -8670
rect 15325 -8790 15445 -8670
rect 15500 -8790 15620 -8670
rect 15665 -8790 15785 -8670
rect 15830 -8790 15950 -8670
rect 15995 -8790 16115 -8670
rect 16170 -8790 16290 -8670
rect 16335 -8790 16455 -8670
rect 16500 -8790 16620 -8670
rect 16665 -8790 16785 -8670
rect 16840 -8790 16960 -8670
rect 17005 -8790 17125 -8670
rect 17170 -8790 17290 -8670
rect 17335 -8790 17455 -8670
rect 17510 -8790 17630 -8670
rect 17675 -8790 17795 -8670
rect 17840 -8790 17960 -8670
rect 18005 -8790 18125 -8670
rect 18180 -8790 18300 -8670
rect 12820 -8955 12940 -8835
rect 12985 -8955 13105 -8835
rect 13150 -8955 13270 -8835
rect 13315 -8955 13435 -8835
rect 13490 -8955 13610 -8835
rect 13655 -8955 13775 -8835
rect 13820 -8955 13940 -8835
rect 13985 -8955 14105 -8835
rect 14160 -8955 14280 -8835
rect 14325 -8955 14445 -8835
rect 14490 -8955 14610 -8835
rect 14655 -8955 14775 -8835
rect 14830 -8955 14950 -8835
rect 14995 -8955 15115 -8835
rect 15160 -8955 15280 -8835
rect 15325 -8955 15445 -8835
rect 15500 -8955 15620 -8835
rect 15665 -8955 15785 -8835
rect 15830 -8955 15950 -8835
rect 15995 -8955 16115 -8835
rect 16170 -8955 16290 -8835
rect 16335 -8955 16455 -8835
rect 16500 -8955 16620 -8835
rect 16665 -8955 16785 -8835
rect 16840 -8955 16960 -8835
rect 17005 -8955 17125 -8835
rect 17170 -8955 17290 -8835
rect 17335 -8955 17455 -8835
rect 17510 -8955 17630 -8835
rect 17675 -8955 17795 -8835
rect 17840 -8955 17960 -8835
rect 18005 -8955 18125 -8835
rect 18180 -8955 18300 -8835
rect 12820 -9120 12940 -9000
rect 12985 -9120 13105 -9000
rect 13150 -9120 13270 -9000
rect 13315 -9120 13435 -9000
rect 13490 -9120 13610 -9000
rect 13655 -9120 13775 -9000
rect 13820 -9120 13940 -9000
rect 13985 -9120 14105 -9000
rect 14160 -9120 14280 -9000
rect 14325 -9120 14445 -9000
rect 14490 -9120 14610 -9000
rect 14655 -9120 14775 -9000
rect 14830 -9120 14950 -9000
rect 14995 -9120 15115 -9000
rect 15160 -9120 15280 -9000
rect 15325 -9120 15445 -9000
rect 15500 -9120 15620 -9000
rect 15665 -9120 15785 -9000
rect 15830 -9120 15950 -9000
rect 15995 -9120 16115 -9000
rect 16170 -9120 16290 -9000
rect 16335 -9120 16455 -9000
rect 16500 -9120 16620 -9000
rect 16665 -9120 16785 -9000
rect 16840 -9120 16960 -9000
rect 17005 -9120 17125 -9000
rect 17170 -9120 17290 -9000
rect 17335 -9120 17455 -9000
rect 17510 -9120 17630 -9000
rect 17675 -9120 17795 -9000
rect 17840 -9120 17960 -9000
rect 18005 -9120 18125 -9000
rect 18180 -9120 18300 -9000
rect 12820 -9295 12940 -9175
rect 12985 -9295 13105 -9175
rect 13150 -9295 13270 -9175
rect 13315 -9295 13435 -9175
rect 13490 -9295 13610 -9175
rect 13655 -9295 13775 -9175
rect 13820 -9295 13940 -9175
rect 13985 -9295 14105 -9175
rect 14160 -9295 14280 -9175
rect 14325 -9295 14445 -9175
rect 14490 -9295 14610 -9175
rect 14655 -9295 14775 -9175
rect 14830 -9295 14950 -9175
rect 14995 -9295 15115 -9175
rect 15160 -9295 15280 -9175
rect 15325 -9295 15445 -9175
rect 15500 -9295 15620 -9175
rect 15665 -9295 15785 -9175
rect 15830 -9295 15950 -9175
rect 15995 -9295 16115 -9175
rect 16170 -9295 16290 -9175
rect 16335 -9295 16455 -9175
rect 16500 -9295 16620 -9175
rect 16665 -9295 16785 -9175
rect 16840 -9295 16960 -9175
rect 17005 -9295 17125 -9175
rect 17170 -9295 17290 -9175
rect 17335 -9295 17455 -9175
rect 17510 -9295 17630 -9175
rect 17675 -9295 17795 -9175
rect 17840 -9295 17960 -9175
rect 18005 -9295 18125 -9175
rect 18180 -9295 18300 -9175
rect 12820 -9460 12940 -9340
rect 12985 -9460 13105 -9340
rect 13150 -9460 13270 -9340
rect 13315 -9460 13435 -9340
rect 13490 -9460 13610 -9340
rect 13655 -9460 13775 -9340
rect 13820 -9460 13940 -9340
rect 13985 -9460 14105 -9340
rect 14160 -9460 14280 -9340
rect 14325 -9460 14445 -9340
rect 14490 -9460 14610 -9340
rect 14655 -9460 14775 -9340
rect 14830 -9460 14950 -9340
rect 14995 -9460 15115 -9340
rect 15160 -9460 15280 -9340
rect 15325 -9460 15445 -9340
rect 15500 -9460 15620 -9340
rect 15665 -9460 15785 -9340
rect 15830 -9460 15950 -9340
rect 15995 -9460 16115 -9340
rect 16170 -9460 16290 -9340
rect 16335 -9460 16455 -9340
rect 16500 -9460 16620 -9340
rect 16665 -9460 16785 -9340
rect 16840 -9460 16960 -9340
rect 17005 -9460 17125 -9340
rect 17170 -9460 17290 -9340
rect 17335 -9460 17455 -9340
rect 17510 -9460 17630 -9340
rect 17675 -9460 17795 -9340
rect 17840 -9460 17960 -9340
rect 18005 -9460 18125 -9340
rect 18180 -9460 18300 -9340
rect 12820 -9625 12940 -9505
rect 12985 -9625 13105 -9505
rect 13150 -9625 13270 -9505
rect 13315 -9625 13435 -9505
rect 13490 -9625 13610 -9505
rect 13655 -9625 13775 -9505
rect 13820 -9625 13940 -9505
rect 13985 -9625 14105 -9505
rect 14160 -9625 14280 -9505
rect 14325 -9625 14445 -9505
rect 14490 -9625 14610 -9505
rect 14655 -9625 14775 -9505
rect 14830 -9625 14950 -9505
rect 14995 -9625 15115 -9505
rect 15160 -9625 15280 -9505
rect 15325 -9625 15445 -9505
rect 15500 -9625 15620 -9505
rect 15665 -9625 15785 -9505
rect 15830 -9625 15950 -9505
rect 15995 -9625 16115 -9505
rect 16170 -9625 16290 -9505
rect 16335 -9625 16455 -9505
rect 16500 -9625 16620 -9505
rect 16665 -9625 16785 -9505
rect 16840 -9625 16960 -9505
rect 17005 -9625 17125 -9505
rect 17170 -9625 17290 -9505
rect 17335 -9625 17455 -9505
rect 17510 -9625 17630 -9505
rect 17675 -9625 17795 -9505
rect 17840 -9625 17960 -9505
rect 18005 -9625 18125 -9505
rect 18180 -9625 18300 -9505
rect 12820 -9790 12940 -9670
rect 12985 -9790 13105 -9670
rect 13150 -9790 13270 -9670
rect 13315 -9790 13435 -9670
rect 13490 -9790 13610 -9670
rect 13655 -9790 13775 -9670
rect 13820 -9790 13940 -9670
rect 13985 -9790 14105 -9670
rect 14160 -9790 14280 -9670
rect 14325 -9790 14445 -9670
rect 14490 -9790 14610 -9670
rect 14655 -9790 14775 -9670
rect 14830 -9790 14950 -9670
rect 14995 -9790 15115 -9670
rect 15160 -9790 15280 -9670
rect 15325 -9790 15445 -9670
rect 15500 -9790 15620 -9670
rect 15665 -9790 15785 -9670
rect 15830 -9790 15950 -9670
rect 15995 -9790 16115 -9670
rect 16170 -9790 16290 -9670
rect 16335 -9790 16455 -9670
rect 16500 -9790 16620 -9670
rect 16665 -9790 16785 -9670
rect 16840 -9790 16960 -9670
rect 17005 -9790 17125 -9670
rect 17170 -9790 17290 -9670
rect 17335 -9790 17455 -9670
rect 17510 -9790 17630 -9670
rect 17675 -9790 17795 -9670
rect 17840 -9790 17960 -9670
rect 18005 -9790 18125 -9670
rect 18180 -9790 18300 -9670
rect 18510 -4430 18630 -4310
rect 18675 -4430 18795 -4310
rect 18840 -4430 18960 -4310
rect 19005 -4430 19125 -4310
rect 19180 -4430 19300 -4310
rect 19345 -4430 19465 -4310
rect 19510 -4430 19630 -4310
rect 19675 -4430 19795 -4310
rect 19850 -4430 19970 -4310
rect 20015 -4430 20135 -4310
rect 20180 -4430 20300 -4310
rect 20345 -4430 20465 -4310
rect 20520 -4430 20640 -4310
rect 20685 -4430 20805 -4310
rect 20850 -4430 20970 -4310
rect 21015 -4430 21135 -4310
rect 21190 -4430 21310 -4310
rect 21355 -4430 21475 -4310
rect 21520 -4430 21640 -4310
rect 21685 -4430 21805 -4310
rect 21860 -4430 21980 -4310
rect 22025 -4430 22145 -4310
rect 22190 -4430 22310 -4310
rect 22355 -4430 22475 -4310
rect 22530 -4430 22650 -4310
rect 22695 -4430 22815 -4310
rect 22860 -4430 22980 -4310
rect 23025 -4430 23145 -4310
rect 23200 -4430 23320 -4310
rect 23365 -4430 23485 -4310
rect 23530 -4430 23650 -4310
rect 23695 -4430 23815 -4310
rect 23870 -4430 23990 -4310
rect 18510 -4605 18630 -4485
rect 18675 -4605 18795 -4485
rect 18840 -4605 18960 -4485
rect 19005 -4605 19125 -4485
rect 19180 -4605 19300 -4485
rect 19345 -4605 19465 -4485
rect 19510 -4605 19630 -4485
rect 19675 -4605 19795 -4485
rect 19850 -4605 19970 -4485
rect 20015 -4605 20135 -4485
rect 20180 -4605 20300 -4485
rect 20345 -4605 20465 -4485
rect 20520 -4605 20640 -4485
rect 20685 -4605 20805 -4485
rect 20850 -4605 20970 -4485
rect 21015 -4605 21135 -4485
rect 21190 -4605 21310 -4485
rect 21355 -4605 21475 -4485
rect 21520 -4605 21640 -4485
rect 21685 -4605 21805 -4485
rect 21860 -4605 21980 -4485
rect 22025 -4605 22145 -4485
rect 22190 -4605 22310 -4485
rect 22355 -4605 22475 -4485
rect 22530 -4605 22650 -4485
rect 22695 -4605 22815 -4485
rect 22860 -4605 22980 -4485
rect 23025 -4605 23145 -4485
rect 23200 -4605 23320 -4485
rect 23365 -4605 23485 -4485
rect 23530 -4605 23650 -4485
rect 23695 -4605 23815 -4485
rect 23870 -4605 23990 -4485
rect 18510 -4770 18630 -4650
rect 18675 -4770 18795 -4650
rect 18840 -4770 18960 -4650
rect 19005 -4770 19125 -4650
rect 19180 -4770 19300 -4650
rect 19345 -4770 19465 -4650
rect 19510 -4770 19630 -4650
rect 19675 -4770 19795 -4650
rect 19850 -4770 19970 -4650
rect 20015 -4770 20135 -4650
rect 20180 -4770 20300 -4650
rect 20345 -4770 20465 -4650
rect 20520 -4770 20640 -4650
rect 20685 -4770 20805 -4650
rect 20850 -4770 20970 -4650
rect 21015 -4770 21135 -4650
rect 21190 -4770 21310 -4650
rect 21355 -4770 21475 -4650
rect 21520 -4770 21640 -4650
rect 21685 -4770 21805 -4650
rect 21860 -4770 21980 -4650
rect 22025 -4770 22145 -4650
rect 22190 -4770 22310 -4650
rect 22355 -4770 22475 -4650
rect 22530 -4770 22650 -4650
rect 22695 -4770 22815 -4650
rect 22860 -4770 22980 -4650
rect 23025 -4770 23145 -4650
rect 23200 -4770 23320 -4650
rect 23365 -4770 23485 -4650
rect 23530 -4770 23650 -4650
rect 23695 -4770 23815 -4650
rect 23870 -4770 23990 -4650
rect 18510 -4935 18630 -4815
rect 18675 -4935 18795 -4815
rect 18840 -4935 18960 -4815
rect 19005 -4935 19125 -4815
rect 19180 -4935 19300 -4815
rect 19345 -4935 19465 -4815
rect 19510 -4935 19630 -4815
rect 19675 -4935 19795 -4815
rect 19850 -4935 19970 -4815
rect 20015 -4935 20135 -4815
rect 20180 -4935 20300 -4815
rect 20345 -4935 20465 -4815
rect 20520 -4935 20640 -4815
rect 20685 -4935 20805 -4815
rect 20850 -4935 20970 -4815
rect 21015 -4935 21135 -4815
rect 21190 -4935 21310 -4815
rect 21355 -4935 21475 -4815
rect 21520 -4935 21640 -4815
rect 21685 -4935 21805 -4815
rect 21860 -4935 21980 -4815
rect 22025 -4935 22145 -4815
rect 22190 -4935 22310 -4815
rect 22355 -4935 22475 -4815
rect 22530 -4935 22650 -4815
rect 22695 -4935 22815 -4815
rect 22860 -4935 22980 -4815
rect 23025 -4935 23145 -4815
rect 23200 -4935 23320 -4815
rect 23365 -4935 23485 -4815
rect 23530 -4935 23650 -4815
rect 23695 -4935 23815 -4815
rect 23870 -4935 23990 -4815
rect 18510 -5100 18630 -4980
rect 18675 -5100 18795 -4980
rect 18840 -5100 18960 -4980
rect 19005 -5100 19125 -4980
rect 19180 -5100 19300 -4980
rect 19345 -5100 19465 -4980
rect 19510 -5100 19630 -4980
rect 19675 -5100 19795 -4980
rect 19850 -5100 19970 -4980
rect 20015 -5100 20135 -4980
rect 20180 -5100 20300 -4980
rect 20345 -5100 20465 -4980
rect 20520 -5100 20640 -4980
rect 20685 -5100 20805 -4980
rect 20850 -5100 20970 -4980
rect 21015 -5100 21135 -4980
rect 21190 -5100 21310 -4980
rect 21355 -5100 21475 -4980
rect 21520 -5100 21640 -4980
rect 21685 -5100 21805 -4980
rect 21860 -5100 21980 -4980
rect 22025 -5100 22145 -4980
rect 22190 -5100 22310 -4980
rect 22355 -5100 22475 -4980
rect 22530 -5100 22650 -4980
rect 22695 -5100 22815 -4980
rect 22860 -5100 22980 -4980
rect 23025 -5100 23145 -4980
rect 23200 -5100 23320 -4980
rect 23365 -5100 23485 -4980
rect 23530 -5100 23650 -4980
rect 23695 -5100 23815 -4980
rect 23870 -5100 23990 -4980
rect 18510 -5275 18630 -5155
rect 18675 -5275 18795 -5155
rect 18840 -5275 18960 -5155
rect 19005 -5275 19125 -5155
rect 19180 -5275 19300 -5155
rect 19345 -5275 19465 -5155
rect 19510 -5275 19630 -5155
rect 19675 -5275 19795 -5155
rect 19850 -5275 19970 -5155
rect 20015 -5275 20135 -5155
rect 20180 -5275 20300 -5155
rect 20345 -5275 20465 -5155
rect 20520 -5275 20640 -5155
rect 20685 -5275 20805 -5155
rect 20850 -5275 20970 -5155
rect 21015 -5275 21135 -5155
rect 21190 -5275 21310 -5155
rect 21355 -5275 21475 -5155
rect 21520 -5275 21640 -5155
rect 21685 -5275 21805 -5155
rect 21860 -5275 21980 -5155
rect 22025 -5275 22145 -5155
rect 22190 -5275 22310 -5155
rect 22355 -5275 22475 -5155
rect 22530 -5275 22650 -5155
rect 22695 -5275 22815 -5155
rect 22860 -5275 22980 -5155
rect 23025 -5275 23145 -5155
rect 23200 -5275 23320 -5155
rect 23365 -5275 23485 -5155
rect 23530 -5275 23650 -5155
rect 23695 -5275 23815 -5155
rect 23870 -5275 23990 -5155
rect 18510 -5440 18630 -5320
rect 18675 -5440 18795 -5320
rect 18840 -5440 18960 -5320
rect 19005 -5440 19125 -5320
rect 19180 -5440 19300 -5320
rect 19345 -5440 19465 -5320
rect 19510 -5440 19630 -5320
rect 19675 -5440 19795 -5320
rect 19850 -5440 19970 -5320
rect 20015 -5440 20135 -5320
rect 20180 -5440 20300 -5320
rect 20345 -5440 20465 -5320
rect 20520 -5440 20640 -5320
rect 20685 -5440 20805 -5320
rect 20850 -5440 20970 -5320
rect 21015 -5440 21135 -5320
rect 21190 -5440 21310 -5320
rect 21355 -5440 21475 -5320
rect 21520 -5440 21640 -5320
rect 21685 -5440 21805 -5320
rect 21860 -5440 21980 -5320
rect 22025 -5440 22145 -5320
rect 22190 -5440 22310 -5320
rect 22355 -5440 22475 -5320
rect 22530 -5440 22650 -5320
rect 22695 -5440 22815 -5320
rect 22860 -5440 22980 -5320
rect 23025 -5440 23145 -5320
rect 23200 -5440 23320 -5320
rect 23365 -5440 23485 -5320
rect 23530 -5440 23650 -5320
rect 23695 -5440 23815 -5320
rect 23870 -5440 23990 -5320
rect 18510 -5605 18630 -5485
rect 18675 -5605 18795 -5485
rect 18840 -5605 18960 -5485
rect 19005 -5605 19125 -5485
rect 19180 -5605 19300 -5485
rect 19345 -5605 19465 -5485
rect 19510 -5605 19630 -5485
rect 19675 -5605 19795 -5485
rect 19850 -5605 19970 -5485
rect 20015 -5605 20135 -5485
rect 20180 -5605 20300 -5485
rect 20345 -5605 20465 -5485
rect 20520 -5605 20640 -5485
rect 20685 -5605 20805 -5485
rect 20850 -5605 20970 -5485
rect 21015 -5605 21135 -5485
rect 21190 -5605 21310 -5485
rect 21355 -5605 21475 -5485
rect 21520 -5605 21640 -5485
rect 21685 -5605 21805 -5485
rect 21860 -5605 21980 -5485
rect 22025 -5605 22145 -5485
rect 22190 -5605 22310 -5485
rect 22355 -5605 22475 -5485
rect 22530 -5605 22650 -5485
rect 22695 -5605 22815 -5485
rect 22860 -5605 22980 -5485
rect 23025 -5605 23145 -5485
rect 23200 -5605 23320 -5485
rect 23365 -5605 23485 -5485
rect 23530 -5605 23650 -5485
rect 23695 -5605 23815 -5485
rect 23870 -5605 23990 -5485
rect 18510 -5770 18630 -5650
rect 18675 -5770 18795 -5650
rect 18840 -5770 18960 -5650
rect 19005 -5770 19125 -5650
rect 19180 -5770 19300 -5650
rect 19345 -5770 19465 -5650
rect 19510 -5770 19630 -5650
rect 19675 -5770 19795 -5650
rect 19850 -5770 19970 -5650
rect 20015 -5770 20135 -5650
rect 20180 -5770 20300 -5650
rect 20345 -5770 20465 -5650
rect 20520 -5770 20640 -5650
rect 20685 -5770 20805 -5650
rect 20850 -5770 20970 -5650
rect 21015 -5770 21135 -5650
rect 21190 -5770 21310 -5650
rect 21355 -5770 21475 -5650
rect 21520 -5770 21640 -5650
rect 21685 -5770 21805 -5650
rect 21860 -5770 21980 -5650
rect 22025 -5770 22145 -5650
rect 22190 -5770 22310 -5650
rect 22355 -5770 22475 -5650
rect 22530 -5770 22650 -5650
rect 22695 -5770 22815 -5650
rect 22860 -5770 22980 -5650
rect 23025 -5770 23145 -5650
rect 23200 -5770 23320 -5650
rect 23365 -5770 23485 -5650
rect 23530 -5770 23650 -5650
rect 23695 -5770 23815 -5650
rect 23870 -5770 23990 -5650
rect 18510 -5945 18630 -5825
rect 18675 -5945 18795 -5825
rect 18840 -5945 18960 -5825
rect 19005 -5945 19125 -5825
rect 19180 -5945 19300 -5825
rect 19345 -5945 19465 -5825
rect 19510 -5945 19630 -5825
rect 19675 -5945 19795 -5825
rect 19850 -5945 19970 -5825
rect 20015 -5945 20135 -5825
rect 20180 -5945 20300 -5825
rect 20345 -5945 20465 -5825
rect 20520 -5945 20640 -5825
rect 20685 -5945 20805 -5825
rect 20850 -5945 20970 -5825
rect 21015 -5945 21135 -5825
rect 21190 -5945 21310 -5825
rect 21355 -5945 21475 -5825
rect 21520 -5945 21640 -5825
rect 21685 -5945 21805 -5825
rect 21860 -5945 21980 -5825
rect 22025 -5945 22145 -5825
rect 22190 -5945 22310 -5825
rect 22355 -5945 22475 -5825
rect 22530 -5945 22650 -5825
rect 22695 -5945 22815 -5825
rect 22860 -5945 22980 -5825
rect 23025 -5945 23145 -5825
rect 23200 -5945 23320 -5825
rect 23365 -5945 23485 -5825
rect 23530 -5945 23650 -5825
rect 23695 -5945 23815 -5825
rect 23870 -5945 23990 -5825
rect 18510 -6110 18630 -5990
rect 18675 -6110 18795 -5990
rect 18840 -6110 18960 -5990
rect 19005 -6110 19125 -5990
rect 19180 -6110 19300 -5990
rect 19345 -6110 19465 -5990
rect 19510 -6110 19630 -5990
rect 19675 -6110 19795 -5990
rect 19850 -6110 19970 -5990
rect 20015 -6110 20135 -5990
rect 20180 -6110 20300 -5990
rect 20345 -6110 20465 -5990
rect 20520 -6110 20640 -5990
rect 20685 -6110 20805 -5990
rect 20850 -6110 20970 -5990
rect 21015 -6110 21135 -5990
rect 21190 -6110 21310 -5990
rect 21355 -6110 21475 -5990
rect 21520 -6110 21640 -5990
rect 21685 -6110 21805 -5990
rect 21860 -6110 21980 -5990
rect 22025 -6110 22145 -5990
rect 22190 -6110 22310 -5990
rect 22355 -6110 22475 -5990
rect 22530 -6110 22650 -5990
rect 22695 -6110 22815 -5990
rect 22860 -6110 22980 -5990
rect 23025 -6110 23145 -5990
rect 23200 -6110 23320 -5990
rect 23365 -6110 23485 -5990
rect 23530 -6110 23650 -5990
rect 23695 -6110 23815 -5990
rect 23870 -6110 23990 -5990
rect 18510 -6275 18630 -6155
rect 18675 -6275 18795 -6155
rect 18840 -6275 18960 -6155
rect 19005 -6275 19125 -6155
rect 19180 -6275 19300 -6155
rect 19345 -6275 19465 -6155
rect 19510 -6275 19630 -6155
rect 19675 -6275 19795 -6155
rect 19850 -6275 19970 -6155
rect 20015 -6275 20135 -6155
rect 20180 -6275 20300 -6155
rect 20345 -6275 20465 -6155
rect 20520 -6275 20640 -6155
rect 20685 -6275 20805 -6155
rect 20850 -6275 20970 -6155
rect 21015 -6275 21135 -6155
rect 21190 -6275 21310 -6155
rect 21355 -6275 21475 -6155
rect 21520 -6275 21640 -6155
rect 21685 -6275 21805 -6155
rect 21860 -6275 21980 -6155
rect 22025 -6275 22145 -6155
rect 22190 -6275 22310 -6155
rect 22355 -6275 22475 -6155
rect 22530 -6275 22650 -6155
rect 22695 -6275 22815 -6155
rect 22860 -6275 22980 -6155
rect 23025 -6275 23145 -6155
rect 23200 -6275 23320 -6155
rect 23365 -6275 23485 -6155
rect 23530 -6275 23650 -6155
rect 23695 -6275 23815 -6155
rect 23870 -6275 23990 -6155
rect 18510 -6440 18630 -6320
rect 18675 -6440 18795 -6320
rect 18840 -6440 18960 -6320
rect 19005 -6440 19125 -6320
rect 19180 -6440 19300 -6320
rect 19345 -6440 19465 -6320
rect 19510 -6440 19630 -6320
rect 19675 -6440 19795 -6320
rect 19850 -6440 19970 -6320
rect 20015 -6440 20135 -6320
rect 20180 -6440 20300 -6320
rect 20345 -6440 20465 -6320
rect 20520 -6440 20640 -6320
rect 20685 -6440 20805 -6320
rect 20850 -6440 20970 -6320
rect 21015 -6440 21135 -6320
rect 21190 -6440 21310 -6320
rect 21355 -6440 21475 -6320
rect 21520 -6440 21640 -6320
rect 21685 -6440 21805 -6320
rect 21860 -6440 21980 -6320
rect 22025 -6440 22145 -6320
rect 22190 -6440 22310 -6320
rect 22355 -6440 22475 -6320
rect 22530 -6440 22650 -6320
rect 22695 -6440 22815 -6320
rect 22860 -6440 22980 -6320
rect 23025 -6440 23145 -6320
rect 23200 -6440 23320 -6320
rect 23365 -6440 23485 -6320
rect 23530 -6440 23650 -6320
rect 23695 -6440 23815 -6320
rect 23870 -6440 23990 -6320
rect 18510 -6615 18630 -6495
rect 18675 -6615 18795 -6495
rect 18840 -6615 18960 -6495
rect 19005 -6615 19125 -6495
rect 19180 -6615 19300 -6495
rect 19345 -6615 19465 -6495
rect 19510 -6615 19630 -6495
rect 19675 -6615 19795 -6495
rect 19850 -6615 19970 -6495
rect 20015 -6615 20135 -6495
rect 20180 -6615 20300 -6495
rect 20345 -6615 20465 -6495
rect 20520 -6615 20640 -6495
rect 20685 -6615 20805 -6495
rect 20850 -6615 20970 -6495
rect 21015 -6615 21135 -6495
rect 21190 -6615 21310 -6495
rect 21355 -6615 21475 -6495
rect 21520 -6615 21640 -6495
rect 21685 -6615 21805 -6495
rect 21860 -6615 21980 -6495
rect 22025 -6615 22145 -6495
rect 22190 -6615 22310 -6495
rect 22355 -6615 22475 -6495
rect 22530 -6615 22650 -6495
rect 22695 -6615 22815 -6495
rect 22860 -6615 22980 -6495
rect 23025 -6615 23145 -6495
rect 23200 -6615 23320 -6495
rect 23365 -6615 23485 -6495
rect 23530 -6615 23650 -6495
rect 23695 -6615 23815 -6495
rect 23870 -6615 23990 -6495
rect 18510 -6780 18630 -6660
rect 18675 -6780 18795 -6660
rect 18840 -6780 18960 -6660
rect 19005 -6780 19125 -6660
rect 19180 -6780 19300 -6660
rect 19345 -6780 19465 -6660
rect 19510 -6780 19630 -6660
rect 19675 -6780 19795 -6660
rect 19850 -6780 19970 -6660
rect 20015 -6780 20135 -6660
rect 20180 -6780 20300 -6660
rect 20345 -6780 20465 -6660
rect 20520 -6780 20640 -6660
rect 20685 -6780 20805 -6660
rect 20850 -6780 20970 -6660
rect 21015 -6780 21135 -6660
rect 21190 -6780 21310 -6660
rect 21355 -6780 21475 -6660
rect 21520 -6780 21640 -6660
rect 21685 -6780 21805 -6660
rect 21860 -6780 21980 -6660
rect 22025 -6780 22145 -6660
rect 22190 -6780 22310 -6660
rect 22355 -6780 22475 -6660
rect 22530 -6780 22650 -6660
rect 22695 -6780 22815 -6660
rect 22860 -6780 22980 -6660
rect 23025 -6780 23145 -6660
rect 23200 -6780 23320 -6660
rect 23365 -6780 23485 -6660
rect 23530 -6780 23650 -6660
rect 23695 -6780 23815 -6660
rect 23870 -6780 23990 -6660
rect 18510 -6945 18630 -6825
rect 18675 -6945 18795 -6825
rect 18840 -6945 18960 -6825
rect 19005 -6945 19125 -6825
rect 19180 -6945 19300 -6825
rect 19345 -6945 19465 -6825
rect 19510 -6945 19630 -6825
rect 19675 -6945 19795 -6825
rect 19850 -6945 19970 -6825
rect 20015 -6945 20135 -6825
rect 20180 -6945 20300 -6825
rect 20345 -6945 20465 -6825
rect 20520 -6945 20640 -6825
rect 20685 -6945 20805 -6825
rect 20850 -6945 20970 -6825
rect 21015 -6945 21135 -6825
rect 21190 -6945 21310 -6825
rect 21355 -6945 21475 -6825
rect 21520 -6945 21640 -6825
rect 21685 -6945 21805 -6825
rect 21860 -6945 21980 -6825
rect 22025 -6945 22145 -6825
rect 22190 -6945 22310 -6825
rect 22355 -6945 22475 -6825
rect 22530 -6945 22650 -6825
rect 22695 -6945 22815 -6825
rect 22860 -6945 22980 -6825
rect 23025 -6945 23145 -6825
rect 23200 -6945 23320 -6825
rect 23365 -6945 23485 -6825
rect 23530 -6945 23650 -6825
rect 23695 -6945 23815 -6825
rect 23870 -6945 23990 -6825
rect 18510 -7110 18630 -6990
rect 18675 -7110 18795 -6990
rect 18840 -7110 18960 -6990
rect 19005 -7110 19125 -6990
rect 19180 -7110 19300 -6990
rect 19345 -7110 19465 -6990
rect 19510 -7110 19630 -6990
rect 19675 -7110 19795 -6990
rect 19850 -7110 19970 -6990
rect 20015 -7110 20135 -6990
rect 20180 -7110 20300 -6990
rect 20345 -7110 20465 -6990
rect 20520 -7110 20640 -6990
rect 20685 -7110 20805 -6990
rect 20850 -7110 20970 -6990
rect 21015 -7110 21135 -6990
rect 21190 -7110 21310 -6990
rect 21355 -7110 21475 -6990
rect 21520 -7110 21640 -6990
rect 21685 -7110 21805 -6990
rect 21860 -7110 21980 -6990
rect 22025 -7110 22145 -6990
rect 22190 -7110 22310 -6990
rect 22355 -7110 22475 -6990
rect 22530 -7110 22650 -6990
rect 22695 -7110 22815 -6990
rect 22860 -7110 22980 -6990
rect 23025 -7110 23145 -6990
rect 23200 -7110 23320 -6990
rect 23365 -7110 23485 -6990
rect 23530 -7110 23650 -6990
rect 23695 -7110 23815 -6990
rect 23870 -7110 23990 -6990
rect 18510 -7285 18630 -7165
rect 18675 -7285 18795 -7165
rect 18840 -7285 18960 -7165
rect 19005 -7285 19125 -7165
rect 19180 -7285 19300 -7165
rect 19345 -7285 19465 -7165
rect 19510 -7285 19630 -7165
rect 19675 -7285 19795 -7165
rect 19850 -7285 19970 -7165
rect 20015 -7285 20135 -7165
rect 20180 -7285 20300 -7165
rect 20345 -7285 20465 -7165
rect 20520 -7285 20640 -7165
rect 20685 -7285 20805 -7165
rect 20850 -7285 20970 -7165
rect 21015 -7285 21135 -7165
rect 21190 -7285 21310 -7165
rect 21355 -7285 21475 -7165
rect 21520 -7285 21640 -7165
rect 21685 -7285 21805 -7165
rect 21860 -7285 21980 -7165
rect 22025 -7285 22145 -7165
rect 22190 -7285 22310 -7165
rect 22355 -7285 22475 -7165
rect 22530 -7285 22650 -7165
rect 22695 -7285 22815 -7165
rect 22860 -7285 22980 -7165
rect 23025 -7285 23145 -7165
rect 23200 -7285 23320 -7165
rect 23365 -7285 23485 -7165
rect 23530 -7285 23650 -7165
rect 23695 -7285 23815 -7165
rect 23870 -7285 23990 -7165
rect 18510 -7450 18630 -7330
rect 18675 -7450 18795 -7330
rect 18840 -7450 18960 -7330
rect 19005 -7450 19125 -7330
rect 19180 -7450 19300 -7330
rect 19345 -7450 19465 -7330
rect 19510 -7450 19630 -7330
rect 19675 -7450 19795 -7330
rect 19850 -7450 19970 -7330
rect 20015 -7450 20135 -7330
rect 20180 -7450 20300 -7330
rect 20345 -7450 20465 -7330
rect 20520 -7450 20640 -7330
rect 20685 -7450 20805 -7330
rect 20850 -7450 20970 -7330
rect 21015 -7450 21135 -7330
rect 21190 -7450 21310 -7330
rect 21355 -7450 21475 -7330
rect 21520 -7450 21640 -7330
rect 21685 -7450 21805 -7330
rect 21860 -7450 21980 -7330
rect 22025 -7450 22145 -7330
rect 22190 -7450 22310 -7330
rect 22355 -7450 22475 -7330
rect 22530 -7450 22650 -7330
rect 22695 -7450 22815 -7330
rect 22860 -7450 22980 -7330
rect 23025 -7450 23145 -7330
rect 23200 -7450 23320 -7330
rect 23365 -7450 23485 -7330
rect 23530 -7450 23650 -7330
rect 23695 -7450 23815 -7330
rect 23870 -7450 23990 -7330
rect 18510 -7615 18630 -7495
rect 18675 -7615 18795 -7495
rect 18840 -7615 18960 -7495
rect 19005 -7615 19125 -7495
rect 19180 -7615 19300 -7495
rect 19345 -7615 19465 -7495
rect 19510 -7615 19630 -7495
rect 19675 -7615 19795 -7495
rect 19850 -7615 19970 -7495
rect 20015 -7615 20135 -7495
rect 20180 -7615 20300 -7495
rect 20345 -7615 20465 -7495
rect 20520 -7615 20640 -7495
rect 20685 -7615 20805 -7495
rect 20850 -7615 20970 -7495
rect 21015 -7615 21135 -7495
rect 21190 -7615 21310 -7495
rect 21355 -7615 21475 -7495
rect 21520 -7615 21640 -7495
rect 21685 -7615 21805 -7495
rect 21860 -7615 21980 -7495
rect 22025 -7615 22145 -7495
rect 22190 -7615 22310 -7495
rect 22355 -7615 22475 -7495
rect 22530 -7615 22650 -7495
rect 22695 -7615 22815 -7495
rect 22860 -7615 22980 -7495
rect 23025 -7615 23145 -7495
rect 23200 -7615 23320 -7495
rect 23365 -7615 23485 -7495
rect 23530 -7615 23650 -7495
rect 23695 -7615 23815 -7495
rect 23870 -7615 23990 -7495
rect 18510 -7780 18630 -7660
rect 18675 -7780 18795 -7660
rect 18840 -7780 18960 -7660
rect 19005 -7780 19125 -7660
rect 19180 -7780 19300 -7660
rect 19345 -7780 19465 -7660
rect 19510 -7780 19630 -7660
rect 19675 -7780 19795 -7660
rect 19850 -7780 19970 -7660
rect 20015 -7780 20135 -7660
rect 20180 -7780 20300 -7660
rect 20345 -7780 20465 -7660
rect 20520 -7780 20640 -7660
rect 20685 -7780 20805 -7660
rect 20850 -7780 20970 -7660
rect 21015 -7780 21135 -7660
rect 21190 -7780 21310 -7660
rect 21355 -7780 21475 -7660
rect 21520 -7780 21640 -7660
rect 21685 -7780 21805 -7660
rect 21860 -7780 21980 -7660
rect 22025 -7780 22145 -7660
rect 22190 -7780 22310 -7660
rect 22355 -7780 22475 -7660
rect 22530 -7780 22650 -7660
rect 22695 -7780 22815 -7660
rect 22860 -7780 22980 -7660
rect 23025 -7780 23145 -7660
rect 23200 -7780 23320 -7660
rect 23365 -7780 23485 -7660
rect 23530 -7780 23650 -7660
rect 23695 -7780 23815 -7660
rect 23870 -7780 23990 -7660
rect 18510 -7955 18630 -7835
rect 18675 -7955 18795 -7835
rect 18840 -7955 18960 -7835
rect 19005 -7955 19125 -7835
rect 19180 -7955 19300 -7835
rect 19345 -7955 19465 -7835
rect 19510 -7955 19630 -7835
rect 19675 -7955 19795 -7835
rect 19850 -7955 19970 -7835
rect 20015 -7955 20135 -7835
rect 20180 -7955 20300 -7835
rect 20345 -7955 20465 -7835
rect 20520 -7955 20640 -7835
rect 20685 -7955 20805 -7835
rect 20850 -7955 20970 -7835
rect 21015 -7955 21135 -7835
rect 21190 -7955 21310 -7835
rect 21355 -7955 21475 -7835
rect 21520 -7955 21640 -7835
rect 21685 -7955 21805 -7835
rect 21860 -7955 21980 -7835
rect 22025 -7955 22145 -7835
rect 22190 -7955 22310 -7835
rect 22355 -7955 22475 -7835
rect 22530 -7955 22650 -7835
rect 22695 -7955 22815 -7835
rect 22860 -7955 22980 -7835
rect 23025 -7955 23145 -7835
rect 23200 -7955 23320 -7835
rect 23365 -7955 23485 -7835
rect 23530 -7955 23650 -7835
rect 23695 -7955 23815 -7835
rect 23870 -7955 23990 -7835
rect 18510 -8120 18630 -8000
rect 18675 -8120 18795 -8000
rect 18840 -8120 18960 -8000
rect 19005 -8120 19125 -8000
rect 19180 -8120 19300 -8000
rect 19345 -8120 19465 -8000
rect 19510 -8120 19630 -8000
rect 19675 -8120 19795 -8000
rect 19850 -8120 19970 -8000
rect 20015 -8120 20135 -8000
rect 20180 -8120 20300 -8000
rect 20345 -8120 20465 -8000
rect 20520 -8120 20640 -8000
rect 20685 -8120 20805 -8000
rect 20850 -8120 20970 -8000
rect 21015 -8120 21135 -8000
rect 21190 -8120 21310 -8000
rect 21355 -8120 21475 -8000
rect 21520 -8120 21640 -8000
rect 21685 -8120 21805 -8000
rect 21860 -8120 21980 -8000
rect 22025 -8120 22145 -8000
rect 22190 -8120 22310 -8000
rect 22355 -8120 22475 -8000
rect 22530 -8120 22650 -8000
rect 22695 -8120 22815 -8000
rect 22860 -8120 22980 -8000
rect 23025 -8120 23145 -8000
rect 23200 -8120 23320 -8000
rect 23365 -8120 23485 -8000
rect 23530 -8120 23650 -8000
rect 23695 -8120 23815 -8000
rect 23870 -8120 23990 -8000
rect 18510 -8285 18630 -8165
rect 18675 -8285 18795 -8165
rect 18840 -8285 18960 -8165
rect 19005 -8285 19125 -8165
rect 19180 -8285 19300 -8165
rect 19345 -8285 19465 -8165
rect 19510 -8285 19630 -8165
rect 19675 -8285 19795 -8165
rect 19850 -8285 19970 -8165
rect 20015 -8285 20135 -8165
rect 20180 -8285 20300 -8165
rect 20345 -8285 20465 -8165
rect 20520 -8285 20640 -8165
rect 20685 -8285 20805 -8165
rect 20850 -8285 20970 -8165
rect 21015 -8285 21135 -8165
rect 21190 -8285 21310 -8165
rect 21355 -8285 21475 -8165
rect 21520 -8285 21640 -8165
rect 21685 -8285 21805 -8165
rect 21860 -8285 21980 -8165
rect 22025 -8285 22145 -8165
rect 22190 -8285 22310 -8165
rect 22355 -8285 22475 -8165
rect 22530 -8285 22650 -8165
rect 22695 -8285 22815 -8165
rect 22860 -8285 22980 -8165
rect 23025 -8285 23145 -8165
rect 23200 -8285 23320 -8165
rect 23365 -8285 23485 -8165
rect 23530 -8285 23650 -8165
rect 23695 -8285 23815 -8165
rect 23870 -8285 23990 -8165
rect 18510 -8450 18630 -8330
rect 18675 -8450 18795 -8330
rect 18840 -8450 18960 -8330
rect 19005 -8450 19125 -8330
rect 19180 -8450 19300 -8330
rect 19345 -8450 19465 -8330
rect 19510 -8450 19630 -8330
rect 19675 -8450 19795 -8330
rect 19850 -8450 19970 -8330
rect 20015 -8450 20135 -8330
rect 20180 -8450 20300 -8330
rect 20345 -8450 20465 -8330
rect 20520 -8450 20640 -8330
rect 20685 -8450 20805 -8330
rect 20850 -8450 20970 -8330
rect 21015 -8450 21135 -8330
rect 21190 -8450 21310 -8330
rect 21355 -8450 21475 -8330
rect 21520 -8450 21640 -8330
rect 21685 -8450 21805 -8330
rect 21860 -8450 21980 -8330
rect 22025 -8450 22145 -8330
rect 22190 -8450 22310 -8330
rect 22355 -8450 22475 -8330
rect 22530 -8450 22650 -8330
rect 22695 -8450 22815 -8330
rect 22860 -8450 22980 -8330
rect 23025 -8450 23145 -8330
rect 23200 -8450 23320 -8330
rect 23365 -8450 23485 -8330
rect 23530 -8450 23650 -8330
rect 23695 -8450 23815 -8330
rect 23870 -8450 23990 -8330
rect 18510 -8625 18630 -8505
rect 18675 -8625 18795 -8505
rect 18840 -8625 18960 -8505
rect 19005 -8625 19125 -8505
rect 19180 -8625 19300 -8505
rect 19345 -8625 19465 -8505
rect 19510 -8625 19630 -8505
rect 19675 -8625 19795 -8505
rect 19850 -8625 19970 -8505
rect 20015 -8625 20135 -8505
rect 20180 -8625 20300 -8505
rect 20345 -8625 20465 -8505
rect 20520 -8625 20640 -8505
rect 20685 -8625 20805 -8505
rect 20850 -8625 20970 -8505
rect 21015 -8625 21135 -8505
rect 21190 -8625 21310 -8505
rect 21355 -8625 21475 -8505
rect 21520 -8625 21640 -8505
rect 21685 -8625 21805 -8505
rect 21860 -8625 21980 -8505
rect 22025 -8625 22145 -8505
rect 22190 -8625 22310 -8505
rect 22355 -8625 22475 -8505
rect 22530 -8625 22650 -8505
rect 22695 -8625 22815 -8505
rect 22860 -8625 22980 -8505
rect 23025 -8625 23145 -8505
rect 23200 -8625 23320 -8505
rect 23365 -8625 23485 -8505
rect 23530 -8625 23650 -8505
rect 23695 -8625 23815 -8505
rect 23870 -8625 23990 -8505
rect 18510 -8790 18630 -8670
rect 18675 -8790 18795 -8670
rect 18840 -8790 18960 -8670
rect 19005 -8790 19125 -8670
rect 19180 -8790 19300 -8670
rect 19345 -8790 19465 -8670
rect 19510 -8790 19630 -8670
rect 19675 -8790 19795 -8670
rect 19850 -8790 19970 -8670
rect 20015 -8790 20135 -8670
rect 20180 -8790 20300 -8670
rect 20345 -8790 20465 -8670
rect 20520 -8790 20640 -8670
rect 20685 -8790 20805 -8670
rect 20850 -8790 20970 -8670
rect 21015 -8790 21135 -8670
rect 21190 -8790 21310 -8670
rect 21355 -8790 21475 -8670
rect 21520 -8790 21640 -8670
rect 21685 -8790 21805 -8670
rect 21860 -8790 21980 -8670
rect 22025 -8790 22145 -8670
rect 22190 -8790 22310 -8670
rect 22355 -8790 22475 -8670
rect 22530 -8790 22650 -8670
rect 22695 -8790 22815 -8670
rect 22860 -8790 22980 -8670
rect 23025 -8790 23145 -8670
rect 23200 -8790 23320 -8670
rect 23365 -8790 23485 -8670
rect 23530 -8790 23650 -8670
rect 23695 -8790 23815 -8670
rect 23870 -8790 23990 -8670
rect 18510 -8955 18630 -8835
rect 18675 -8955 18795 -8835
rect 18840 -8955 18960 -8835
rect 19005 -8955 19125 -8835
rect 19180 -8955 19300 -8835
rect 19345 -8955 19465 -8835
rect 19510 -8955 19630 -8835
rect 19675 -8955 19795 -8835
rect 19850 -8955 19970 -8835
rect 20015 -8955 20135 -8835
rect 20180 -8955 20300 -8835
rect 20345 -8955 20465 -8835
rect 20520 -8955 20640 -8835
rect 20685 -8955 20805 -8835
rect 20850 -8955 20970 -8835
rect 21015 -8955 21135 -8835
rect 21190 -8955 21310 -8835
rect 21355 -8955 21475 -8835
rect 21520 -8955 21640 -8835
rect 21685 -8955 21805 -8835
rect 21860 -8955 21980 -8835
rect 22025 -8955 22145 -8835
rect 22190 -8955 22310 -8835
rect 22355 -8955 22475 -8835
rect 22530 -8955 22650 -8835
rect 22695 -8955 22815 -8835
rect 22860 -8955 22980 -8835
rect 23025 -8955 23145 -8835
rect 23200 -8955 23320 -8835
rect 23365 -8955 23485 -8835
rect 23530 -8955 23650 -8835
rect 23695 -8955 23815 -8835
rect 23870 -8955 23990 -8835
rect 18510 -9120 18630 -9000
rect 18675 -9120 18795 -9000
rect 18840 -9120 18960 -9000
rect 19005 -9120 19125 -9000
rect 19180 -9120 19300 -9000
rect 19345 -9120 19465 -9000
rect 19510 -9120 19630 -9000
rect 19675 -9120 19795 -9000
rect 19850 -9120 19970 -9000
rect 20015 -9120 20135 -9000
rect 20180 -9120 20300 -9000
rect 20345 -9120 20465 -9000
rect 20520 -9120 20640 -9000
rect 20685 -9120 20805 -9000
rect 20850 -9120 20970 -9000
rect 21015 -9120 21135 -9000
rect 21190 -9120 21310 -9000
rect 21355 -9120 21475 -9000
rect 21520 -9120 21640 -9000
rect 21685 -9120 21805 -9000
rect 21860 -9120 21980 -9000
rect 22025 -9120 22145 -9000
rect 22190 -9120 22310 -9000
rect 22355 -9120 22475 -9000
rect 22530 -9120 22650 -9000
rect 22695 -9120 22815 -9000
rect 22860 -9120 22980 -9000
rect 23025 -9120 23145 -9000
rect 23200 -9120 23320 -9000
rect 23365 -9120 23485 -9000
rect 23530 -9120 23650 -9000
rect 23695 -9120 23815 -9000
rect 23870 -9120 23990 -9000
rect 18510 -9295 18630 -9175
rect 18675 -9295 18795 -9175
rect 18840 -9295 18960 -9175
rect 19005 -9295 19125 -9175
rect 19180 -9295 19300 -9175
rect 19345 -9295 19465 -9175
rect 19510 -9295 19630 -9175
rect 19675 -9295 19795 -9175
rect 19850 -9295 19970 -9175
rect 20015 -9295 20135 -9175
rect 20180 -9295 20300 -9175
rect 20345 -9295 20465 -9175
rect 20520 -9295 20640 -9175
rect 20685 -9295 20805 -9175
rect 20850 -9295 20970 -9175
rect 21015 -9295 21135 -9175
rect 21190 -9295 21310 -9175
rect 21355 -9295 21475 -9175
rect 21520 -9295 21640 -9175
rect 21685 -9295 21805 -9175
rect 21860 -9295 21980 -9175
rect 22025 -9295 22145 -9175
rect 22190 -9295 22310 -9175
rect 22355 -9295 22475 -9175
rect 22530 -9295 22650 -9175
rect 22695 -9295 22815 -9175
rect 22860 -9295 22980 -9175
rect 23025 -9295 23145 -9175
rect 23200 -9295 23320 -9175
rect 23365 -9295 23485 -9175
rect 23530 -9295 23650 -9175
rect 23695 -9295 23815 -9175
rect 23870 -9295 23990 -9175
rect 18510 -9460 18630 -9340
rect 18675 -9460 18795 -9340
rect 18840 -9460 18960 -9340
rect 19005 -9460 19125 -9340
rect 19180 -9460 19300 -9340
rect 19345 -9460 19465 -9340
rect 19510 -9460 19630 -9340
rect 19675 -9460 19795 -9340
rect 19850 -9460 19970 -9340
rect 20015 -9460 20135 -9340
rect 20180 -9460 20300 -9340
rect 20345 -9460 20465 -9340
rect 20520 -9460 20640 -9340
rect 20685 -9460 20805 -9340
rect 20850 -9460 20970 -9340
rect 21015 -9460 21135 -9340
rect 21190 -9460 21310 -9340
rect 21355 -9460 21475 -9340
rect 21520 -9460 21640 -9340
rect 21685 -9460 21805 -9340
rect 21860 -9460 21980 -9340
rect 22025 -9460 22145 -9340
rect 22190 -9460 22310 -9340
rect 22355 -9460 22475 -9340
rect 22530 -9460 22650 -9340
rect 22695 -9460 22815 -9340
rect 22860 -9460 22980 -9340
rect 23025 -9460 23145 -9340
rect 23200 -9460 23320 -9340
rect 23365 -9460 23485 -9340
rect 23530 -9460 23650 -9340
rect 23695 -9460 23815 -9340
rect 23870 -9460 23990 -9340
rect 18510 -9625 18630 -9505
rect 18675 -9625 18795 -9505
rect 18840 -9625 18960 -9505
rect 19005 -9625 19125 -9505
rect 19180 -9625 19300 -9505
rect 19345 -9625 19465 -9505
rect 19510 -9625 19630 -9505
rect 19675 -9625 19795 -9505
rect 19850 -9625 19970 -9505
rect 20015 -9625 20135 -9505
rect 20180 -9625 20300 -9505
rect 20345 -9625 20465 -9505
rect 20520 -9625 20640 -9505
rect 20685 -9625 20805 -9505
rect 20850 -9625 20970 -9505
rect 21015 -9625 21135 -9505
rect 21190 -9625 21310 -9505
rect 21355 -9625 21475 -9505
rect 21520 -9625 21640 -9505
rect 21685 -9625 21805 -9505
rect 21860 -9625 21980 -9505
rect 22025 -9625 22145 -9505
rect 22190 -9625 22310 -9505
rect 22355 -9625 22475 -9505
rect 22530 -9625 22650 -9505
rect 22695 -9625 22815 -9505
rect 22860 -9625 22980 -9505
rect 23025 -9625 23145 -9505
rect 23200 -9625 23320 -9505
rect 23365 -9625 23485 -9505
rect 23530 -9625 23650 -9505
rect 23695 -9625 23815 -9505
rect 23870 -9625 23990 -9505
rect 18510 -9790 18630 -9670
rect 18675 -9790 18795 -9670
rect 18840 -9790 18960 -9670
rect 19005 -9790 19125 -9670
rect 19180 -9790 19300 -9670
rect 19345 -9790 19465 -9670
rect 19510 -9790 19630 -9670
rect 19675 -9790 19795 -9670
rect 19850 -9790 19970 -9670
rect 20015 -9790 20135 -9670
rect 20180 -9790 20300 -9670
rect 20345 -9790 20465 -9670
rect 20520 -9790 20640 -9670
rect 20685 -9790 20805 -9670
rect 20850 -9790 20970 -9670
rect 21015 -9790 21135 -9670
rect 21190 -9790 21310 -9670
rect 21355 -9790 21475 -9670
rect 21520 -9790 21640 -9670
rect 21685 -9790 21805 -9670
rect 21860 -9790 21980 -9670
rect 22025 -9790 22145 -9670
rect 22190 -9790 22310 -9670
rect 22355 -9790 22475 -9670
rect 22530 -9790 22650 -9670
rect 22695 -9790 22815 -9670
rect 22860 -9790 22980 -9670
rect 23025 -9790 23145 -9670
rect 23200 -9790 23320 -9670
rect 23365 -9790 23485 -9670
rect 23530 -9790 23650 -9670
rect 23695 -9790 23815 -9670
rect 23870 -9790 23990 -9670
rect 24200 -4430 24320 -4310
rect 24365 -4430 24485 -4310
rect 24530 -4430 24650 -4310
rect 24695 -4430 24815 -4310
rect 24870 -4430 24990 -4310
rect 25035 -4430 25155 -4310
rect 25200 -4430 25320 -4310
rect 25365 -4430 25485 -4310
rect 25540 -4430 25660 -4310
rect 25705 -4430 25825 -4310
rect 25870 -4430 25990 -4310
rect 26035 -4430 26155 -4310
rect 26210 -4430 26330 -4310
rect 26375 -4430 26495 -4310
rect 26540 -4430 26660 -4310
rect 26705 -4430 26825 -4310
rect 26880 -4430 27000 -4310
rect 27045 -4430 27165 -4310
rect 27210 -4430 27330 -4310
rect 27375 -4430 27495 -4310
rect 27550 -4430 27670 -4310
rect 27715 -4430 27835 -4310
rect 27880 -4430 28000 -4310
rect 28045 -4430 28165 -4310
rect 28220 -4430 28340 -4310
rect 28385 -4430 28505 -4310
rect 28550 -4430 28670 -4310
rect 28715 -4430 28835 -4310
rect 28890 -4430 29010 -4310
rect 29055 -4430 29175 -4310
rect 29220 -4430 29340 -4310
rect 29385 -4430 29505 -4310
rect 29560 -4430 29680 -4310
rect 24200 -4605 24320 -4485
rect 24365 -4605 24485 -4485
rect 24530 -4605 24650 -4485
rect 24695 -4605 24815 -4485
rect 24870 -4605 24990 -4485
rect 25035 -4605 25155 -4485
rect 25200 -4605 25320 -4485
rect 25365 -4605 25485 -4485
rect 25540 -4605 25660 -4485
rect 25705 -4605 25825 -4485
rect 25870 -4605 25990 -4485
rect 26035 -4605 26155 -4485
rect 26210 -4605 26330 -4485
rect 26375 -4605 26495 -4485
rect 26540 -4605 26660 -4485
rect 26705 -4605 26825 -4485
rect 26880 -4605 27000 -4485
rect 27045 -4605 27165 -4485
rect 27210 -4605 27330 -4485
rect 27375 -4605 27495 -4485
rect 27550 -4605 27670 -4485
rect 27715 -4605 27835 -4485
rect 27880 -4605 28000 -4485
rect 28045 -4605 28165 -4485
rect 28220 -4605 28340 -4485
rect 28385 -4605 28505 -4485
rect 28550 -4605 28670 -4485
rect 28715 -4605 28835 -4485
rect 28890 -4605 29010 -4485
rect 29055 -4605 29175 -4485
rect 29220 -4605 29340 -4485
rect 29385 -4605 29505 -4485
rect 29560 -4605 29680 -4485
rect 24200 -4770 24320 -4650
rect 24365 -4770 24485 -4650
rect 24530 -4770 24650 -4650
rect 24695 -4770 24815 -4650
rect 24870 -4770 24990 -4650
rect 25035 -4770 25155 -4650
rect 25200 -4770 25320 -4650
rect 25365 -4770 25485 -4650
rect 25540 -4770 25660 -4650
rect 25705 -4770 25825 -4650
rect 25870 -4770 25990 -4650
rect 26035 -4770 26155 -4650
rect 26210 -4770 26330 -4650
rect 26375 -4770 26495 -4650
rect 26540 -4770 26660 -4650
rect 26705 -4770 26825 -4650
rect 26880 -4770 27000 -4650
rect 27045 -4770 27165 -4650
rect 27210 -4770 27330 -4650
rect 27375 -4770 27495 -4650
rect 27550 -4770 27670 -4650
rect 27715 -4770 27835 -4650
rect 27880 -4770 28000 -4650
rect 28045 -4770 28165 -4650
rect 28220 -4770 28340 -4650
rect 28385 -4770 28505 -4650
rect 28550 -4770 28670 -4650
rect 28715 -4770 28835 -4650
rect 28890 -4770 29010 -4650
rect 29055 -4770 29175 -4650
rect 29220 -4770 29340 -4650
rect 29385 -4770 29505 -4650
rect 29560 -4770 29680 -4650
rect 24200 -4935 24320 -4815
rect 24365 -4935 24485 -4815
rect 24530 -4935 24650 -4815
rect 24695 -4935 24815 -4815
rect 24870 -4935 24990 -4815
rect 25035 -4935 25155 -4815
rect 25200 -4935 25320 -4815
rect 25365 -4935 25485 -4815
rect 25540 -4935 25660 -4815
rect 25705 -4935 25825 -4815
rect 25870 -4935 25990 -4815
rect 26035 -4935 26155 -4815
rect 26210 -4935 26330 -4815
rect 26375 -4935 26495 -4815
rect 26540 -4935 26660 -4815
rect 26705 -4935 26825 -4815
rect 26880 -4935 27000 -4815
rect 27045 -4935 27165 -4815
rect 27210 -4935 27330 -4815
rect 27375 -4935 27495 -4815
rect 27550 -4935 27670 -4815
rect 27715 -4935 27835 -4815
rect 27880 -4935 28000 -4815
rect 28045 -4935 28165 -4815
rect 28220 -4935 28340 -4815
rect 28385 -4935 28505 -4815
rect 28550 -4935 28670 -4815
rect 28715 -4935 28835 -4815
rect 28890 -4935 29010 -4815
rect 29055 -4935 29175 -4815
rect 29220 -4935 29340 -4815
rect 29385 -4935 29505 -4815
rect 29560 -4935 29680 -4815
rect 24200 -5100 24320 -4980
rect 24365 -5100 24485 -4980
rect 24530 -5100 24650 -4980
rect 24695 -5100 24815 -4980
rect 24870 -5100 24990 -4980
rect 25035 -5100 25155 -4980
rect 25200 -5100 25320 -4980
rect 25365 -5100 25485 -4980
rect 25540 -5100 25660 -4980
rect 25705 -5100 25825 -4980
rect 25870 -5100 25990 -4980
rect 26035 -5100 26155 -4980
rect 26210 -5100 26330 -4980
rect 26375 -5100 26495 -4980
rect 26540 -5100 26660 -4980
rect 26705 -5100 26825 -4980
rect 26880 -5100 27000 -4980
rect 27045 -5100 27165 -4980
rect 27210 -5100 27330 -4980
rect 27375 -5100 27495 -4980
rect 27550 -5100 27670 -4980
rect 27715 -5100 27835 -4980
rect 27880 -5100 28000 -4980
rect 28045 -5100 28165 -4980
rect 28220 -5100 28340 -4980
rect 28385 -5100 28505 -4980
rect 28550 -5100 28670 -4980
rect 28715 -5100 28835 -4980
rect 28890 -5100 29010 -4980
rect 29055 -5100 29175 -4980
rect 29220 -5100 29340 -4980
rect 29385 -5100 29505 -4980
rect 29560 -5100 29680 -4980
rect 24200 -5275 24320 -5155
rect 24365 -5275 24485 -5155
rect 24530 -5275 24650 -5155
rect 24695 -5275 24815 -5155
rect 24870 -5275 24990 -5155
rect 25035 -5275 25155 -5155
rect 25200 -5275 25320 -5155
rect 25365 -5275 25485 -5155
rect 25540 -5275 25660 -5155
rect 25705 -5275 25825 -5155
rect 25870 -5275 25990 -5155
rect 26035 -5275 26155 -5155
rect 26210 -5275 26330 -5155
rect 26375 -5275 26495 -5155
rect 26540 -5275 26660 -5155
rect 26705 -5275 26825 -5155
rect 26880 -5275 27000 -5155
rect 27045 -5275 27165 -5155
rect 27210 -5275 27330 -5155
rect 27375 -5275 27495 -5155
rect 27550 -5275 27670 -5155
rect 27715 -5275 27835 -5155
rect 27880 -5275 28000 -5155
rect 28045 -5275 28165 -5155
rect 28220 -5275 28340 -5155
rect 28385 -5275 28505 -5155
rect 28550 -5275 28670 -5155
rect 28715 -5275 28835 -5155
rect 28890 -5275 29010 -5155
rect 29055 -5275 29175 -5155
rect 29220 -5275 29340 -5155
rect 29385 -5275 29505 -5155
rect 29560 -5275 29680 -5155
rect 24200 -5440 24320 -5320
rect 24365 -5440 24485 -5320
rect 24530 -5440 24650 -5320
rect 24695 -5440 24815 -5320
rect 24870 -5440 24990 -5320
rect 25035 -5440 25155 -5320
rect 25200 -5440 25320 -5320
rect 25365 -5440 25485 -5320
rect 25540 -5440 25660 -5320
rect 25705 -5440 25825 -5320
rect 25870 -5440 25990 -5320
rect 26035 -5440 26155 -5320
rect 26210 -5440 26330 -5320
rect 26375 -5440 26495 -5320
rect 26540 -5440 26660 -5320
rect 26705 -5440 26825 -5320
rect 26880 -5440 27000 -5320
rect 27045 -5440 27165 -5320
rect 27210 -5440 27330 -5320
rect 27375 -5440 27495 -5320
rect 27550 -5440 27670 -5320
rect 27715 -5440 27835 -5320
rect 27880 -5440 28000 -5320
rect 28045 -5440 28165 -5320
rect 28220 -5440 28340 -5320
rect 28385 -5440 28505 -5320
rect 28550 -5440 28670 -5320
rect 28715 -5440 28835 -5320
rect 28890 -5440 29010 -5320
rect 29055 -5440 29175 -5320
rect 29220 -5440 29340 -5320
rect 29385 -5440 29505 -5320
rect 29560 -5440 29680 -5320
rect 24200 -5605 24320 -5485
rect 24365 -5605 24485 -5485
rect 24530 -5605 24650 -5485
rect 24695 -5605 24815 -5485
rect 24870 -5605 24990 -5485
rect 25035 -5605 25155 -5485
rect 25200 -5605 25320 -5485
rect 25365 -5605 25485 -5485
rect 25540 -5605 25660 -5485
rect 25705 -5605 25825 -5485
rect 25870 -5605 25990 -5485
rect 26035 -5605 26155 -5485
rect 26210 -5605 26330 -5485
rect 26375 -5605 26495 -5485
rect 26540 -5605 26660 -5485
rect 26705 -5605 26825 -5485
rect 26880 -5605 27000 -5485
rect 27045 -5605 27165 -5485
rect 27210 -5605 27330 -5485
rect 27375 -5605 27495 -5485
rect 27550 -5605 27670 -5485
rect 27715 -5605 27835 -5485
rect 27880 -5605 28000 -5485
rect 28045 -5605 28165 -5485
rect 28220 -5605 28340 -5485
rect 28385 -5605 28505 -5485
rect 28550 -5605 28670 -5485
rect 28715 -5605 28835 -5485
rect 28890 -5605 29010 -5485
rect 29055 -5605 29175 -5485
rect 29220 -5605 29340 -5485
rect 29385 -5605 29505 -5485
rect 29560 -5605 29680 -5485
rect 24200 -5770 24320 -5650
rect 24365 -5770 24485 -5650
rect 24530 -5770 24650 -5650
rect 24695 -5770 24815 -5650
rect 24870 -5770 24990 -5650
rect 25035 -5770 25155 -5650
rect 25200 -5770 25320 -5650
rect 25365 -5770 25485 -5650
rect 25540 -5770 25660 -5650
rect 25705 -5770 25825 -5650
rect 25870 -5770 25990 -5650
rect 26035 -5770 26155 -5650
rect 26210 -5770 26330 -5650
rect 26375 -5770 26495 -5650
rect 26540 -5770 26660 -5650
rect 26705 -5770 26825 -5650
rect 26880 -5770 27000 -5650
rect 27045 -5770 27165 -5650
rect 27210 -5770 27330 -5650
rect 27375 -5770 27495 -5650
rect 27550 -5770 27670 -5650
rect 27715 -5770 27835 -5650
rect 27880 -5770 28000 -5650
rect 28045 -5770 28165 -5650
rect 28220 -5770 28340 -5650
rect 28385 -5770 28505 -5650
rect 28550 -5770 28670 -5650
rect 28715 -5770 28835 -5650
rect 28890 -5770 29010 -5650
rect 29055 -5770 29175 -5650
rect 29220 -5770 29340 -5650
rect 29385 -5770 29505 -5650
rect 29560 -5770 29680 -5650
rect 24200 -5945 24320 -5825
rect 24365 -5945 24485 -5825
rect 24530 -5945 24650 -5825
rect 24695 -5945 24815 -5825
rect 24870 -5945 24990 -5825
rect 25035 -5945 25155 -5825
rect 25200 -5945 25320 -5825
rect 25365 -5945 25485 -5825
rect 25540 -5945 25660 -5825
rect 25705 -5945 25825 -5825
rect 25870 -5945 25990 -5825
rect 26035 -5945 26155 -5825
rect 26210 -5945 26330 -5825
rect 26375 -5945 26495 -5825
rect 26540 -5945 26660 -5825
rect 26705 -5945 26825 -5825
rect 26880 -5945 27000 -5825
rect 27045 -5945 27165 -5825
rect 27210 -5945 27330 -5825
rect 27375 -5945 27495 -5825
rect 27550 -5945 27670 -5825
rect 27715 -5945 27835 -5825
rect 27880 -5945 28000 -5825
rect 28045 -5945 28165 -5825
rect 28220 -5945 28340 -5825
rect 28385 -5945 28505 -5825
rect 28550 -5945 28670 -5825
rect 28715 -5945 28835 -5825
rect 28890 -5945 29010 -5825
rect 29055 -5945 29175 -5825
rect 29220 -5945 29340 -5825
rect 29385 -5945 29505 -5825
rect 29560 -5945 29680 -5825
rect 24200 -6110 24320 -5990
rect 24365 -6110 24485 -5990
rect 24530 -6110 24650 -5990
rect 24695 -6110 24815 -5990
rect 24870 -6110 24990 -5990
rect 25035 -6110 25155 -5990
rect 25200 -6110 25320 -5990
rect 25365 -6110 25485 -5990
rect 25540 -6110 25660 -5990
rect 25705 -6110 25825 -5990
rect 25870 -6110 25990 -5990
rect 26035 -6110 26155 -5990
rect 26210 -6110 26330 -5990
rect 26375 -6110 26495 -5990
rect 26540 -6110 26660 -5990
rect 26705 -6110 26825 -5990
rect 26880 -6110 27000 -5990
rect 27045 -6110 27165 -5990
rect 27210 -6110 27330 -5990
rect 27375 -6110 27495 -5990
rect 27550 -6110 27670 -5990
rect 27715 -6110 27835 -5990
rect 27880 -6110 28000 -5990
rect 28045 -6110 28165 -5990
rect 28220 -6110 28340 -5990
rect 28385 -6110 28505 -5990
rect 28550 -6110 28670 -5990
rect 28715 -6110 28835 -5990
rect 28890 -6110 29010 -5990
rect 29055 -6110 29175 -5990
rect 29220 -6110 29340 -5990
rect 29385 -6110 29505 -5990
rect 29560 -6110 29680 -5990
rect 24200 -6275 24320 -6155
rect 24365 -6275 24485 -6155
rect 24530 -6275 24650 -6155
rect 24695 -6275 24815 -6155
rect 24870 -6275 24990 -6155
rect 25035 -6275 25155 -6155
rect 25200 -6275 25320 -6155
rect 25365 -6275 25485 -6155
rect 25540 -6275 25660 -6155
rect 25705 -6275 25825 -6155
rect 25870 -6275 25990 -6155
rect 26035 -6275 26155 -6155
rect 26210 -6275 26330 -6155
rect 26375 -6275 26495 -6155
rect 26540 -6275 26660 -6155
rect 26705 -6275 26825 -6155
rect 26880 -6275 27000 -6155
rect 27045 -6275 27165 -6155
rect 27210 -6275 27330 -6155
rect 27375 -6275 27495 -6155
rect 27550 -6275 27670 -6155
rect 27715 -6275 27835 -6155
rect 27880 -6275 28000 -6155
rect 28045 -6275 28165 -6155
rect 28220 -6275 28340 -6155
rect 28385 -6275 28505 -6155
rect 28550 -6275 28670 -6155
rect 28715 -6275 28835 -6155
rect 28890 -6275 29010 -6155
rect 29055 -6275 29175 -6155
rect 29220 -6275 29340 -6155
rect 29385 -6275 29505 -6155
rect 29560 -6275 29680 -6155
rect 24200 -6440 24320 -6320
rect 24365 -6440 24485 -6320
rect 24530 -6440 24650 -6320
rect 24695 -6440 24815 -6320
rect 24870 -6440 24990 -6320
rect 25035 -6440 25155 -6320
rect 25200 -6440 25320 -6320
rect 25365 -6440 25485 -6320
rect 25540 -6440 25660 -6320
rect 25705 -6440 25825 -6320
rect 25870 -6440 25990 -6320
rect 26035 -6440 26155 -6320
rect 26210 -6440 26330 -6320
rect 26375 -6440 26495 -6320
rect 26540 -6440 26660 -6320
rect 26705 -6440 26825 -6320
rect 26880 -6440 27000 -6320
rect 27045 -6440 27165 -6320
rect 27210 -6440 27330 -6320
rect 27375 -6440 27495 -6320
rect 27550 -6440 27670 -6320
rect 27715 -6440 27835 -6320
rect 27880 -6440 28000 -6320
rect 28045 -6440 28165 -6320
rect 28220 -6440 28340 -6320
rect 28385 -6440 28505 -6320
rect 28550 -6440 28670 -6320
rect 28715 -6440 28835 -6320
rect 28890 -6440 29010 -6320
rect 29055 -6440 29175 -6320
rect 29220 -6440 29340 -6320
rect 29385 -6440 29505 -6320
rect 29560 -6440 29680 -6320
rect 24200 -6615 24320 -6495
rect 24365 -6615 24485 -6495
rect 24530 -6615 24650 -6495
rect 24695 -6615 24815 -6495
rect 24870 -6615 24990 -6495
rect 25035 -6615 25155 -6495
rect 25200 -6615 25320 -6495
rect 25365 -6615 25485 -6495
rect 25540 -6615 25660 -6495
rect 25705 -6615 25825 -6495
rect 25870 -6615 25990 -6495
rect 26035 -6615 26155 -6495
rect 26210 -6615 26330 -6495
rect 26375 -6615 26495 -6495
rect 26540 -6615 26660 -6495
rect 26705 -6615 26825 -6495
rect 26880 -6615 27000 -6495
rect 27045 -6615 27165 -6495
rect 27210 -6615 27330 -6495
rect 27375 -6615 27495 -6495
rect 27550 -6615 27670 -6495
rect 27715 -6615 27835 -6495
rect 27880 -6615 28000 -6495
rect 28045 -6615 28165 -6495
rect 28220 -6615 28340 -6495
rect 28385 -6615 28505 -6495
rect 28550 -6615 28670 -6495
rect 28715 -6615 28835 -6495
rect 28890 -6615 29010 -6495
rect 29055 -6615 29175 -6495
rect 29220 -6615 29340 -6495
rect 29385 -6615 29505 -6495
rect 29560 -6615 29680 -6495
rect 24200 -6780 24320 -6660
rect 24365 -6780 24485 -6660
rect 24530 -6780 24650 -6660
rect 24695 -6780 24815 -6660
rect 24870 -6780 24990 -6660
rect 25035 -6780 25155 -6660
rect 25200 -6780 25320 -6660
rect 25365 -6780 25485 -6660
rect 25540 -6780 25660 -6660
rect 25705 -6780 25825 -6660
rect 25870 -6780 25990 -6660
rect 26035 -6780 26155 -6660
rect 26210 -6780 26330 -6660
rect 26375 -6780 26495 -6660
rect 26540 -6780 26660 -6660
rect 26705 -6780 26825 -6660
rect 26880 -6780 27000 -6660
rect 27045 -6780 27165 -6660
rect 27210 -6780 27330 -6660
rect 27375 -6780 27495 -6660
rect 27550 -6780 27670 -6660
rect 27715 -6780 27835 -6660
rect 27880 -6780 28000 -6660
rect 28045 -6780 28165 -6660
rect 28220 -6780 28340 -6660
rect 28385 -6780 28505 -6660
rect 28550 -6780 28670 -6660
rect 28715 -6780 28835 -6660
rect 28890 -6780 29010 -6660
rect 29055 -6780 29175 -6660
rect 29220 -6780 29340 -6660
rect 29385 -6780 29505 -6660
rect 29560 -6780 29680 -6660
rect 24200 -6945 24320 -6825
rect 24365 -6945 24485 -6825
rect 24530 -6945 24650 -6825
rect 24695 -6945 24815 -6825
rect 24870 -6945 24990 -6825
rect 25035 -6945 25155 -6825
rect 25200 -6945 25320 -6825
rect 25365 -6945 25485 -6825
rect 25540 -6945 25660 -6825
rect 25705 -6945 25825 -6825
rect 25870 -6945 25990 -6825
rect 26035 -6945 26155 -6825
rect 26210 -6945 26330 -6825
rect 26375 -6945 26495 -6825
rect 26540 -6945 26660 -6825
rect 26705 -6945 26825 -6825
rect 26880 -6945 27000 -6825
rect 27045 -6945 27165 -6825
rect 27210 -6945 27330 -6825
rect 27375 -6945 27495 -6825
rect 27550 -6945 27670 -6825
rect 27715 -6945 27835 -6825
rect 27880 -6945 28000 -6825
rect 28045 -6945 28165 -6825
rect 28220 -6945 28340 -6825
rect 28385 -6945 28505 -6825
rect 28550 -6945 28670 -6825
rect 28715 -6945 28835 -6825
rect 28890 -6945 29010 -6825
rect 29055 -6945 29175 -6825
rect 29220 -6945 29340 -6825
rect 29385 -6945 29505 -6825
rect 29560 -6945 29680 -6825
rect 24200 -7110 24320 -6990
rect 24365 -7110 24485 -6990
rect 24530 -7110 24650 -6990
rect 24695 -7110 24815 -6990
rect 24870 -7110 24990 -6990
rect 25035 -7110 25155 -6990
rect 25200 -7110 25320 -6990
rect 25365 -7110 25485 -6990
rect 25540 -7110 25660 -6990
rect 25705 -7110 25825 -6990
rect 25870 -7110 25990 -6990
rect 26035 -7110 26155 -6990
rect 26210 -7110 26330 -6990
rect 26375 -7110 26495 -6990
rect 26540 -7110 26660 -6990
rect 26705 -7110 26825 -6990
rect 26880 -7110 27000 -6990
rect 27045 -7110 27165 -6990
rect 27210 -7110 27330 -6990
rect 27375 -7110 27495 -6990
rect 27550 -7110 27670 -6990
rect 27715 -7110 27835 -6990
rect 27880 -7110 28000 -6990
rect 28045 -7110 28165 -6990
rect 28220 -7110 28340 -6990
rect 28385 -7110 28505 -6990
rect 28550 -7110 28670 -6990
rect 28715 -7110 28835 -6990
rect 28890 -7110 29010 -6990
rect 29055 -7110 29175 -6990
rect 29220 -7110 29340 -6990
rect 29385 -7110 29505 -6990
rect 29560 -7110 29680 -6990
rect 24200 -7285 24320 -7165
rect 24365 -7285 24485 -7165
rect 24530 -7285 24650 -7165
rect 24695 -7285 24815 -7165
rect 24870 -7285 24990 -7165
rect 25035 -7285 25155 -7165
rect 25200 -7285 25320 -7165
rect 25365 -7285 25485 -7165
rect 25540 -7285 25660 -7165
rect 25705 -7285 25825 -7165
rect 25870 -7285 25990 -7165
rect 26035 -7285 26155 -7165
rect 26210 -7285 26330 -7165
rect 26375 -7285 26495 -7165
rect 26540 -7285 26660 -7165
rect 26705 -7285 26825 -7165
rect 26880 -7285 27000 -7165
rect 27045 -7285 27165 -7165
rect 27210 -7285 27330 -7165
rect 27375 -7285 27495 -7165
rect 27550 -7285 27670 -7165
rect 27715 -7285 27835 -7165
rect 27880 -7285 28000 -7165
rect 28045 -7285 28165 -7165
rect 28220 -7285 28340 -7165
rect 28385 -7285 28505 -7165
rect 28550 -7285 28670 -7165
rect 28715 -7285 28835 -7165
rect 28890 -7285 29010 -7165
rect 29055 -7285 29175 -7165
rect 29220 -7285 29340 -7165
rect 29385 -7285 29505 -7165
rect 29560 -7285 29680 -7165
rect 24200 -7450 24320 -7330
rect 24365 -7450 24485 -7330
rect 24530 -7450 24650 -7330
rect 24695 -7450 24815 -7330
rect 24870 -7450 24990 -7330
rect 25035 -7450 25155 -7330
rect 25200 -7450 25320 -7330
rect 25365 -7450 25485 -7330
rect 25540 -7450 25660 -7330
rect 25705 -7450 25825 -7330
rect 25870 -7450 25990 -7330
rect 26035 -7450 26155 -7330
rect 26210 -7450 26330 -7330
rect 26375 -7450 26495 -7330
rect 26540 -7450 26660 -7330
rect 26705 -7450 26825 -7330
rect 26880 -7450 27000 -7330
rect 27045 -7450 27165 -7330
rect 27210 -7450 27330 -7330
rect 27375 -7450 27495 -7330
rect 27550 -7450 27670 -7330
rect 27715 -7450 27835 -7330
rect 27880 -7450 28000 -7330
rect 28045 -7450 28165 -7330
rect 28220 -7450 28340 -7330
rect 28385 -7450 28505 -7330
rect 28550 -7450 28670 -7330
rect 28715 -7450 28835 -7330
rect 28890 -7450 29010 -7330
rect 29055 -7450 29175 -7330
rect 29220 -7450 29340 -7330
rect 29385 -7450 29505 -7330
rect 29560 -7450 29680 -7330
rect 24200 -7615 24320 -7495
rect 24365 -7615 24485 -7495
rect 24530 -7615 24650 -7495
rect 24695 -7615 24815 -7495
rect 24870 -7615 24990 -7495
rect 25035 -7615 25155 -7495
rect 25200 -7615 25320 -7495
rect 25365 -7615 25485 -7495
rect 25540 -7615 25660 -7495
rect 25705 -7615 25825 -7495
rect 25870 -7615 25990 -7495
rect 26035 -7615 26155 -7495
rect 26210 -7615 26330 -7495
rect 26375 -7615 26495 -7495
rect 26540 -7615 26660 -7495
rect 26705 -7615 26825 -7495
rect 26880 -7615 27000 -7495
rect 27045 -7615 27165 -7495
rect 27210 -7615 27330 -7495
rect 27375 -7615 27495 -7495
rect 27550 -7615 27670 -7495
rect 27715 -7615 27835 -7495
rect 27880 -7615 28000 -7495
rect 28045 -7615 28165 -7495
rect 28220 -7615 28340 -7495
rect 28385 -7615 28505 -7495
rect 28550 -7615 28670 -7495
rect 28715 -7615 28835 -7495
rect 28890 -7615 29010 -7495
rect 29055 -7615 29175 -7495
rect 29220 -7615 29340 -7495
rect 29385 -7615 29505 -7495
rect 29560 -7615 29680 -7495
rect 24200 -7780 24320 -7660
rect 24365 -7780 24485 -7660
rect 24530 -7780 24650 -7660
rect 24695 -7780 24815 -7660
rect 24870 -7780 24990 -7660
rect 25035 -7780 25155 -7660
rect 25200 -7780 25320 -7660
rect 25365 -7780 25485 -7660
rect 25540 -7780 25660 -7660
rect 25705 -7780 25825 -7660
rect 25870 -7780 25990 -7660
rect 26035 -7780 26155 -7660
rect 26210 -7780 26330 -7660
rect 26375 -7780 26495 -7660
rect 26540 -7780 26660 -7660
rect 26705 -7780 26825 -7660
rect 26880 -7780 27000 -7660
rect 27045 -7780 27165 -7660
rect 27210 -7780 27330 -7660
rect 27375 -7780 27495 -7660
rect 27550 -7780 27670 -7660
rect 27715 -7780 27835 -7660
rect 27880 -7780 28000 -7660
rect 28045 -7780 28165 -7660
rect 28220 -7780 28340 -7660
rect 28385 -7780 28505 -7660
rect 28550 -7780 28670 -7660
rect 28715 -7780 28835 -7660
rect 28890 -7780 29010 -7660
rect 29055 -7780 29175 -7660
rect 29220 -7780 29340 -7660
rect 29385 -7780 29505 -7660
rect 29560 -7780 29680 -7660
rect 24200 -7955 24320 -7835
rect 24365 -7955 24485 -7835
rect 24530 -7955 24650 -7835
rect 24695 -7955 24815 -7835
rect 24870 -7955 24990 -7835
rect 25035 -7955 25155 -7835
rect 25200 -7955 25320 -7835
rect 25365 -7955 25485 -7835
rect 25540 -7955 25660 -7835
rect 25705 -7955 25825 -7835
rect 25870 -7955 25990 -7835
rect 26035 -7955 26155 -7835
rect 26210 -7955 26330 -7835
rect 26375 -7955 26495 -7835
rect 26540 -7955 26660 -7835
rect 26705 -7955 26825 -7835
rect 26880 -7955 27000 -7835
rect 27045 -7955 27165 -7835
rect 27210 -7955 27330 -7835
rect 27375 -7955 27495 -7835
rect 27550 -7955 27670 -7835
rect 27715 -7955 27835 -7835
rect 27880 -7955 28000 -7835
rect 28045 -7955 28165 -7835
rect 28220 -7955 28340 -7835
rect 28385 -7955 28505 -7835
rect 28550 -7955 28670 -7835
rect 28715 -7955 28835 -7835
rect 28890 -7955 29010 -7835
rect 29055 -7955 29175 -7835
rect 29220 -7955 29340 -7835
rect 29385 -7955 29505 -7835
rect 29560 -7955 29680 -7835
rect 24200 -8120 24320 -8000
rect 24365 -8120 24485 -8000
rect 24530 -8120 24650 -8000
rect 24695 -8120 24815 -8000
rect 24870 -8120 24990 -8000
rect 25035 -8120 25155 -8000
rect 25200 -8120 25320 -8000
rect 25365 -8120 25485 -8000
rect 25540 -8120 25660 -8000
rect 25705 -8120 25825 -8000
rect 25870 -8120 25990 -8000
rect 26035 -8120 26155 -8000
rect 26210 -8120 26330 -8000
rect 26375 -8120 26495 -8000
rect 26540 -8120 26660 -8000
rect 26705 -8120 26825 -8000
rect 26880 -8120 27000 -8000
rect 27045 -8120 27165 -8000
rect 27210 -8120 27330 -8000
rect 27375 -8120 27495 -8000
rect 27550 -8120 27670 -8000
rect 27715 -8120 27835 -8000
rect 27880 -8120 28000 -8000
rect 28045 -8120 28165 -8000
rect 28220 -8120 28340 -8000
rect 28385 -8120 28505 -8000
rect 28550 -8120 28670 -8000
rect 28715 -8120 28835 -8000
rect 28890 -8120 29010 -8000
rect 29055 -8120 29175 -8000
rect 29220 -8120 29340 -8000
rect 29385 -8120 29505 -8000
rect 29560 -8120 29680 -8000
rect 24200 -8285 24320 -8165
rect 24365 -8285 24485 -8165
rect 24530 -8285 24650 -8165
rect 24695 -8285 24815 -8165
rect 24870 -8285 24990 -8165
rect 25035 -8285 25155 -8165
rect 25200 -8285 25320 -8165
rect 25365 -8285 25485 -8165
rect 25540 -8285 25660 -8165
rect 25705 -8285 25825 -8165
rect 25870 -8285 25990 -8165
rect 26035 -8285 26155 -8165
rect 26210 -8285 26330 -8165
rect 26375 -8285 26495 -8165
rect 26540 -8285 26660 -8165
rect 26705 -8285 26825 -8165
rect 26880 -8285 27000 -8165
rect 27045 -8285 27165 -8165
rect 27210 -8285 27330 -8165
rect 27375 -8285 27495 -8165
rect 27550 -8285 27670 -8165
rect 27715 -8285 27835 -8165
rect 27880 -8285 28000 -8165
rect 28045 -8285 28165 -8165
rect 28220 -8285 28340 -8165
rect 28385 -8285 28505 -8165
rect 28550 -8285 28670 -8165
rect 28715 -8285 28835 -8165
rect 28890 -8285 29010 -8165
rect 29055 -8285 29175 -8165
rect 29220 -8285 29340 -8165
rect 29385 -8285 29505 -8165
rect 29560 -8285 29680 -8165
rect 24200 -8450 24320 -8330
rect 24365 -8450 24485 -8330
rect 24530 -8450 24650 -8330
rect 24695 -8450 24815 -8330
rect 24870 -8450 24990 -8330
rect 25035 -8450 25155 -8330
rect 25200 -8450 25320 -8330
rect 25365 -8450 25485 -8330
rect 25540 -8450 25660 -8330
rect 25705 -8450 25825 -8330
rect 25870 -8450 25990 -8330
rect 26035 -8450 26155 -8330
rect 26210 -8450 26330 -8330
rect 26375 -8450 26495 -8330
rect 26540 -8450 26660 -8330
rect 26705 -8450 26825 -8330
rect 26880 -8450 27000 -8330
rect 27045 -8450 27165 -8330
rect 27210 -8450 27330 -8330
rect 27375 -8450 27495 -8330
rect 27550 -8450 27670 -8330
rect 27715 -8450 27835 -8330
rect 27880 -8450 28000 -8330
rect 28045 -8450 28165 -8330
rect 28220 -8450 28340 -8330
rect 28385 -8450 28505 -8330
rect 28550 -8450 28670 -8330
rect 28715 -8450 28835 -8330
rect 28890 -8450 29010 -8330
rect 29055 -8450 29175 -8330
rect 29220 -8450 29340 -8330
rect 29385 -8450 29505 -8330
rect 29560 -8450 29680 -8330
rect 24200 -8625 24320 -8505
rect 24365 -8625 24485 -8505
rect 24530 -8625 24650 -8505
rect 24695 -8625 24815 -8505
rect 24870 -8625 24990 -8505
rect 25035 -8625 25155 -8505
rect 25200 -8625 25320 -8505
rect 25365 -8625 25485 -8505
rect 25540 -8625 25660 -8505
rect 25705 -8625 25825 -8505
rect 25870 -8625 25990 -8505
rect 26035 -8625 26155 -8505
rect 26210 -8625 26330 -8505
rect 26375 -8625 26495 -8505
rect 26540 -8625 26660 -8505
rect 26705 -8625 26825 -8505
rect 26880 -8625 27000 -8505
rect 27045 -8625 27165 -8505
rect 27210 -8625 27330 -8505
rect 27375 -8625 27495 -8505
rect 27550 -8625 27670 -8505
rect 27715 -8625 27835 -8505
rect 27880 -8625 28000 -8505
rect 28045 -8625 28165 -8505
rect 28220 -8625 28340 -8505
rect 28385 -8625 28505 -8505
rect 28550 -8625 28670 -8505
rect 28715 -8625 28835 -8505
rect 28890 -8625 29010 -8505
rect 29055 -8625 29175 -8505
rect 29220 -8625 29340 -8505
rect 29385 -8625 29505 -8505
rect 29560 -8625 29680 -8505
rect 24200 -8790 24320 -8670
rect 24365 -8790 24485 -8670
rect 24530 -8790 24650 -8670
rect 24695 -8790 24815 -8670
rect 24870 -8790 24990 -8670
rect 25035 -8790 25155 -8670
rect 25200 -8790 25320 -8670
rect 25365 -8790 25485 -8670
rect 25540 -8790 25660 -8670
rect 25705 -8790 25825 -8670
rect 25870 -8790 25990 -8670
rect 26035 -8790 26155 -8670
rect 26210 -8790 26330 -8670
rect 26375 -8790 26495 -8670
rect 26540 -8790 26660 -8670
rect 26705 -8790 26825 -8670
rect 26880 -8790 27000 -8670
rect 27045 -8790 27165 -8670
rect 27210 -8790 27330 -8670
rect 27375 -8790 27495 -8670
rect 27550 -8790 27670 -8670
rect 27715 -8790 27835 -8670
rect 27880 -8790 28000 -8670
rect 28045 -8790 28165 -8670
rect 28220 -8790 28340 -8670
rect 28385 -8790 28505 -8670
rect 28550 -8790 28670 -8670
rect 28715 -8790 28835 -8670
rect 28890 -8790 29010 -8670
rect 29055 -8790 29175 -8670
rect 29220 -8790 29340 -8670
rect 29385 -8790 29505 -8670
rect 29560 -8790 29680 -8670
rect 24200 -8955 24320 -8835
rect 24365 -8955 24485 -8835
rect 24530 -8955 24650 -8835
rect 24695 -8955 24815 -8835
rect 24870 -8955 24990 -8835
rect 25035 -8955 25155 -8835
rect 25200 -8955 25320 -8835
rect 25365 -8955 25485 -8835
rect 25540 -8955 25660 -8835
rect 25705 -8955 25825 -8835
rect 25870 -8955 25990 -8835
rect 26035 -8955 26155 -8835
rect 26210 -8955 26330 -8835
rect 26375 -8955 26495 -8835
rect 26540 -8955 26660 -8835
rect 26705 -8955 26825 -8835
rect 26880 -8955 27000 -8835
rect 27045 -8955 27165 -8835
rect 27210 -8955 27330 -8835
rect 27375 -8955 27495 -8835
rect 27550 -8955 27670 -8835
rect 27715 -8955 27835 -8835
rect 27880 -8955 28000 -8835
rect 28045 -8955 28165 -8835
rect 28220 -8955 28340 -8835
rect 28385 -8955 28505 -8835
rect 28550 -8955 28670 -8835
rect 28715 -8955 28835 -8835
rect 28890 -8955 29010 -8835
rect 29055 -8955 29175 -8835
rect 29220 -8955 29340 -8835
rect 29385 -8955 29505 -8835
rect 29560 -8955 29680 -8835
rect 24200 -9120 24320 -9000
rect 24365 -9120 24485 -9000
rect 24530 -9120 24650 -9000
rect 24695 -9120 24815 -9000
rect 24870 -9120 24990 -9000
rect 25035 -9120 25155 -9000
rect 25200 -9120 25320 -9000
rect 25365 -9120 25485 -9000
rect 25540 -9120 25660 -9000
rect 25705 -9120 25825 -9000
rect 25870 -9120 25990 -9000
rect 26035 -9120 26155 -9000
rect 26210 -9120 26330 -9000
rect 26375 -9120 26495 -9000
rect 26540 -9120 26660 -9000
rect 26705 -9120 26825 -9000
rect 26880 -9120 27000 -9000
rect 27045 -9120 27165 -9000
rect 27210 -9120 27330 -9000
rect 27375 -9120 27495 -9000
rect 27550 -9120 27670 -9000
rect 27715 -9120 27835 -9000
rect 27880 -9120 28000 -9000
rect 28045 -9120 28165 -9000
rect 28220 -9120 28340 -9000
rect 28385 -9120 28505 -9000
rect 28550 -9120 28670 -9000
rect 28715 -9120 28835 -9000
rect 28890 -9120 29010 -9000
rect 29055 -9120 29175 -9000
rect 29220 -9120 29340 -9000
rect 29385 -9120 29505 -9000
rect 29560 -9120 29680 -9000
rect 24200 -9295 24320 -9175
rect 24365 -9295 24485 -9175
rect 24530 -9295 24650 -9175
rect 24695 -9295 24815 -9175
rect 24870 -9295 24990 -9175
rect 25035 -9295 25155 -9175
rect 25200 -9295 25320 -9175
rect 25365 -9295 25485 -9175
rect 25540 -9295 25660 -9175
rect 25705 -9295 25825 -9175
rect 25870 -9295 25990 -9175
rect 26035 -9295 26155 -9175
rect 26210 -9295 26330 -9175
rect 26375 -9295 26495 -9175
rect 26540 -9295 26660 -9175
rect 26705 -9295 26825 -9175
rect 26880 -9295 27000 -9175
rect 27045 -9295 27165 -9175
rect 27210 -9295 27330 -9175
rect 27375 -9295 27495 -9175
rect 27550 -9295 27670 -9175
rect 27715 -9295 27835 -9175
rect 27880 -9295 28000 -9175
rect 28045 -9295 28165 -9175
rect 28220 -9295 28340 -9175
rect 28385 -9295 28505 -9175
rect 28550 -9295 28670 -9175
rect 28715 -9295 28835 -9175
rect 28890 -9295 29010 -9175
rect 29055 -9295 29175 -9175
rect 29220 -9295 29340 -9175
rect 29385 -9295 29505 -9175
rect 29560 -9295 29680 -9175
rect 24200 -9460 24320 -9340
rect 24365 -9460 24485 -9340
rect 24530 -9460 24650 -9340
rect 24695 -9460 24815 -9340
rect 24870 -9460 24990 -9340
rect 25035 -9460 25155 -9340
rect 25200 -9460 25320 -9340
rect 25365 -9460 25485 -9340
rect 25540 -9460 25660 -9340
rect 25705 -9460 25825 -9340
rect 25870 -9460 25990 -9340
rect 26035 -9460 26155 -9340
rect 26210 -9460 26330 -9340
rect 26375 -9460 26495 -9340
rect 26540 -9460 26660 -9340
rect 26705 -9460 26825 -9340
rect 26880 -9460 27000 -9340
rect 27045 -9460 27165 -9340
rect 27210 -9460 27330 -9340
rect 27375 -9460 27495 -9340
rect 27550 -9460 27670 -9340
rect 27715 -9460 27835 -9340
rect 27880 -9460 28000 -9340
rect 28045 -9460 28165 -9340
rect 28220 -9460 28340 -9340
rect 28385 -9460 28505 -9340
rect 28550 -9460 28670 -9340
rect 28715 -9460 28835 -9340
rect 28890 -9460 29010 -9340
rect 29055 -9460 29175 -9340
rect 29220 -9460 29340 -9340
rect 29385 -9460 29505 -9340
rect 29560 -9460 29680 -9340
rect 24200 -9625 24320 -9505
rect 24365 -9625 24485 -9505
rect 24530 -9625 24650 -9505
rect 24695 -9625 24815 -9505
rect 24870 -9625 24990 -9505
rect 25035 -9625 25155 -9505
rect 25200 -9625 25320 -9505
rect 25365 -9625 25485 -9505
rect 25540 -9625 25660 -9505
rect 25705 -9625 25825 -9505
rect 25870 -9625 25990 -9505
rect 26035 -9625 26155 -9505
rect 26210 -9625 26330 -9505
rect 26375 -9625 26495 -9505
rect 26540 -9625 26660 -9505
rect 26705 -9625 26825 -9505
rect 26880 -9625 27000 -9505
rect 27045 -9625 27165 -9505
rect 27210 -9625 27330 -9505
rect 27375 -9625 27495 -9505
rect 27550 -9625 27670 -9505
rect 27715 -9625 27835 -9505
rect 27880 -9625 28000 -9505
rect 28045 -9625 28165 -9505
rect 28220 -9625 28340 -9505
rect 28385 -9625 28505 -9505
rect 28550 -9625 28670 -9505
rect 28715 -9625 28835 -9505
rect 28890 -9625 29010 -9505
rect 29055 -9625 29175 -9505
rect 29220 -9625 29340 -9505
rect 29385 -9625 29505 -9505
rect 29560 -9625 29680 -9505
rect 24200 -9790 24320 -9670
rect 24365 -9790 24485 -9670
rect 24530 -9790 24650 -9670
rect 24695 -9790 24815 -9670
rect 24870 -9790 24990 -9670
rect 25035 -9790 25155 -9670
rect 25200 -9790 25320 -9670
rect 25365 -9790 25485 -9670
rect 25540 -9790 25660 -9670
rect 25705 -9790 25825 -9670
rect 25870 -9790 25990 -9670
rect 26035 -9790 26155 -9670
rect 26210 -9790 26330 -9670
rect 26375 -9790 26495 -9670
rect 26540 -9790 26660 -9670
rect 26705 -9790 26825 -9670
rect 26880 -9790 27000 -9670
rect 27045 -9790 27165 -9670
rect 27210 -9790 27330 -9670
rect 27375 -9790 27495 -9670
rect 27550 -9790 27670 -9670
rect 27715 -9790 27835 -9670
rect 27880 -9790 28000 -9670
rect 28045 -9790 28165 -9670
rect 28220 -9790 28340 -9670
rect 28385 -9790 28505 -9670
rect 28550 -9790 28670 -9670
rect 28715 -9790 28835 -9670
rect 28890 -9790 29010 -9670
rect 29055 -9790 29175 -9670
rect 29220 -9790 29340 -9670
rect 29385 -9790 29505 -9670
rect 29560 -9790 29680 -9670
rect 7130 -10210 7250 -10090
rect 7305 -10210 7425 -10090
rect 7470 -10210 7590 -10090
rect 7635 -10210 7755 -10090
rect 7800 -10210 7920 -10090
rect 7975 -10210 8095 -10090
rect 8140 -10210 8260 -10090
rect 8305 -10210 8425 -10090
rect 8470 -10210 8590 -10090
rect 8645 -10210 8765 -10090
rect 8810 -10210 8930 -10090
rect 8975 -10210 9095 -10090
rect 9140 -10210 9260 -10090
rect 9315 -10210 9435 -10090
rect 9480 -10210 9600 -10090
rect 9645 -10210 9765 -10090
rect 9810 -10210 9930 -10090
rect 9985 -10210 10105 -10090
rect 10150 -10210 10270 -10090
rect 10315 -10210 10435 -10090
rect 10480 -10210 10600 -10090
rect 10655 -10210 10775 -10090
rect 10820 -10210 10940 -10090
rect 10985 -10210 11105 -10090
rect 11150 -10210 11270 -10090
rect 11325 -10210 11445 -10090
rect 11490 -10210 11610 -10090
rect 11655 -10210 11775 -10090
rect 11820 -10210 11940 -10090
rect 11995 -10210 12115 -10090
rect 12160 -10210 12280 -10090
rect 12325 -10210 12445 -10090
rect 12490 -10210 12610 -10090
rect 7130 -10375 7250 -10255
rect 7305 -10375 7425 -10255
rect 7470 -10375 7590 -10255
rect 7635 -10375 7755 -10255
rect 7800 -10375 7920 -10255
rect 7975 -10375 8095 -10255
rect 8140 -10375 8260 -10255
rect 8305 -10375 8425 -10255
rect 8470 -10375 8590 -10255
rect 8645 -10375 8765 -10255
rect 8810 -10375 8930 -10255
rect 8975 -10375 9095 -10255
rect 9140 -10375 9260 -10255
rect 9315 -10375 9435 -10255
rect 9480 -10375 9600 -10255
rect 9645 -10375 9765 -10255
rect 9810 -10375 9930 -10255
rect 9985 -10375 10105 -10255
rect 10150 -10375 10270 -10255
rect 10315 -10375 10435 -10255
rect 10480 -10375 10600 -10255
rect 10655 -10375 10775 -10255
rect 10820 -10375 10940 -10255
rect 10985 -10375 11105 -10255
rect 11150 -10375 11270 -10255
rect 11325 -10375 11445 -10255
rect 11490 -10375 11610 -10255
rect 11655 -10375 11775 -10255
rect 11820 -10375 11940 -10255
rect 11995 -10375 12115 -10255
rect 12160 -10375 12280 -10255
rect 12325 -10375 12445 -10255
rect 12490 -10375 12610 -10255
rect 7130 -10540 7250 -10420
rect 7305 -10540 7425 -10420
rect 7470 -10540 7590 -10420
rect 7635 -10540 7755 -10420
rect 7800 -10540 7920 -10420
rect 7975 -10540 8095 -10420
rect 8140 -10540 8260 -10420
rect 8305 -10540 8425 -10420
rect 8470 -10540 8590 -10420
rect 8645 -10540 8765 -10420
rect 8810 -10540 8930 -10420
rect 8975 -10540 9095 -10420
rect 9140 -10540 9260 -10420
rect 9315 -10540 9435 -10420
rect 9480 -10540 9600 -10420
rect 9645 -10540 9765 -10420
rect 9810 -10540 9930 -10420
rect 9985 -10540 10105 -10420
rect 10150 -10540 10270 -10420
rect 10315 -10540 10435 -10420
rect 10480 -10540 10600 -10420
rect 10655 -10540 10775 -10420
rect 10820 -10540 10940 -10420
rect 10985 -10540 11105 -10420
rect 11150 -10540 11270 -10420
rect 11325 -10540 11445 -10420
rect 11490 -10540 11610 -10420
rect 11655 -10540 11775 -10420
rect 11820 -10540 11940 -10420
rect 11995 -10540 12115 -10420
rect 12160 -10540 12280 -10420
rect 12325 -10540 12445 -10420
rect 12490 -10540 12610 -10420
rect 7130 -10705 7250 -10585
rect 7305 -10705 7425 -10585
rect 7470 -10705 7590 -10585
rect 7635 -10705 7755 -10585
rect 7800 -10705 7920 -10585
rect 7975 -10705 8095 -10585
rect 8140 -10705 8260 -10585
rect 8305 -10705 8425 -10585
rect 8470 -10705 8590 -10585
rect 8645 -10705 8765 -10585
rect 8810 -10705 8930 -10585
rect 8975 -10705 9095 -10585
rect 9140 -10705 9260 -10585
rect 9315 -10705 9435 -10585
rect 9480 -10705 9600 -10585
rect 9645 -10705 9765 -10585
rect 9810 -10705 9930 -10585
rect 9985 -10705 10105 -10585
rect 10150 -10705 10270 -10585
rect 10315 -10705 10435 -10585
rect 10480 -10705 10600 -10585
rect 10655 -10705 10775 -10585
rect 10820 -10705 10940 -10585
rect 10985 -10705 11105 -10585
rect 11150 -10705 11270 -10585
rect 11325 -10705 11445 -10585
rect 11490 -10705 11610 -10585
rect 11655 -10705 11775 -10585
rect 11820 -10705 11940 -10585
rect 11995 -10705 12115 -10585
rect 12160 -10705 12280 -10585
rect 12325 -10705 12445 -10585
rect 12490 -10705 12610 -10585
rect 7130 -10880 7250 -10760
rect 7305 -10880 7425 -10760
rect 7470 -10880 7590 -10760
rect 7635 -10880 7755 -10760
rect 7800 -10880 7920 -10760
rect 7975 -10880 8095 -10760
rect 8140 -10880 8260 -10760
rect 8305 -10880 8425 -10760
rect 8470 -10880 8590 -10760
rect 8645 -10880 8765 -10760
rect 8810 -10880 8930 -10760
rect 8975 -10880 9095 -10760
rect 9140 -10880 9260 -10760
rect 9315 -10880 9435 -10760
rect 9480 -10880 9600 -10760
rect 9645 -10880 9765 -10760
rect 9810 -10880 9930 -10760
rect 9985 -10880 10105 -10760
rect 10150 -10880 10270 -10760
rect 10315 -10880 10435 -10760
rect 10480 -10880 10600 -10760
rect 10655 -10880 10775 -10760
rect 10820 -10880 10940 -10760
rect 10985 -10880 11105 -10760
rect 11150 -10880 11270 -10760
rect 11325 -10880 11445 -10760
rect 11490 -10880 11610 -10760
rect 11655 -10880 11775 -10760
rect 11820 -10880 11940 -10760
rect 11995 -10880 12115 -10760
rect 12160 -10880 12280 -10760
rect 12325 -10880 12445 -10760
rect 12490 -10880 12610 -10760
rect 7130 -11045 7250 -10925
rect 7305 -11045 7425 -10925
rect 7470 -11045 7590 -10925
rect 7635 -11045 7755 -10925
rect 7800 -11045 7920 -10925
rect 7975 -11045 8095 -10925
rect 8140 -11045 8260 -10925
rect 8305 -11045 8425 -10925
rect 8470 -11045 8590 -10925
rect 8645 -11045 8765 -10925
rect 8810 -11045 8930 -10925
rect 8975 -11045 9095 -10925
rect 9140 -11045 9260 -10925
rect 9315 -11045 9435 -10925
rect 9480 -11045 9600 -10925
rect 9645 -11045 9765 -10925
rect 9810 -11045 9930 -10925
rect 9985 -11045 10105 -10925
rect 10150 -11045 10270 -10925
rect 10315 -11045 10435 -10925
rect 10480 -11045 10600 -10925
rect 10655 -11045 10775 -10925
rect 10820 -11045 10940 -10925
rect 10985 -11045 11105 -10925
rect 11150 -11045 11270 -10925
rect 11325 -11045 11445 -10925
rect 11490 -11045 11610 -10925
rect 11655 -11045 11775 -10925
rect 11820 -11045 11940 -10925
rect 11995 -11045 12115 -10925
rect 12160 -11045 12280 -10925
rect 12325 -11045 12445 -10925
rect 12490 -11045 12610 -10925
rect 7130 -11210 7250 -11090
rect 7305 -11210 7425 -11090
rect 7470 -11210 7590 -11090
rect 7635 -11210 7755 -11090
rect 7800 -11210 7920 -11090
rect 7975 -11210 8095 -11090
rect 8140 -11210 8260 -11090
rect 8305 -11210 8425 -11090
rect 8470 -11210 8590 -11090
rect 8645 -11210 8765 -11090
rect 8810 -11210 8930 -11090
rect 8975 -11210 9095 -11090
rect 9140 -11210 9260 -11090
rect 9315 -11210 9435 -11090
rect 9480 -11210 9600 -11090
rect 9645 -11210 9765 -11090
rect 9810 -11210 9930 -11090
rect 9985 -11210 10105 -11090
rect 10150 -11210 10270 -11090
rect 10315 -11210 10435 -11090
rect 10480 -11210 10600 -11090
rect 10655 -11210 10775 -11090
rect 10820 -11210 10940 -11090
rect 10985 -11210 11105 -11090
rect 11150 -11210 11270 -11090
rect 11325 -11210 11445 -11090
rect 11490 -11210 11610 -11090
rect 11655 -11210 11775 -11090
rect 11820 -11210 11940 -11090
rect 11995 -11210 12115 -11090
rect 12160 -11210 12280 -11090
rect 12325 -11210 12445 -11090
rect 12490 -11210 12610 -11090
rect 7130 -11375 7250 -11255
rect 7305 -11375 7425 -11255
rect 7470 -11375 7590 -11255
rect 7635 -11375 7755 -11255
rect 7800 -11375 7920 -11255
rect 7975 -11375 8095 -11255
rect 8140 -11375 8260 -11255
rect 8305 -11375 8425 -11255
rect 8470 -11375 8590 -11255
rect 8645 -11375 8765 -11255
rect 8810 -11375 8930 -11255
rect 8975 -11375 9095 -11255
rect 9140 -11375 9260 -11255
rect 9315 -11375 9435 -11255
rect 9480 -11375 9600 -11255
rect 9645 -11375 9765 -11255
rect 9810 -11375 9930 -11255
rect 9985 -11375 10105 -11255
rect 10150 -11375 10270 -11255
rect 10315 -11375 10435 -11255
rect 10480 -11375 10600 -11255
rect 10655 -11375 10775 -11255
rect 10820 -11375 10940 -11255
rect 10985 -11375 11105 -11255
rect 11150 -11375 11270 -11255
rect 11325 -11375 11445 -11255
rect 11490 -11375 11610 -11255
rect 11655 -11375 11775 -11255
rect 11820 -11375 11940 -11255
rect 11995 -11375 12115 -11255
rect 12160 -11375 12280 -11255
rect 12325 -11375 12445 -11255
rect 12490 -11375 12610 -11255
rect 7130 -11550 7250 -11430
rect 7305 -11550 7425 -11430
rect 7470 -11550 7590 -11430
rect 7635 -11550 7755 -11430
rect 7800 -11550 7920 -11430
rect 7975 -11550 8095 -11430
rect 8140 -11550 8260 -11430
rect 8305 -11550 8425 -11430
rect 8470 -11550 8590 -11430
rect 8645 -11550 8765 -11430
rect 8810 -11550 8930 -11430
rect 8975 -11550 9095 -11430
rect 9140 -11550 9260 -11430
rect 9315 -11550 9435 -11430
rect 9480 -11550 9600 -11430
rect 9645 -11550 9765 -11430
rect 9810 -11550 9930 -11430
rect 9985 -11550 10105 -11430
rect 10150 -11550 10270 -11430
rect 10315 -11550 10435 -11430
rect 10480 -11550 10600 -11430
rect 10655 -11550 10775 -11430
rect 10820 -11550 10940 -11430
rect 10985 -11550 11105 -11430
rect 11150 -11550 11270 -11430
rect 11325 -11550 11445 -11430
rect 11490 -11550 11610 -11430
rect 11655 -11550 11775 -11430
rect 11820 -11550 11940 -11430
rect 11995 -11550 12115 -11430
rect 12160 -11550 12280 -11430
rect 12325 -11550 12445 -11430
rect 12490 -11550 12610 -11430
rect 7130 -11715 7250 -11595
rect 7305 -11715 7425 -11595
rect 7470 -11715 7590 -11595
rect 7635 -11715 7755 -11595
rect 7800 -11715 7920 -11595
rect 7975 -11715 8095 -11595
rect 8140 -11715 8260 -11595
rect 8305 -11715 8425 -11595
rect 8470 -11715 8590 -11595
rect 8645 -11715 8765 -11595
rect 8810 -11715 8930 -11595
rect 8975 -11715 9095 -11595
rect 9140 -11715 9260 -11595
rect 9315 -11715 9435 -11595
rect 9480 -11715 9600 -11595
rect 9645 -11715 9765 -11595
rect 9810 -11715 9930 -11595
rect 9985 -11715 10105 -11595
rect 10150 -11715 10270 -11595
rect 10315 -11715 10435 -11595
rect 10480 -11715 10600 -11595
rect 10655 -11715 10775 -11595
rect 10820 -11715 10940 -11595
rect 10985 -11715 11105 -11595
rect 11150 -11715 11270 -11595
rect 11325 -11715 11445 -11595
rect 11490 -11715 11610 -11595
rect 11655 -11715 11775 -11595
rect 11820 -11715 11940 -11595
rect 11995 -11715 12115 -11595
rect 12160 -11715 12280 -11595
rect 12325 -11715 12445 -11595
rect 12490 -11715 12610 -11595
rect 7130 -11880 7250 -11760
rect 7305 -11880 7425 -11760
rect 7470 -11880 7590 -11760
rect 7635 -11880 7755 -11760
rect 7800 -11880 7920 -11760
rect 7975 -11880 8095 -11760
rect 8140 -11880 8260 -11760
rect 8305 -11880 8425 -11760
rect 8470 -11880 8590 -11760
rect 8645 -11880 8765 -11760
rect 8810 -11880 8930 -11760
rect 8975 -11880 9095 -11760
rect 9140 -11880 9260 -11760
rect 9315 -11880 9435 -11760
rect 9480 -11880 9600 -11760
rect 9645 -11880 9765 -11760
rect 9810 -11880 9930 -11760
rect 9985 -11880 10105 -11760
rect 10150 -11880 10270 -11760
rect 10315 -11880 10435 -11760
rect 10480 -11880 10600 -11760
rect 10655 -11880 10775 -11760
rect 10820 -11880 10940 -11760
rect 10985 -11880 11105 -11760
rect 11150 -11880 11270 -11760
rect 11325 -11880 11445 -11760
rect 11490 -11880 11610 -11760
rect 11655 -11880 11775 -11760
rect 11820 -11880 11940 -11760
rect 11995 -11880 12115 -11760
rect 12160 -11880 12280 -11760
rect 12325 -11880 12445 -11760
rect 12490 -11880 12610 -11760
rect 7130 -12045 7250 -11925
rect 7305 -12045 7425 -11925
rect 7470 -12045 7590 -11925
rect 7635 -12045 7755 -11925
rect 7800 -12045 7920 -11925
rect 7975 -12045 8095 -11925
rect 8140 -12045 8260 -11925
rect 8305 -12045 8425 -11925
rect 8470 -12045 8590 -11925
rect 8645 -12045 8765 -11925
rect 8810 -12045 8930 -11925
rect 8975 -12045 9095 -11925
rect 9140 -12045 9260 -11925
rect 9315 -12045 9435 -11925
rect 9480 -12045 9600 -11925
rect 9645 -12045 9765 -11925
rect 9810 -12045 9930 -11925
rect 9985 -12045 10105 -11925
rect 10150 -12045 10270 -11925
rect 10315 -12045 10435 -11925
rect 10480 -12045 10600 -11925
rect 10655 -12045 10775 -11925
rect 10820 -12045 10940 -11925
rect 10985 -12045 11105 -11925
rect 11150 -12045 11270 -11925
rect 11325 -12045 11445 -11925
rect 11490 -12045 11610 -11925
rect 11655 -12045 11775 -11925
rect 11820 -12045 11940 -11925
rect 11995 -12045 12115 -11925
rect 12160 -12045 12280 -11925
rect 12325 -12045 12445 -11925
rect 12490 -12045 12610 -11925
rect 7130 -12220 7250 -12100
rect 7305 -12220 7425 -12100
rect 7470 -12220 7590 -12100
rect 7635 -12220 7755 -12100
rect 7800 -12220 7920 -12100
rect 7975 -12220 8095 -12100
rect 8140 -12220 8260 -12100
rect 8305 -12220 8425 -12100
rect 8470 -12220 8590 -12100
rect 8645 -12220 8765 -12100
rect 8810 -12220 8930 -12100
rect 8975 -12220 9095 -12100
rect 9140 -12220 9260 -12100
rect 9315 -12220 9435 -12100
rect 9480 -12220 9600 -12100
rect 9645 -12220 9765 -12100
rect 9810 -12220 9930 -12100
rect 9985 -12220 10105 -12100
rect 10150 -12220 10270 -12100
rect 10315 -12220 10435 -12100
rect 10480 -12220 10600 -12100
rect 10655 -12220 10775 -12100
rect 10820 -12220 10940 -12100
rect 10985 -12220 11105 -12100
rect 11150 -12220 11270 -12100
rect 11325 -12220 11445 -12100
rect 11490 -12220 11610 -12100
rect 11655 -12220 11775 -12100
rect 11820 -12220 11940 -12100
rect 11995 -12220 12115 -12100
rect 12160 -12220 12280 -12100
rect 12325 -12220 12445 -12100
rect 12490 -12220 12610 -12100
rect 7130 -12385 7250 -12265
rect 7305 -12385 7425 -12265
rect 7470 -12385 7590 -12265
rect 7635 -12385 7755 -12265
rect 7800 -12385 7920 -12265
rect 7975 -12385 8095 -12265
rect 8140 -12385 8260 -12265
rect 8305 -12385 8425 -12265
rect 8470 -12385 8590 -12265
rect 8645 -12385 8765 -12265
rect 8810 -12385 8930 -12265
rect 8975 -12385 9095 -12265
rect 9140 -12385 9260 -12265
rect 9315 -12385 9435 -12265
rect 9480 -12385 9600 -12265
rect 9645 -12385 9765 -12265
rect 9810 -12385 9930 -12265
rect 9985 -12385 10105 -12265
rect 10150 -12385 10270 -12265
rect 10315 -12385 10435 -12265
rect 10480 -12385 10600 -12265
rect 10655 -12385 10775 -12265
rect 10820 -12385 10940 -12265
rect 10985 -12385 11105 -12265
rect 11150 -12385 11270 -12265
rect 11325 -12385 11445 -12265
rect 11490 -12385 11610 -12265
rect 11655 -12385 11775 -12265
rect 11820 -12385 11940 -12265
rect 11995 -12385 12115 -12265
rect 12160 -12385 12280 -12265
rect 12325 -12385 12445 -12265
rect 12490 -12385 12610 -12265
rect 7130 -12550 7250 -12430
rect 7305 -12550 7425 -12430
rect 7470 -12550 7590 -12430
rect 7635 -12550 7755 -12430
rect 7800 -12550 7920 -12430
rect 7975 -12550 8095 -12430
rect 8140 -12550 8260 -12430
rect 8305 -12550 8425 -12430
rect 8470 -12550 8590 -12430
rect 8645 -12550 8765 -12430
rect 8810 -12550 8930 -12430
rect 8975 -12550 9095 -12430
rect 9140 -12550 9260 -12430
rect 9315 -12550 9435 -12430
rect 9480 -12550 9600 -12430
rect 9645 -12550 9765 -12430
rect 9810 -12550 9930 -12430
rect 9985 -12550 10105 -12430
rect 10150 -12550 10270 -12430
rect 10315 -12550 10435 -12430
rect 10480 -12550 10600 -12430
rect 10655 -12550 10775 -12430
rect 10820 -12550 10940 -12430
rect 10985 -12550 11105 -12430
rect 11150 -12550 11270 -12430
rect 11325 -12550 11445 -12430
rect 11490 -12550 11610 -12430
rect 11655 -12550 11775 -12430
rect 11820 -12550 11940 -12430
rect 11995 -12550 12115 -12430
rect 12160 -12550 12280 -12430
rect 12325 -12550 12445 -12430
rect 12490 -12550 12610 -12430
rect 7130 -12715 7250 -12595
rect 7305 -12715 7425 -12595
rect 7470 -12715 7590 -12595
rect 7635 -12715 7755 -12595
rect 7800 -12715 7920 -12595
rect 7975 -12715 8095 -12595
rect 8140 -12715 8260 -12595
rect 8305 -12715 8425 -12595
rect 8470 -12715 8590 -12595
rect 8645 -12715 8765 -12595
rect 8810 -12715 8930 -12595
rect 8975 -12715 9095 -12595
rect 9140 -12715 9260 -12595
rect 9315 -12715 9435 -12595
rect 9480 -12715 9600 -12595
rect 9645 -12715 9765 -12595
rect 9810 -12715 9930 -12595
rect 9985 -12715 10105 -12595
rect 10150 -12715 10270 -12595
rect 10315 -12715 10435 -12595
rect 10480 -12715 10600 -12595
rect 10655 -12715 10775 -12595
rect 10820 -12715 10940 -12595
rect 10985 -12715 11105 -12595
rect 11150 -12715 11270 -12595
rect 11325 -12715 11445 -12595
rect 11490 -12715 11610 -12595
rect 11655 -12715 11775 -12595
rect 11820 -12715 11940 -12595
rect 11995 -12715 12115 -12595
rect 12160 -12715 12280 -12595
rect 12325 -12715 12445 -12595
rect 12490 -12715 12610 -12595
rect 7130 -12890 7250 -12770
rect 7305 -12890 7425 -12770
rect 7470 -12890 7590 -12770
rect 7635 -12890 7755 -12770
rect 7800 -12890 7920 -12770
rect 7975 -12890 8095 -12770
rect 8140 -12890 8260 -12770
rect 8305 -12890 8425 -12770
rect 8470 -12890 8590 -12770
rect 8645 -12890 8765 -12770
rect 8810 -12890 8930 -12770
rect 8975 -12890 9095 -12770
rect 9140 -12890 9260 -12770
rect 9315 -12890 9435 -12770
rect 9480 -12890 9600 -12770
rect 9645 -12890 9765 -12770
rect 9810 -12890 9930 -12770
rect 9985 -12890 10105 -12770
rect 10150 -12890 10270 -12770
rect 10315 -12890 10435 -12770
rect 10480 -12890 10600 -12770
rect 10655 -12890 10775 -12770
rect 10820 -12890 10940 -12770
rect 10985 -12890 11105 -12770
rect 11150 -12890 11270 -12770
rect 11325 -12890 11445 -12770
rect 11490 -12890 11610 -12770
rect 11655 -12890 11775 -12770
rect 11820 -12890 11940 -12770
rect 11995 -12890 12115 -12770
rect 12160 -12890 12280 -12770
rect 12325 -12890 12445 -12770
rect 12490 -12890 12610 -12770
rect 7130 -13055 7250 -12935
rect 7305 -13055 7425 -12935
rect 7470 -13055 7590 -12935
rect 7635 -13055 7755 -12935
rect 7800 -13055 7920 -12935
rect 7975 -13055 8095 -12935
rect 8140 -13055 8260 -12935
rect 8305 -13055 8425 -12935
rect 8470 -13055 8590 -12935
rect 8645 -13055 8765 -12935
rect 8810 -13055 8930 -12935
rect 8975 -13055 9095 -12935
rect 9140 -13055 9260 -12935
rect 9315 -13055 9435 -12935
rect 9480 -13055 9600 -12935
rect 9645 -13055 9765 -12935
rect 9810 -13055 9930 -12935
rect 9985 -13055 10105 -12935
rect 10150 -13055 10270 -12935
rect 10315 -13055 10435 -12935
rect 10480 -13055 10600 -12935
rect 10655 -13055 10775 -12935
rect 10820 -13055 10940 -12935
rect 10985 -13055 11105 -12935
rect 11150 -13055 11270 -12935
rect 11325 -13055 11445 -12935
rect 11490 -13055 11610 -12935
rect 11655 -13055 11775 -12935
rect 11820 -13055 11940 -12935
rect 11995 -13055 12115 -12935
rect 12160 -13055 12280 -12935
rect 12325 -13055 12445 -12935
rect 12490 -13055 12610 -12935
rect 7130 -13220 7250 -13100
rect 7305 -13220 7425 -13100
rect 7470 -13220 7590 -13100
rect 7635 -13220 7755 -13100
rect 7800 -13220 7920 -13100
rect 7975 -13220 8095 -13100
rect 8140 -13220 8260 -13100
rect 8305 -13220 8425 -13100
rect 8470 -13220 8590 -13100
rect 8645 -13220 8765 -13100
rect 8810 -13220 8930 -13100
rect 8975 -13220 9095 -13100
rect 9140 -13220 9260 -13100
rect 9315 -13220 9435 -13100
rect 9480 -13220 9600 -13100
rect 9645 -13220 9765 -13100
rect 9810 -13220 9930 -13100
rect 9985 -13220 10105 -13100
rect 10150 -13220 10270 -13100
rect 10315 -13220 10435 -13100
rect 10480 -13220 10600 -13100
rect 10655 -13220 10775 -13100
rect 10820 -13220 10940 -13100
rect 10985 -13220 11105 -13100
rect 11150 -13220 11270 -13100
rect 11325 -13220 11445 -13100
rect 11490 -13220 11610 -13100
rect 11655 -13220 11775 -13100
rect 11820 -13220 11940 -13100
rect 11995 -13220 12115 -13100
rect 12160 -13220 12280 -13100
rect 12325 -13220 12445 -13100
rect 12490 -13220 12610 -13100
rect 7130 -13385 7250 -13265
rect 7305 -13385 7425 -13265
rect 7470 -13385 7590 -13265
rect 7635 -13385 7755 -13265
rect 7800 -13385 7920 -13265
rect 7975 -13385 8095 -13265
rect 8140 -13385 8260 -13265
rect 8305 -13385 8425 -13265
rect 8470 -13385 8590 -13265
rect 8645 -13385 8765 -13265
rect 8810 -13385 8930 -13265
rect 8975 -13385 9095 -13265
rect 9140 -13385 9260 -13265
rect 9315 -13385 9435 -13265
rect 9480 -13385 9600 -13265
rect 9645 -13385 9765 -13265
rect 9810 -13385 9930 -13265
rect 9985 -13385 10105 -13265
rect 10150 -13385 10270 -13265
rect 10315 -13385 10435 -13265
rect 10480 -13385 10600 -13265
rect 10655 -13385 10775 -13265
rect 10820 -13385 10940 -13265
rect 10985 -13385 11105 -13265
rect 11150 -13385 11270 -13265
rect 11325 -13385 11445 -13265
rect 11490 -13385 11610 -13265
rect 11655 -13385 11775 -13265
rect 11820 -13385 11940 -13265
rect 11995 -13385 12115 -13265
rect 12160 -13385 12280 -13265
rect 12325 -13385 12445 -13265
rect 12490 -13385 12610 -13265
rect 7130 -13560 7250 -13440
rect 7305 -13560 7425 -13440
rect 7470 -13560 7590 -13440
rect 7635 -13560 7755 -13440
rect 7800 -13560 7920 -13440
rect 7975 -13560 8095 -13440
rect 8140 -13560 8260 -13440
rect 8305 -13560 8425 -13440
rect 8470 -13560 8590 -13440
rect 8645 -13560 8765 -13440
rect 8810 -13560 8930 -13440
rect 8975 -13560 9095 -13440
rect 9140 -13560 9260 -13440
rect 9315 -13560 9435 -13440
rect 9480 -13560 9600 -13440
rect 9645 -13560 9765 -13440
rect 9810 -13560 9930 -13440
rect 9985 -13560 10105 -13440
rect 10150 -13560 10270 -13440
rect 10315 -13560 10435 -13440
rect 10480 -13560 10600 -13440
rect 10655 -13560 10775 -13440
rect 10820 -13560 10940 -13440
rect 10985 -13560 11105 -13440
rect 11150 -13560 11270 -13440
rect 11325 -13560 11445 -13440
rect 11490 -13560 11610 -13440
rect 11655 -13560 11775 -13440
rect 11820 -13560 11940 -13440
rect 11995 -13560 12115 -13440
rect 12160 -13560 12280 -13440
rect 12325 -13560 12445 -13440
rect 12490 -13560 12610 -13440
rect 7130 -13725 7250 -13605
rect 7305 -13725 7425 -13605
rect 7470 -13725 7590 -13605
rect 7635 -13725 7755 -13605
rect 7800 -13725 7920 -13605
rect 7975 -13725 8095 -13605
rect 8140 -13725 8260 -13605
rect 8305 -13725 8425 -13605
rect 8470 -13725 8590 -13605
rect 8645 -13725 8765 -13605
rect 8810 -13725 8930 -13605
rect 8975 -13725 9095 -13605
rect 9140 -13725 9260 -13605
rect 9315 -13725 9435 -13605
rect 9480 -13725 9600 -13605
rect 9645 -13725 9765 -13605
rect 9810 -13725 9930 -13605
rect 9985 -13725 10105 -13605
rect 10150 -13725 10270 -13605
rect 10315 -13725 10435 -13605
rect 10480 -13725 10600 -13605
rect 10655 -13725 10775 -13605
rect 10820 -13725 10940 -13605
rect 10985 -13725 11105 -13605
rect 11150 -13725 11270 -13605
rect 11325 -13725 11445 -13605
rect 11490 -13725 11610 -13605
rect 11655 -13725 11775 -13605
rect 11820 -13725 11940 -13605
rect 11995 -13725 12115 -13605
rect 12160 -13725 12280 -13605
rect 12325 -13725 12445 -13605
rect 12490 -13725 12610 -13605
rect 7130 -13890 7250 -13770
rect 7305 -13890 7425 -13770
rect 7470 -13890 7590 -13770
rect 7635 -13890 7755 -13770
rect 7800 -13890 7920 -13770
rect 7975 -13890 8095 -13770
rect 8140 -13890 8260 -13770
rect 8305 -13890 8425 -13770
rect 8470 -13890 8590 -13770
rect 8645 -13890 8765 -13770
rect 8810 -13890 8930 -13770
rect 8975 -13890 9095 -13770
rect 9140 -13890 9260 -13770
rect 9315 -13890 9435 -13770
rect 9480 -13890 9600 -13770
rect 9645 -13890 9765 -13770
rect 9810 -13890 9930 -13770
rect 9985 -13890 10105 -13770
rect 10150 -13890 10270 -13770
rect 10315 -13890 10435 -13770
rect 10480 -13890 10600 -13770
rect 10655 -13890 10775 -13770
rect 10820 -13890 10940 -13770
rect 10985 -13890 11105 -13770
rect 11150 -13890 11270 -13770
rect 11325 -13890 11445 -13770
rect 11490 -13890 11610 -13770
rect 11655 -13890 11775 -13770
rect 11820 -13890 11940 -13770
rect 11995 -13890 12115 -13770
rect 12160 -13890 12280 -13770
rect 12325 -13890 12445 -13770
rect 12490 -13890 12610 -13770
rect 7130 -14055 7250 -13935
rect 7305 -14055 7425 -13935
rect 7470 -14055 7590 -13935
rect 7635 -14055 7755 -13935
rect 7800 -14055 7920 -13935
rect 7975 -14055 8095 -13935
rect 8140 -14055 8260 -13935
rect 8305 -14055 8425 -13935
rect 8470 -14055 8590 -13935
rect 8645 -14055 8765 -13935
rect 8810 -14055 8930 -13935
rect 8975 -14055 9095 -13935
rect 9140 -14055 9260 -13935
rect 9315 -14055 9435 -13935
rect 9480 -14055 9600 -13935
rect 9645 -14055 9765 -13935
rect 9810 -14055 9930 -13935
rect 9985 -14055 10105 -13935
rect 10150 -14055 10270 -13935
rect 10315 -14055 10435 -13935
rect 10480 -14055 10600 -13935
rect 10655 -14055 10775 -13935
rect 10820 -14055 10940 -13935
rect 10985 -14055 11105 -13935
rect 11150 -14055 11270 -13935
rect 11325 -14055 11445 -13935
rect 11490 -14055 11610 -13935
rect 11655 -14055 11775 -13935
rect 11820 -14055 11940 -13935
rect 11995 -14055 12115 -13935
rect 12160 -14055 12280 -13935
rect 12325 -14055 12445 -13935
rect 12490 -14055 12610 -13935
rect 7130 -14230 7250 -14110
rect 7305 -14230 7425 -14110
rect 7470 -14230 7590 -14110
rect 7635 -14230 7755 -14110
rect 7800 -14230 7920 -14110
rect 7975 -14230 8095 -14110
rect 8140 -14230 8260 -14110
rect 8305 -14230 8425 -14110
rect 8470 -14230 8590 -14110
rect 8645 -14230 8765 -14110
rect 8810 -14230 8930 -14110
rect 8975 -14230 9095 -14110
rect 9140 -14230 9260 -14110
rect 9315 -14230 9435 -14110
rect 9480 -14230 9600 -14110
rect 9645 -14230 9765 -14110
rect 9810 -14230 9930 -14110
rect 9985 -14230 10105 -14110
rect 10150 -14230 10270 -14110
rect 10315 -14230 10435 -14110
rect 10480 -14230 10600 -14110
rect 10655 -14230 10775 -14110
rect 10820 -14230 10940 -14110
rect 10985 -14230 11105 -14110
rect 11150 -14230 11270 -14110
rect 11325 -14230 11445 -14110
rect 11490 -14230 11610 -14110
rect 11655 -14230 11775 -14110
rect 11820 -14230 11940 -14110
rect 11995 -14230 12115 -14110
rect 12160 -14230 12280 -14110
rect 12325 -14230 12445 -14110
rect 12490 -14230 12610 -14110
rect 7130 -14395 7250 -14275
rect 7305 -14395 7425 -14275
rect 7470 -14395 7590 -14275
rect 7635 -14395 7755 -14275
rect 7800 -14395 7920 -14275
rect 7975 -14395 8095 -14275
rect 8140 -14395 8260 -14275
rect 8305 -14395 8425 -14275
rect 8470 -14395 8590 -14275
rect 8645 -14395 8765 -14275
rect 8810 -14395 8930 -14275
rect 8975 -14395 9095 -14275
rect 9140 -14395 9260 -14275
rect 9315 -14395 9435 -14275
rect 9480 -14395 9600 -14275
rect 9645 -14395 9765 -14275
rect 9810 -14395 9930 -14275
rect 9985 -14395 10105 -14275
rect 10150 -14395 10270 -14275
rect 10315 -14395 10435 -14275
rect 10480 -14395 10600 -14275
rect 10655 -14395 10775 -14275
rect 10820 -14395 10940 -14275
rect 10985 -14395 11105 -14275
rect 11150 -14395 11270 -14275
rect 11325 -14395 11445 -14275
rect 11490 -14395 11610 -14275
rect 11655 -14395 11775 -14275
rect 11820 -14395 11940 -14275
rect 11995 -14395 12115 -14275
rect 12160 -14395 12280 -14275
rect 12325 -14395 12445 -14275
rect 12490 -14395 12610 -14275
rect 7130 -14560 7250 -14440
rect 7305 -14560 7425 -14440
rect 7470 -14560 7590 -14440
rect 7635 -14560 7755 -14440
rect 7800 -14560 7920 -14440
rect 7975 -14560 8095 -14440
rect 8140 -14560 8260 -14440
rect 8305 -14560 8425 -14440
rect 8470 -14560 8590 -14440
rect 8645 -14560 8765 -14440
rect 8810 -14560 8930 -14440
rect 8975 -14560 9095 -14440
rect 9140 -14560 9260 -14440
rect 9315 -14560 9435 -14440
rect 9480 -14560 9600 -14440
rect 9645 -14560 9765 -14440
rect 9810 -14560 9930 -14440
rect 9985 -14560 10105 -14440
rect 10150 -14560 10270 -14440
rect 10315 -14560 10435 -14440
rect 10480 -14560 10600 -14440
rect 10655 -14560 10775 -14440
rect 10820 -14560 10940 -14440
rect 10985 -14560 11105 -14440
rect 11150 -14560 11270 -14440
rect 11325 -14560 11445 -14440
rect 11490 -14560 11610 -14440
rect 11655 -14560 11775 -14440
rect 11820 -14560 11940 -14440
rect 11995 -14560 12115 -14440
rect 12160 -14560 12280 -14440
rect 12325 -14560 12445 -14440
rect 12490 -14560 12610 -14440
rect 7130 -14725 7250 -14605
rect 7305 -14725 7425 -14605
rect 7470 -14725 7590 -14605
rect 7635 -14725 7755 -14605
rect 7800 -14725 7920 -14605
rect 7975 -14725 8095 -14605
rect 8140 -14725 8260 -14605
rect 8305 -14725 8425 -14605
rect 8470 -14725 8590 -14605
rect 8645 -14725 8765 -14605
rect 8810 -14725 8930 -14605
rect 8975 -14725 9095 -14605
rect 9140 -14725 9260 -14605
rect 9315 -14725 9435 -14605
rect 9480 -14725 9600 -14605
rect 9645 -14725 9765 -14605
rect 9810 -14725 9930 -14605
rect 9985 -14725 10105 -14605
rect 10150 -14725 10270 -14605
rect 10315 -14725 10435 -14605
rect 10480 -14725 10600 -14605
rect 10655 -14725 10775 -14605
rect 10820 -14725 10940 -14605
rect 10985 -14725 11105 -14605
rect 11150 -14725 11270 -14605
rect 11325 -14725 11445 -14605
rect 11490 -14725 11610 -14605
rect 11655 -14725 11775 -14605
rect 11820 -14725 11940 -14605
rect 11995 -14725 12115 -14605
rect 12160 -14725 12280 -14605
rect 12325 -14725 12445 -14605
rect 12490 -14725 12610 -14605
rect 7130 -14900 7250 -14780
rect 7305 -14900 7425 -14780
rect 7470 -14900 7590 -14780
rect 7635 -14900 7755 -14780
rect 7800 -14900 7920 -14780
rect 7975 -14900 8095 -14780
rect 8140 -14900 8260 -14780
rect 8305 -14900 8425 -14780
rect 8470 -14900 8590 -14780
rect 8645 -14900 8765 -14780
rect 8810 -14900 8930 -14780
rect 8975 -14900 9095 -14780
rect 9140 -14900 9260 -14780
rect 9315 -14900 9435 -14780
rect 9480 -14900 9600 -14780
rect 9645 -14900 9765 -14780
rect 9810 -14900 9930 -14780
rect 9985 -14900 10105 -14780
rect 10150 -14900 10270 -14780
rect 10315 -14900 10435 -14780
rect 10480 -14900 10600 -14780
rect 10655 -14900 10775 -14780
rect 10820 -14900 10940 -14780
rect 10985 -14900 11105 -14780
rect 11150 -14900 11270 -14780
rect 11325 -14900 11445 -14780
rect 11490 -14900 11610 -14780
rect 11655 -14900 11775 -14780
rect 11820 -14900 11940 -14780
rect 11995 -14900 12115 -14780
rect 12160 -14900 12280 -14780
rect 12325 -14900 12445 -14780
rect 12490 -14900 12610 -14780
rect 7130 -15065 7250 -14945
rect 7305 -15065 7425 -14945
rect 7470 -15065 7590 -14945
rect 7635 -15065 7755 -14945
rect 7800 -15065 7920 -14945
rect 7975 -15065 8095 -14945
rect 8140 -15065 8260 -14945
rect 8305 -15065 8425 -14945
rect 8470 -15065 8590 -14945
rect 8645 -15065 8765 -14945
rect 8810 -15065 8930 -14945
rect 8975 -15065 9095 -14945
rect 9140 -15065 9260 -14945
rect 9315 -15065 9435 -14945
rect 9480 -15065 9600 -14945
rect 9645 -15065 9765 -14945
rect 9810 -15065 9930 -14945
rect 9985 -15065 10105 -14945
rect 10150 -15065 10270 -14945
rect 10315 -15065 10435 -14945
rect 10480 -15065 10600 -14945
rect 10655 -15065 10775 -14945
rect 10820 -15065 10940 -14945
rect 10985 -15065 11105 -14945
rect 11150 -15065 11270 -14945
rect 11325 -15065 11445 -14945
rect 11490 -15065 11610 -14945
rect 11655 -15065 11775 -14945
rect 11820 -15065 11940 -14945
rect 11995 -15065 12115 -14945
rect 12160 -15065 12280 -14945
rect 12325 -15065 12445 -14945
rect 12490 -15065 12610 -14945
rect 7130 -15230 7250 -15110
rect 7305 -15230 7425 -15110
rect 7470 -15230 7590 -15110
rect 7635 -15230 7755 -15110
rect 7800 -15230 7920 -15110
rect 7975 -15230 8095 -15110
rect 8140 -15230 8260 -15110
rect 8305 -15230 8425 -15110
rect 8470 -15230 8590 -15110
rect 8645 -15230 8765 -15110
rect 8810 -15230 8930 -15110
rect 8975 -15230 9095 -15110
rect 9140 -15230 9260 -15110
rect 9315 -15230 9435 -15110
rect 9480 -15230 9600 -15110
rect 9645 -15230 9765 -15110
rect 9810 -15230 9930 -15110
rect 9985 -15230 10105 -15110
rect 10150 -15230 10270 -15110
rect 10315 -15230 10435 -15110
rect 10480 -15230 10600 -15110
rect 10655 -15230 10775 -15110
rect 10820 -15230 10940 -15110
rect 10985 -15230 11105 -15110
rect 11150 -15230 11270 -15110
rect 11325 -15230 11445 -15110
rect 11490 -15230 11610 -15110
rect 11655 -15230 11775 -15110
rect 11820 -15230 11940 -15110
rect 11995 -15230 12115 -15110
rect 12160 -15230 12280 -15110
rect 12325 -15230 12445 -15110
rect 12490 -15230 12610 -15110
rect 7130 -15395 7250 -15275
rect 7305 -15395 7425 -15275
rect 7470 -15395 7590 -15275
rect 7635 -15395 7755 -15275
rect 7800 -15395 7920 -15275
rect 7975 -15395 8095 -15275
rect 8140 -15395 8260 -15275
rect 8305 -15395 8425 -15275
rect 8470 -15395 8590 -15275
rect 8645 -15395 8765 -15275
rect 8810 -15395 8930 -15275
rect 8975 -15395 9095 -15275
rect 9140 -15395 9260 -15275
rect 9315 -15395 9435 -15275
rect 9480 -15395 9600 -15275
rect 9645 -15395 9765 -15275
rect 9810 -15395 9930 -15275
rect 9985 -15395 10105 -15275
rect 10150 -15395 10270 -15275
rect 10315 -15395 10435 -15275
rect 10480 -15395 10600 -15275
rect 10655 -15395 10775 -15275
rect 10820 -15395 10940 -15275
rect 10985 -15395 11105 -15275
rect 11150 -15395 11270 -15275
rect 11325 -15395 11445 -15275
rect 11490 -15395 11610 -15275
rect 11655 -15395 11775 -15275
rect 11820 -15395 11940 -15275
rect 11995 -15395 12115 -15275
rect 12160 -15395 12280 -15275
rect 12325 -15395 12445 -15275
rect 12490 -15395 12610 -15275
rect 7130 -15570 7250 -15450
rect 7305 -15570 7425 -15450
rect 7470 -15570 7590 -15450
rect 7635 -15570 7755 -15450
rect 7800 -15570 7920 -15450
rect 7975 -15570 8095 -15450
rect 8140 -15570 8260 -15450
rect 8305 -15570 8425 -15450
rect 8470 -15570 8590 -15450
rect 8645 -15570 8765 -15450
rect 8810 -15570 8930 -15450
rect 8975 -15570 9095 -15450
rect 9140 -15570 9260 -15450
rect 9315 -15570 9435 -15450
rect 9480 -15570 9600 -15450
rect 9645 -15570 9765 -15450
rect 9810 -15570 9930 -15450
rect 9985 -15570 10105 -15450
rect 10150 -15570 10270 -15450
rect 10315 -15570 10435 -15450
rect 10480 -15570 10600 -15450
rect 10655 -15570 10775 -15450
rect 10820 -15570 10940 -15450
rect 10985 -15570 11105 -15450
rect 11150 -15570 11270 -15450
rect 11325 -15570 11445 -15450
rect 11490 -15570 11610 -15450
rect 11655 -15570 11775 -15450
rect 11820 -15570 11940 -15450
rect 11995 -15570 12115 -15450
rect 12160 -15570 12280 -15450
rect 12325 -15570 12445 -15450
rect 12490 -15570 12610 -15450
rect 12820 -10210 12940 -10090
rect 12995 -10210 13115 -10090
rect 13160 -10210 13280 -10090
rect 13325 -10210 13445 -10090
rect 13490 -10210 13610 -10090
rect 13665 -10210 13785 -10090
rect 13830 -10210 13950 -10090
rect 13995 -10210 14115 -10090
rect 14160 -10210 14280 -10090
rect 14335 -10210 14455 -10090
rect 14500 -10210 14620 -10090
rect 14665 -10210 14785 -10090
rect 14830 -10210 14950 -10090
rect 15005 -10210 15125 -10090
rect 15170 -10210 15290 -10090
rect 15335 -10210 15455 -10090
rect 15500 -10210 15620 -10090
rect 15675 -10210 15795 -10090
rect 15840 -10210 15960 -10090
rect 16005 -10210 16125 -10090
rect 16170 -10210 16290 -10090
rect 16345 -10210 16465 -10090
rect 16510 -10210 16630 -10090
rect 16675 -10210 16795 -10090
rect 16840 -10210 16960 -10090
rect 17015 -10210 17135 -10090
rect 17180 -10210 17300 -10090
rect 17345 -10210 17465 -10090
rect 17510 -10210 17630 -10090
rect 17685 -10210 17805 -10090
rect 17850 -10210 17970 -10090
rect 18015 -10210 18135 -10090
rect 18180 -10210 18300 -10090
rect 12820 -10375 12940 -10255
rect 12995 -10375 13115 -10255
rect 13160 -10375 13280 -10255
rect 13325 -10375 13445 -10255
rect 13490 -10375 13610 -10255
rect 13665 -10375 13785 -10255
rect 13830 -10375 13950 -10255
rect 13995 -10375 14115 -10255
rect 14160 -10375 14280 -10255
rect 14335 -10375 14455 -10255
rect 14500 -10375 14620 -10255
rect 14665 -10375 14785 -10255
rect 14830 -10375 14950 -10255
rect 15005 -10375 15125 -10255
rect 15170 -10375 15290 -10255
rect 15335 -10375 15455 -10255
rect 15500 -10375 15620 -10255
rect 15675 -10375 15795 -10255
rect 15840 -10375 15960 -10255
rect 16005 -10375 16125 -10255
rect 16170 -10375 16290 -10255
rect 16345 -10375 16465 -10255
rect 16510 -10375 16630 -10255
rect 16675 -10375 16795 -10255
rect 16840 -10375 16960 -10255
rect 17015 -10375 17135 -10255
rect 17180 -10375 17300 -10255
rect 17345 -10375 17465 -10255
rect 17510 -10375 17630 -10255
rect 17685 -10375 17805 -10255
rect 17850 -10375 17970 -10255
rect 18015 -10375 18135 -10255
rect 18180 -10375 18300 -10255
rect 12820 -10540 12940 -10420
rect 12995 -10540 13115 -10420
rect 13160 -10540 13280 -10420
rect 13325 -10540 13445 -10420
rect 13490 -10540 13610 -10420
rect 13665 -10540 13785 -10420
rect 13830 -10540 13950 -10420
rect 13995 -10540 14115 -10420
rect 14160 -10540 14280 -10420
rect 14335 -10540 14455 -10420
rect 14500 -10540 14620 -10420
rect 14665 -10540 14785 -10420
rect 14830 -10540 14950 -10420
rect 15005 -10540 15125 -10420
rect 15170 -10540 15290 -10420
rect 15335 -10540 15455 -10420
rect 15500 -10540 15620 -10420
rect 15675 -10540 15795 -10420
rect 15840 -10540 15960 -10420
rect 16005 -10540 16125 -10420
rect 16170 -10540 16290 -10420
rect 16345 -10540 16465 -10420
rect 16510 -10540 16630 -10420
rect 16675 -10540 16795 -10420
rect 16840 -10540 16960 -10420
rect 17015 -10540 17135 -10420
rect 17180 -10540 17300 -10420
rect 17345 -10540 17465 -10420
rect 17510 -10540 17630 -10420
rect 17685 -10540 17805 -10420
rect 17850 -10540 17970 -10420
rect 18015 -10540 18135 -10420
rect 18180 -10540 18300 -10420
rect 12820 -10705 12940 -10585
rect 12995 -10705 13115 -10585
rect 13160 -10705 13280 -10585
rect 13325 -10705 13445 -10585
rect 13490 -10705 13610 -10585
rect 13665 -10705 13785 -10585
rect 13830 -10705 13950 -10585
rect 13995 -10705 14115 -10585
rect 14160 -10705 14280 -10585
rect 14335 -10705 14455 -10585
rect 14500 -10705 14620 -10585
rect 14665 -10705 14785 -10585
rect 14830 -10705 14950 -10585
rect 15005 -10705 15125 -10585
rect 15170 -10705 15290 -10585
rect 15335 -10705 15455 -10585
rect 15500 -10705 15620 -10585
rect 15675 -10705 15795 -10585
rect 15840 -10705 15960 -10585
rect 16005 -10705 16125 -10585
rect 16170 -10705 16290 -10585
rect 16345 -10705 16465 -10585
rect 16510 -10705 16630 -10585
rect 16675 -10705 16795 -10585
rect 16840 -10705 16960 -10585
rect 17015 -10705 17135 -10585
rect 17180 -10705 17300 -10585
rect 17345 -10705 17465 -10585
rect 17510 -10705 17630 -10585
rect 17685 -10705 17805 -10585
rect 17850 -10705 17970 -10585
rect 18015 -10705 18135 -10585
rect 18180 -10705 18300 -10585
rect 12820 -10880 12940 -10760
rect 12995 -10880 13115 -10760
rect 13160 -10880 13280 -10760
rect 13325 -10880 13445 -10760
rect 13490 -10880 13610 -10760
rect 13665 -10880 13785 -10760
rect 13830 -10880 13950 -10760
rect 13995 -10880 14115 -10760
rect 14160 -10880 14280 -10760
rect 14335 -10880 14455 -10760
rect 14500 -10880 14620 -10760
rect 14665 -10880 14785 -10760
rect 14830 -10880 14950 -10760
rect 15005 -10880 15125 -10760
rect 15170 -10880 15290 -10760
rect 15335 -10880 15455 -10760
rect 15500 -10880 15620 -10760
rect 15675 -10880 15795 -10760
rect 15840 -10880 15960 -10760
rect 16005 -10880 16125 -10760
rect 16170 -10880 16290 -10760
rect 16345 -10880 16465 -10760
rect 16510 -10880 16630 -10760
rect 16675 -10880 16795 -10760
rect 16840 -10880 16960 -10760
rect 17015 -10880 17135 -10760
rect 17180 -10880 17300 -10760
rect 17345 -10880 17465 -10760
rect 17510 -10880 17630 -10760
rect 17685 -10880 17805 -10760
rect 17850 -10880 17970 -10760
rect 18015 -10880 18135 -10760
rect 18180 -10880 18300 -10760
rect 12820 -11045 12940 -10925
rect 12995 -11045 13115 -10925
rect 13160 -11045 13280 -10925
rect 13325 -11045 13445 -10925
rect 13490 -11045 13610 -10925
rect 13665 -11045 13785 -10925
rect 13830 -11045 13950 -10925
rect 13995 -11045 14115 -10925
rect 14160 -11045 14280 -10925
rect 14335 -11045 14455 -10925
rect 14500 -11045 14620 -10925
rect 14665 -11045 14785 -10925
rect 14830 -11045 14950 -10925
rect 15005 -11045 15125 -10925
rect 15170 -11045 15290 -10925
rect 15335 -11045 15455 -10925
rect 15500 -11045 15620 -10925
rect 15675 -11045 15795 -10925
rect 15840 -11045 15960 -10925
rect 16005 -11045 16125 -10925
rect 16170 -11045 16290 -10925
rect 16345 -11045 16465 -10925
rect 16510 -11045 16630 -10925
rect 16675 -11045 16795 -10925
rect 16840 -11045 16960 -10925
rect 17015 -11045 17135 -10925
rect 17180 -11045 17300 -10925
rect 17345 -11045 17465 -10925
rect 17510 -11045 17630 -10925
rect 17685 -11045 17805 -10925
rect 17850 -11045 17970 -10925
rect 18015 -11045 18135 -10925
rect 18180 -11045 18300 -10925
rect 12820 -11210 12940 -11090
rect 12995 -11210 13115 -11090
rect 13160 -11210 13280 -11090
rect 13325 -11210 13445 -11090
rect 13490 -11210 13610 -11090
rect 13665 -11210 13785 -11090
rect 13830 -11210 13950 -11090
rect 13995 -11210 14115 -11090
rect 14160 -11210 14280 -11090
rect 14335 -11210 14455 -11090
rect 14500 -11210 14620 -11090
rect 14665 -11210 14785 -11090
rect 14830 -11210 14950 -11090
rect 15005 -11210 15125 -11090
rect 15170 -11210 15290 -11090
rect 15335 -11210 15455 -11090
rect 15500 -11210 15620 -11090
rect 15675 -11210 15795 -11090
rect 15840 -11210 15960 -11090
rect 16005 -11210 16125 -11090
rect 16170 -11210 16290 -11090
rect 16345 -11210 16465 -11090
rect 16510 -11210 16630 -11090
rect 16675 -11210 16795 -11090
rect 16840 -11210 16960 -11090
rect 17015 -11210 17135 -11090
rect 17180 -11210 17300 -11090
rect 17345 -11210 17465 -11090
rect 17510 -11210 17630 -11090
rect 17685 -11210 17805 -11090
rect 17850 -11210 17970 -11090
rect 18015 -11210 18135 -11090
rect 18180 -11210 18300 -11090
rect 12820 -11375 12940 -11255
rect 12995 -11375 13115 -11255
rect 13160 -11375 13280 -11255
rect 13325 -11375 13445 -11255
rect 13490 -11375 13610 -11255
rect 13665 -11375 13785 -11255
rect 13830 -11375 13950 -11255
rect 13995 -11375 14115 -11255
rect 14160 -11375 14280 -11255
rect 14335 -11375 14455 -11255
rect 14500 -11375 14620 -11255
rect 14665 -11375 14785 -11255
rect 14830 -11375 14950 -11255
rect 15005 -11375 15125 -11255
rect 15170 -11375 15290 -11255
rect 15335 -11375 15455 -11255
rect 15500 -11375 15620 -11255
rect 15675 -11375 15795 -11255
rect 15840 -11375 15960 -11255
rect 16005 -11375 16125 -11255
rect 16170 -11375 16290 -11255
rect 16345 -11375 16465 -11255
rect 16510 -11375 16630 -11255
rect 16675 -11375 16795 -11255
rect 16840 -11375 16960 -11255
rect 17015 -11375 17135 -11255
rect 17180 -11375 17300 -11255
rect 17345 -11375 17465 -11255
rect 17510 -11375 17630 -11255
rect 17685 -11375 17805 -11255
rect 17850 -11375 17970 -11255
rect 18015 -11375 18135 -11255
rect 18180 -11375 18300 -11255
rect 12820 -11550 12940 -11430
rect 12995 -11550 13115 -11430
rect 13160 -11550 13280 -11430
rect 13325 -11550 13445 -11430
rect 13490 -11550 13610 -11430
rect 13665 -11550 13785 -11430
rect 13830 -11550 13950 -11430
rect 13995 -11550 14115 -11430
rect 14160 -11550 14280 -11430
rect 14335 -11550 14455 -11430
rect 14500 -11550 14620 -11430
rect 14665 -11550 14785 -11430
rect 14830 -11550 14950 -11430
rect 15005 -11550 15125 -11430
rect 15170 -11550 15290 -11430
rect 15335 -11550 15455 -11430
rect 15500 -11550 15620 -11430
rect 15675 -11550 15795 -11430
rect 15840 -11550 15960 -11430
rect 16005 -11550 16125 -11430
rect 16170 -11550 16290 -11430
rect 16345 -11550 16465 -11430
rect 16510 -11550 16630 -11430
rect 16675 -11550 16795 -11430
rect 16840 -11550 16960 -11430
rect 17015 -11550 17135 -11430
rect 17180 -11550 17300 -11430
rect 17345 -11550 17465 -11430
rect 17510 -11550 17630 -11430
rect 17685 -11550 17805 -11430
rect 17850 -11550 17970 -11430
rect 18015 -11550 18135 -11430
rect 18180 -11550 18300 -11430
rect 12820 -11715 12940 -11595
rect 12995 -11715 13115 -11595
rect 13160 -11715 13280 -11595
rect 13325 -11715 13445 -11595
rect 13490 -11715 13610 -11595
rect 13665 -11715 13785 -11595
rect 13830 -11715 13950 -11595
rect 13995 -11715 14115 -11595
rect 14160 -11715 14280 -11595
rect 14335 -11715 14455 -11595
rect 14500 -11715 14620 -11595
rect 14665 -11715 14785 -11595
rect 14830 -11715 14950 -11595
rect 15005 -11715 15125 -11595
rect 15170 -11715 15290 -11595
rect 15335 -11715 15455 -11595
rect 15500 -11715 15620 -11595
rect 15675 -11715 15795 -11595
rect 15840 -11715 15960 -11595
rect 16005 -11715 16125 -11595
rect 16170 -11715 16290 -11595
rect 16345 -11715 16465 -11595
rect 16510 -11715 16630 -11595
rect 16675 -11715 16795 -11595
rect 16840 -11715 16960 -11595
rect 17015 -11715 17135 -11595
rect 17180 -11715 17300 -11595
rect 17345 -11715 17465 -11595
rect 17510 -11715 17630 -11595
rect 17685 -11715 17805 -11595
rect 17850 -11715 17970 -11595
rect 18015 -11715 18135 -11595
rect 18180 -11715 18300 -11595
rect 12820 -11880 12940 -11760
rect 12995 -11880 13115 -11760
rect 13160 -11880 13280 -11760
rect 13325 -11880 13445 -11760
rect 13490 -11880 13610 -11760
rect 13665 -11880 13785 -11760
rect 13830 -11880 13950 -11760
rect 13995 -11880 14115 -11760
rect 14160 -11880 14280 -11760
rect 14335 -11880 14455 -11760
rect 14500 -11880 14620 -11760
rect 14665 -11880 14785 -11760
rect 14830 -11880 14950 -11760
rect 15005 -11880 15125 -11760
rect 15170 -11880 15290 -11760
rect 15335 -11880 15455 -11760
rect 15500 -11880 15620 -11760
rect 15675 -11880 15795 -11760
rect 15840 -11880 15960 -11760
rect 16005 -11880 16125 -11760
rect 16170 -11880 16290 -11760
rect 16345 -11880 16465 -11760
rect 16510 -11880 16630 -11760
rect 16675 -11880 16795 -11760
rect 16840 -11880 16960 -11760
rect 17015 -11880 17135 -11760
rect 17180 -11880 17300 -11760
rect 17345 -11880 17465 -11760
rect 17510 -11880 17630 -11760
rect 17685 -11880 17805 -11760
rect 17850 -11880 17970 -11760
rect 18015 -11880 18135 -11760
rect 18180 -11880 18300 -11760
rect 12820 -12045 12940 -11925
rect 12995 -12045 13115 -11925
rect 13160 -12045 13280 -11925
rect 13325 -12045 13445 -11925
rect 13490 -12045 13610 -11925
rect 13665 -12045 13785 -11925
rect 13830 -12045 13950 -11925
rect 13995 -12045 14115 -11925
rect 14160 -12045 14280 -11925
rect 14335 -12045 14455 -11925
rect 14500 -12045 14620 -11925
rect 14665 -12045 14785 -11925
rect 14830 -12045 14950 -11925
rect 15005 -12045 15125 -11925
rect 15170 -12045 15290 -11925
rect 15335 -12045 15455 -11925
rect 15500 -12045 15620 -11925
rect 15675 -12045 15795 -11925
rect 15840 -12045 15960 -11925
rect 16005 -12045 16125 -11925
rect 16170 -12045 16290 -11925
rect 16345 -12045 16465 -11925
rect 16510 -12045 16630 -11925
rect 16675 -12045 16795 -11925
rect 16840 -12045 16960 -11925
rect 17015 -12045 17135 -11925
rect 17180 -12045 17300 -11925
rect 17345 -12045 17465 -11925
rect 17510 -12045 17630 -11925
rect 17685 -12045 17805 -11925
rect 17850 -12045 17970 -11925
rect 18015 -12045 18135 -11925
rect 18180 -12045 18300 -11925
rect 12820 -12220 12940 -12100
rect 12995 -12220 13115 -12100
rect 13160 -12220 13280 -12100
rect 13325 -12220 13445 -12100
rect 13490 -12220 13610 -12100
rect 13665 -12220 13785 -12100
rect 13830 -12220 13950 -12100
rect 13995 -12220 14115 -12100
rect 14160 -12220 14280 -12100
rect 14335 -12220 14455 -12100
rect 14500 -12220 14620 -12100
rect 14665 -12220 14785 -12100
rect 14830 -12220 14950 -12100
rect 15005 -12220 15125 -12100
rect 15170 -12220 15290 -12100
rect 15335 -12220 15455 -12100
rect 15500 -12220 15620 -12100
rect 15675 -12220 15795 -12100
rect 15840 -12220 15960 -12100
rect 16005 -12220 16125 -12100
rect 16170 -12220 16290 -12100
rect 16345 -12220 16465 -12100
rect 16510 -12220 16630 -12100
rect 16675 -12220 16795 -12100
rect 16840 -12220 16960 -12100
rect 17015 -12220 17135 -12100
rect 17180 -12220 17300 -12100
rect 17345 -12220 17465 -12100
rect 17510 -12220 17630 -12100
rect 17685 -12220 17805 -12100
rect 17850 -12220 17970 -12100
rect 18015 -12220 18135 -12100
rect 18180 -12220 18300 -12100
rect 12820 -12385 12940 -12265
rect 12995 -12385 13115 -12265
rect 13160 -12385 13280 -12265
rect 13325 -12385 13445 -12265
rect 13490 -12385 13610 -12265
rect 13665 -12385 13785 -12265
rect 13830 -12385 13950 -12265
rect 13995 -12385 14115 -12265
rect 14160 -12385 14280 -12265
rect 14335 -12385 14455 -12265
rect 14500 -12385 14620 -12265
rect 14665 -12385 14785 -12265
rect 14830 -12385 14950 -12265
rect 15005 -12385 15125 -12265
rect 15170 -12385 15290 -12265
rect 15335 -12385 15455 -12265
rect 15500 -12385 15620 -12265
rect 15675 -12385 15795 -12265
rect 15840 -12385 15960 -12265
rect 16005 -12385 16125 -12265
rect 16170 -12385 16290 -12265
rect 16345 -12385 16465 -12265
rect 16510 -12385 16630 -12265
rect 16675 -12385 16795 -12265
rect 16840 -12385 16960 -12265
rect 17015 -12385 17135 -12265
rect 17180 -12385 17300 -12265
rect 17345 -12385 17465 -12265
rect 17510 -12385 17630 -12265
rect 17685 -12385 17805 -12265
rect 17850 -12385 17970 -12265
rect 18015 -12385 18135 -12265
rect 18180 -12385 18300 -12265
rect 12820 -12550 12940 -12430
rect 12995 -12550 13115 -12430
rect 13160 -12550 13280 -12430
rect 13325 -12550 13445 -12430
rect 13490 -12550 13610 -12430
rect 13665 -12550 13785 -12430
rect 13830 -12550 13950 -12430
rect 13995 -12550 14115 -12430
rect 14160 -12550 14280 -12430
rect 14335 -12550 14455 -12430
rect 14500 -12550 14620 -12430
rect 14665 -12550 14785 -12430
rect 14830 -12550 14950 -12430
rect 15005 -12550 15125 -12430
rect 15170 -12550 15290 -12430
rect 15335 -12550 15455 -12430
rect 15500 -12550 15620 -12430
rect 15675 -12550 15795 -12430
rect 15840 -12550 15960 -12430
rect 16005 -12550 16125 -12430
rect 16170 -12550 16290 -12430
rect 16345 -12550 16465 -12430
rect 16510 -12550 16630 -12430
rect 16675 -12550 16795 -12430
rect 16840 -12550 16960 -12430
rect 17015 -12550 17135 -12430
rect 17180 -12550 17300 -12430
rect 17345 -12550 17465 -12430
rect 17510 -12550 17630 -12430
rect 17685 -12550 17805 -12430
rect 17850 -12550 17970 -12430
rect 18015 -12550 18135 -12430
rect 18180 -12550 18300 -12430
rect 12820 -12715 12940 -12595
rect 12995 -12715 13115 -12595
rect 13160 -12715 13280 -12595
rect 13325 -12715 13445 -12595
rect 13490 -12715 13610 -12595
rect 13665 -12715 13785 -12595
rect 13830 -12715 13950 -12595
rect 13995 -12715 14115 -12595
rect 14160 -12715 14280 -12595
rect 14335 -12715 14455 -12595
rect 14500 -12715 14620 -12595
rect 14665 -12715 14785 -12595
rect 14830 -12715 14950 -12595
rect 15005 -12715 15125 -12595
rect 15170 -12715 15290 -12595
rect 15335 -12715 15455 -12595
rect 15500 -12715 15620 -12595
rect 15675 -12715 15795 -12595
rect 15840 -12715 15960 -12595
rect 16005 -12715 16125 -12595
rect 16170 -12715 16290 -12595
rect 16345 -12715 16465 -12595
rect 16510 -12715 16630 -12595
rect 16675 -12715 16795 -12595
rect 16840 -12715 16960 -12595
rect 17015 -12715 17135 -12595
rect 17180 -12715 17300 -12595
rect 17345 -12715 17465 -12595
rect 17510 -12715 17630 -12595
rect 17685 -12715 17805 -12595
rect 17850 -12715 17970 -12595
rect 18015 -12715 18135 -12595
rect 18180 -12715 18300 -12595
rect 12820 -12890 12940 -12770
rect 12995 -12890 13115 -12770
rect 13160 -12890 13280 -12770
rect 13325 -12890 13445 -12770
rect 13490 -12890 13610 -12770
rect 13665 -12890 13785 -12770
rect 13830 -12890 13950 -12770
rect 13995 -12890 14115 -12770
rect 14160 -12890 14280 -12770
rect 14335 -12890 14455 -12770
rect 14500 -12890 14620 -12770
rect 14665 -12890 14785 -12770
rect 14830 -12890 14950 -12770
rect 15005 -12890 15125 -12770
rect 15170 -12890 15290 -12770
rect 15335 -12890 15455 -12770
rect 15500 -12890 15620 -12770
rect 15675 -12890 15795 -12770
rect 15840 -12890 15960 -12770
rect 16005 -12890 16125 -12770
rect 16170 -12890 16290 -12770
rect 16345 -12890 16465 -12770
rect 16510 -12890 16630 -12770
rect 16675 -12890 16795 -12770
rect 16840 -12890 16960 -12770
rect 17015 -12890 17135 -12770
rect 17180 -12890 17300 -12770
rect 17345 -12890 17465 -12770
rect 17510 -12890 17630 -12770
rect 17685 -12890 17805 -12770
rect 17850 -12890 17970 -12770
rect 18015 -12890 18135 -12770
rect 18180 -12890 18300 -12770
rect 12820 -13055 12940 -12935
rect 12995 -13055 13115 -12935
rect 13160 -13055 13280 -12935
rect 13325 -13055 13445 -12935
rect 13490 -13055 13610 -12935
rect 13665 -13055 13785 -12935
rect 13830 -13055 13950 -12935
rect 13995 -13055 14115 -12935
rect 14160 -13055 14280 -12935
rect 14335 -13055 14455 -12935
rect 14500 -13055 14620 -12935
rect 14665 -13055 14785 -12935
rect 14830 -13055 14950 -12935
rect 15005 -13055 15125 -12935
rect 15170 -13055 15290 -12935
rect 15335 -13055 15455 -12935
rect 15500 -13055 15620 -12935
rect 15675 -13055 15795 -12935
rect 15840 -13055 15960 -12935
rect 16005 -13055 16125 -12935
rect 16170 -13055 16290 -12935
rect 16345 -13055 16465 -12935
rect 16510 -13055 16630 -12935
rect 16675 -13055 16795 -12935
rect 16840 -13055 16960 -12935
rect 17015 -13055 17135 -12935
rect 17180 -13055 17300 -12935
rect 17345 -13055 17465 -12935
rect 17510 -13055 17630 -12935
rect 17685 -13055 17805 -12935
rect 17850 -13055 17970 -12935
rect 18015 -13055 18135 -12935
rect 18180 -13055 18300 -12935
rect 12820 -13220 12940 -13100
rect 12995 -13220 13115 -13100
rect 13160 -13220 13280 -13100
rect 13325 -13220 13445 -13100
rect 13490 -13220 13610 -13100
rect 13665 -13220 13785 -13100
rect 13830 -13220 13950 -13100
rect 13995 -13220 14115 -13100
rect 14160 -13220 14280 -13100
rect 14335 -13220 14455 -13100
rect 14500 -13220 14620 -13100
rect 14665 -13220 14785 -13100
rect 14830 -13220 14950 -13100
rect 15005 -13220 15125 -13100
rect 15170 -13220 15290 -13100
rect 15335 -13220 15455 -13100
rect 15500 -13220 15620 -13100
rect 15675 -13220 15795 -13100
rect 15840 -13220 15960 -13100
rect 16005 -13220 16125 -13100
rect 16170 -13220 16290 -13100
rect 16345 -13220 16465 -13100
rect 16510 -13220 16630 -13100
rect 16675 -13220 16795 -13100
rect 16840 -13220 16960 -13100
rect 17015 -13220 17135 -13100
rect 17180 -13220 17300 -13100
rect 17345 -13220 17465 -13100
rect 17510 -13220 17630 -13100
rect 17685 -13220 17805 -13100
rect 17850 -13220 17970 -13100
rect 18015 -13220 18135 -13100
rect 18180 -13220 18300 -13100
rect 12820 -13385 12940 -13265
rect 12995 -13385 13115 -13265
rect 13160 -13385 13280 -13265
rect 13325 -13385 13445 -13265
rect 13490 -13385 13610 -13265
rect 13665 -13385 13785 -13265
rect 13830 -13385 13950 -13265
rect 13995 -13385 14115 -13265
rect 14160 -13385 14280 -13265
rect 14335 -13385 14455 -13265
rect 14500 -13385 14620 -13265
rect 14665 -13385 14785 -13265
rect 14830 -13385 14950 -13265
rect 15005 -13385 15125 -13265
rect 15170 -13385 15290 -13265
rect 15335 -13385 15455 -13265
rect 15500 -13385 15620 -13265
rect 15675 -13385 15795 -13265
rect 15840 -13385 15960 -13265
rect 16005 -13385 16125 -13265
rect 16170 -13385 16290 -13265
rect 16345 -13385 16465 -13265
rect 16510 -13385 16630 -13265
rect 16675 -13385 16795 -13265
rect 16840 -13385 16960 -13265
rect 17015 -13385 17135 -13265
rect 17180 -13385 17300 -13265
rect 17345 -13385 17465 -13265
rect 17510 -13385 17630 -13265
rect 17685 -13385 17805 -13265
rect 17850 -13385 17970 -13265
rect 18015 -13385 18135 -13265
rect 18180 -13385 18300 -13265
rect 12820 -13560 12940 -13440
rect 12995 -13560 13115 -13440
rect 13160 -13560 13280 -13440
rect 13325 -13560 13445 -13440
rect 13490 -13560 13610 -13440
rect 13665 -13560 13785 -13440
rect 13830 -13560 13950 -13440
rect 13995 -13560 14115 -13440
rect 14160 -13560 14280 -13440
rect 14335 -13560 14455 -13440
rect 14500 -13560 14620 -13440
rect 14665 -13560 14785 -13440
rect 14830 -13560 14950 -13440
rect 15005 -13560 15125 -13440
rect 15170 -13560 15290 -13440
rect 15335 -13560 15455 -13440
rect 15500 -13560 15620 -13440
rect 15675 -13560 15795 -13440
rect 15840 -13560 15960 -13440
rect 16005 -13560 16125 -13440
rect 16170 -13560 16290 -13440
rect 16345 -13560 16465 -13440
rect 16510 -13560 16630 -13440
rect 16675 -13560 16795 -13440
rect 16840 -13560 16960 -13440
rect 17015 -13560 17135 -13440
rect 17180 -13560 17300 -13440
rect 17345 -13560 17465 -13440
rect 17510 -13560 17630 -13440
rect 17685 -13560 17805 -13440
rect 17850 -13560 17970 -13440
rect 18015 -13560 18135 -13440
rect 18180 -13560 18300 -13440
rect 12820 -13725 12940 -13605
rect 12995 -13725 13115 -13605
rect 13160 -13725 13280 -13605
rect 13325 -13725 13445 -13605
rect 13490 -13725 13610 -13605
rect 13665 -13725 13785 -13605
rect 13830 -13725 13950 -13605
rect 13995 -13725 14115 -13605
rect 14160 -13725 14280 -13605
rect 14335 -13725 14455 -13605
rect 14500 -13725 14620 -13605
rect 14665 -13725 14785 -13605
rect 14830 -13725 14950 -13605
rect 15005 -13725 15125 -13605
rect 15170 -13725 15290 -13605
rect 15335 -13725 15455 -13605
rect 15500 -13725 15620 -13605
rect 15675 -13725 15795 -13605
rect 15840 -13725 15960 -13605
rect 16005 -13725 16125 -13605
rect 16170 -13725 16290 -13605
rect 16345 -13725 16465 -13605
rect 16510 -13725 16630 -13605
rect 16675 -13725 16795 -13605
rect 16840 -13725 16960 -13605
rect 17015 -13725 17135 -13605
rect 17180 -13725 17300 -13605
rect 17345 -13725 17465 -13605
rect 17510 -13725 17630 -13605
rect 17685 -13725 17805 -13605
rect 17850 -13725 17970 -13605
rect 18015 -13725 18135 -13605
rect 18180 -13725 18300 -13605
rect 12820 -13890 12940 -13770
rect 12995 -13890 13115 -13770
rect 13160 -13890 13280 -13770
rect 13325 -13890 13445 -13770
rect 13490 -13890 13610 -13770
rect 13665 -13890 13785 -13770
rect 13830 -13890 13950 -13770
rect 13995 -13890 14115 -13770
rect 14160 -13890 14280 -13770
rect 14335 -13890 14455 -13770
rect 14500 -13890 14620 -13770
rect 14665 -13890 14785 -13770
rect 14830 -13890 14950 -13770
rect 15005 -13890 15125 -13770
rect 15170 -13890 15290 -13770
rect 15335 -13890 15455 -13770
rect 15500 -13890 15620 -13770
rect 15675 -13890 15795 -13770
rect 15840 -13890 15960 -13770
rect 16005 -13890 16125 -13770
rect 16170 -13890 16290 -13770
rect 16345 -13890 16465 -13770
rect 16510 -13890 16630 -13770
rect 16675 -13890 16795 -13770
rect 16840 -13890 16960 -13770
rect 17015 -13890 17135 -13770
rect 17180 -13890 17300 -13770
rect 17345 -13890 17465 -13770
rect 17510 -13890 17630 -13770
rect 17685 -13890 17805 -13770
rect 17850 -13890 17970 -13770
rect 18015 -13890 18135 -13770
rect 18180 -13890 18300 -13770
rect 12820 -14055 12940 -13935
rect 12995 -14055 13115 -13935
rect 13160 -14055 13280 -13935
rect 13325 -14055 13445 -13935
rect 13490 -14055 13610 -13935
rect 13665 -14055 13785 -13935
rect 13830 -14055 13950 -13935
rect 13995 -14055 14115 -13935
rect 14160 -14055 14280 -13935
rect 14335 -14055 14455 -13935
rect 14500 -14055 14620 -13935
rect 14665 -14055 14785 -13935
rect 14830 -14055 14950 -13935
rect 15005 -14055 15125 -13935
rect 15170 -14055 15290 -13935
rect 15335 -14055 15455 -13935
rect 15500 -14055 15620 -13935
rect 15675 -14055 15795 -13935
rect 15840 -14055 15960 -13935
rect 16005 -14055 16125 -13935
rect 16170 -14055 16290 -13935
rect 16345 -14055 16465 -13935
rect 16510 -14055 16630 -13935
rect 16675 -14055 16795 -13935
rect 16840 -14055 16960 -13935
rect 17015 -14055 17135 -13935
rect 17180 -14055 17300 -13935
rect 17345 -14055 17465 -13935
rect 17510 -14055 17630 -13935
rect 17685 -14055 17805 -13935
rect 17850 -14055 17970 -13935
rect 18015 -14055 18135 -13935
rect 18180 -14055 18300 -13935
rect 12820 -14230 12940 -14110
rect 12995 -14230 13115 -14110
rect 13160 -14230 13280 -14110
rect 13325 -14230 13445 -14110
rect 13490 -14230 13610 -14110
rect 13665 -14230 13785 -14110
rect 13830 -14230 13950 -14110
rect 13995 -14230 14115 -14110
rect 14160 -14230 14280 -14110
rect 14335 -14230 14455 -14110
rect 14500 -14230 14620 -14110
rect 14665 -14230 14785 -14110
rect 14830 -14230 14950 -14110
rect 15005 -14230 15125 -14110
rect 15170 -14230 15290 -14110
rect 15335 -14230 15455 -14110
rect 15500 -14230 15620 -14110
rect 15675 -14230 15795 -14110
rect 15840 -14230 15960 -14110
rect 16005 -14230 16125 -14110
rect 16170 -14230 16290 -14110
rect 16345 -14230 16465 -14110
rect 16510 -14230 16630 -14110
rect 16675 -14230 16795 -14110
rect 16840 -14230 16960 -14110
rect 17015 -14230 17135 -14110
rect 17180 -14230 17300 -14110
rect 17345 -14230 17465 -14110
rect 17510 -14230 17630 -14110
rect 17685 -14230 17805 -14110
rect 17850 -14230 17970 -14110
rect 18015 -14230 18135 -14110
rect 18180 -14230 18300 -14110
rect 12820 -14395 12940 -14275
rect 12995 -14395 13115 -14275
rect 13160 -14395 13280 -14275
rect 13325 -14395 13445 -14275
rect 13490 -14395 13610 -14275
rect 13665 -14395 13785 -14275
rect 13830 -14395 13950 -14275
rect 13995 -14395 14115 -14275
rect 14160 -14395 14280 -14275
rect 14335 -14395 14455 -14275
rect 14500 -14395 14620 -14275
rect 14665 -14395 14785 -14275
rect 14830 -14395 14950 -14275
rect 15005 -14395 15125 -14275
rect 15170 -14395 15290 -14275
rect 15335 -14395 15455 -14275
rect 15500 -14395 15620 -14275
rect 15675 -14395 15795 -14275
rect 15840 -14395 15960 -14275
rect 16005 -14395 16125 -14275
rect 16170 -14395 16290 -14275
rect 16345 -14395 16465 -14275
rect 16510 -14395 16630 -14275
rect 16675 -14395 16795 -14275
rect 16840 -14395 16960 -14275
rect 17015 -14395 17135 -14275
rect 17180 -14395 17300 -14275
rect 17345 -14395 17465 -14275
rect 17510 -14395 17630 -14275
rect 17685 -14395 17805 -14275
rect 17850 -14395 17970 -14275
rect 18015 -14395 18135 -14275
rect 18180 -14395 18300 -14275
rect 12820 -14560 12940 -14440
rect 12995 -14560 13115 -14440
rect 13160 -14560 13280 -14440
rect 13325 -14560 13445 -14440
rect 13490 -14560 13610 -14440
rect 13665 -14560 13785 -14440
rect 13830 -14560 13950 -14440
rect 13995 -14560 14115 -14440
rect 14160 -14560 14280 -14440
rect 14335 -14560 14455 -14440
rect 14500 -14560 14620 -14440
rect 14665 -14560 14785 -14440
rect 14830 -14560 14950 -14440
rect 15005 -14560 15125 -14440
rect 15170 -14560 15290 -14440
rect 15335 -14560 15455 -14440
rect 15500 -14560 15620 -14440
rect 15675 -14560 15795 -14440
rect 15840 -14560 15960 -14440
rect 16005 -14560 16125 -14440
rect 16170 -14560 16290 -14440
rect 16345 -14560 16465 -14440
rect 16510 -14560 16630 -14440
rect 16675 -14560 16795 -14440
rect 16840 -14560 16960 -14440
rect 17015 -14560 17135 -14440
rect 17180 -14560 17300 -14440
rect 17345 -14560 17465 -14440
rect 17510 -14560 17630 -14440
rect 17685 -14560 17805 -14440
rect 17850 -14560 17970 -14440
rect 18015 -14560 18135 -14440
rect 18180 -14560 18300 -14440
rect 12820 -14725 12940 -14605
rect 12995 -14725 13115 -14605
rect 13160 -14725 13280 -14605
rect 13325 -14725 13445 -14605
rect 13490 -14725 13610 -14605
rect 13665 -14725 13785 -14605
rect 13830 -14725 13950 -14605
rect 13995 -14725 14115 -14605
rect 14160 -14725 14280 -14605
rect 14335 -14725 14455 -14605
rect 14500 -14725 14620 -14605
rect 14665 -14725 14785 -14605
rect 14830 -14725 14950 -14605
rect 15005 -14725 15125 -14605
rect 15170 -14725 15290 -14605
rect 15335 -14725 15455 -14605
rect 15500 -14725 15620 -14605
rect 15675 -14725 15795 -14605
rect 15840 -14725 15960 -14605
rect 16005 -14725 16125 -14605
rect 16170 -14725 16290 -14605
rect 16345 -14725 16465 -14605
rect 16510 -14725 16630 -14605
rect 16675 -14725 16795 -14605
rect 16840 -14725 16960 -14605
rect 17015 -14725 17135 -14605
rect 17180 -14725 17300 -14605
rect 17345 -14725 17465 -14605
rect 17510 -14725 17630 -14605
rect 17685 -14725 17805 -14605
rect 17850 -14725 17970 -14605
rect 18015 -14725 18135 -14605
rect 18180 -14725 18300 -14605
rect 12820 -14900 12940 -14780
rect 12995 -14900 13115 -14780
rect 13160 -14900 13280 -14780
rect 13325 -14900 13445 -14780
rect 13490 -14900 13610 -14780
rect 13665 -14900 13785 -14780
rect 13830 -14900 13950 -14780
rect 13995 -14900 14115 -14780
rect 14160 -14900 14280 -14780
rect 14335 -14900 14455 -14780
rect 14500 -14900 14620 -14780
rect 14665 -14900 14785 -14780
rect 14830 -14900 14950 -14780
rect 15005 -14900 15125 -14780
rect 15170 -14900 15290 -14780
rect 15335 -14900 15455 -14780
rect 15500 -14900 15620 -14780
rect 15675 -14900 15795 -14780
rect 15840 -14900 15960 -14780
rect 16005 -14900 16125 -14780
rect 16170 -14900 16290 -14780
rect 16345 -14900 16465 -14780
rect 16510 -14900 16630 -14780
rect 16675 -14900 16795 -14780
rect 16840 -14900 16960 -14780
rect 17015 -14900 17135 -14780
rect 17180 -14900 17300 -14780
rect 17345 -14900 17465 -14780
rect 17510 -14900 17630 -14780
rect 17685 -14900 17805 -14780
rect 17850 -14900 17970 -14780
rect 18015 -14900 18135 -14780
rect 18180 -14900 18300 -14780
rect 12820 -15065 12940 -14945
rect 12995 -15065 13115 -14945
rect 13160 -15065 13280 -14945
rect 13325 -15065 13445 -14945
rect 13490 -15065 13610 -14945
rect 13665 -15065 13785 -14945
rect 13830 -15065 13950 -14945
rect 13995 -15065 14115 -14945
rect 14160 -15065 14280 -14945
rect 14335 -15065 14455 -14945
rect 14500 -15065 14620 -14945
rect 14665 -15065 14785 -14945
rect 14830 -15065 14950 -14945
rect 15005 -15065 15125 -14945
rect 15170 -15065 15290 -14945
rect 15335 -15065 15455 -14945
rect 15500 -15065 15620 -14945
rect 15675 -15065 15795 -14945
rect 15840 -15065 15960 -14945
rect 16005 -15065 16125 -14945
rect 16170 -15065 16290 -14945
rect 16345 -15065 16465 -14945
rect 16510 -15065 16630 -14945
rect 16675 -15065 16795 -14945
rect 16840 -15065 16960 -14945
rect 17015 -15065 17135 -14945
rect 17180 -15065 17300 -14945
rect 17345 -15065 17465 -14945
rect 17510 -15065 17630 -14945
rect 17685 -15065 17805 -14945
rect 17850 -15065 17970 -14945
rect 18015 -15065 18135 -14945
rect 18180 -15065 18300 -14945
rect 12820 -15230 12940 -15110
rect 12995 -15230 13115 -15110
rect 13160 -15230 13280 -15110
rect 13325 -15230 13445 -15110
rect 13490 -15230 13610 -15110
rect 13665 -15230 13785 -15110
rect 13830 -15230 13950 -15110
rect 13995 -15230 14115 -15110
rect 14160 -15230 14280 -15110
rect 14335 -15230 14455 -15110
rect 14500 -15230 14620 -15110
rect 14665 -15230 14785 -15110
rect 14830 -15230 14950 -15110
rect 15005 -15230 15125 -15110
rect 15170 -15230 15290 -15110
rect 15335 -15230 15455 -15110
rect 15500 -15230 15620 -15110
rect 15675 -15230 15795 -15110
rect 15840 -15230 15960 -15110
rect 16005 -15230 16125 -15110
rect 16170 -15230 16290 -15110
rect 16345 -15230 16465 -15110
rect 16510 -15230 16630 -15110
rect 16675 -15230 16795 -15110
rect 16840 -15230 16960 -15110
rect 17015 -15230 17135 -15110
rect 17180 -15230 17300 -15110
rect 17345 -15230 17465 -15110
rect 17510 -15230 17630 -15110
rect 17685 -15230 17805 -15110
rect 17850 -15230 17970 -15110
rect 18015 -15230 18135 -15110
rect 18180 -15230 18300 -15110
rect 12820 -15395 12940 -15275
rect 12995 -15395 13115 -15275
rect 13160 -15395 13280 -15275
rect 13325 -15395 13445 -15275
rect 13490 -15395 13610 -15275
rect 13665 -15395 13785 -15275
rect 13830 -15395 13950 -15275
rect 13995 -15395 14115 -15275
rect 14160 -15395 14280 -15275
rect 14335 -15395 14455 -15275
rect 14500 -15395 14620 -15275
rect 14665 -15395 14785 -15275
rect 14830 -15395 14950 -15275
rect 15005 -15395 15125 -15275
rect 15170 -15395 15290 -15275
rect 15335 -15395 15455 -15275
rect 15500 -15395 15620 -15275
rect 15675 -15395 15795 -15275
rect 15840 -15395 15960 -15275
rect 16005 -15395 16125 -15275
rect 16170 -15395 16290 -15275
rect 16345 -15395 16465 -15275
rect 16510 -15395 16630 -15275
rect 16675 -15395 16795 -15275
rect 16840 -15395 16960 -15275
rect 17015 -15395 17135 -15275
rect 17180 -15395 17300 -15275
rect 17345 -15395 17465 -15275
rect 17510 -15395 17630 -15275
rect 17685 -15395 17805 -15275
rect 17850 -15395 17970 -15275
rect 18015 -15395 18135 -15275
rect 18180 -15395 18300 -15275
rect 12820 -15570 12940 -15450
rect 12995 -15570 13115 -15450
rect 13160 -15570 13280 -15450
rect 13325 -15570 13445 -15450
rect 13490 -15570 13610 -15450
rect 13665 -15570 13785 -15450
rect 13830 -15570 13950 -15450
rect 13995 -15570 14115 -15450
rect 14160 -15570 14280 -15450
rect 14335 -15570 14455 -15450
rect 14500 -15570 14620 -15450
rect 14665 -15570 14785 -15450
rect 14830 -15570 14950 -15450
rect 15005 -15570 15125 -15450
rect 15170 -15570 15290 -15450
rect 15335 -15570 15455 -15450
rect 15500 -15570 15620 -15450
rect 15675 -15570 15795 -15450
rect 15840 -15570 15960 -15450
rect 16005 -15570 16125 -15450
rect 16170 -15570 16290 -15450
rect 16345 -15570 16465 -15450
rect 16510 -15570 16630 -15450
rect 16675 -15570 16795 -15450
rect 16840 -15570 16960 -15450
rect 17015 -15570 17135 -15450
rect 17180 -15570 17300 -15450
rect 17345 -15570 17465 -15450
rect 17510 -15570 17630 -15450
rect 17685 -15570 17805 -15450
rect 17850 -15570 17970 -15450
rect 18015 -15570 18135 -15450
rect 18180 -15570 18300 -15450
rect 18510 -10210 18630 -10090
rect 18685 -10210 18805 -10090
rect 18850 -10210 18970 -10090
rect 19015 -10210 19135 -10090
rect 19180 -10210 19300 -10090
rect 19355 -10210 19475 -10090
rect 19520 -10210 19640 -10090
rect 19685 -10210 19805 -10090
rect 19850 -10210 19970 -10090
rect 20025 -10210 20145 -10090
rect 20190 -10210 20310 -10090
rect 20355 -10210 20475 -10090
rect 20520 -10210 20640 -10090
rect 20695 -10210 20815 -10090
rect 20860 -10210 20980 -10090
rect 21025 -10210 21145 -10090
rect 21190 -10210 21310 -10090
rect 21365 -10210 21485 -10090
rect 21530 -10210 21650 -10090
rect 21695 -10210 21815 -10090
rect 21860 -10210 21980 -10090
rect 22035 -10210 22155 -10090
rect 22200 -10210 22320 -10090
rect 22365 -10210 22485 -10090
rect 22530 -10210 22650 -10090
rect 22705 -10210 22825 -10090
rect 22870 -10210 22990 -10090
rect 23035 -10210 23155 -10090
rect 23200 -10210 23320 -10090
rect 23375 -10210 23495 -10090
rect 23540 -10210 23660 -10090
rect 23705 -10210 23825 -10090
rect 23870 -10210 23990 -10090
rect 18510 -10375 18630 -10255
rect 18685 -10375 18805 -10255
rect 18850 -10375 18970 -10255
rect 19015 -10375 19135 -10255
rect 19180 -10375 19300 -10255
rect 19355 -10375 19475 -10255
rect 19520 -10375 19640 -10255
rect 19685 -10375 19805 -10255
rect 19850 -10375 19970 -10255
rect 20025 -10375 20145 -10255
rect 20190 -10375 20310 -10255
rect 20355 -10375 20475 -10255
rect 20520 -10375 20640 -10255
rect 20695 -10375 20815 -10255
rect 20860 -10375 20980 -10255
rect 21025 -10375 21145 -10255
rect 21190 -10375 21310 -10255
rect 21365 -10375 21485 -10255
rect 21530 -10375 21650 -10255
rect 21695 -10375 21815 -10255
rect 21860 -10375 21980 -10255
rect 22035 -10375 22155 -10255
rect 22200 -10375 22320 -10255
rect 22365 -10375 22485 -10255
rect 22530 -10375 22650 -10255
rect 22705 -10375 22825 -10255
rect 22870 -10375 22990 -10255
rect 23035 -10375 23155 -10255
rect 23200 -10375 23320 -10255
rect 23375 -10375 23495 -10255
rect 23540 -10375 23660 -10255
rect 23705 -10375 23825 -10255
rect 23870 -10375 23990 -10255
rect 18510 -10540 18630 -10420
rect 18685 -10540 18805 -10420
rect 18850 -10540 18970 -10420
rect 19015 -10540 19135 -10420
rect 19180 -10540 19300 -10420
rect 19355 -10540 19475 -10420
rect 19520 -10540 19640 -10420
rect 19685 -10540 19805 -10420
rect 19850 -10540 19970 -10420
rect 20025 -10540 20145 -10420
rect 20190 -10540 20310 -10420
rect 20355 -10540 20475 -10420
rect 20520 -10540 20640 -10420
rect 20695 -10540 20815 -10420
rect 20860 -10540 20980 -10420
rect 21025 -10540 21145 -10420
rect 21190 -10540 21310 -10420
rect 21365 -10540 21485 -10420
rect 21530 -10540 21650 -10420
rect 21695 -10540 21815 -10420
rect 21860 -10540 21980 -10420
rect 22035 -10540 22155 -10420
rect 22200 -10540 22320 -10420
rect 22365 -10540 22485 -10420
rect 22530 -10540 22650 -10420
rect 22705 -10540 22825 -10420
rect 22870 -10540 22990 -10420
rect 23035 -10540 23155 -10420
rect 23200 -10540 23320 -10420
rect 23375 -10540 23495 -10420
rect 23540 -10540 23660 -10420
rect 23705 -10540 23825 -10420
rect 23870 -10540 23990 -10420
rect 18510 -10705 18630 -10585
rect 18685 -10705 18805 -10585
rect 18850 -10705 18970 -10585
rect 19015 -10705 19135 -10585
rect 19180 -10705 19300 -10585
rect 19355 -10705 19475 -10585
rect 19520 -10705 19640 -10585
rect 19685 -10705 19805 -10585
rect 19850 -10705 19970 -10585
rect 20025 -10705 20145 -10585
rect 20190 -10705 20310 -10585
rect 20355 -10705 20475 -10585
rect 20520 -10705 20640 -10585
rect 20695 -10705 20815 -10585
rect 20860 -10705 20980 -10585
rect 21025 -10705 21145 -10585
rect 21190 -10705 21310 -10585
rect 21365 -10705 21485 -10585
rect 21530 -10705 21650 -10585
rect 21695 -10705 21815 -10585
rect 21860 -10705 21980 -10585
rect 22035 -10705 22155 -10585
rect 22200 -10705 22320 -10585
rect 22365 -10705 22485 -10585
rect 22530 -10705 22650 -10585
rect 22705 -10705 22825 -10585
rect 22870 -10705 22990 -10585
rect 23035 -10705 23155 -10585
rect 23200 -10705 23320 -10585
rect 23375 -10705 23495 -10585
rect 23540 -10705 23660 -10585
rect 23705 -10705 23825 -10585
rect 23870 -10705 23990 -10585
rect 18510 -10880 18630 -10760
rect 18685 -10880 18805 -10760
rect 18850 -10880 18970 -10760
rect 19015 -10880 19135 -10760
rect 19180 -10880 19300 -10760
rect 19355 -10880 19475 -10760
rect 19520 -10880 19640 -10760
rect 19685 -10880 19805 -10760
rect 19850 -10880 19970 -10760
rect 20025 -10880 20145 -10760
rect 20190 -10880 20310 -10760
rect 20355 -10880 20475 -10760
rect 20520 -10880 20640 -10760
rect 20695 -10880 20815 -10760
rect 20860 -10880 20980 -10760
rect 21025 -10880 21145 -10760
rect 21190 -10880 21310 -10760
rect 21365 -10880 21485 -10760
rect 21530 -10880 21650 -10760
rect 21695 -10880 21815 -10760
rect 21860 -10880 21980 -10760
rect 22035 -10880 22155 -10760
rect 22200 -10880 22320 -10760
rect 22365 -10880 22485 -10760
rect 22530 -10880 22650 -10760
rect 22705 -10880 22825 -10760
rect 22870 -10880 22990 -10760
rect 23035 -10880 23155 -10760
rect 23200 -10880 23320 -10760
rect 23375 -10880 23495 -10760
rect 23540 -10880 23660 -10760
rect 23705 -10880 23825 -10760
rect 23870 -10880 23990 -10760
rect 18510 -11045 18630 -10925
rect 18685 -11045 18805 -10925
rect 18850 -11045 18970 -10925
rect 19015 -11045 19135 -10925
rect 19180 -11045 19300 -10925
rect 19355 -11045 19475 -10925
rect 19520 -11045 19640 -10925
rect 19685 -11045 19805 -10925
rect 19850 -11045 19970 -10925
rect 20025 -11045 20145 -10925
rect 20190 -11045 20310 -10925
rect 20355 -11045 20475 -10925
rect 20520 -11045 20640 -10925
rect 20695 -11045 20815 -10925
rect 20860 -11045 20980 -10925
rect 21025 -11045 21145 -10925
rect 21190 -11045 21310 -10925
rect 21365 -11045 21485 -10925
rect 21530 -11045 21650 -10925
rect 21695 -11045 21815 -10925
rect 21860 -11045 21980 -10925
rect 22035 -11045 22155 -10925
rect 22200 -11045 22320 -10925
rect 22365 -11045 22485 -10925
rect 22530 -11045 22650 -10925
rect 22705 -11045 22825 -10925
rect 22870 -11045 22990 -10925
rect 23035 -11045 23155 -10925
rect 23200 -11045 23320 -10925
rect 23375 -11045 23495 -10925
rect 23540 -11045 23660 -10925
rect 23705 -11045 23825 -10925
rect 23870 -11045 23990 -10925
rect 18510 -11210 18630 -11090
rect 18685 -11210 18805 -11090
rect 18850 -11210 18970 -11090
rect 19015 -11210 19135 -11090
rect 19180 -11210 19300 -11090
rect 19355 -11210 19475 -11090
rect 19520 -11210 19640 -11090
rect 19685 -11210 19805 -11090
rect 19850 -11210 19970 -11090
rect 20025 -11210 20145 -11090
rect 20190 -11210 20310 -11090
rect 20355 -11210 20475 -11090
rect 20520 -11210 20640 -11090
rect 20695 -11210 20815 -11090
rect 20860 -11210 20980 -11090
rect 21025 -11210 21145 -11090
rect 21190 -11210 21310 -11090
rect 21365 -11210 21485 -11090
rect 21530 -11210 21650 -11090
rect 21695 -11210 21815 -11090
rect 21860 -11210 21980 -11090
rect 22035 -11210 22155 -11090
rect 22200 -11210 22320 -11090
rect 22365 -11210 22485 -11090
rect 22530 -11210 22650 -11090
rect 22705 -11210 22825 -11090
rect 22870 -11210 22990 -11090
rect 23035 -11210 23155 -11090
rect 23200 -11210 23320 -11090
rect 23375 -11210 23495 -11090
rect 23540 -11210 23660 -11090
rect 23705 -11210 23825 -11090
rect 23870 -11210 23990 -11090
rect 18510 -11375 18630 -11255
rect 18685 -11375 18805 -11255
rect 18850 -11375 18970 -11255
rect 19015 -11375 19135 -11255
rect 19180 -11375 19300 -11255
rect 19355 -11375 19475 -11255
rect 19520 -11375 19640 -11255
rect 19685 -11375 19805 -11255
rect 19850 -11375 19970 -11255
rect 20025 -11375 20145 -11255
rect 20190 -11375 20310 -11255
rect 20355 -11375 20475 -11255
rect 20520 -11375 20640 -11255
rect 20695 -11375 20815 -11255
rect 20860 -11375 20980 -11255
rect 21025 -11375 21145 -11255
rect 21190 -11375 21310 -11255
rect 21365 -11375 21485 -11255
rect 21530 -11375 21650 -11255
rect 21695 -11375 21815 -11255
rect 21860 -11375 21980 -11255
rect 22035 -11375 22155 -11255
rect 22200 -11375 22320 -11255
rect 22365 -11375 22485 -11255
rect 22530 -11375 22650 -11255
rect 22705 -11375 22825 -11255
rect 22870 -11375 22990 -11255
rect 23035 -11375 23155 -11255
rect 23200 -11375 23320 -11255
rect 23375 -11375 23495 -11255
rect 23540 -11375 23660 -11255
rect 23705 -11375 23825 -11255
rect 23870 -11375 23990 -11255
rect 18510 -11550 18630 -11430
rect 18685 -11550 18805 -11430
rect 18850 -11550 18970 -11430
rect 19015 -11550 19135 -11430
rect 19180 -11550 19300 -11430
rect 19355 -11550 19475 -11430
rect 19520 -11550 19640 -11430
rect 19685 -11550 19805 -11430
rect 19850 -11550 19970 -11430
rect 20025 -11550 20145 -11430
rect 20190 -11550 20310 -11430
rect 20355 -11550 20475 -11430
rect 20520 -11550 20640 -11430
rect 20695 -11550 20815 -11430
rect 20860 -11550 20980 -11430
rect 21025 -11550 21145 -11430
rect 21190 -11550 21310 -11430
rect 21365 -11550 21485 -11430
rect 21530 -11550 21650 -11430
rect 21695 -11550 21815 -11430
rect 21860 -11550 21980 -11430
rect 22035 -11550 22155 -11430
rect 22200 -11550 22320 -11430
rect 22365 -11550 22485 -11430
rect 22530 -11550 22650 -11430
rect 22705 -11550 22825 -11430
rect 22870 -11550 22990 -11430
rect 23035 -11550 23155 -11430
rect 23200 -11550 23320 -11430
rect 23375 -11550 23495 -11430
rect 23540 -11550 23660 -11430
rect 23705 -11550 23825 -11430
rect 23870 -11550 23990 -11430
rect 18510 -11715 18630 -11595
rect 18685 -11715 18805 -11595
rect 18850 -11715 18970 -11595
rect 19015 -11715 19135 -11595
rect 19180 -11715 19300 -11595
rect 19355 -11715 19475 -11595
rect 19520 -11715 19640 -11595
rect 19685 -11715 19805 -11595
rect 19850 -11715 19970 -11595
rect 20025 -11715 20145 -11595
rect 20190 -11715 20310 -11595
rect 20355 -11715 20475 -11595
rect 20520 -11715 20640 -11595
rect 20695 -11715 20815 -11595
rect 20860 -11715 20980 -11595
rect 21025 -11715 21145 -11595
rect 21190 -11715 21310 -11595
rect 21365 -11715 21485 -11595
rect 21530 -11715 21650 -11595
rect 21695 -11715 21815 -11595
rect 21860 -11715 21980 -11595
rect 22035 -11715 22155 -11595
rect 22200 -11715 22320 -11595
rect 22365 -11715 22485 -11595
rect 22530 -11715 22650 -11595
rect 22705 -11715 22825 -11595
rect 22870 -11715 22990 -11595
rect 23035 -11715 23155 -11595
rect 23200 -11715 23320 -11595
rect 23375 -11715 23495 -11595
rect 23540 -11715 23660 -11595
rect 23705 -11715 23825 -11595
rect 23870 -11715 23990 -11595
rect 18510 -11880 18630 -11760
rect 18685 -11880 18805 -11760
rect 18850 -11880 18970 -11760
rect 19015 -11880 19135 -11760
rect 19180 -11880 19300 -11760
rect 19355 -11880 19475 -11760
rect 19520 -11880 19640 -11760
rect 19685 -11880 19805 -11760
rect 19850 -11880 19970 -11760
rect 20025 -11880 20145 -11760
rect 20190 -11880 20310 -11760
rect 20355 -11880 20475 -11760
rect 20520 -11880 20640 -11760
rect 20695 -11880 20815 -11760
rect 20860 -11880 20980 -11760
rect 21025 -11880 21145 -11760
rect 21190 -11880 21310 -11760
rect 21365 -11880 21485 -11760
rect 21530 -11880 21650 -11760
rect 21695 -11880 21815 -11760
rect 21860 -11880 21980 -11760
rect 22035 -11880 22155 -11760
rect 22200 -11880 22320 -11760
rect 22365 -11880 22485 -11760
rect 22530 -11880 22650 -11760
rect 22705 -11880 22825 -11760
rect 22870 -11880 22990 -11760
rect 23035 -11880 23155 -11760
rect 23200 -11880 23320 -11760
rect 23375 -11880 23495 -11760
rect 23540 -11880 23660 -11760
rect 23705 -11880 23825 -11760
rect 23870 -11880 23990 -11760
rect 18510 -12045 18630 -11925
rect 18685 -12045 18805 -11925
rect 18850 -12045 18970 -11925
rect 19015 -12045 19135 -11925
rect 19180 -12045 19300 -11925
rect 19355 -12045 19475 -11925
rect 19520 -12045 19640 -11925
rect 19685 -12045 19805 -11925
rect 19850 -12045 19970 -11925
rect 20025 -12045 20145 -11925
rect 20190 -12045 20310 -11925
rect 20355 -12045 20475 -11925
rect 20520 -12045 20640 -11925
rect 20695 -12045 20815 -11925
rect 20860 -12045 20980 -11925
rect 21025 -12045 21145 -11925
rect 21190 -12045 21310 -11925
rect 21365 -12045 21485 -11925
rect 21530 -12045 21650 -11925
rect 21695 -12045 21815 -11925
rect 21860 -12045 21980 -11925
rect 22035 -12045 22155 -11925
rect 22200 -12045 22320 -11925
rect 22365 -12045 22485 -11925
rect 22530 -12045 22650 -11925
rect 22705 -12045 22825 -11925
rect 22870 -12045 22990 -11925
rect 23035 -12045 23155 -11925
rect 23200 -12045 23320 -11925
rect 23375 -12045 23495 -11925
rect 23540 -12045 23660 -11925
rect 23705 -12045 23825 -11925
rect 23870 -12045 23990 -11925
rect 18510 -12220 18630 -12100
rect 18685 -12220 18805 -12100
rect 18850 -12220 18970 -12100
rect 19015 -12220 19135 -12100
rect 19180 -12220 19300 -12100
rect 19355 -12220 19475 -12100
rect 19520 -12220 19640 -12100
rect 19685 -12220 19805 -12100
rect 19850 -12220 19970 -12100
rect 20025 -12220 20145 -12100
rect 20190 -12220 20310 -12100
rect 20355 -12220 20475 -12100
rect 20520 -12220 20640 -12100
rect 20695 -12220 20815 -12100
rect 20860 -12220 20980 -12100
rect 21025 -12220 21145 -12100
rect 21190 -12220 21310 -12100
rect 21365 -12220 21485 -12100
rect 21530 -12220 21650 -12100
rect 21695 -12220 21815 -12100
rect 21860 -12220 21980 -12100
rect 22035 -12220 22155 -12100
rect 22200 -12220 22320 -12100
rect 22365 -12220 22485 -12100
rect 22530 -12220 22650 -12100
rect 22705 -12220 22825 -12100
rect 22870 -12220 22990 -12100
rect 23035 -12220 23155 -12100
rect 23200 -12220 23320 -12100
rect 23375 -12220 23495 -12100
rect 23540 -12220 23660 -12100
rect 23705 -12220 23825 -12100
rect 23870 -12220 23990 -12100
rect 18510 -12385 18630 -12265
rect 18685 -12385 18805 -12265
rect 18850 -12385 18970 -12265
rect 19015 -12385 19135 -12265
rect 19180 -12385 19300 -12265
rect 19355 -12385 19475 -12265
rect 19520 -12385 19640 -12265
rect 19685 -12385 19805 -12265
rect 19850 -12385 19970 -12265
rect 20025 -12385 20145 -12265
rect 20190 -12385 20310 -12265
rect 20355 -12385 20475 -12265
rect 20520 -12385 20640 -12265
rect 20695 -12385 20815 -12265
rect 20860 -12385 20980 -12265
rect 21025 -12385 21145 -12265
rect 21190 -12385 21310 -12265
rect 21365 -12385 21485 -12265
rect 21530 -12385 21650 -12265
rect 21695 -12385 21815 -12265
rect 21860 -12385 21980 -12265
rect 22035 -12385 22155 -12265
rect 22200 -12385 22320 -12265
rect 22365 -12385 22485 -12265
rect 22530 -12385 22650 -12265
rect 22705 -12385 22825 -12265
rect 22870 -12385 22990 -12265
rect 23035 -12385 23155 -12265
rect 23200 -12385 23320 -12265
rect 23375 -12385 23495 -12265
rect 23540 -12385 23660 -12265
rect 23705 -12385 23825 -12265
rect 23870 -12385 23990 -12265
rect 18510 -12550 18630 -12430
rect 18685 -12550 18805 -12430
rect 18850 -12550 18970 -12430
rect 19015 -12550 19135 -12430
rect 19180 -12550 19300 -12430
rect 19355 -12550 19475 -12430
rect 19520 -12550 19640 -12430
rect 19685 -12550 19805 -12430
rect 19850 -12550 19970 -12430
rect 20025 -12550 20145 -12430
rect 20190 -12550 20310 -12430
rect 20355 -12550 20475 -12430
rect 20520 -12550 20640 -12430
rect 20695 -12550 20815 -12430
rect 20860 -12550 20980 -12430
rect 21025 -12550 21145 -12430
rect 21190 -12550 21310 -12430
rect 21365 -12550 21485 -12430
rect 21530 -12550 21650 -12430
rect 21695 -12550 21815 -12430
rect 21860 -12550 21980 -12430
rect 22035 -12550 22155 -12430
rect 22200 -12550 22320 -12430
rect 22365 -12550 22485 -12430
rect 22530 -12550 22650 -12430
rect 22705 -12550 22825 -12430
rect 22870 -12550 22990 -12430
rect 23035 -12550 23155 -12430
rect 23200 -12550 23320 -12430
rect 23375 -12550 23495 -12430
rect 23540 -12550 23660 -12430
rect 23705 -12550 23825 -12430
rect 23870 -12550 23990 -12430
rect 18510 -12715 18630 -12595
rect 18685 -12715 18805 -12595
rect 18850 -12715 18970 -12595
rect 19015 -12715 19135 -12595
rect 19180 -12715 19300 -12595
rect 19355 -12715 19475 -12595
rect 19520 -12715 19640 -12595
rect 19685 -12715 19805 -12595
rect 19850 -12715 19970 -12595
rect 20025 -12715 20145 -12595
rect 20190 -12715 20310 -12595
rect 20355 -12715 20475 -12595
rect 20520 -12715 20640 -12595
rect 20695 -12715 20815 -12595
rect 20860 -12715 20980 -12595
rect 21025 -12715 21145 -12595
rect 21190 -12715 21310 -12595
rect 21365 -12715 21485 -12595
rect 21530 -12715 21650 -12595
rect 21695 -12715 21815 -12595
rect 21860 -12715 21980 -12595
rect 22035 -12715 22155 -12595
rect 22200 -12715 22320 -12595
rect 22365 -12715 22485 -12595
rect 22530 -12715 22650 -12595
rect 22705 -12715 22825 -12595
rect 22870 -12715 22990 -12595
rect 23035 -12715 23155 -12595
rect 23200 -12715 23320 -12595
rect 23375 -12715 23495 -12595
rect 23540 -12715 23660 -12595
rect 23705 -12715 23825 -12595
rect 23870 -12715 23990 -12595
rect 18510 -12890 18630 -12770
rect 18685 -12890 18805 -12770
rect 18850 -12890 18970 -12770
rect 19015 -12890 19135 -12770
rect 19180 -12890 19300 -12770
rect 19355 -12890 19475 -12770
rect 19520 -12890 19640 -12770
rect 19685 -12890 19805 -12770
rect 19850 -12890 19970 -12770
rect 20025 -12890 20145 -12770
rect 20190 -12890 20310 -12770
rect 20355 -12890 20475 -12770
rect 20520 -12890 20640 -12770
rect 20695 -12890 20815 -12770
rect 20860 -12890 20980 -12770
rect 21025 -12890 21145 -12770
rect 21190 -12890 21310 -12770
rect 21365 -12890 21485 -12770
rect 21530 -12890 21650 -12770
rect 21695 -12890 21815 -12770
rect 21860 -12890 21980 -12770
rect 22035 -12890 22155 -12770
rect 22200 -12890 22320 -12770
rect 22365 -12890 22485 -12770
rect 22530 -12890 22650 -12770
rect 22705 -12890 22825 -12770
rect 22870 -12890 22990 -12770
rect 23035 -12890 23155 -12770
rect 23200 -12890 23320 -12770
rect 23375 -12890 23495 -12770
rect 23540 -12890 23660 -12770
rect 23705 -12890 23825 -12770
rect 23870 -12890 23990 -12770
rect 18510 -13055 18630 -12935
rect 18685 -13055 18805 -12935
rect 18850 -13055 18970 -12935
rect 19015 -13055 19135 -12935
rect 19180 -13055 19300 -12935
rect 19355 -13055 19475 -12935
rect 19520 -13055 19640 -12935
rect 19685 -13055 19805 -12935
rect 19850 -13055 19970 -12935
rect 20025 -13055 20145 -12935
rect 20190 -13055 20310 -12935
rect 20355 -13055 20475 -12935
rect 20520 -13055 20640 -12935
rect 20695 -13055 20815 -12935
rect 20860 -13055 20980 -12935
rect 21025 -13055 21145 -12935
rect 21190 -13055 21310 -12935
rect 21365 -13055 21485 -12935
rect 21530 -13055 21650 -12935
rect 21695 -13055 21815 -12935
rect 21860 -13055 21980 -12935
rect 22035 -13055 22155 -12935
rect 22200 -13055 22320 -12935
rect 22365 -13055 22485 -12935
rect 22530 -13055 22650 -12935
rect 22705 -13055 22825 -12935
rect 22870 -13055 22990 -12935
rect 23035 -13055 23155 -12935
rect 23200 -13055 23320 -12935
rect 23375 -13055 23495 -12935
rect 23540 -13055 23660 -12935
rect 23705 -13055 23825 -12935
rect 23870 -13055 23990 -12935
rect 18510 -13220 18630 -13100
rect 18685 -13220 18805 -13100
rect 18850 -13220 18970 -13100
rect 19015 -13220 19135 -13100
rect 19180 -13220 19300 -13100
rect 19355 -13220 19475 -13100
rect 19520 -13220 19640 -13100
rect 19685 -13220 19805 -13100
rect 19850 -13220 19970 -13100
rect 20025 -13220 20145 -13100
rect 20190 -13220 20310 -13100
rect 20355 -13220 20475 -13100
rect 20520 -13220 20640 -13100
rect 20695 -13220 20815 -13100
rect 20860 -13220 20980 -13100
rect 21025 -13220 21145 -13100
rect 21190 -13220 21310 -13100
rect 21365 -13220 21485 -13100
rect 21530 -13220 21650 -13100
rect 21695 -13220 21815 -13100
rect 21860 -13220 21980 -13100
rect 22035 -13220 22155 -13100
rect 22200 -13220 22320 -13100
rect 22365 -13220 22485 -13100
rect 22530 -13220 22650 -13100
rect 22705 -13220 22825 -13100
rect 22870 -13220 22990 -13100
rect 23035 -13220 23155 -13100
rect 23200 -13220 23320 -13100
rect 23375 -13220 23495 -13100
rect 23540 -13220 23660 -13100
rect 23705 -13220 23825 -13100
rect 23870 -13220 23990 -13100
rect 18510 -13385 18630 -13265
rect 18685 -13385 18805 -13265
rect 18850 -13385 18970 -13265
rect 19015 -13385 19135 -13265
rect 19180 -13385 19300 -13265
rect 19355 -13385 19475 -13265
rect 19520 -13385 19640 -13265
rect 19685 -13385 19805 -13265
rect 19850 -13385 19970 -13265
rect 20025 -13385 20145 -13265
rect 20190 -13385 20310 -13265
rect 20355 -13385 20475 -13265
rect 20520 -13385 20640 -13265
rect 20695 -13385 20815 -13265
rect 20860 -13385 20980 -13265
rect 21025 -13385 21145 -13265
rect 21190 -13385 21310 -13265
rect 21365 -13385 21485 -13265
rect 21530 -13385 21650 -13265
rect 21695 -13385 21815 -13265
rect 21860 -13385 21980 -13265
rect 22035 -13385 22155 -13265
rect 22200 -13385 22320 -13265
rect 22365 -13385 22485 -13265
rect 22530 -13385 22650 -13265
rect 22705 -13385 22825 -13265
rect 22870 -13385 22990 -13265
rect 23035 -13385 23155 -13265
rect 23200 -13385 23320 -13265
rect 23375 -13385 23495 -13265
rect 23540 -13385 23660 -13265
rect 23705 -13385 23825 -13265
rect 23870 -13385 23990 -13265
rect 18510 -13560 18630 -13440
rect 18685 -13560 18805 -13440
rect 18850 -13560 18970 -13440
rect 19015 -13560 19135 -13440
rect 19180 -13560 19300 -13440
rect 19355 -13560 19475 -13440
rect 19520 -13560 19640 -13440
rect 19685 -13560 19805 -13440
rect 19850 -13560 19970 -13440
rect 20025 -13560 20145 -13440
rect 20190 -13560 20310 -13440
rect 20355 -13560 20475 -13440
rect 20520 -13560 20640 -13440
rect 20695 -13560 20815 -13440
rect 20860 -13560 20980 -13440
rect 21025 -13560 21145 -13440
rect 21190 -13560 21310 -13440
rect 21365 -13560 21485 -13440
rect 21530 -13560 21650 -13440
rect 21695 -13560 21815 -13440
rect 21860 -13560 21980 -13440
rect 22035 -13560 22155 -13440
rect 22200 -13560 22320 -13440
rect 22365 -13560 22485 -13440
rect 22530 -13560 22650 -13440
rect 22705 -13560 22825 -13440
rect 22870 -13560 22990 -13440
rect 23035 -13560 23155 -13440
rect 23200 -13560 23320 -13440
rect 23375 -13560 23495 -13440
rect 23540 -13560 23660 -13440
rect 23705 -13560 23825 -13440
rect 23870 -13560 23990 -13440
rect 18510 -13725 18630 -13605
rect 18685 -13725 18805 -13605
rect 18850 -13725 18970 -13605
rect 19015 -13725 19135 -13605
rect 19180 -13725 19300 -13605
rect 19355 -13725 19475 -13605
rect 19520 -13725 19640 -13605
rect 19685 -13725 19805 -13605
rect 19850 -13725 19970 -13605
rect 20025 -13725 20145 -13605
rect 20190 -13725 20310 -13605
rect 20355 -13725 20475 -13605
rect 20520 -13725 20640 -13605
rect 20695 -13725 20815 -13605
rect 20860 -13725 20980 -13605
rect 21025 -13725 21145 -13605
rect 21190 -13725 21310 -13605
rect 21365 -13725 21485 -13605
rect 21530 -13725 21650 -13605
rect 21695 -13725 21815 -13605
rect 21860 -13725 21980 -13605
rect 22035 -13725 22155 -13605
rect 22200 -13725 22320 -13605
rect 22365 -13725 22485 -13605
rect 22530 -13725 22650 -13605
rect 22705 -13725 22825 -13605
rect 22870 -13725 22990 -13605
rect 23035 -13725 23155 -13605
rect 23200 -13725 23320 -13605
rect 23375 -13725 23495 -13605
rect 23540 -13725 23660 -13605
rect 23705 -13725 23825 -13605
rect 23870 -13725 23990 -13605
rect 18510 -13890 18630 -13770
rect 18685 -13890 18805 -13770
rect 18850 -13890 18970 -13770
rect 19015 -13890 19135 -13770
rect 19180 -13890 19300 -13770
rect 19355 -13890 19475 -13770
rect 19520 -13890 19640 -13770
rect 19685 -13890 19805 -13770
rect 19850 -13890 19970 -13770
rect 20025 -13890 20145 -13770
rect 20190 -13890 20310 -13770
rect 20355 -13890 20475 -13770
rect 20520 -13890 20640 -13770
rect 20695 -13890 20815 -13770
rect 20860 -13890 20980 -13770
rect 21025 -13890 21145 -13770
rect 21190 -13890 21310 -13770
rect 21365 -13890 21485 -13770
rect 21530 -13890 21650 -13770
rect 21695 -13890 21815 -13770
rect 21860 -13890 21980 -13770
rect 22035 -13890 22155 -13770
rect 22200 -13890 22320 -13770
rect 22365 -13890 22485 -13770
rect 22530 -13890 22650 -13770
rect 22705 -13890 22825 -13770
rect 22870 -13890 22990 -13770
rect 23035 -13890 23155 -13770
rect 23200 -13890 23320 -13770
rect 23375 -13890 23495 -13770
rect 23540 -13890 23660 -13770
rect 23705 -13890 23825 -13770
rect 23870 -13890 23990 -13770
rect 18510 -14055 18630 -13935
rect 18685 -14055 18805 -13935
rect 18850 -14055 18970 -13935
rect 19015 -14055 19135 -13935
rect 19180 -14055 19300 -13935
rect 19355 -14055 19475 -13935
rect 19520 -14055 19640 -13935
rect 19685 -14055 19805 -13935
rect 19850 -14055 19970 -13935
rect 20025 -14055 20145 -13935
rect 20190 -14055 20310 -13935
rect 20355 -14055 20475 -13935
rect 20520 -14055 20640 -13935
rect 20695 -14055 20815 -13935
rect 20860 -14055 20980 -13935
rect 21025 -14055 21145 -13935
rect 21190 -14055 21310 -13935
rect 21365 -14055 21485 -13935
rect 21530 -14055 21650 -13935
rect 21695 -14055 21815 -13935
rect 21860 -14055 21980 -13935
rect 22035 -14055 22155 -13935
rect 22200 -14055 22320 -13935
rect 22365 -14055 22485 -13935
rect 22530 -14055 22650 -13935
rect 22705 -14055 22825 -13935
rect 22870 -14055 22990 -13935
rect 23035 -14055 23155 -13935
rect 23200 -14055 23320 -13935
rect 23375 -14055 23495 -13935
rect 23540 -14055 23660 -13935
rect 23705 -14055 23825 -13935
rect 23870 -14055 23990 -13935
rect 18510 -14230 18630 -14110
rect 18685 -14230 18805 -14110
rect 18850 -14230 18970 -14110
rect 19015 -14230 19135 -14110
rect 19180 -14230 19300 -14110
rect 19355 -14230 19475 -14110
rect 19520 -14230 19640 -14110
rect 19685 -14230 19805 -14110
rect 19850 -14230 19970 -14110
rect 20025 -14230 20145 -14110
rect 20190 -14230 20310 -14110
rect 20355 -14230 20475 -14110
rect 20520 -14230 20640 -14110
rect 20695 -14230 20815 -14110
rect 20860 -14230 20980 -14110
rect 21025 -14230 21145 -14110
rect 21190 -14230 21310 -14110
rect 21365 -14230 21485 -14110
rect 21530 -14230 21650 -14110
rect 21695 -14230 21815 -14110
rect 21860 -14230 21980 -14110
rect 22035 -14230 22155 -14110
rect 22200 -14230 22320 -14110
rect 22365 -14230 22485 -14110
rect 22530 -14230 22650 -14110
rect 22705 -14230 22825 -14110
rect 22870 -14230 22990 -14110
rect 23035 -14230 23155 -14110
rect 23200 -14230 23320 -14110
rect 23375 -14230 23495 -14110
rect 23540 -14230 23660 -14110
rect 23705 -14230 23825 -14110
rect 23870 -14230 23990 -14110
rect 18510 -14395 18630 -14275
rect 18685 -14395 18805 -14275
rect 18850 -14395 18970 -14275
rect 19015 -14395 19135 -14275
rect 19180 -14395 19300 -14275
rect 19355 -14395 19475 -14275
rect 19520 -14395 19640 -14275
rect 19685 -14395 19805 -14275
rect 19850 -14395 19970 -14275
rect 20025 -14395 20145 -14275
rect 20190 -14395 20310 -14275
rect 20355 -14395 20475 -14275
rect 20520 -14395 20640 -14275
rect 20695 -14395 20815 -14275
rect 20860 -14395 20980 -14275
rect 21025 -14395 21145 -14275
rect 21190 -14395 21310 -14275
rect 21365 -14395 21485 -14275
rect 21530 -14395 21650 -14275
rect 21695 -14395 21815 -14275
rect 21860 -14395 21980 -14275
rect 22035 -14395 22155 -14275
rect 22200 -14395 22320 -14275
rect 22365 -14395 22485 -14275
rect 22530 -14395 22650 -14275
rect 22705 -14395 22825 -14275
rect 22870 -14395 22990 -14275
rect 23035 -14395 23155 -14275
rect 23200 -14395 23320 -14275
rect 23375 -14395 23495 -14275
rect 23540 -14395 23660 -14275
rect 23705 -14395 23825 -14275
rect 23870 -14395 23990 -14275
rect 18510 -14560 18630 -14440
rect 18685 -14560 18805 -14440
rect 18850 -14560 18970 -14440
rect 19015 -14560 19135 -14440
rect 19180 -14560 19300 -14440
rect 19355 -14560 19475 -14440
rect 19520 -14560 19640 -14440
rect 19685 -14560 19805 -14440
rect 19850 -14560 19970 -14440
rect 20025 -14560 20145 -14440
rect 20190 -14560 20310 -14440
rect 20355 -14560 20475 -14440
rect 20520 -14560 20640 -14440
rect 20695 -14560 20815 -14440
rect 20860 -14560 20980 -14440
rect 21025 -14560 21145 -14440
rect 21190 -14560 21310 -14440
rect 21365 -14560 21485 -14440
rect 21530 -14560 21650 -14440
rect 21695 -14560 21815 -14440
rect 21860 -14560 21980 -14440
rect 22035 -14560 22155 -14440
rect 22200 -14560 22320 -14440
rect 22365 -14560 22485 -14440
rect 22530 -14560 22650 -14440
rect 22705 -14560 22825 -14440
rect 22870 -14560 22990 -14440
rect 23035 -14560 23155 -14440
rect 23200 -14560 23320 -14440
rect 23375 -14560 23495 -14440
rect 23540 -14560 23660 -14440
rect 23705 -14560 23825 -14440
rect 23870 -14560 23990 -14440
rect 18510 -14725 18630 -14605
rect 18685 -14725 18805 -14605
rect 18850 -14725 18970 -14605
rect 19015 -14725 19135 -14605
rect 19180 -14725 19300 -14605
rect 19355 -14725 19475 -14605
rect 19520 -14725 19640 -14605
rect 19685 -14725 19805 -14605
rect 19850 -14725 19970 -14605
rect 20025 -14725 20145 -14605
rect 20190 -14725 20310 -14605
rect 20355 -14725 20475 -14605
rect 20520 -14725 20640 -14605
rect 20695 -14725 20815 -14605
rect 20860 -14725 20980 -14605
rect 21025 -14725 21145 -14605
rect 21190 -14725 21310 -14605
rect 21365 -14725 21485 -14605
rect 21530 -14725 21650 -14605
rect 21695 -14725 21815 -14605
rect 21860 -14725 21980 -14605
rect 22035 -14725 22155 -14605
rect 22200 -14725 22320 -14605
rect 22365 -14725 22485 -14605
rect 22530 -14725 22650 -14605
rect 22705 -14725 22825 -14605
rect 22870 -14725 22990 -14605
rect 23035 -14725 23155 -14605
rect 23200 -14725 23320 -14605
rect 23375 -14725 23495 -14605
rect 23540 -14725 23660 -14605
rect 23705 -14725 23825 -14605
rect 23870 -14725 23990 -14605
rect 18510 -14900 18630 -14780
rect 18685 -14900 18805 -14780
rect 18850 -14900 18970 -14780
rect 19015 -14900 19135 -14780
rect 19180 -14900 19300 -14780
rect 19355 -14900 19475 -14780
rect 19520 -14900 19640 -14780
rect 19685 -14900 19805 -14780
rect 19850 -14900 19970 -14780
rect 20025 -14900 20145 -14780
rect 20190 -14900 20310 -14780
rect 20355 -14900 20475 -14780
rect 20520 -14900 20640 -14780
rect 20695 -14900 20815 -14780
rect 20860 -14900 20980 -14780
rect 21025 -14900 21145 -14780
rect 21190 -14900 21310 -14780
rect 21365 -14900 21485 -14780
rect 21530 -14900 21650 -14780
rect 21695 -14900 21815 -14780
rect 21860 -14900 21980 -14780
rect 22035 -14900 22155 -14780
rect 22200 -14900 22320 -14780
rect 22365 -14900 22485 -14780
rect 22530 -14900 22650 -14780
rect 22705 -14900 22825 -14780
rect 22870 -14900 22990 -14780
rect 23035 -14900 23155 -14780
rect 23200 -14900 23320 -14780
rect 23375 -14900 23495 -14780
rect 23540 -14900 23660 -14780
rect 23705 -14900 23825 -14780
rect 23870 -14900 23990 -14780
rect 18510 -15065 18630 -14945
rect 18685 -15065 18805 -14945
rect 18850 -15065 18970 -14945
rect 19015 -15065 19135 -14945
rect 19180 -15065 19300 -14945
rect 19355 -15065 19475 -14945
rect 19520 -15065 19640 -14945
rect 19685 -15065 19805 -14945
rect 19850 -15065 19970 -14945
rect 20025 -15065 20145 -14945
rect 20190 -15065 20310 -14945
rect 20355 -15065 20475 -14945
rect 20520 -15065 20640 -14945
rect 20695 -15065 20815 -14945
rect 20860 -15065 20980 -14945
rect 21025 -15065 21145 -14945
rect 21190 -15065 21310 -14945
rect 21365 -15065 21485 -14945
rect 21530 -15065 21650 -14945
rect 21695 -15065 21815 -14945
rect 21860 -15065 21980 -14945
rect 22035 -15065 22155 -14945
rect 22200 -15065 22320 -14945
rect 22365 -15065 22485 -14945
rect 22530 -15065 22650 -14945
rect 22705 -15065 22825 -14945
rect 22870 -15065 22990 -14945
rect 23035 -15065 23155 -14945
rect 23200 -15065 23320 -14945
rect 23375 -15065 23495 -14945
rect 23540 -15065 23660 -14945
rect 23705 -15065 23825 -14945
rect 23870 -15065 23990 -14945
rect 18510 -15230 18630 -15110
rect 18685 -15230 18805 -15110
rect 18850 -15230 18970 -15110
rect 19015 -15230 19135 -15110
rect 19180 -15230 19300 -15110
rect 19355 -15230 19475 -15110
rect 19520 -15230 19640 -15110
rect 19685 -15230 19805 -15110
rect 19850 -15230 19970 -15110
rect 20025 -15230 20145 -15110
rect 20190 -15230 20310 -15110
rect 20355 -15230 20475 -15110
rect 20520 -15230 20640 -15110
rect 20695 -15230 20815 -15110
rect 20860 -15230 20980 -15110
rect 21025 -15230 21145 -15110
rect 21190 -15230 21310 -15110
rect 21365 -15230 21485 -15110
rect 21530 -15230 21650 -15110
rect 21695 -15230 21815 -15110
rect 21860 -15230 21980 -15110
rect 22035 -15230 22155 -15110
rect 22200 -15230 22320 -15110
rect 22365 -15230 22485 -15110
rect 22530 -15230 22650 -15110
rect 22705 -15230 22825 -15110
rect 22870 -15230 22990 -15110
rect 23035 -15230 23155 -15110
rect 23200 -15230 23320 -15110
rect 23375 -15230 23495 -15110
rect 23540 -15230 23660 -15110
rect 23705 -15230 23825 -15110
rect 23870 -15230 23990 -15110
rect 18510 -15395 18630 -15275
rect 18685 -15395 18805 -15275
rect 18850 -15395 18970 -15275
rect 19015 -15395 19135 -15275
rect 19180 -15395 19300 -15275
rect 19355 -15395 19475 -15275
rect 19520 -15395 19640 -15275
rect 19685 -15395 19805 -15275
rect 19850 -15395 19970 -15275
rect 20025 -15395 20145 -15275
rect 20190 -15395 20310 -15275
rect 20355 -15395 20475 -15275
rect 20520 -15395 20640 -15275
rect 20695 -15395 20815 -15275
rect 20860 -15395 20980 -15275
rect 21025 -15395 21145 -15275
rect 21190 -15395 21310 -15275
rect 21365 -15395 21485 -15275
rect 21530 -15395 21650 -15275
rect 21695 -15395 21815 -15275
rect 21860 -15395 21980 -15275
rect 22035 -15395 22155 -15275
rect 22200 -15395 22320 -15275
rect 22365 -15395 22485 -15275
rect 22530 -15395 22650 -15275
rect 22705 -15395 22825 -15275
rect 22870 -15395 22990 -15275
rect 23035 -15395 23155 -15275
rect 23200 -15395 23320 -15275
rect 23375 -15395 23495 -15275
rect 23540 -15395 23660 -15275
rect 23705 -15395 23825 -15275
rect 23870 -15395 23990 -15275
rect 18510 -15570 18630 -15450
rect 18685 -15570 18805 -15450
rect 18850 -15570 18970 -15450
rect 19015 -15570 19135 -15450
rect 19180 -15570 19300 -15450
rect 19355 -15570 19475 -15450
rect 19520 -15570 19640 -15450
rect 19685 -15570 19805 -15450
rect 19850 -15570 19970 -15450
rect 20025 -15570 20145 -15450
rect 20190 -15570 20310 -15450
rect 20355 -15570 20475 -15450
rect 20520 -15570 20640 -15450
rect 20695 -15570 20815 -15450
rect 20860 -15570 20980 -15450
rect 21025 -15570 21145 -15450
rect 21190 -15570 21310 -15450
rect 21365 -15570 21485 -15450
rect 21530 -15570 21650 -15450
rect 21695 -15570 21815 -15450
rect 21860 -15570 21980 -15450
rect 22035 -15570 22155 -15450
rect 22200 -15570 22320 -15450
rect 22365 -15570 22485 -15450
rect 22530 -15570 22650 -15450
rect 22705 -15570 22825 -15450
rect 22870 -15570 22990 -15450
rect 23035 -15570 23155 -15450
rect 23200 -15570 23320 -15450
rect 23375 -15570 23495 -15450
rect 23540 -15570 23660 -15450
rect 23705 -15570 23825 -15450
rect 23870 -15570 23990 -15450
rect 24200 -10210 24320 -10090
rect 24375 -10210 24495 -10090
rect 24540 -10210 24660 -10090
rect 24705 -10210 24825 -10090
rect 24870 -10210 24990 -10090
rect 25045 -10210 25165 -10090
rect 25210 -10210 25330 -10090
rect 25375 -10210 25495 -10090
rect 25540 -10210 25660 -10090
rect 25715 -10210 25835 -10090
rect 25880 -10210 26000 -10090
rect 26045 -10210 26165 -10090
rect 26210 -10210 26330 -10090
rect 26385 -10210 26505 -10090
rect 26550 -10210 26670 -10090
rect 26715 -10210 26835 -10090
rect 26880 -10210 27000 -10090
rect 27055 -10210 27175 -10090
rect 27220 -10210 27340 -10090
rect 27385 -10210 27505 -10090
rect 27550 -10210 27670 -10090
rect 27725 -10210 27845 -10090
rect 27890 -10210 28010 -10090
rect 28055 -10210 28175 -10090
rect 28220 -10210 28340 -10090
rect 28395 -10210 28515 -10090
rect 28560 -10210 28680 -10090
rect 28725 -10210 28845 -10090
rect 28890 -10210 29010 -10090
rect 29065 -10210 29185 -10090
rect 29230 -10210 29350 -10090
rect 29395 -10210 29515 -10090
rect 29560 -10210 29680 -10090
rect 24200 -10375 24320 -10255
rect 24375 -10375 24495 -10255
rect 24540 -10375 24660 -10255
rect 24705 -10375 24825 -10255
rect 24870 -10375 24990 -10255
rect 25045 -10375 25165 -10255
rect 25210 -10375 25330 -10255
rect 25375 -10375 25495 -10255
rect 25540 -10375 25660 -10255
rect 25715 -10375 25835 -10255
rect 25880 -10375 26000 -10255
rect 26045 -10375 26165 -10255
rect 26210 -10375 26330 -10255
rect 26385 -10375 26505 -10255
rect 26550 -10375 26670 -10255
rect 26715 -10375 26835 -10255
rect 26880 -10375 27000 -10255
rect 27055 -10375 27175 -10255
rect 27220 -10375 27340 -10255
rect 27385 -10375 27505 -10255
rect 27550 -10375 27670 -10255
rect 27725 -10375 27845 -10255
rect 27890 -10375 28010 -10255
rect 28055 -10375 28175 -10255
rect 28220 -10375 28340 -10255
rect 28395 -10375 28515 -10255
rect 28560 -10375 28680 -10255
rect 28725 -10375 28845 -10255
rect 28890 -10375 29010 -10255
rect 29065 -10375 29185 -10255
rect 29230 -10375 29350 -10255
rect 29395 -10375 29515 -10255
rect 29560 -10375 29680 -10255
rect 24200 -10540 24320 -10420
rect 24375 -10540 24495 -10420
rect 24540 -10540 24660 -10420
rect 24705 -10540 24825 -10420
rect 24870 -10540 24990 -10420
rect 25045 -10540 25165 -10420
rect 25210 -10540 25330 -10420
rect 25375 -10540 25495 -10420
rect 25540 -10540 25660 -10420
rect 25715 -10540 25835 -10420
rect 25880 -10540 26000 -10420
rect 26045 -10540 26165 -10420
rect 26210 -10540 26330 -10420
rect 26385 -10540 26505 -10420
rect 26550 -10540 26670 -10420
rect 26715 -10540 26835 -10420
rect 26880 -10540 27000 -10420
rect 27055 -10540 27175 -10420
rect 27220 -10540 27340 -10420
rect 27385 -10540 27505 -10420
rect 27550 -10540 27670 -10420
rect 27725 -10540 27845 -10420
rect 27890 -10540 28010 -10420
rect 28055 -10540 28175 -10420
rect 28220 -10540 28340 -10420
rect 28395 -10540 28515 -10420
rect 28560 -10540 28680 -10420
rect 28725 -10540 28845 -10420
rect 28890 -10540 29010 -10420
rect 29065 -10540 29185 -10420
rect 29230 -10540 29350 -10420
rect 29395 -10540 29515 -10420
rect 29560 -10540 29680 -10420
rect 24200 -10705 24320 -10585
rect 24375 -10705 24495 -10585
rect 24540 -10705 24660 -10585
rect 24705 -10705 24825 -10585
rect 24870 -10705 24990 -10585
rect 25045 -10705 25165 -10585
rect 25210 -10705 25330 -10585
rect 25375 -10705 25495 -10585
rect 25540 -10705 25660 -10585
rect 25715 -10705 25835 -10585
rect 25880 -10705 26000 -10585
rect 26045 -10705 26165 -10585
rect 26210 -10705 26330 -10585
rect 26385 -10705 26505 -10585
rect 26550 -10705 26670 -10585
rect 26715 -10705 26835 -10585
rect 26880 -10705 27000 -10585
rect 27055 -10705 27175 -10585
rect 27220 -10705 27340 -10585
rect 27385 -10705 27505 -10585
rect 27550 -10705 27670 -10585
rect 27725 -10705 27845 -10585
rect 27890 -10705 28010 -10585
rect 28055 -10705 28175 -10585
rect 28220 -10705 28340 -10585
rect 28395 -10705 28515 -10585
rect 28560 -10705 28680 -10585
rect 28725 -10705 28845 -10585
rect 28890 -10705 29010 -10585
rect 29065 -10705 29185 -10585
rect 29230 -10705 29350 -10585
rect 29395 -10705 29515 -10585
rect 29560 -10705 29680 -10585
rect 24200 -10880 24320 -10760
rect 24375 -10880 24495 -10760
rect 24540 -10880 24660 -10760
rect 24705 -10880 24825 -10760
rect 24870 -10880 24990 -10760
rect 25045 -10880 25165 -10760
rect 25210 -10880 25330 -10760
rect 25375 -10880 25495 -10760
rect 25540 -10880 25660 -10760
rect 25715 -10880 25835 -10760
rect 25880 -10880 26000 -10760
rect 26045 -10880 26165 -10760
rect 26210 -10880 26330 -10760
rect 26385 -10880 26505 -10760
rect 26550 -10880 26670 -10760
rect 26715 -10880 26835 -10760
rect 26880 -10880 27000 -10760
rect 27055 -10880 27175 -10760
rect 27220 -10880 27340 -10760
rect 27385 -10880 27505 -10760
rect 27550 -10880 27670 -10760
rect 27725 -10880 27845 -10760
rect 27890 -10880 28010 -10760
rect 28055 -10880 28175 -10760
rect 28220 -10880 28340 -10760
rect 28395 -10880 28515 -10760
rect 28560 -10880 28680 -10760
rect 28725 -10880 28845 -10760
rect 28890 -10880 29010 -10760
rect 29065 -10880 29185 -10760
rect 29230 -10880 29350 -10760
rect 29395 -10880 29515 -10760
rect 29560 -10880 29680 -10760
rect 24200 -11045 24320 -10925
rect 24375 -11045 24495 -10925
rect 24540 -11045 24660 -10925
rect 24705 -11045 24825 -10925
rect 24870 -11045 24990 -10925
rect 25045 -11045 25165 -10925
rect 25210 -11045 25330 -10925
rect 25375 -11045 25495 -10925
rect 25540 -11045 25660 -10925
rect 25715 -11045 25835 -10925
rect 25880 -11045 26000 -10925
rect 26045 -11045 26165 -10925
rect 26210 -11045 26330 -10925
rect 26385 -11045 26505 -10925
rect 26550 -11045 26670 -10925
rect 26715 -11045 26835 -10925
rect 26880 -11045 27000 -10925
rect 27055 -11045 27175 -10925
rect 27220 -11045 27340 -10925
rect 27385 -11045 27505 -10925
rect 27550 -11045 27670 -10925
rect 27725 -11045 27845 -10925
rect 27890 -11045 28010 -10925
rect 28055 -11045 28175 -10925
rect 28220 -11045 28340 -10925
rect 28395 -11045 28515 -10925
rect 28560 -11045 28680 -10925
rect 28725 -11045 28845 -10925
rect 28890 -11045 29010 -10925
rect 29065 -11045 29185 -10925
rect 29230 -11045 29350 -10925
rect 29395 -11045 29515 -10925
rect 29560 -11045 29680 -10925
rect 24200 -11210 24320 -11090
rect 24375 -11210 24495 -11090
rect 24540 -11210 24660 -11090
rect 24705 -11210 24825 -11090
rect 24870 -11210 24990 -11090
rect 25045 -11210 25165 -11090
rect 25210 -11210 25330 -11090
rect 25375 -11210 25495 -11090
rect 25540 -11210 25660 -11090
rect 25715 -11210 25835 -11090
rect 25880 -11210 26000 -11090
rect 26045 -11210 26165 -11090
rect 26210 -11210 26330 -11090
rect 26385 -11210 26505 -11090
rect 26550 -11210 26670 -11090
rect 26715 -11210 26835 -11090
rect 26880 -11210 27000 -11090
rect 27055 -11210 27175 -11090
rect 27220 -11210 27340 -11090
rect 27385 -11210 27505 -11090
rect 27550 -11210 27670 -11090
rect 27725 -11210 27845 -11090
rect 27890 -11210 28010 -11090
rect 28055 -11210 28175 -11090
rect 28220 -11210 28340 -11090
rect 28395 -11210 28515 -11090
rect 28560 -11210 28680 -11090
rect 28725 -11210 28845 -11090
rect 28890 -11210 29010 -11090
rect 29065 -11210 29185 -11090
rect 29230 -11210 29350 -11090
rect 29395 -11210 29515 -11090
rect 29560 -11210 29680 -11090
rect 24200 -11375 24320 -11255
rect 24375 -11375 24495 -11255
rect 24540 -11375 24660 -11255
rect 24705 -11375 24825 -11255
rect 24870 -11375 24990 -11255
rect 25045 -11375 25165 -11255
rect 25210 -11375 25330 -11255
rect 25375 -11375 25495 -11255
rect 25540 -11375 25660 -11255
rect 25715 -11375 25835 -11255
rect 25880 -11375 26000 -11255
rect 26045 -11375 26165 -11255
rect 26210 -11375 26330 -11255
rect 26385 -11375 26505 -11255
rect 26550 -11375 26670 -11255
rect 26715 -11375 26835 -11255
rect 26880 -11375 27000 -11255
rect 27055 -11375 27175 -11255
rect 27220 -11375 27340 -11255
rect 27385 -11375 27505 -11255
rect 27550 -11375 27670 -11255
rect 27725 -11375 27845 -11255
rect 27890 -11375 28010 -11255
rect 28055 -11375 28175 -11255
rect 28220 -11375 28340 -11255
rect 28395 -11375 28515 -11255
rect 28560 -11375 28680 -11255
rect 28725 -11375 28845 -11255
rect 28890 -11375 29010 -11255
rect 29065 -11375 29185 -11255
rect 29230 -11375 29350 -11255
rect 29395 -11375 29515 -11255
rect 29560 -11375 29680 -11255
rect 24200 -11550 24320 -11430
rect 24375 -11550 24495 -11430
rect 24540 -11550 24660 -11430
rect 24705 -11550 24825 -11430
rect 24870 -11550 24990 -11430
rect 25045 -11550 25165 -11430
rect 25210 -11550 25330 -11430
rect 25375 -11550 25495 -11430
rect 25540 -11550 25660 -11430
rect 25715 -11550 25835 -11430
rect 25880 -11550 26000 -11430
rect 26045 -11550 26165 -11430
rect 26210 -11550 26330 -11430
rect 26385 -11550 26505 -11430
rect 26550 -11550 26670 -11430
rect 26715 -11550 26835 -11430
rect 26880 -11550 27000 -11430
rect 27055 -11550 27175 -11430
rect 27220 -11550 27340 -11430
rect 27385 -11550 27505 -11430
rect 27550 -11550 27670 -11430
rect 27725 -11550 27845 -11430
rect 27890 -11550 28010 -11430
rect 28055 -11550 28175 -11430
rect 28220 -11550 28340 -11430
rect 28395 -11550 28515 -11430
rect 28560 -11550 28680 -11430
rect 28725 -11550 28845 -11430
rect 28890 -11550 29010 -11430
rect 29065 -11550 29185 -11430
rect 29230 -11550 29350 -11430
rect 29395 -11550 29515 -11430
rect 29560 -11550 29680 -11430
rect 24200 -11715 24320 -11595
rect 24375 -11715 24495 -11595
rect 24540 -11715 24660 -11595
rect 24705 -11715 24825 -11595
rect 24870 -11715 24990 -11595
rect 25045 -11715 25165 -11595
rect 25210 -11715 25330 -11595
rect 25375 -11715 25495 -11595
rect 25540 -11715 25660 -11595
rect 25715 -11715 25835 -11595
rect 25880 -11715 26000 -11595
rect 26045 -11715 26165 -11595
rect 26210 -11715 26330 -11595
rect 26385 -11715 26505 -11595
rect 26550 -11715 26670 -11595
rect 26715 -11715 26835 -11595
rect 26880 -11715 27000 -11595
rect 27055 -11715 27175 -11595
rect 27220 -11715 27340 -11595
rect 27385 -11715 27505 -11595
rect 27550 -11715 27670 -11595
rect 27725 -11715 27845 -11595
rect 27890 -11715 28010 -11595
rect 28055 -11715 28175 -11595
rect 28220 -11715 28340 -11595
rect 28395 -11715 28515 -11595
rect 28560 -11715 28680 -11595
rect 28725 -11715 28845 -11595
rect 28890 -11715 29010 -11595
rect 29065 -11715 29185 -11595
rect 29230 -11715 29350 -11595
rect 29395 -11715 29515 -11595
rect 29560 -11715 29680 -11595
rect 24200 -11880 24320 -11760
rect 24375 -11880 24495 -11760
rect 24540 -11880 24660 -11760
rect 24705 -11880 24825 -11760
rect 24870 -11880 24990 -11760
rect 25045 -11880 25165 -11760
rect 25210 -11880 25330 -11760
rect 25375 -11880 25495 -11760
rect 25540 -11880 25660 -11760
rect 25715 -11880 25835 -11760
rect 25880 -11880 26000 -11760
rect 26045 -11880 26165 -11760
rect 26210 -11880 26330 -11760
rect 26385 -11880 26505 -11760
rect 26550 -11880 26670 -11760
rect 26715 -11880 26835 -11760
rect 26880 -11880 27000 -11760
rect 27055 -11880 27175 -11760
rect 27220 -11880 27340 -11760
rect 27385 -11880 27505 -11760
rect 27550 -11880 27670 -11760
rect 27725 -11880 27845 -11760
rect 27890 -11880 28010 -11760
rect 28055 -11880 28175 -11760
rect 28220 -11880 28340 -11760
rect 28395 -11880 28515 -11760
rect 28560 -11880 28680 -11760
rect 28725 -11880 28845 -11760
rect 28890 -11880 29010 -11760
rect 29065 -11880 29185 -11760
rect 29230 -11880 29350 -11760
rect 29395 -11880 29515 -11760
rect 29560 -11880 29680 -11760
rect 24200 -12045 24320 -11925
rect 24375 -12045 24495 -11925
rect 24540 -12045 24660 -11925
rect 24705 -12045 24825 -11925
rect 24870 -12045 24990 -11925
rect 25045 -12045 25165 -11925
rect 25210 -12045 25330 -11925
rect 25375 -12045 25495 -11925
rect 25540 -12045 25660 -11925
rect 25715 -12045 25835 -11925
rect 25880 -12045 26000 -11925
rect 26045 -12045 26165 -11925
rect 26210 -12045 26330 -11925
rect 26385 -12045 26505 -11925
rect 26550 -12045 26670 -11925
rect 26715 -12045 26835 -11925
rect 26880 -12045 27000 -11925
rect 27055 -12045 27175 -11925
rect 27220 -12045 27340 -11925
rect 27385 -12045 27505 -11925
rect 27550 -12045 27670 -11925
rect 27725 -12045 27845 -11925
rect 27890 -12045 28010 -11925
rect 28055 -12045 28175 -11925
rect 28220 -12045 28340 -11925
rect 28395 -12045 28515 -11925
rect 28560 -12045 28680 -11925
rect 28725 -12045 28845 -11925
rect 28890 -12045 29010 -11925
rect 29065 -12045 29185 -11925
rect 29230 -12045 29350 -11925
rect 29395 -12045 29515 -11925
rect 29560 -12045 29680 -11925
rect 24200 -12220 24320 -12100
rect 24375 -12220 24495 -12100
rect 24540 -12220 24660 -12100
rect 24705 -12220 24825 -12100
rect 24870 -12220 24990 -12100
rect 25045 -12220 25165 -12100
rect 25210 -12220 25330 -12100
rect 25375 -12220 25495 -12100
rect 25540 -12220 25660 -12100
rect 25715 -12220 25835 -12100
rect 25880 -12220 26000 -12100
rect 26045 -12220 26165 -12100
rect 26210 -12220 26330 -12100
rect 26385 -12220 26505 -12100
rect 26550 -12220 26670 -12100
rect 26715 -12220 26835 -12100
rect 26880 -12220 27000 -12100
rect 27055 -12220 27175 -12100
rect 27220 -12220 27340 -12100
rect 27385 -12220 27505 -12100
rect 27550 -12220 27670 -12100
rect 27725 -12220 27845 -12100
rect 27890 -12220 28010 -12100
rect 28055 -12220 28175 -12100
rect 28220 -12220 28340 -12100
rect 28395 -12220 28515 -12100
rect 28560 -12220 28680 -12100
rect 28725 -12220 28845 -12100
rect 28890 -12220 29010 -12100
rect 29065 -12220 29185 -12100
rect 29230 -12220 29350 -12100
rect 29395 -12220 29515 -12100
rect 29560 -12220 29680 -12100
rect 24200 -12385 24320 -12265
rect 24375 -12385 24495 -12265
rect 24540 -12385 24660 -12265
rect 24705 -12385 24825 -12265
rect 24870 -12385 24990 -12265
rect 25045 -12385 25165 -12265
rect 25210 -12385 25330 -12265
rect 25375 -12385 25495 -12265
rect 25540 -12385 25660 -12265
rect 25715 -12385 25835 -12265
rect 25880 -12385 26000 -12265
rect 26045 -12385 26165 -12265
rect 26210 -12385 26330 -12265
rect 26385 -12385 26505 -12265
rect 26550 -12385 26670 -12265
rect 26715 -12385 26835 -12265
rect 26880 -12385 27000 -12265
rect 27055 -12385 27175 -12265
rect 27220 -12385 27340 -12265
rect 27385 -12385 27505 -12265
rect 27550 -12385 27670 -12265
rect 27725 -12385 27845 -12265
rect 27890 -12385 28010 -12265
rect 28055 -12385 28175 -12265
rect 28220 -12385 28340 -12265
rect 28395 -12385 28515 -12265
rect 28560 -12385 28680 -12265
rect 28725 -12385 28845 -12265
rect 28890 -12385 29010 -12265
rect 29065 -12385 29185 -12265
rect 29230 -12385 29350 -12265
rect 29395 -12385 29515 -12265
rect 29560 -12385 29680 -12265
rect 24200 -12550 24320 -12430
rect 24375 -12550 24495 -12430
rect 24540 -12550 24660 -12430
rect 24705 -12550 24825 -12430
rect 24870 -12550 24990 -12430
rect 25045 -12550 25165 -12430
rect 25210 -12550 25330 -12430
rect 25375 -12550 25495 -12430
rect 25540 -12550 25660 -12430
rect 25715 -12550 25835 -12430
rect 25880 -12550 26000 -12430
rect 26045 -12550 26165 -12430
rect 26210 -12550 26330 -12430
rect 26385 -12550 26505 -12430
rect 26550 -12550 26670 -12430
rect 26715 -12550 26835 -12430
rect 26880 -12550 27000 -12430
rect 27055 -12550 27175 -12430
rect 27220 -12550 27340 -12430
rect 27385 -12550 27505 -12430
rect 27550 -12550 27670 -12430
rect 27725 -12550 27845 -12430
rect 27890 -12550 28010 -12430
rect 28055 -12550 28175 -12430
rect 28220 -12550 28340 -12430
rect 28395 -12550 28515 -12430
rect 28560 -12550 28680 -12430
rect 28725 -12550 28845 -12430
rect 28890 -12550 29010 -12430
rect 29065 -12550 29185 -12430
rect 29230 -12550 29350 -12430
rect 29395 -12550 29515 -12430
rect 29560 -12550 29680 -12430
rect 24200 -12715 24320 -12595
rect 24375 -12715 24495 -12595
rect 24540 -12715 24660 -12595
rect 24705 -12715 24825 -12595
rect 24870 -12715 24990 -12595
rect 25045 -12715 25165 -12595
rect 25210 -12715 25330 -12595
rect 25375 -12715 25495 -12595
rect 25540 -12715 25660 -12595
rect 25715 -12715 25835 -12595
rect 25880 -12715 26000 -12595
rect 26045 -12715 26165 -12595
rect 26210 -12715 26330 -12595
rect 26385 -12715 26505 -12595
rect 26550 -12715 26670 -12595
rect 26715 -12715 26835 -12595
rect 26880 -12715 27000 -12595
rect 27055 -12715 27175 -12595
rect 27220 -12715 27340 -12595
rect 27385 -12715 27505 -12595
rect 27550 -12715 27670 -12595
rect 27725 -12715 27845 -12595
rect 27890 -12715 28010 -12595
rect 28055 -12715 28175 -12595
rect 28220 -12715 28340 -12595
rect 28395 -12715 28515 -12595
rect 28560 -12715 28680 -12595
rect 28725 -12715 28845 -12595
rect 28890 -12715 29010 -12595
rect 29065 -12715 29185 -12595
rect 29230 -12715 29350 -12595
rect 29395 -12715 29515 -12595
rect 29560 -12715 29680 -12595
rect 24200 -12890 24320 -12770
rect 24375 -12890 24495 -12770
rect 24540 -12890 24660 -12770
rect 24705 -12890 24825 -12770
rect 24870 -12890 24990 -12770
rect 25045 -12890 25165 -12770
rect 25210 -12890 25330 -12770
rect 25375 -12890 25495 -12770
rect 25540 -12890 25660 -12770
rect 25715 -12890 25835 -12770
rect 25880 -12890 26000 -12770
rect 26045 -12890 26165 -12770
rect 26210 -12890 26330 -12770
rect 26385 -12890 26505 -12770
rect 26550 -12890 26670 -12770
rect 26715 -12890 26835 -12770
rect 26880 -12890 27000 -12770
rect 27055 -12890 27175 -12770
rect 27220 -12890 27340 -12770
rect 27385 -12890 27505 -12770
rect 27550 -12890 27670 -12770
rect 27725 -12890 27845 -12770
rect 27890 -12890 28010 -12770
rect 28055 -12890 28175 -12770
rect 28220 -12890 28340 -12770
rect 28395 -12890 28515 -12770
rect 28560 -12890 28680 -12770
rect 28725 -12890 28845 -12770
rect 28890 -12890 29010 -12770
rect 29065 -12890 29185 -12770
rect 29230 -12890 29350 -12770
rect 29395 -12890 29515 -12770
rect 29560 -12890 29680 -12770
rect 24200 -13055 24320 -12935
rect 24375 -13055 24495 -12935
rect 24540 -13055 24660 -12935
rect 24705 -13055 24825 -12935
rect 24870 -13055 24990 -12935
rect 25045 -13055 25165 -12935
rect 25210 -13055 25330 -12935
rect 25375 -13055 25495 -12935
rect 25540 -13055 25660 -12935
rect 25715 -13055 25835 -12935
rect 25880 -13055 26000 -12935
rect 26045 -13055 26165 -12935
rect 26210 -13055 26330 -12935
rect 26385 -13055 26505 -12935
rect 26550 -13055 26670 -12935
rect 26715 -13055 26835 -12935
rect 26880 -13055 27000 -12935
rect 27055 -13055 27175 -12935
rect 27220 -13055 27340 -12935
rect 27385 -13055 27505 -12935
rect 27550 -13055 27670 -12935
rect 27725 -13055 27845 -12935
rect 27890 -13055 28010 -12935
rect 28055 -13055 28175 -12935
rect 28220 -13055 28340 -12935
rect 28395 -13055 28515 -12935
rect 28560 -13055 28680 -12935
rect 28725 -13055 28845 -12935
rect 28890 -13055 29010 -12935
rect 29065 -13055 29185 -12935
rect 29230 -13055 29350 -12935
rect 29395 -13055 29515 -12935
rect 29560 -13055 29680 -12935
rect 24200 -13220 24320 -13100
rect 24375 -13220 24495 -13100
rect 24540 -13220 24660 -13100
rect 24705 -13220 24825 -13100
rect 24870 -13220 24990 -13100
rect 25045 -13220 25165 -13100
rect 25210 -13220 25330 -13100
rect 25375 -13220 25495 -13100
rect 25540 -13220 25660 -13100
rect 25715 -13220 25835 -13100
rect 25880 -13220 26000 -13100
rect 26045 -13220 26165 -13100
rect 26210 -13220 26330 -13100
rect 26385 -13220 26505 -13100
rect 26550 -13220 26670 -13100
rect 26715 -13220 26835 -13100
rect 26880 -13220 27000 -13100
rect 27055 -13220 27175 -13100
rect 27220 -13220 27340 -13100
rect 27385 -13220 27505 -13100
rect 27550 -13220 27670 -13100
rect 27725 -13220 27845 -13100
rect 27890 -13220 28010 -13100
rect 28055 -13220 28175 -13100
rect 28220 -13220 28340 -13100
rect 28395 -13220 28515 -13100
rect 28560 -13220 28680 -13100
rect 28725 -13220 28845 -13100
rect 28890 -13220 29010 -13100
rect 29065 -13220 29185 -13100
rect 29230 -13220 29350 -13100
rect 29395 -13220 29515 -13100
rect 29560 -13220 29680 -13100
rect 24200 -13385 24320 -13265
rect 24375 -13385 24495 -13265
rect 24540 -13385 24660 -13265
rect 24705 -13385 24825 -13265
rect 24870 -13385 24990 -13265
rect 25045 -13385 25165 -13265
rect 25210 -13385 25330 -13265
rect 25375 -13385 25495 -13265
rect 25540 -13385 25660 -13265
rect 25715 -13385 25835 -13265
rect 25880 -13385 26000 -13265
rect 26045 -13385 26165 -13265
rect 26210 -13385 26330 -13265
rect 26385 -13385 26505 -13265
rect 26550 -13385 26670 -13265
rect 26715 -13385 26835 -13265
rect 26880 -13385 27000 -13265
rect 27055 -13385 27175 -13265
rect 27220 -13385 27340 -13265
rect 27385 -13385 27505 -13265
rect 27550 -13385 27670 -13265
rect 27725 -13385 27845 -13265
rect 27890 -13385 28010 -13265
rect 28055 -13385 28175 -13265
rect 28220 -13385 28340 -13265
rect 28395 -13385 28515 -13265
rect 28560 -13385 28680 -13265
rect 28725 -13385 28845 -13265
rect 28890 -13385 29010 -13265
rect 29065 -13385 29185 -13265
rect 29230 -13385 29350 -13265
rect 29395 -13385 29515 -13265
rect 29560 -13385 29680 -13265
rect 24200 -13560 24320 -13440
rect 24375 -13560 24495 -13440
rect 24540 -13560 24660 -13440
rect 24705 -13560 24825 -13440
rect 24870 -13560 24990 -13440
rect 25045 -13560 25165 -13440
rect 25210 -13560 25330 -13440
rect 25375 -13560 25495 -13440
rect 25540 -13560 25660 -13440
rect 25715 -13560 25835 -13440
rect 25880 -13560 26000 -13440
rect 26045 -13560 26165 -13440
rect 26210 -13560 26330 -13440
rect 26385 -13560 26505 -13440
rect 26550 -13560 26670 -13440
rect 26715 -13560 26835 -13440
rect 26880 -13560 27000 -13440
rect 27055 -13560 27175 -13440
rect 27220 -13560 27340 -13440
rect 27385 -13560 27505 -13440
rect 27550 -13560 27670 -13440
rect 27725 -13560 27845 -13440
rect 27890 -13560 28010 -13440
rect 28055 -13560 28175 -13440
rect 28220 -13560 28340 -13440
rect 28395 -13560 28515 -13440
rect 28560 -13560 28680 -13440
rect 28725 -13560 28845 -13440
rect 28890 -13560 29010 -13440
rect 29065 -13560 29185 -13440
rect 29230 -13560 29350 -13440
rect 29395 -13560 29515 -13440
rect 29560 -13560 29680 -13440
rect 24200 -13725 24320 -13605
rect 24375 -13725 24495 -13605
rect 24540 -13725 24660 -13605
rect 24705 -13725 24825 -13605
rect 24870 -13725 24990 -13605
rect 25045 -13725 25165 -13605
rect 25210 -13725 25330 -13605
rect 25375 -13725 25495 -13605
rect 25540 -13725 25660 -13605
rect 25715 -13725 25835 -13605
rect 25880 -13725 26000 -13605
rect 26045 -13725 26165 -13605
rect 26210 -13725 26330 -13605
rect 26385 -13725 26505 -13605
rect 26550 -13725 26670 -13605
rect 26715 -13725 26835 -13605
rect 26880 -13725 27000 -13605
rect 27055 -13725 27175 -13605
rect 27220 -13725 27340 -13605
rect 27385 -13725 27505 -13605
rect 27550 -13725 27670 -13605
rect 27725 -13725 27845 -13605
rect 27890 -13725 28010 -13605
rect 28055 -13725 28175 -13605
rect 28220 -13725 28340 -13605
rect 28395 -13725 28515 -13605
rect 28560 -13725 28680 -13605
rect 28725 -13725 28845 -13605
rect 28890 -13725 29010 -13605
rect 29065 -13725 29185 -13605
rect 29230 -13725 29350 -13605
rect 29395 -13725 29515 -13605
rect 29560 -13725 29680 -13605
rect 24200 -13890 24320 -13770
rect 24375 -13890 24495 -13770
rect 24540 -13890 24660 -13770
rect 24705 -13890 24825 -13770
rect 24870 -13890 24990 -13770
rect 25045 -13890 25165 -13770
rect 25210 -13890 25330 -13770
rect 25375 -13890 25495 -13770
rect 25540 -13890 25660 -13770
rect 25715 -13890 25835 -13770
rect 25880 -13890 26000 -13770
rect 26045 -13890 26165 -13770
rect 26210 -13890 26330 -13770
rect 26385 -13890 26505 -13770
rect 26550 -13890 26670 -13770
rect 26715 -13890 26835 -13770
rect 26880 -13890 27000 -13770
rect 27055 -13890 27175 -13770
rect 27220 -13890 27340 -13770
rect 27385 -13890 27505 -13770
rect 27550 -13890 27670 -13770
rect 27725 -13890 27845 -13770
rect 27890 -13890 28010 -13770
rect 28055 -13890 28175 -13770
rect 28220 -13890 28340 -13770
rect 28395 -13890 28515 -13770
rect 28560 -13890 28680 -13770
rect 28725 -13890 28845 -13770
rect 28890 -13890 29010 -13770
rect 29065 -13890 29185 -13770
rect 29230 -13890 29350 -13770
rect 29395 -13890 29515 -13770
rect 29560 -13890 29680 -13770
rect 24200 -14055 24320 -13935
rect 24375 -14055 24495 -13935
rect 24540 -14055 24660 -13935
rect 24705 -14055 24825 -13935
rect 24870 -14055 24990 -13935
rect 25045 -14055 25165 -13935
rect 25210 -14055 25330 -13935
rect 25375 -14055 25495 -13935
rect 25540 -14055 25660 -13935
rect 25715 -14055 25835 -13935
rect 25880 -14055 26000 -13935
rect 26045 -14055 26165 -13935
rect 26210 -14055 26330 -13935
rect 26385 -14055 26505 -13935
rect 26550 -14055 26670 -13935
rect 26715 -14055 26835 -13935
rect 26880 -14055 27000 -13935
rect 27055 -14055 27175 -13935
rect 27220 -14055 27340 -13935
rect 27385 -14055 27505 -13935
rect 27550 -14055 27670 -13935
rect 27725 -14055 27845 -13935
rect 27890 -14055 28010 -13935
rect 28055 -14055 28175 -13935
rect 28220 -14055 28340 -13935
rect 28395 -14055 28515 -13935
rect 28560 -14055 28680 -13935
rect 28725 -14055 28845 -13935
rect 28890 -14055 29010 -13935
rect 29065 -14055 29185 -13935
rect 29230 -14055 29350 -13935
rect 29395 -14055 29515 -13935
rect 29560 -14055 29680 -13935
rect 24200 -14230 24320 -14110
rect 24375 -14230 24495 -14110
rect 24540 -14230 24660 -14110
rect 24705 -14230 24825 -14110
rect 24870 -14230 24990 -14110
rect 25045 -14230 25165 -14110
rect 25210 -14230 25330 -14110
rect 25375 -14230 25495 -14110
rect 25540 -14230 25660 -14110
rect 25715 -14230 25835 -14110
rect 25880 -14230 26000 -14110
rect 26045 -14230 26165 -14110
rect 26210 -14230 26330 -14110
rect 26385 -14230 26505 -14110
rect 26550 -14230 26670 -14110
rect 26715 -14230 26835 -14110
rect 26880 -14230 27000 -14110
rect 27055 -14230 27175 -14110
rect 27220 -14230 27340 -14110
rect 27385 -14230 27505 -14110
rect 27550 -14230 27670 -14110
rect 27725 -14230 27845 -14110
rect 27890 -14230 28010 -14110
rect 28055 -14230 28175 -14110
rect 28220 -14230 28340 -14110
rect 28395 -14230 28515 -14110
rect 28560 -14230 28680 -14110
rect 28725 -14230 28845 -14110
rect 28890 -14230 29010 -14110
rect 29065 -14230 29185 -14110
rect 29230 -14230 29350 -14110
rect 29395 -14230 29515 -14110
rect 29560 -14230 29680 -14110
rect 24200 -14395 24320 -14275
rect 24375 -14395 24495 -14275
rect 24540 -14395 24660 -14275
rect 24705 -14395 24825 -14275
rect 24870 -14395 24990 -14275
rect 25045 -14395 25165 -14275
rect 25210 -14395 25330 -14275
rect 25375 -14395 25495 -14275
rect 25540 -14395 25660 -14275
rect 25715 -14395 25835 -14275
rect 25880 -14395 26000 -14275
rect 26045 -14395 26165 -14275
rect 26210 -14395 26330 -14275
rect 26385 -14395 26505 -14275
rect 26550 -14395 26670 -14275
rect 26715 -14395 26835 -14275
rect 26880 -14395 27000 -14275
rect 27055 -14395 27175 -14275
rect 27220 -14395 27340 -14275
rect 27385 -14395 27505 -14275
rect 27550 -14395 27670 -14275
rect 27725 -14395 27845 -14275
rect 27890 -14395 28010 -14275
rect 28055 -14395 28175 -14275
rect 28220 -14395 28340 -14275
rect 28395 -14395 28515 -14275
rect 28560 -14395 28680 -14275
rect 28725 -14395 28845 -14275
rect 28890 -14395 29010 -14275
rect 29065 -14395 29185 -14275
rect 29230 -14395 29350 -14275
rect 29395 -14395 29515 -14275
rect 29560 -14395 29680 -14275
rect 24200 -14560 24320 -14440
rect 24375 -14560 24495 -14440
rect 24540 -14560 24660 -14440
rect 24705 -14560 24825 -14440
rect 24870 -14560 24990 -14440
rect 25045 -14560 25165 -14440
rect 25210 -14560 25330 -14440
rect 25375 -14560 25495 -14440
rect 25540 -14560 25660 -14440
rect 25715 -14560 25835 -14440
rect 25880 -14560 26000 -14440
rect 26045 -14560 26165 -14440
rect 26210 -14560 26330 -14440
rect 26385 -14560 26505 -14440
rect 26550 -14560 26670 -14440
rect 26715 -14560 26835 -14440
rect 26880 -14560 27000 -14440
rect 27055 -14560 27175 -14440
rect 27220 -14560 27340 -14440
rect 27385 -14560 27505 -14440
rect 27550 -14560 27670 -14440
rect 27725 -14560 27845 -14440
rect 27890 -14560 28010 -14440
rect 28055 -14560 28175 -14440
rect 28220 -14560 28340 -14440
rect 28395 -14560 28515 -14440
rect 28560 -14560 28680 -14440
rect 28725 -14560 28845 -14440
rect 28890 -14560 29010 -14440
rect 29065 -14560 29185 -14440
rect 29230 -14560 29350 -14440
rect 29395 -14560 29515 -14440
rect 29560 -14560 29680 -14440
rect 24200 -14725 24320 -14605
rect 24375 -14725 24495 -14605
rect 24540 -14725 24660 -14605
rect 24705 -14725 24825 -14605
rect 24870 -14725 24990 -14605
rect 25045 -14725 25165 -14605
rect 25210 -14725 25330 -14605
rect 25375 -14725 25495 -14605
rect 25540 -14725 25660 -14605
rect 25715 -14725 25835 -14605
rect 25880 -14725 26000 -14605
rect 26045 -14725 26165 -14605
rect 26210 -14725 26330 -14605
rect 26385 -14725 26505 -14605
rect 26550 -14725 26670 -14605
rect 26715 -14725 26835 -14605
rect 26880 -14725 27000 -14605
rect 27055 -14725 27175 -14605
rect 27220 -14725 27340 -14605
rect 27385 -14725 27505 -14605
rect 27550 -14725 27670 -14605
rect 27725 -14725 27845 -14605
rect 27890 -14725 28010 -14605
rect 28055 -14725 28175 -14605
rect 28220 -14725 28340 -14605
rect 28395 -14725 28515 -14605
rect 28560 -14725 28680 -14605
rect 28725 -14725 28845 -14605
rect 28890 -14725 29010 -14605
rect 29065 -14725 29185 -14605
rect 29230 -14725 29350 -14605
rect 29395 -14725 29515 -14605
rect 29560 -14725 29680 -14605
rect 24200 -14900 24320 -14780
rect 24375 -14900 24495 -14780
rect 24540 -14900 24660 -14780
rect 24705 -14900 24825 -14780
rect 24870 -14900 24990 -14780
rect 25045 -14900 25165 -14780
rect 25210 -14900 25330 -14780
rect 25375 -14900 25495 -14780
rect 25540 -14900 25660 -14780
rect 25715 -14900 25835 -14780
rect 25880 -14900 26000 -14780
rect 26045 -14900 26165 -14780
rect 26210 -14900 26330 -14780
rect 26385 -14900 26505 -14780
rect 26550 -14900 26670 -14780
rect 26715 -14900 26835 -14780
rect 26880 -14900 27000 -14780
rect 27055 -14900 27175 -14780
rect 27220 -14900 27340 -14780
rect 27385 -14900 27505 -14780
rect 27550 -14900 27670 -14780
rect 27725 -14900 27845 -14780
rect 27890 -14900 28010 -14780
rect 28055 -14900 28175 -14780
rect 28220 -14900 28340 -14780
rect 28395 -14900 28515 -14780
rect 28560 -14900 28680 -14780
rect 28725 -14900 28845 -14780
rect 28890 -14900 29010 -14780
rect 29065 -14900 29185 -14780
rect 29230 -14900 29350 -14780
rect 29395 -14900 29515 -14780
rect 29560 -14900 29680 -14780
rect 24200 -15065 24320 -14945
rect 24375 -15065 24495 -14945
rect 24540 -15065 24660 -14945
rect 24705 -15065 24825 -14945
rect 24870 -15065 24990 -14945
rect 25045 -15065 25165 -14945
rect 25210 -15065 25330 -14945
rect 25375 -15065 25495 -14945
rect 25540 -15065 25660 -14945
rect 25715 -15065 25835 -14945
rect 25880 -15065 26000 -14945
rect 26045 -15065 26165 -14945
rect 26210 -15065 26330 -14945
rect 26385 -15065 26505 -14945
rect 26550 -15065 26670 -14945
rect 26715 -15065 26835 -14945
rect 26880 -15065 27000 -14945
rect 27055 -15065 27175 -14945
rect 27220 -15065 27340 -14945
rect 27385 -15065 27505 -14945
rect 27550 -15065 27670 -14945
rect 27725 -15065 27845 -14945
rect 27890 -15065 28010 -14945
rect 28055 -15065 28175 -14945
rect 28220 -15065 28340 -14945
rect 28395 -15065 28515 -14945
rect 28560 -15065 28680 -14945
rect 28725 -15065 28845 -14945
rect 28890 -15065 29010 -14945
rect 29065 -15065 29185 -14945
rect 29230 -15065 29350 -14945
rect 29395 -15065 29515 -14945
rect 29560 -15065 29680 -14945
rect 24200 -15230 24320 -15110
rect 24375 -15230 24495 -15110
rect 24540 -15230 24660 -15110
rect 24705 -15230 24825 -15110
rect 24870 -15230 24990 -15110
rect 25045 -15230 25165 -15110
rect 25210 -15230 25330 -15110
rect 25375 -15230 25495 -15110
rect 25540 -15230 25660 -15110
rect 25715 -15230 25835 -15110
rect 25880 -15230 26000 -15110
rect 26045 -15230 26165 -15110
rect 26210 -15230 26330 -15110
rect 26385 -15230 26505 -15110
rect 26550 -15230 26670 -15110
rect 26715 -15230 26835 -15110
rect 26880 -15230 27000 -15110
rect 27055 -15230 27175 -15110
rect 27220 -15230 27340 -15110
rect 27385 -15230 27505 -15110
rect 27550 -15230 27670 -15110
rect 27725 -15230 27845 -15110
rect 27890 -15230 28010 -15110
rect 28055 -15230 28175 -15110
rect 28220 -15230 28340 -15110
rect 28395 -15230 28515 -15110
rect 28560 -15230 28680 -15110
rect 28725 -15230 28845 -15110
rect 28890 -15230 29010 -15110
rect 29065 -15230 29185 -15110
rect 29230 -15230 29350 -15110
rect 29395 -15230 29515 -15110
rect 29560 -15230 29680 -15110
rect 24200 -15395 24320 -15275
rect 24375 -15395 24495 -15275
rect 24540 -15395 24660 -15275
rect 24705 -15395 24825 -15275
rect 24870 -15395 24990 -15275
rect 25045 -15395 25165 -15275
rect 25210 -15395 25330 -15275
rect 25375 -15395 25495 -15275
rect 25540 -15395 25660 -15275
rect 25715 -15395 25835 -15275
rect 25880 -15395 26000 -15275
rect 26045 -15395 26165 -15275
rect 26210 -15395 26330 -15275
rect 26385 -15395 26505 -15275
rect 26550 -15395 26670 -15275
rect 26715 -15395 26835 -15275
rect 26880 -15395 27000 -15275
rect 27055 -15395 27175 -15275
rect 27220 -15395 27340 -15275
rect 27385 -15395 27505 -15275
rect 27550 -15395 27670 -15275
rect 27725 -15395 27845 -15275
rect 27890 -15395 28010 -15275
rect 28055 -15395 28175 -15275
rect 28220 -15395 28340 -15275
rect 28395 -15395 28515 -15275
rect 28560 -15395 28680 -15275
rect 28725 -15395 28845 -15275
rect 28890 -15395 29010 -15275
rect 29065 -15395 29185 -15275
rect 29230 -15395 29350 -15275
rect 29395 -15395 29515 -15275
rect 29560 -15395 29680 -15275
rect 24200 -15570 24320 -15450
rect 24375 -15570 24495 -15450
rect 24540 -15570 24660 -15450
rect 24705 -15570 24825 -15450
rect 24870 -15570 24990 -15450
rect 25045 -15570 25165 -15450
rect 25210 -15570 25330 -15450
rect 25375 -15570 25495 -15450
rect 25540 -15570 25660 -15450
rect 25715 -15570 25835 -15450
rect 25880 -15570 26000 -15450
rect 26045 -15570 26165 -15450
rect 26210 -15570 26330 -15450
rect 26385 -15570 26505 -15450
rect 26550 -15570 26670 -15450
rect 26715 -15570 26835 -15450
rect 26880 -15570 27000 -15450
rect 27055 -15570 27175 -15450
rect 27220 -15570 27340 -15450
rect 27385 -15570 27505 -15450
rect 27550 -15570 27670 -15450
rect 27725 -15570 27845 -15450
rect 27890 -15570 28010 -15450
rect 28055 -15570 28175 -15450
rect 28220 -15570 28340 -15450
rect 28395 -15570 28515 -15450
rect 28560 -15570 28680 -15450
rect 28725 -15570 28845 -15450
rect 28890 -15570 29010 -15450
rect 29065 -15570 29185 -15450
rect 29230 -15570 29350 -15450
rect 29395 -15570 29515 -15450
rect 29560 -15570 29680 -15450
<< metal4 >>
rect 7105 7160 29705 7185
rect 7105 7040 7130 7160
rect 7250 7040 7295 7160
rect 7415 7040 7460 7160
rect 7580 7040 7625 7160
rect 7745 7040 7800 7160
rect 7920 7040 7965 7160
rect 8085 7040 8130 7160
rect 8250 7040 8295 7160
rect 8415 7040 8470 7160
rect 8590 7040 8635 7160
rect 8755 7040 8800 7160
rect 8920 7040 8965 7160
rect 9085 7040 9140 7160
rect 9260 7040 9305 7160
rect 9425 7040 9470 7160
rect 9590 7040 9635 7160
rect 9755 7040 9810 7160
rect 9930 7040 9975 7160
rect 10095 7040 10140 7160
rect 10260 7040 10305 7160
rect 10425 7040 10480 7160
rect 10600 7040 10645 7160
rect 10765 7040 10810 7160
rect 10930 7040 10975 7160
rect 11095 7040 11150 7160
rect 11270 7040 11315 7160
rect 11435 7040 11480 7160
rect 11600 7040 11645 7160
rect 11765 7040 11820 7160
rect 11940 7040 11985 7160
rect 12105 7040 12150 7160
rect 12270 7040 12315 7160
rect 12435 7040 12490 7160
rect 12610 7125 12820 7160
rect 12610 7040 12635 7125
rect 7105 6985 12635 7040
rect 7105 6865 7130 6985
rect 7250 6865 7295 6985
rect 7415 6865 7460 6985
rect 7580 6865 7625 6985
rect 7745 6865 7800 6985
rect 7920 6865 7965 6985
rect 8085 6865 8130 6985
rect 8250 6865 8295 6985
rect 8415 6865 8470 6985
rect 8590 6865 8635 6985
rect 8755 6865 8800 6985
rect 8920 6865 8965 6985
rect 9085 6865 9140 6985
rect 9260 6865 9305 6985
rect 9425 6865 9470 6985
rect 9590 6865 9635 6985
rect 9755 6865 9810 6985
rect 9930 6865 9975 6985
rect 10095 6865 10140 6985
rect 10260 6865 10305 6985
rect 10425 6865 10480 6985
rect 10600 6865 10645 6985
rect 10765 6865 10810 6985
rect 10930 6865 10975 6985
rect 11095 6865 11150 6985
rect 11270 6865 11315 6985
rect 11435 6865 11480 6985
rect 11600 6865 11645 6985
rect 11765 6865 11820 6985
rect 11940 6865 11985 6985
rect 12105 6865 12150 6985
rect 12270 6865 12315 6985
rect 12435 6865 12490 6985
rect 12610 6865 12635 6985
rect 7105 6820 12635 6865
rect 7105 6700 7130 6820
rect 7250 6700 7295 6820
rect 7415 6700 7460 6820
rect 7580 6700 7625 6820
rect 7745 6700 7800 6820
rect 7920 6700 7965 6820
rect 8085 6700 8130 6820
rect 8250 6700 8295 6820
rect 8415 6700 8470 6820
rect 8590 6700 8635 6820
rect 8755 6700 8800 6820
rect 8920 6700 8965 6820
rect 9085 6700 9140 6820
rect 9260 6700 9305 6820
rect 9425 6700 9470 6820
rect 9590 6700 9635 6820
rect 9755 6700 9810 6820
rect 9930 6700 9975 6820
rect 10095 6700 10140 6820
rect 10260 6700 10305 6820
rect 10425 6700 10480 6820
rect 10600 6700 10645 6820
rect 10765 6700 10810 6820
rect 10930 6700 10975 6820
rect 11095 6700 11150 6820
rect 11270 6700 11315 6820
rect 11435 6700 11480 6820
rect 11600 6700 11645 6820
rect 11765 6700 11820 6820
rect 11940 6700 11985 6820
rect 12105 6700 12150 6820
rect 12270 6700 12315 6820
rect 12435 6700 12490 6820
rect 12610 6700 12635 6820
rect 7105 6655 12635 6700
rect 7105 6535 7130 6655
rect 7250 6535 7295 6655
rect 7415 6535 7460 6655
rect 7580 6535 7625 6655
rect 7745 6535 7800 6655
rect 7920 6535 7965 6655
rect 8085 6535 8130 6655
rect 8250 6535 8295 6655
rect 8415 6535 8470 6655
rect 8590 6535 8635 6655
rect 8755 6535 8800 6655
rect 8920 6535 8965 6655
rect 9085 6535 9140 6655
rect 9260 6535 9305 6655
rect 9425 6535 9470 6655
rect 9590 6535 9635 6655
rect 9755 6535 9810 6655
rect 9930 6535 9975 6655
rect 10095 6535 10140 6655
rect 10260 6535 10305 6655
rect 10425 6535 10480 6655
rect 10600 6535 10645 6655
rect 10765 6535 10810 6655
rect 10930 6535 10975 6655
rect 11095 6535 11150 6655
rect 11270 6535 11315 6655
rect 11435 6535 11480 6655
rect 11600 6535 11645 6655
rect 11765 6535 11820 6655
rect 11940 6535 11985 6655
rect 12105 6535 12150 6655
rect 12270 6535 12315 6655
rect 12435 6535 12490 6655
rect 12610 6535 12635 6655
rect 7105 6490 12635 6535
rect 7105 6370 7130 6490
rect 7250 6370 7295 6490
rect 7415 6370 7460 6490
rect 7580 6370 7625 6490
rect 7745 6370 7800 6490
rect 7920 6370 7965 6490
rect 8085 6370 8130 6490
rect 8250 6370 8295 6490
rect 8415 6370 8470 6490
rect 8590 6370 8635 6490
rect 8755 6370 8800 6490
rect 8920 6370 8965 6490
rect 9085 6370 9140 6490
rect 9260 6370 9305 6490
rect 9425 6370 9470 6490
rect 9590 6370 9635 6490
rect 9755 6370 9810 6490
rect 9930 6370 9975 6490
rect 10095 6370 10140 6490
rect 10260 6370 10305 6490
rect 10425 6370 10480 6490
rect 10600 6370 10645 6490
rect 10765 6370 10810 6490
rect 10930 6370 10975 6490
rect 11095 6370 11150 6490
rect 11270 6370 11315 6490
rect 11435 6370 11480 6490
rect 11600 6370 11645 6490
rect 11765 6370 11820 6490
rect 11940 6370 11985 6490
rect 12105 6370 12150 6490
rect 12270 6370 12315 6490
rect 12435 6370 12490 6490
rect 12610 6370 12635 6490
rect 7105 6315 12635 6370
rect 7105 6195 7130 6315
rect 7250 6195 7295 6315
rect 7415 6195 7460 6315
rect 7580 6195 7625 6315
rect 7745 6195 7800 6315
rect 7920 6195 7965 6315
rect 8085 6195 8130 6315
rect 8250 6195 8295 6315
rect 8415 6195 8470 6315
rect 8590 6195 8635 6315
rect 8755 6195 8800 6315
rect 8920 6195 8965 6315
rect 9085 6195 9140 6315
rect 9260 6195 9305 6315
rect 9425 6195 9470 6315
rect 9590 6195 9635 6315
rect 9755 6195 9810 6315
rect 9930 6195 9975 6315
rect 10095 6195 10140 6315
rect 10260 6195 10305 6315
rect 10425 6195 10480 6315
rect 10600 6195 10645 6315
rect 10765 6195 10810 6315
rect 10930 6195 10975 6315
rect 11095 6195 11150 6315
rect 11270 6195 11315 6315
rect 11435 6195 11480 6315
rect 11600 6195 11645 6315
rect 11765 6195 11820 6315
rect 11940 6195 11985 6315
rect 12105 6195 12150 6315
rect 12270 6195 12315 6315
rect 12435 6195 12490 6315
rect 12610 6195 12635 6315
rect 7105 6150 12635 6195
rect 7105 6030 7130 6150
rect 7250 6030 7295 6150
rect 7415 6030 7460 6150
rect 7580 6030 7625 6150
rect 7745 6030 7800 6150
rect 7920 6030 7965 6150
rect 8085 6030 8130 6150
rect 8250 6030 8295 6150
rect 8415 6030 8470 6150
rect 8590 6030 8635 6150
rect 8755 6030 8800 6150
rect 8920 6030 8965 6150
rect 9085 6030 9140 6150
rect 9260 6030 9305 6150
rect 9425 6030 9470 6150
rect 9590 6030 9635 6150
rect 9755 6030 9810 6150
rect 9930 6030 9975 6150
rect 10095 6030 10140 6150
rect 10260 6030 10305 6150
rect 10425 6030 10480 6150
rect 10600 6030 10645 6150
rect 10765 6030 10810 6150
rect 10930 6030 10975 6150
rect 11095 6030 11150 6150
rect 11270 6030 11315 6150
rect 11435 6030 11480 6150
rect 11600 6030 11645 6150
rect 11765 6030 11820 6150
rect 11940 6030 11985 6150
rect 12105 6030 12150 6150
rect 12270 6030 12315 6150
rect 12435 6030 12490 6150
rect 12610 6030 12635 6150
rect 7105 5985 12635 6030
rect 7105 5865 7130 5985
rect 7250 5865 7295 5985
rect 7415 5865 7460 5985
rect 7580 5865 7625 5985
rect 7745 5865 7800 5985
rect 7920 5865 7965 5985
rect 8085 5865 8130 5985
rect 8250 5865 8295 5985
rect 8415 5865 8470 5985
rect 8590 5865 8635 5985
rect 8755 5865 8800 5985
rect 8920 5865 8965 5985
rect 9085 5865 9140 5985
rect 9260 5865 9305 5985
rect 9425 5865 9470 5985
rect 9590 5865 9635 5985
rect 9755 5865 9810 5985
rect 9930 5865 9975 5985
rect 10095 5865 10140 5985
rect 10260 5865 10305 5985
rect 10425 5865 10480 5985
rect 10600 5865 10645 5985
rect 10765 5865 10810 5985
rect 10930 5865 10975 5985
rect 11095 5865 11150 5985
rect 11270 5865 11315 5985
rect 11435 5865 11480 5985
rect 11600 5865 11645 5985
rect 11765 5865 11820 5985
rect 11940 5865 11985 5985
rect 12105 5865 12150 5985
rect 12270 5865 12315 5985
rect 12435 5865 12490 5985
rect 12610 5865 12635 5985
rect 7105 5820 12635 5865
rect 7105 5700 7130 5820
rect 7250 5700 7295 5820
rect 7415 5700 7460 5820
rect 7580 5700 7625 5820
rect 7745 5700 7800 5820
rect 7920 5700 7965 5820
rect 8085 5700 8130 5820
rect 8250 5700 8295 5820
rect 8415 5700 8470 5820
rect 8590 5700 8635 5820
rect 8755 5700 8800 5820
rect 8920 5700 8965 5820
rect 9085 5700 9140 5820
rect 9260 5700 9305 5820
rect 9425 5700 9470 5820
rect 9590 5700 9635 5820
rect 9755 5700 9810 5820
rect 9930 5700 9975 5820
rect 10095 5700 10140 5820
rect 10260 5700 10305 5820
rect 10425 5700 10480 5820
rect 10600 5700 10645 5820
rect 10765 5700 10810 5820
rect 10930 5700 10975 5820
rect 11095 5700 11150 5820
rect 11270 5700 11315 5820
rect 11435 5700 11480 5820
rect 11600 5700 11645 5820
rect 11765 5700 11820 5820
rect 11940 5700 11985 5820
rect 12105 5700 12150 5820
rect 12270 5700 12315 5820
rect 12435 5700 12490 5820
rect 12610 5700 12635 5820
rect 7105 5645 12635 5700
rect 7105 5525 7130 5645
rect 7250 5525 7295 5645
rect 7415 5525 7460 5645
rect 7580 5525 7625 5645
rect 7745 5525 7800 5645
rect 7920 5525 7965 5645
rect 8085 5525 8130 5645
rect 8250 5525 8295 5645
rect 8415 5525 8470 5645
rect 8590 5525 8635 5645
rect 8755 5525 8800 5645
rect 8920 5525 8965 5645
rect 9085 5525 9140 5645
rect 9260 5525 9305 5645
rect 9425 5525 9470 5645
rect 9590 5525 9635 5645
rect 9755 5525 9810 5645
rect 9930 5525 9975 5645
rect 10095 5525 10140 5645
rect 10260 5525 10305 5645
rect 10425 5525 10480 5645
rect 10600 5525 10645 5645
rect 10765 5525 10810 5645
rect 10930 5525 10975 5645
rect 11095 5525 11150 5645
rect 11270 5525 11315 5645
rect 11435 5525 11480 5645
rect 11600 5525 11645 5645
rect 11765 5525 11820 5645
rect 11940 5525 11985 5645
rect 12105 5525 12150 5645
rect 12270 5525 12315 5645
rect 12435 5525 12490 5645
rect 12610 5525 12635 5645
rect 7105 5480 12635 5525
rect 7105 5360 7130 5480
rect 7250 5360 7295 5480
rect 7415 5360 7460 5480
rect 7580 5360 7625 5480
rect 7745 5360 7800 5480
rect 7920 5360 7965 5480
rect 8085 5360 8130 5480
rect 8250 5360 8295 5480
rect 8415 5360 8470 5480
rect 8590 5360 8635 5480
rect 8755 5360 8800 5480
rect 8920 5360 8965 5480
rect 9085 5360 9140 5480
rect 9260 5360 9305 5480
rect 9425 5360 9470 5480
rect 9590 5360 9635 5480
rect 9755 5360 9810 5480
rect 9930 5360 9975 5480
rect 10095 5360 10140 5480
rect 10260 5360 10305 5480
rect 10425 5360 10480 5480
rect 10600 5360 10645 5480
rect 10765 5360 10810 5480
rect 10930 5360 10975 5480
rect 11095 5360 11150 5480
rect 11270 5360 11315 5480
rect 11435 5360 11480 5480
rect 11600 5360 11645 5480
rect 11765 5360 11820 5480
rect 11940 5360 11985 5480
rect 12105 5360 12150 5480
rect 12270 5360 12315 5480
rect 12435 5360 12490 5480
rect 12610 5360 12635 5480
rect 7105 5315 12635 5360
rect 7105 5195 7130 5315
rect 7250 5195 7295 5315
rect 7415 5195 7460 5315
rect 7580 5195 7625 5315
rect 7745 5195 7800 5315
rect 7920 5195 7965 5315
rect 8085 5195 8130 5315
rect 8250 5195 8295 5315
rect 8415 5195 8470 5315
rect 8590 5195 8635 5315
rect 8755 5195 8800 5315
rect 8920 5195 8965 5315
rect 9085 5195 9140 5315
rect 9260 5195 9305 5315
rect 9425 5195 9470 5315
rect 9590 5195 9635 5315
rect 9755 5195 9810 5315
rect 9930 5195 9975 5315
rect 10095 5195 10140 5315
rect 10260 5195 10305 5315
rect 10425 5195 10480 5315
rect 10600 5195 10645 5315
rect 10765 5195 10810 5315
rect 10930 5195 10975 5315
rect 11095 5195 11150 5315
rect 11270 5195 11315 5315
rect 11435 5195 11480 5315
rect 11600 5195 11645 5315
rect 11765 5195 11820 5315
rect 11940 5195 11985 5315
rect 12105 5195 12150 5315
rect 12270 5195 12315 5315
rect 12435 5195 12490 5315
rect 12610 5195 12635 5315
rect 7105 5150 12635 5195
rect 7105 5030 7130 5150
rect 7250 5030 7295 5150
rect 7415 5030 7460 5150
rect 7580 5030 7625 5150
rect 7745 5030 7800 5150
rect 7920 5030 7965 5150
rect 8085 5030 8130 5150
rect 8250 5030 8295 5150
rect 8415 5030 8470 5150
rect 8590 5030 8635 5150
rect 8755 5030 8800 5150
rect 8920 5030 8965 5150
rect 9085 5030 9140 5150
rect 9260 5030 9305 5150
rect 9425 5030 9470 5150
rect 9590 5030 9635 5150
rect 9755 5030 9810 5150
rect 9930 5030 9975 5150
rect 10095 5030 10140 5150
rect 10260 5030 10305 5150
rect 10425 5030 10480 5150
rect 10600 5030 10645 5150
rect 10765 5030 10810 5150
rect 10930 5030 10975 5150
rect 11095 5030 11150 5150
rect 11270 5030 11315 5150
rect 11435 5030 11480 5150
rect 11600 5030 11645 5150
rect 11765 5030 11820 5150
rect 11940 5030 11985 5150
rect 12105 5030 12150 5150
rect 12270 5030 12315 5150
rect 12435 5030 12490 5150
rect 12610 5030 12635 5150
rect 7105 4975 12635 5030
rect 7105 4855 7130 4975
rect 7250 4855 7295 4975
rect 7415 4855 7460 4975
rect 7580 4855 7625 4975
rect 7745 4855 7800 4975
rect 7920 4855 7965 4975
rect 8085 4855 8130 4975
rect 8250 4855 8295 4975
rect 8415 4855 8470 4975
rect 8590 4855 8635 4975
rect 8755 4855 8800 4975
rect 8920 4855 8965 4975
rect 9085 4855 9140 4975
rect 9260 4855 9305 4975
rect 9425 4855 9470 4975
rect 9590 4855 9635 4975
rect 9755 4855 9810 4975
rect 9930 4855 9975 4975
rect 10095 4855 10140 4975
rect 10260 4855 10305 4975
rect 10425 4855 10480 4975
rect 10600 4855 10645 4975
rect 10765 4855 10810 4975
rect 10930 4855 10975 4975
rect 11095 4855 11150 4975
rect 11270 4855 11315 4975
rect 11435 4855 11480 4975
rect 11600 4855 11645 4975
rect 11765 4855 11820 4975
rect 11940 4855 11985 4975
rect 12105 4855 12150 4975
rect 12270 4855 12315 4975
rect 12435 4855 12490 4975
rect 12610 4855 12635 4975
rect 7105 4810 12635 4855
rect 7105 4690 7130 4810
rect 7250 4690 7295 4810
rect 7415 4690 7460 4810
rect 7580 4690 7625 4810
rect 7745 4690 7800 4810
rect 7920 4690 7965 4810
rect 8085 4690 8130 4810
rect 8250 4690 8295 4810
rect 8415 4690 8470 4810
rect 8590 4690 8635 4810
rect 8755 4690 8800 4810
rect 8920 4690 8965 4810
rect 9085 4690 9140 4810
rect 9260 4690 9305 4810
rect 9425 4690 9470 4810
rect 9590 4690 9635 4810
rect 9755 4690 9810 4810
rect 9930 4690 9975 4810
rect 10095 4690 10140 4810
rect 10260 4690 10305 4810
rect 10425 4690 10480 4810
rect 10600 4690 10645 4810
rect 10765 4690 10810 4810
rect 10930 4690 10975 4810
rect 11095 4690 11150 4810
rect 11270 4690 11315 4810
rect 11435 4690 11480 4810
rect 11600 4690 11645 4810
rect 11765 4690 11820 4810
rect 11940 4690 11985 4810
rect 12105 4690 12150 4810
rect 12270 4690 12315 4810
rect 12435 4690 12490 4810
rect 12610 4690 12635 4810
rect 7105 4645 12635 4690
rect 7105 4525 7130 4645
rect 7250 4525 7295 4645
rect 7415 4525 7460 4645
rect 7580 4525 7625 4645
rect 7745 4525 7800 4645
rect 7920 4525 7965 4645
rect 8085 4525 8130 4645
rect 8250 4525 8295 4645
rect 8415 4525 8470 4645
rect 8590 4525 8635 4645
rect 8755 4525 8800 4645
rect 8920 4525 8965 4645
rect 9085 4525 9140 4645
rect 9260 4525 9305 4645
rect 9425 4525 9470 4645
rect 9590 4525 9635 4645
rect 9755 4525 9810 4645
rect 9930 4525 9975 4645
rect 10095 4525 10140 4645
rect 10260 4525 10305 4645
rect 10425 4525 10480 4645
rect 10600 4525 10645 4645
rect 10765 4525 10810 4645
rect 10930 4525 10975 4645
rect 11095 4525 11150 4645
rect 11270 4525 11315 4645
rect 11435 4525 11480 4645
rect 11600 4525 11645 4645
rect 11765 4525 11820 4645
rect 11940 4525 11985 4645
rect 12105 4525 12150 4645
rect 12270 4525 12315 4645
rect 12435 4525 12490 4645
rect 12610 4525 12635 4645
rect 7105 4480 12635 4525
rect 7105 4360 7130 4480
rect 7250 4360 7295 4480
rect 7415 4360 7460 4480
rect 7580 4360 7625 4480
rect 7745 4360 7800 4480
rect 7920 4360 7965 4480
rect 8085 4360 8130 4480
rect 8250 4360 8295 4480
rect 8415 4360 8470 4480
rect 8590 4360 8635 4480
rect 8755 4360 8800 4480
rect 8920 4360 8965 4480
rect 9085 4360 9140 4480
rect 9260 4360 9305 4480
rect 9425 4360 9470 4480
rect 9590 4360 9635 4480
rect 9755 4360 9810 4480
rect 9930 4360 9975 4480
rect 10095 4360 10140 4480
rect 10260 4360 10305 4480
rect 10425 4360 10480 4480
rect 10600 4360 10645 4480
rect 10765 4360 10810 4480
rect 10930 4360 10975 4480
rect 11095 4360 11150 4480
rect 11270 4360 11315 4480
rect 11435 4360 11480 4480
rect 11600 4360 11645 4480
rect 11765 4360 11820 4480
rect 11940 4360 11985 4480
rect 12105 4360 12150 4480
rect 12270 4360 12315 4480
rect 12435 4360 12490 4480
rect 12610 4360 12635 4480
rect 7105 4305 12635 4360
rect 7105 4185 7130 4305
rect 7250 4185 7295 4305
rect 7415 4185 7460 4305
rect 7580 4185 7625 4305
rect 7745 4185 7800 4305
rect 7920 4185 7965 4305
rect 8085 4185 8130 4305
rect 8250 4185 8295 4305
rect 8415 4185 8470 4305
rect 8590 4185 8635 4305
rect 8755 4185 8800 4305
rect 8920 4185 8965 4305
rect 9085 4185 9140 4305
rect 9260 4185 9305 4305
rect 9425 4185 9470 4305
rect 9590 4185 9635 4305
rect 9755 4185 9810 4305
rect 9930 4185 9975 4305
rect 10095 4185 10140 4305
rect 10260 4185 10305 4305
rect 10425 4185 10480 4305
rect 10600 4185 10645 4305
rect 10765 4185 10810 4305
rect 10930 4185 10975 4305
rect 11095 4185 11150 4305
rect 11270 4185 11315 4305
rect 11435 4185 11480 4305
rect 11600 4185 11645 4305
rect 11765 4185 11820 4305
rect 11940 4185 11985 4305
rect 12105 4185 12150 4305
rect 12270 4185 12315 4305
rect 12435 4185 12490 4305
rect 12610 4185 12635 4305
rect 7105 4140 12635 4185
rect 7105 4020 7130 4140
rect 7250 4020 7295 4140
rect 7415 4020 7460 4140
rect 7580 4020 7625 4140
rect 7745 4020 7800 4140
rect 7920 4020 7965 4140
rect 8085 4020 8130 4140
rect 8250 4020 8295 4140
rect 8415 4020 8470 4140
rect 8590 4020 8635 4140
rect 8755 4020 8800 4140
rect 8920 4020 8965 4140
rect 9085 4020 9140 4140
rect 9260 4020 9305 4140
rect 9425 4020 9470 4140
rect 9590 4020 9635 4140
rect 9755 4020 9810 4140
rect 9930 4020 9975 4140
rect 10095 4020 10140 4140
rect 10260 4020 10305 4140
rect 10425 4020 10480 4140
rect 10600 4020 10645 4140
rect 10765 4020 10810 4140
rect 10930 4020 10975 4140
rect 11095 4020 11150 4140
rect 11270 4020 11315 4140
rect 11435 4020 11480 4140
rect 11600 4020 11645 4140
rect 11765 4020 11820 4140
rect 11940 4020 11985 4140
rect 12105 4020 12150 4140
rect 12270 4020 12315 4140
rect 12435 4020 12490 4140
rect 12610 4020 12635 4140
rect 7105 3975 12635 4020
rect 7105 3855 7130 3975
rect 7250 3855 7295 3975
rect 7415 3855 7460 3975
rect 7580 3855 7625 3975
rect 7745 3855 7800 3975
rect 7920 3855 7965 3975
rect 8085 3855 8130 3975
rect 8250 3855 8295 3975
rect 8415 3855 8470 3975
rect 8590 3855 8635 3975
rect 8755 3855 8800 3975
rect 8920 3855 8965 3975
rect 9085 3855 9140 3975
rect 9260 3855 9305 3975
rect 9425 3855 9470 3975
rect 9590 3855 9635 3975
rect 9755 3855 9810 3975
rect 9930 3855 9975 3975
rect 10095 3855 10140 3975
rect 10260 3855 10305 3975
rect 10425 3855 10480 3975
rect 10600 3855 10645 3975
rect 10765 3855 10810 3975
rect 10930 3855 10975 3975
rect 11095 3855 11150 3975
rect 11270 3855 11315 3975
rect 11435 3855 11480 3975
rect 11600 3855 11645 3975
rect 11765 3855 11820 3975
rect 11940 3855 11985 3975
rect 12105 3855 12150 3975
rect 12270 3855 12315 3975
rect 12435 3855 12490 3975
rect 12610 3855 12635 3975
rect 7105 3810 12635 3855
rect 7105 3690 7130 3810
rect 7250 3690 7295 3810
rect 7415 3690 7460 3810
rect 7580 3690 7625 3810
rect 7745 3690 7800 3810
rect 7920 3690 7965 3810
rect 8085 3690 8130 3810
rect 8250 3690 8295 3810
rect 8415 3690 8470 3810
rect 8590 3690 8635 3810
rect 8755 3690 8800 3810
rect 8920 3690 8965 3810
rect 9085 3690 9140 3810
rect 9260 3690 9305 3810
rect 9425 3690 9470 3810
rect 9590 3690 9635 3810
rect 9755 3690 9810 3810
rect 9930 3690 9975 3810
rect 10095 3690 10140 3810
rect 10260 3690 10305 3810
rect 10425 3690 10480 3810
rect 10600 3690 10645 3810
rect 10765 3690 10810 3810
rect 10930 3690 10975 3810
rect 11095 3690 11150 3810
rect 11270 3690 11315 3810
rect 11435 3690 11480 3810
rect 11600 3690 11645 3810
rect 11765 3690 11820 3810
rect 11940 3690 11985 3810
rect 12105 3690 12150 3810
rect 12270 3690 12315 3810
rect 12435 3690 12490 3810
rect 12610 3690 12635 3810
rect 7105 3635 12635 3690
rect 7105 3515 7130 3635
rect 7250 3515 7295 3635
rect 7415 3515 7460 3635
rect 7580 3515 7625 3635
rect 7745 3515 7800 3635
rect 7920 3515 7965 3635
rect 8085 3515 8130 3635
rect 8250 3515 8295 3635
rect 8415 3515 8470 3635
rect 8590 3515 8635 3635
rect 8755 3515 8800 3635
rect 8920 3515 8965 3635
rect 9085 3515 9140 3635
rect 9260 3515 9305 3635
rect 9425 3515 9470 3635
rect 9590 3515 9635 3635
rect 9755 3515 9810 3635
rect 9930 3515 9975 3635
rect 10095 3515 10140 3635
rect 10260 3515 10305 3635
rect 10425 3515 10480 3635
rect 10600 3515 10645 3635
rect 10765 3515 10810 3635
rect 10930 3515 10975 3635
rect 11095 3515 11150 3635
rect 11270 3515 11315 3635
rect 11435 3515 11480 3635
rect 11600 3515 11645 3635
rect 11765 3515 11820 3635
rect 11940 3515 11985 3635
rect 12105 3515 12150 3635
rect 12270 3515 12315 3635
rect 12435 3515 12490 3635
rect 12610 3515 12635 3635
rect 7105 3470 12635 3515
rect 7105 3350 7130 3470
rect 7250 3350 7295 3470
rect 7415 3350 7460 3470
rect 7580 3350 7625 3470
rect 7745 3350 7800 3470
rect 7920 3350 7965 3470
rect 8085 3350 8130 3470
rect 8250 3350 8295 3470
rect 8415 3350 8470 3470
rect 8590 3350 8635 3470
rect 8755 3350 8800 3470
rect 8920 3350 8965 3470
rect 9085 3350 9140 3470
rect 9260 3350 9305 3470
rect 9425 3350 9470 3470
rect 9590 3350 9635 3470
rect 9755 3350 9810 3470
rect 9930 3350 9975 3470
rect 10095 3350 10140 3470
rect 10260 3350 10305 3470
rect 10425 3350 10480 3470
rect 10600 3350 10645 3470
rect 10765 3350 10810 3470
rect 10930 3350 10975 3470
rect 11095 3350 11150 3470
rect 11270 3350 11315 3470
rect 11435 3350 11480 3470
rect 11600 3350 11645 3470
rect 11765 3350 11820 3470
rect 11940 3350 11985 3470
rect 12105 3350 12150 3470
rect 12270 3350 12315 3470
rect 12435 3350 12490 3470
rect 12610 3350 12635 3470
rect 7105 3305 12635 3350
rect 7105 3185 7130 3305
rect 7250 3185 7295 3305
rect 7415 3185 7460 3305
rect 7580 3185 7625 3305
rect 7745 3185 7800 3305
rect 7920 3185 7965 3305
rect 8085 3185 8130 3305
rect 8250 3185 8295 3305
rect 8415 3185 8470 3305
rect 8590 3185 8635 3305
rect 8755 3185 8800 3305
rect 8920 3185 8965 3305
rect 9085 3185 9140 3305
rect 9260 3185 9305 3305
rect 9425 3185 9470 3305
rect 9590 3185 9635 3305
rect 9755 3185 9810 3305
rect 9930 3185 9975 3305
rect 10095 3185 10140 3305
rect 10260 3185 10305 3305
rect 10425 3185 10480 3305
rect 10600 3185 10645 3305
rect 10765 3185 10810 3305
rect 10930 3185 10975 3305
rect 11095 3185 11150 3305
rect 11270 3185 11315 3305
rect 11435 3185 11480 3305
rect 11600 3185 11645 3305
rect 11765 3185 11820 3305
rect 11940 3185 11985 3305
rect 12105 3185 12150 3305
rect 12270 3185 12315 3305
rect 12435 3185 12490 3305
rect 12610 3185 12635 3305
rect 7105 3140 12635 3185
rect 7105 3020 7130 3140
rect 7250 3020 7295 3140
rect 7415 3020 7460 3140
rect 7580 3020 7625 3140
rect 7745 3020 7800 3140
rect 7920 3020 7965 3140
rect 8085 3020 8130 3140
rect 8250 3020 8295 3140
rect 8415 3020 8470 3140
rect 8590 3020 8635 3140
rect 8755 3020 8800 3140
rect 8920 3020 8965 3140
rect 9085 3020 9140 3140
rect 9260 3020 9305 3140
rect 9425 3020 9470 3140
rect 9590 3020 9635 3140
rect 9755 3020 9810 3140
rect 9930 3020 9975 3140
rect 10095 3020 10140 3140
rect 10260 3020 10305 3140
rect 10425 3020 10480 3140
rect 10600 3020 10645 3140
rect 10765 3020 10810 3140
rect 10930 3020 10975 3140
rect 11095 3020 11150 3140
rect 11270 3020 11315 3140
rect 11435 3020 11480 3140
rect 11600 3020 11645 3140
rect 11765 3020 11820 3140
rect 11940 3020 11985 3140
rect 12105 3020 12150 3140
rect 12270 3020 12315 3140
rect 12435 3020 12490 3140
rect 12610 3020 12635 3140
rect 7105 2965 12635 3020
rect 7105 2845 7130 2965
rect 7250 2845 7295 2965
rect 7415 2845 7460 2965
rect 7580 2845 7625 2965
rect 7745 2845 7800 2965
rect 7920 2845 7965 2965
rect 8085 2845 8130 2965
rect 8250 2845 8295 2965
rect 8415 2845 8470 2965
rect 8590 2845 8635 2965
rect 8755 2845 8800 2965
rect 8920 2845 8965 2965
rect 9085 2845 9140 2965
rect 9260 2845 9305 2965
rect 9425 2845 9470 2965
rect 9590 2845 9635 2965
rect 9755 2845 9810 2965
rect 9930 2845 9975 2965
rect 10095 2845 10140 2965
rect 10260 2845 10305 2965
rect 10425 2845 10480 2965
rect 10600 2845 10645 2965
rect 10765 2845 10810 2965
rect 10930 2845 10975 2965
rect 11095 2845 11150 2965
rect 11270 2845 11315 2965
rect 11435 2845 11480 2965
rect 11600 2845 11645 2965
rect 11765 2845 11820 2965
rect 11940 2845 11985 2965
rect 12105 2845 12150 2965
rect 12270 2845 12315 2965
rect 12435 2845 12490 2965
rect 12610 2845 12635 2965
rect 7105 2800 12635 2845
rect 7105 2680 7130 2800
rect 7250 2680 7295 2800
rect 7415 2680 7460 2800
rect 7580 2680 7625 2800
rect 7745 2680 7800 2800
rect 7920 2680 7965 2800
rect 8085 2680 8130 2800
rect 8250 2680 8295 2800
rect 8415 2680 8470 2800
rect 8590 2680 8635 2800
rect 8755 2680 8800 2800
rect 8920 2680 8965 2800
rect 9085 2680 9140 2800
rect 9260 2680 9305 2800
rect 9425 2680 9470 2800
rect 9590 2680 9635 2800
rect 9755 2680 9810 2800
rect 9930 2680 9975 2800
rect 10095 2680 10140 2800
rect 10260 2680 10305 2800
rect 10425 2680 10480 2800
rect 10600 2680 10645 2800
rect 10765 2680 10810 2800
rect 10930 2680 10975 2800
rect 11095 2680 11150 2800
rect 11270 2680 11315 2800
rect 11435 2680 11480 2800
rect 11600 2680 11645 2800
rect 11765 2680 11820 2800
rect 11940 2680 11985 2800
rect 12105 2680 12150 2800
rect 12270 2680 12315 2800
rect 12435 2680 12490 2800
rect 12610 2680 12635 2800
rect 7105 2635 12635 2680
rect 7105 2515 7130 2635
rect 7250 2515 7295 2635
rect 7415 2515 7460 2635
rect 7580 2515 7625 2635
rect 7745 2515 7800 2635
rect 7920 2515 7965 2635
rect 8085 2515 8130 2635
rect 8250 2515 8295 2635
rect 8415 2515 8470 2635
rect 8590 2515 8635 2635
rect 8755 2515 8800 2635
rect 8920 2515 8965 2635
rect 9085 2515 9140 2635
rect 9260 2515 9305 2635
rect 9425 2515 9470 2635
rect 9590 2515 9635 2635
rect 9755 2515 9810 2635
rect 9930 2515 9975 2635
rect 10095 2515 10140 2635
rect 10260 2515 10305 2635
rect 10425 2515 10480 2635
rect 10600 2515 10645 2635
rect 10765 2515 10810 2635
rect 10930 2515 10975 2635
rect 11095 2515 11150 2635
rect 11270 2515 11315 2635
rect 11435 2515 11480 2635
rect 11600 2515 11645 2635
rect 11765 2515 11820 2635
rect 11940 2515 11985 2635
rect 12105 2515 12150 2635
rect 12270 2515 12315 2635
rect 12435 2515 12490 2635
rect 12610 2515 12635 2635
rect 7105 2470 12635 2515
rect 7105 2350 7130 2470
rect 7250 2350 7295 2470
rect 7415 2350 7460 2470
rect 7580 2350 7625 2470
rect 7745 2350 7800 2470
rect 7920 2350 7965 2470
rect 8085 2350 8130 2470
rect 8250 2350 8295 2470
rect 8415 2350 8470 2470
rect 8590 2350 8635 2470
rect 8755 2350 8800 2470
rect 8920 2350 8965 2470
rect 9085 2350 9140 2470
rect 9260 2350 9305 2470
rect 9425 2350 9470 2470
rect 9590 2350 9635 2470
rect 9755 2350 9810 2470
rect 9930 2350 9975 2470
rect 10095 2350 10140 2470
rect 10260 2350 10305 2470
rect 10425 2350 10480 2470
rect 10600 2350 10645 2470
rect 10765 2350 10810 2470
rect 10930 2350 10975 2470
rect 11095 2350 11150 2470
rect 11270 2350 11315 2470
rect 11435 2350 11480 2470
rect 11600 2350 11645 2470
rect 11765 2350 11820 2470
rect 11940 2350 11985 2470
rect 12105 2350 12150 2470
rect 12270 2350 12315 2470
rect 12435 2350 12490 2470
rect 12610 2350 12635 2470
rect 7105 2295 12635 2350
rect 7105 2175 7130 2295
rect 7250 2175 7295 2295
rect 7415 2175 7460 2295
rect 7580 2175 7625 2295
rect 7745 2175 7800 2295
rect 7920 2175 7965 2295
rect 8085 2175 8130 2295
rect 8250 2175 8295 2295
rect 8415 2175 8470 2295
rect 8590 2175 8635 2295
rect 8755 2175 8800 2295
rect 8920 2175 8965 2295
rect 9085 2175 9140 2295
rect 9260 2175 9305 2295
rect 9425 2175 9470 2295
rect 9590 2175 9635 2295
rect 9755 2175 9810 2295
rect 9930 2175 9975 2295
rect 10095 2175 10140 2295
rect 10260 2175 10305 2295
rect 10425 2175 10480 2295
rect 10600 2175 10645 2295
rect 10765 2175 10810 2295
rect 10930 2175 10975 2295
rect 11095 2175 11150 2295
rect 11270 2175 11315 2295
rect 11435 2175 11480 2295
rect 11600 2175 11645 2295
rect 11765 2175 11820 2295
rect 11940 2175 11985 2295
rect 12105 2175 12150 2295
rect 12270 2175 12315 2295
rect 12435 2175 12490 2295
rect 12610 2175 12635 2295
rect 7105 2130 12635 2175
rect 7105 2010 7130 2130
rect 7250 2010 7295 2130
rect 7415 2010 7460 2130
rect 7580 2010 7625 2130
rect 7745 2010 7800 2130
rect 7920 2010 7965 2130
rect 8085 2010 8130 2130
rect 8250 2010 8295 2130
rect 8415 2010 8470 2130
rect 8590 2010 8635 2130
rect 8755 2010 8800 2130
rect 8920 2010 8965 2130
rect 9085 2010 9140 2130
rect 9260 2010 9305 2130
rect 9425 2010 9470 2130
rect 9590 2010 9635 2130
rect 9755 2010 9810 2130
rect 9930 2010 9975 2130
rect 10095 2010 10140 2130
rect 10260 2010 10305 2130
rect 10425 2010 10480 2130
rect 10600 2010 10645 2130
rect 10765 2010 10810 2130
rect 10930 2010 10975 2130
rect 11095 2010 11150 2130
rect 11270 2010 11315 2130
rect 11435 2010 11480 2130
rect 11600 2010 11645 2130
rect 11765 2010 11820 2130
rect 11940 2010 11985 2130
rect 12105 2010 12150 2130
rect 12270 2010 12315 2130
rect 12435 2010 12490 2130
rect 12610 2010 12635 2130
rect 7105 1965 12635 2010
rect 7105 1845 7130 1965
rect 7250 1845 7295 1965
rect 7415 1845 7460 1965
rect 7580 1845 7625 1965
rect 7745 1845 7800 1965
rect 7920 1845 7965 1965
rect 8085 1845 8130 1965
rect 8250 1845 8295 1965
rect 8415 1845 8470 1965
rect 8590 1845 8635 1965
rect 8755 1845 8800 1965
rect 8920 1845 8965 1965
rect 9085 1845 9140 1965
rect 9260 1845 9305 1965
rect 9425 1845 9470 1965
rect 9590 1845 9635 1965
rect 9755 1845 9810 1965
rect 9930 1845 9975 1965
rect 10095 1845 10140 1965
rect 10260 1845 10305 1965
rect 10425 1845 10480 1965
rect 10600 1845 10645 1965
rect 10765 1845 10810 1965
rect 10930 1845 10975 1965
rect 11095 1845 11150 1965
rect 11270 1845 11315 1965
rect 11435 1845 11480 1965
rect 11600 1845 11645 1965
rect 11765 1845 11820 1965
rect 11940 1845 11985 1965
rect 12105 1845 12150 1965
rect 12270 1845 12315 1965
rect 12435 1845 12490 1965
rect 12610 1845 12635 1965
rect 7105 1800 12635 1845
rect 7105 1680 7130 1800
rect 7250 1680 7295 1800
rect 7415 1680 7460 1800
rect 7580 1680 7625 1800
rect 7745 1680 7800 1800
rect 7920 1680 7965 1800
rect 8085 1680 8130 1800
rect 8250 1680 8295 1800
rect 8415 1680 8470 1800
rect 8590 1680 8635 1800
rect 8755 1680 8800 1800
rect 8920 1680 8965 1800
rect 9085 1680 9140 1800
rect 9260 1680 9305 1800
rect 9425 1680 9470 1800
rect 9590 1680 9635 1800
rect 9755 1680 9810 1800
rect 9930 1680 9975 1800
rect 10095 1680 10140 1800
rect 10260 1680 10305 1800
rect 10425 1680 10480 1800
rect 10600 1680 10645 1800
rect 10765 1680 10810 1800
rect 10930 1680 10975 1800
rect 11095 1680 11150 1800
rect 11270 1680 11315 1800
rect 11435 1680 11480 1800
rect 11600 1680 11645 1800
rect 11765 1680 11820 1800
rect 11940 1680 11985 1800
rect 12105 1680 12150 1800
rect 12270 1680 12315 1800
rect 12435 1680 12490 1800
rect 12610 1680 12635 1800
rect 7105 1655 12635 1680
rect 12795 7040 12820 7125
rect 12940 7040 12985 7160
rect 13105 7040 13150 7160
rect 13270 7040 13315 7160
rect 13435 7040 13490 7160
rect 13610 7040 13655 7160
rect 13775 7040 13820 7160
rect 13940 7040 13985 7160
rect 14105 7040 14160 7160
rect 14280 7040 14325 7160
rect 14445 7040 14490 7160
rect 14610 7040 14655 7160
rect 14775 7040 14830 7160
rect 14950 7040 14995 7160
rect 15115 7040 15160 7160
rect 15280 7040 15325 7160
rect 15445 7040 15500 7160
rect 15620 7040 15665 7160
rect 15785 7040 15830 7160
rect 15950 7040 15995 7160
rect 16115 7040 16170 7160
rect 16290 7040 16335 7160
rect 16455 7040 16500 7160
rect 16620 7040 16665 7160
rect 16785 7040 16840 7160
rect 16960 7040 17005 7160
rect 17125 7040 17170 7160
rect 17290 7040 17335 7160
rect 17455 7040 17510 7160
rect 17630 7040 17675 7160
rect 17795 7040 17840 7160
rect 17960 7040 18005 7160
rect 18125 7040 18180 7160
rect 18300 7125 18510 7160
rect 18300 7040 18325 7125
rect 12795 6985 18325 7040
rect 12795 6865 12820 6985
rect 12940 6865 12985 6985
rect 13105 6865 13150 6985
rect 13270 6865 13315 6985
rect 13435 6865 13490 6985
rect 13610 6865 13655 6985
rect 13775 6865 13820 6985
rect 13940 6865 13985 6985
rect 14105 6865 14160 6985
rect 14280 6865 14325 6985
rect 14445 6865 14490 6985
rect 14610 6865 14655 6985
rect 14775 6865 14830 6985
rect 14950 6865 14995 6985
rect 15115 6865 15160 6985
rect 15280 6865 15325 6985
rect 15445 6865 15500 6985
rect 15620 6865 15665 6985
rect 15785 6865 15830 6985
rect 15950 6865 15995 6985
rect 16115 6865 16170 6985
rect 16290 6865 16335 6985
rect 16455 6865 16500 6985
rect 16620 6865 16665 6985
rect 16785 6865 16840 6985
rect 16960 6865 17005 6985
rect 17125 6865 17170 6985
rect 17290 6865 17335 6985
rect 17455 6865 17510 6985
rect 17630 6865 17675 6985
rect 17795 6865 17840 6985
rect 17960 6865 18005 6985
rect 18125 6865 18180 6985
rect 18300 6865 18325 6985
rect 12795 6820 18325 6865
rect 12795 6700 12820 6820
rect 12940 6700 12985 6820
rect 13105 6700 13150 6820
rect 13270 6700 13315 6820
rect 13435 6700 13490 6820
rect 13610 6700 13655 6820
rect 13775 6700 13820 6820
rect 13940 6700 13985 6820
rect 14105 6700 14160 6820
rect 14280 6700 14325 6820
rect 14445 6700 14490 6820
rect 14610 6700 14655 6820
rect 14775 6700 14830 6820
rect 14950 6700 14995 6820
rect 15115 6700 15160 6820
rect 15280 6700 15325 6820
rect 15445 6700 15500 6820
rect 15620 6700 15665 6820
rect 15785 6700 15830 6820
rect 15950 6700 15995 6820
rect 16115 6700 16170 6820
rect 16290 6700 16335 6820
rect 16455 6700 16500 6820
rect 16620 6700 16665 6820
rect 16785 6700 16840 6820
rect 16960 6700 17005 6820
rect 17125 6700 17170 6820
rect 17290 6700 17335 6820
rect 17455 6700 17510 6820
rect 17630 6700 17675 6820
rect 17795 6700 17840 6820
rect 17960 6700 18005 6820
rect 18125 6700 18180 6820
rect 18300 6700 18325 6820
rect 12795 6655 18325 6700
rect 12795 6535 12820 6655
rect 12940 6535 12985 6655
rect 13105 6535 13150 6655
rect 13270 6535 13315 6655
rect 13435 6535 13490 6655
rect 13610 6535 13655 6655
rect 13775 6535 13820 6655
rect 13940 6535 13985 6655
rect 14105 6535 14160 6655
rect 14280 6535 14325 6655
rect 14445 6535 14490 6655
rect 14610 6535 14655 6655
rect 14775 6535 14830 6655
rect 14950 6535 14995 6655
rect 15115 6535 15160 6655
rect 15280 6535 15325 6655
rect 15445 6535 15500 6655
rect 15620 6535 15665 6655
rect 15785 6535 15830 6655
rect 15950 6535 15995 6655
rect 16115 6535 16170 6655
rect 16290 6535 16335 6655
rect 16455 6535 16500 6655
rect 16620 6535 16665 6655
rect 16785 6535 16840 6655
rect 16960 6535 17005 6655
rect 17125 6535 17170 6655
rect 17290 6535 17335 6655
rect 17455 6535 17510 6655
rect 17630 6535 17675 6655
rect 17795 6535 17840 6655
rect 17960 6535 18005 6655
rect 18125 6535 18180 6655
rect 18300 6535 18325 6655
rect 12795 6490 18325 6535
rect 12795 6370 12820 6490
rect 12940 6370 12985 6490
rect 13105 6370 13150 6490
rect 13270 6370 13315 6490
rect 13435 6370 13490 6490
rect 13610 6370 13655 6490
rect 13775 6370 13820 6490
rect 13940 6370 13985 6490
rect 14105 6370 14160 6490
rect 14280 6370 14325 6490
rect 14445 6370 14490 6490
rect 14610 6370 14655 6490
rect 14775 6370 14830 6490
rect 14950 6370 14995 6490
rect 15115 6370 15160 6490
rect 15280 6370 15325 6490
rect 15445 6370 15500 6490
rect 15620 6370 15665 6490
rect 15785 6370 15830 6490
rect 15950 6370 15995 6490
rect 16115 6370 16170 6490
rect 16290 6370 16335 6490
rect 16455 6370 16500 6490
rect 16620 6370 16665 6490
rect 16785 6370 16840 6490
rect 16960 6370 17005 6490
rect 17125 6370 17170 6490
rect 17290 6370 17335 6490
rect 17455 6370 17510 6490
rect 17630 6370 17675 6490
rect 17795 6370 17840 6490
rect 17960 6370 18005 6490
rect 18125 6370 18180 6490
rect 18300 6370 18325 6490
rect 12795 6315 18325 6370
rect 12795 6195 12820 6315
rect 12940 6195 12985 6315
rect 13105 6195 13150 6315
rect 13270 6195 13315 6315
rect 13435 6195 13490 6315
rect 13610 6195 13655 6315
rect 13775 6195 13820 6315
rect 13940 6195 13985 6315
rect 14105 6195 14160 6315
rect 14280 6195 14325 6315
rect 14445 6195 14490 6315
rect 14610 6195 14655 6315
rect 14775 6195 14830 6315
rect 14950 6195 14995 6315
rect 15115 6195 15160 6315
rect 15280 6195 15325 6315
rect 15445 6195 15500 6315
rect 15620 6195 15665 6315
rect 15785 6195 15830 6315
rect 15950 6195 15995 6315
rect 16115 6195 16170 6315
rect 16290 6195 16335 6315
rect 16455 6195 16500 6315
rect 16620 6195 16665 6315
rect 16785 6195 16840 6315
rect 16960 6195 17005 6315
rect 17125 6195 17170 6315
rect 17290 6195 17335 6315
rect 17455 6195 17510 6315
rect 17630 6195 17675 6315
rect 17795 6195 17840 6315
rect 17960 6195 18005 6315
rect 18125 6195 18180 6315
rect 18300 6195 18325 6315
rect 12795 6150 18325 6195
rect 12795 6030 12820 6150
rect 12940 6030 12985 6150
rect 13105 6030 13150 6150
rect 13270 6030 13315 6150
rect 13435 6030 13490 6150
rect 13610 6030 13655 6150
rect 13775 6030 13820 6150
rect 13940 6030 13985 6150
rect 14105 6030 14160 6150
rect 14280 6030 14325 6150
rect 14445 6030 14490 6150
rect 14610 6030 14655 6150
rect 14775 6030 14830 6150
rect 14950 6030 14995 6150
rect 15115 6030 15160 6150
rect 15280 6030 15325 6150
rect 15445 6030 15500 6150
rect 15620 6030 15665 6150
rect 15785 6030 15830 6150
rect 15950 6030 15995 6150
rect 16115 6030 16170 6150
rect 16290 6030 16335 6150
rect 16455 6030 16500 6150
rect 16620 6030 16665 6150
rect 16785 6030 16840 6150
rect 16960 6030 17005 6150
rect 17125 6030 17170 6150
rect 17290 6030 17335 6150
rect 17455 6030 17510 6150
rect 17630 6030 17675 6150
rect 17795 6030 17840 6150
rect 17960 6030 18005 6150
rect 18125 6030 18180 6150
rect 18300 6030 18325 6150
rect 12795 5985 18325 6030
rect 12795 5865 12820 5985
rect 12940 5865 12985 5985
rect 13105 5865 13150 5985
rect 13270 5865 13315 5985
rect 13435 5865 13490 5985
rect 13610 5865 13655 5985
rect 13775 5865 13820 5985
rect 13940 5865 13985 5985
rect 14105 5865 14160 5985
rect 14280 5865 14325 5985
rect 14445 5865 14490 5985
rect 14610 5865 14655 5985
rect 14775 5865 14830 5985
rect 14950 5865 14995 5985
rect 15115 5865 15160 5985
rect 15280 5865 15325 5985
rect 15445 5865 15500 5985
rect 15620 5865 15665 5985
rect 15785 5865 15830 5985
rect 15950 5865 15995 5985
rect 16115 5865 16170 5985
rect 16290 5865 16335 5985
rect 16455 5865 16500 5985
rect 16620 5865 16665 5985
rect 16785 5865 16840 5985
rect 16960 5865 17005 5985
rect 17125 5865 17170 5985
rect 17290 5865 17335 5985
rect 17455 5865 17510 5985
rect 17630 5865 17675 5985
rect 17795 5865 17840 5985
rect 17960 5865 18005 5985
rect 18125 5865 18180 5985
rect 18300 5865 18325 5985
rect 12795 5820 18325 5865
rect 12795 5700 12820 5820
rect 12940 5700 12985 5820
rect 13105 5700 13150 5820
rect 13270 5700 13315 5820
rect 13435 5700 13490 5820
rect 13610 5700 13655 5820
rect 13775 5700 13820 5820
rect 13940 5700 13985 5820
rect 14105 5700 14160 5820
rect 14280 5700 14325 5820
rect 14445 5700 14490 5820
rect 14610 5700 14655 5820
rect 14775 5700 14830 5820
rect 14950 5700 14995 5820
rect 15115 5700 15160 5820
rect 15280 5700 15325 5820
rect 15445 5700 15500 5820
rect 15620 5700 15665 5820
rect 15785 5700 15830 5820
rect 15950 5700 15995 5820
rect 16115 5700 16170 5820
rect 16290 5700 16335 5820
rect 16455 5700 16500 5820
rect 16620 5700 16665 5820
rect 16785 5700 16840 5820
rect 16960 5700 17005 5820
rect 17125 5700 17170 5820
rect 17290 5700 17335 5820
rect 17455 5700 17510 5820
rect 17630 5700 17675 5820
rect 17795 5700 17840 5820
rect 17960 5700 18005 5820
rect 18125 5700 18180 5820
rect 18300 5700 18325 5820
rect 12795 5645 18325 5700
rect 12795 5525 12820 5645
rect 12940 5525 12985 5645
rect 13105 5525 13150 5645
rect 13270 5525 13315 5645
rect 13435 5525 13490 5645
rect 13610 5525 13655 5645
rect 13775 5525 13820 5645
rect 13940 5525 13985 5645
rect 14105 5525 14160 5645
rect 14280 5525 14325 5645
rect 14445 5525 14490 5645
rect 14610 5525 14655 5645
rect 14775 5525 14830 5645
rect 14950 5525 14995 5645
rect 15115 5525 15160 5645
rect 15280 5525 15325 5645
rect 15445 5525 15500 5645
rect 15620 5525 15665 5645
rect 15785 5525 15830 5645
rect 15950 5525 15995 5645
rect 16115 5525 16170 5645
rect 16290 5525 16335 5645
rect 16455 5525 16500 5645
rect 16620 5525 16665 5645
rect 16785 5525 16840 5645
rect 16960 5525 17005 5645
rect 17125 5525 17170 5645
rect 17290 5525 17335 5645
rect 17455 5525 17510 5645
rect 17630 5525 17675 5645
rect 17795 5525 17840 5645
rect 17960 5525 18005 5645
rect 18125 5525 18180 5645
rect 18300 5525 18325 5645
rect 12795 5480 18325 5525
rect 12795 5360 12820 5480
rect 12940 5360 12985 5480
rect 13105 5360 13150 5480
rect 13270 5360 13315 5480
rect 13435 5360 13490 5480
rect 13610 5360 13655 5480
rect 13775 5360 13820 5480
rect 13940 5360 13985 5480
rect 14105 5360 14160 5480
rect 14280 5360 14325 5480
rect 14445 5360 14490 5480
rect 14610 5360 14655 5480
rect 14775 5360 14830 5480
rect 14950 5360 14995 5480
rect 15115 5360 15160 5480
rect 15280 5360 15325 5480
rect 15445 5360 15500 5480
rect 15620 5360 15665 5480
rect 15785 5360 15830 5480
rect 15950 5360 15995 5480
rect 16115 5360 16170 5480
rect 16290 5360 16335 5480
rect 16455 5360 16500 5480
rect 16620 5360 16665 5480
rect 16785 5360 16840 5480
rect 16960 5360 17005 5480
rect 17125 5360 17170 5480
rect 17290 5360 17335 5480
rect 17455 5360 17510 5480
rect 17630 5360 17675 5480
rect 17795 5360 17840 5480
rect 17960 5360 18005 5480
rect 18125 5360 18180 5480
rect 18300 5360 18325 5480
rect 12795 5315 18325 5360
rect 12795 5195 12820 5315
rect 12940 5195 12985 5315
rect 13105 5195 13150 5315
rect 13270 5195 13315 5315
rect 13435 5195 13490 5315
rect 13610 5195 13655 5315
rect 13775 5195 13820 5315
rect 13940 5195 13985 5315
rect 14105 5195 14160 5315
rect 14280 5195 14325 5315
rect 14445 5195 14490 5315
rect 14610 5195 14655 5315
rect 14775 5195 14830 5315
rect 14950 5195 14995 5315
rect 15115 5195 15160 5315
rect 15280 5195 15325 5315
rect 15445 5195 15500 5315
rect 15620 5195 15665 5315
rect 15785 5195 15830 5315
rect 15950 5195 15995 5315
rect 16115 5195 16170 5315
rect 16290 5195 16335 5315
rect 16455 5195 16500 5315
rect 16620 5195 16665 5315
rect 16785 5195 16840 5315
rect 16960 5195 17005 5315
rect 17125 5195 17170 5315
rect 17290 5195 17335 5315
rect 17455 5195 17510 5315
rect 17630 5195 17675 5315
rect 17795 5195 17840 5315
rect 17960 5195 18005 5315
rect 18125 5195 18180 5315
rect 18300 5195 18325 5315
rect 12795 5150 18325 5195
rect 12795 5030 12820 5150
rect 12940 5030 12985 5150
rect 13105 5030 13150 5150
rect 13270 5030 13315 5150
rect 13435 5030 13490 5150
rect 13610 5030 13655 5150
rect 13775 5030 13820 5150
rect 13940 5030 13985 5150
rect 14105 5030 14160 5150
rect 14280 5030 14325 5150
rect 14445 5030 14490 5150
rect 14610 5030 14655 5150
rect 14775 5030 14830 5150
rect 14950 5030 14995 5150
rect 15115 5030 15160 5150
rect 15280 5030 15325 5150
rect 15445 5030 15500 5150
rect 15620 5030 15665 5150
rect 15785 5030 15830 5150
rect 15950 5030 15995 5150
rect 16115 5030 16170 5150
rect 16290 5030 16335 5150
rect 16455 5030 16500 5150
rect 16620 5030 16665 5150
rect 16785 5030 16840 5150
rect 16960 5030 17005 5150
rect 17125 5030 17170 5150
rect 17290 5030 17335 5150
rect 17455 5030 17510 5150
rect 17630 5030 17675 5150
rect 17795 5030 17840 5150
rect 17960 5030 18005 5150
rect 18125 5030 18180 5150
rect 18300 5030 18325 5150
rect 12795 4975 18325 5030
rect 12795 4855 12820 4975
rect 12940 4855 12985 4975
rect 13105 4855 13150 4975
rect 13270 4855 13315 4975
rect 13435 4855 13490 4975
rect 13610 4855 13655 4975
rect 13775 4855 13820 4975
rect 13940 4855 13985 4975
rect 14105 4855 14160 4975
rect 14280 4855 14325 4975
rect 14445 4855 14490 4975
rect 14610 4855 14655 4975
rect 14775 4855 14830 4975
rect 14950 4855 14995 4975
rect 15115 4855 15160 4975
rect 15280 4855 15325 4975
rect 15445 4855 15500 4975
rect 15620 4855 15665 4975
rect 15785 4855 15830 4975
rect 15950 4855 15995 4975
rect 16115 4855 16170 4975
rect 16290 4855 16335 4975
rect 16455 4855 16500 4975
rect 16620 4855 16665 4975
rect 16785 4855 16840 4975
rect 16960 4855 17005 4975
rect 17125 4855 17170 4975
rect 17290 4855 17335 4975
rect 17455 4855 17510 4975
rect 17630 4855 17675 4975
rect 17795 4855 17840 4975
rect 17960 4855 18005 4975
rect 18125 4855 18180 4975
rect 18300 4855 18325 4975
rect 12795 4810 18325 4855
rect 12795 4690 12820 4810
rect 12940 4690 12985 4810
rect 13105 4690 13150 4810
rect 13270 4690 13315 4810
rect 13435 4690 13490 4810
rect 13610 4690 13655 4810
rect 13775 4690 13820 4810
rect 13940 4690 13985 4810
rect 14105 4690 14160 4810
rect 14280 4690 14325 4810
rect 14445 4690 14490 4810
rect 14610 4690 14655 4810
rect 14775 4690 14830 4810
rect 14950 4690 14995 4810
rect 15115 4690 15160 4810
rect 15280 4690 15325 4810
rect 15445 4690 15500 4810
rect 15620 4690 15665 4810
rect 15785 4690 15830 4810
rect 15950 4690 15995 4810
rect 16115 4690 16170 4810
rect 16290 4690 16335 4810
rect 16455 4690 16500 4810
rect 16620 4690 16665 4810
rect 16785 4690 16840 4810
rect 16960 4690 17005 4810
rect 17125 4690 17170 4810
rect 17290 4690 17335 4810
rect 17455 4690 17510 4810
rect 17630 4690 17675 4810
rect 17795 4690 17840 4810
rect 17960 4690 18005 4810
rect 18125 4690 18180 4810
rect 18300 4690 18325 4810
rect 12795 4645 18325 4690
rect 12795 4525 12820 4645
rect 12940 4525 12985 4645
rect 13105 4525 13150 4645
rect 13270 4525 13315 4645
rect 13435 4525 13490 4645
rect 13610 4525 13655 4645
rect 13775 4525 13820 4645
rect 13940 4525 13985 4645
rect 14105 4525 14160 4645
rect 14280 4525 14325 4645
rect 14445 4525 14490 4645
rect 14610 4525 14655 4645
rect 14775 4525 14830 4645
rect 14950 4525 14995 4645
rect 15115 4525 15160 4645
rect 15280 4525 15325 4645
rect 15445 4525 15500 4645
rect 15620 4525 15665 4645
rect 15785 4525 15830 4645
rect 15950 4525 15995 4645
rect 16115 4525 16170 4645
rect 16290 4525 16335 4645
rect 16455 4525 16500 4645
rect 16620 4525 16665 4645
rect 16785 4525 16840 4645
rect 16960 4525 17005 4645
rect 17125 4525 17170 4645
rect 17290 4525 17335 4645
rect 17455 4525 17510 4645
rect 17630 4525 17675 4645
rect 17795 4525 17840 4645
rect 17960 4525 18005 4645
rect 18125 4525 18180 4645
rect 18300 4525 18325 4645
rect 12795 4480 18325 4525
rect 12795 4360 12820 4480
rect 12940 4360 12985 4480
rect 13105 4360 13150 4480
rect 13270 4360 13315 4480
rect 13435 4360 13490 4480
rect 13610 4360 13655 4480
rect 13775 4360 13820 4480
rect 13940 4360 13985 4480
rect 14105 4360 14160 4480
rect 14280 4360 14325 4480
rect 14445 4360 14490 4480
rect 14610 4360 14655 4480
rect 14775 4360 14830 4480
rect 14950 4360 14995 4480
rect 15115 4360 15160 4480
rect 15280 4360 15325 4480
rect 15445 4360 15500 4480
rect 15620 4360 15665 4480
rect 15785 4360 15830 4480
rect 15950 4360 15995 4480
rect 16115 4360 16170 4480
rect 16290 4360 16335 4480
rect 16455 4360 16500 4480
rect 16620 4360 16665 4480
rect 16785 4360 16840 4480
rect 16960 4360 17005 4480
rect 17125 4360 17170 4480
rect 17290 4360 17335 4480
rect 17455 4360 17510 4480
rect 17630 4360 17675 4480
rect 17795 4360 17840 4480
rect 17960 4360 18005 4480
rect 18125 4360 18180 4480
rect 18300 4360 18325 4480
rect 12795 4305 18325 4360
rect 12795 4185 12820 4305
rect 12940 4185 12985 4305
rect 13105 4185 13150 4305
rect 13270 4185 13315 4305
rect 13435 4185 13490 4305
rect 13610 4185 13655 4305
rect 13775 4185 13820 4305
rect 13940 4185 13985 4305
rect 14105 4185 14160 4305
rect 14280 4185 14325 4305
rect 14445 4185 14490 4305
rect 14610 4185 14655 4305
rect 14775 4185 14830 4305
rect 14950 4185 14995 4305
rect 15115 4185 15160 4305
rect 15280 4185 15325 4305
rect 15445 4185 15500 4305
rect 15620 4185 15665 4305
rect 15785 4185 15830 4305
rect 15950 4185 15995 4305
rect 16115 4185 16170 4305
rect 16290 4185 16335 4305
rect 16455 4185 16500 4305
rect 16620 4185 16665 4305
rect 16785 4185 16840 4305
rect 16960 4185 17005 4305
rect 17125 4185 17170 4305
rect 17290 4185 17335 4305
rect 17455 4185 17510 4305
rect 17630 4185 17675 4305
rect 17795 4185 17840 4305
rect 17960 4185 18005 4305
rect 18125 4185 18180 4305
rect 18300 4185 18325 4305
rect 12795 4140 18325 4185
rect 12795 4020 12820 4140
rect 12940 4020 12985 4140
rect 13105 4020 13150 4140
rect 13270 4020 13315 4140
rect 13435 4020 13490 4140
rect 13610 4020 13655 4140
rect 13775 4020 13820 4140
rect 13940 4020 13985 4140
rect 14105 4020 14160 4140
rect 14280 4020 14325 4140
rect 14445 4020 14490 4140
rect 14610 4020 14655 4140
rect 14775 4020 14830 4140
rect 14950 4020 14995 4140
rect 15115 4020 15160 4140
rect 15280 4020 15325 4140
rect 15445 4020 15500 4140
rect 15620 4020 15665 4140
rect 15785 4020 15830 4140
rect 15950 4020 15995 4140
rect 16115 4020 16170 4140
rect 16290 4020 16335 4140
rect 16455 4020 16500 4140
rect 16620 4020 16665 4140
rect 16785 4020 16840 4140
rect 16960 4020 17005 4140
rect 17125 4020 17170 4140
rect 17290 4020 17335 4140
rect 17455 4020 17510 4140
rect 17630 4020 17675 4140
rect 17795 4020 17840 4140
rect 17960 4020 18005 4140
rect 18125 4020 18180 4140
rect 18300 4020 18325 4140
rect 12795 3975 18325 4020
rect 12795 3855 12820 3975
rect 12940 3855 12985 3975
rect 13105 3855 13150 3975
rect 13270 3855 13315 3975
rect 13435 3855 13490 3975
rect 13610 3855 13655 3975
rect 13775 3855 13820 3975
rect 13940 3855 13985 3975
rect 14105 3855 14160 3975
rect 14280 3855 14325 3975
rect 14445 3855 14490 3975
rect 14610 3855 14655 3975
rect 14775 3855 14830 3975
rect 14950 3855 14995 3975
rect 15115 3855 15160 3975
rect 15280 3855 15325 3975
rect 15445 3855 15500 3975
rect 15620 3855 15665 3975
rect 15785 3855 15830 3975
rect 15950 3855 15995 3975
rect 16115 3855 16170 3975
rect 16290 3855 16335 3975
rect 16455 3855 16500 3975
rect 16620 3855 16665 3975
rect 16785 3855 16840 3975
rect 16960 3855 17005 3975
rect 17125 3855 17170 3975
rect 17290 3855 17335 3975
rect 17455 3855 17510 3975
rect 17630 3855 17675 3975
rect 17795 3855 17840 3975
rect 17960 3855 18005 3975
rect 18125 3855 18180 3975
rect 18300 3855 18325 3975
rect 12795 3810 18325 3855
rect 12795 3690 12820 3810
rect 12940 3690 12985 3810
rect 13105 3690 13150 3810
rect 13270 3690 13315 3810
rect 13435 3690 13490 3810
rect 13610 3690 13655 3810
rect 13775 3690 13820 3810
rect 13940 3690 13985 3810
rect 14105 3690 14160 3810
rect 14280 3690 14325 3810
rect 14445 3690 14490 3810
rect 14610 3690 14655 3810
rect 14775 3690 14830 3810
rect 14950 3690 14995 3810
rect 15115 3690 15160 3810
rect 15280 3690 15325 3810
rect 15445 3690 15500 3810
rect 15620 3690 15665 3810
rect 15785 3690 15830 3810
rect 15950 3690 15995 3810
rect 16115 3690 16170 3810
rect 16290 3690 16335 3810
rect 16455 3690 16500 3810
rect 16620 3690 16665 3810
rect 16785 3690 16840 3810
rect 16960 3690 17005 3810
rect 17125 3690 17170 3810
rect 17290 3690 17335 3810
rect 17455 3690 17510 3810
rect 17630 3690 17675 3810
rect 17795 3690 17840 3810
rect 17960 3690 18005 3810
rect 18125 3690 18180 3810
rect 18300 3690 18325 3810
rect 12795 3635 18325 3690
rect 12795 3515 12820 3635
rect 12940 3515 12985 3635
rect 13105 3515 13150 3635
rect 13270 3515 13315 3635
rect 13435 3515 13490 3635
rect 13610 3515 13655 3635
rect 13775 3515 13820 3635
rect 13940 3515 13985 3635
rect 14105 3515 14160 3635
rect 14280 3515 14325 3635
rect 14445 3515 14490 3635
rect 14610 3515 14655 3635
rect 14775 3515 14830 3635
rect 14950 3515 14995 3635
rect 15115 3515 15160 3635
rect 15280 3515 15325 3635
rect 15445 3515 15500 3635
rect 15620 3515 15665 3635
rect 15785 3515 15830 3635
rect 15950 3515 15995 3635
rect 16115 3515 16170 3635
rect 16290 3515 16335 3635
rect 16455 3515 16500 3635
rect 16620 3515 16665 3635
rect 16785 3515 16840 3635
rect 16960 3515 17005 3635
rect 17125 3515 17170 3635
rect 17290 3515 17335 3635
rect 17455 3515 17510 3635
rect 17630 3515 17675 3635
rect 17795 3515 17840 3635
rect 17960 3515 18005 3635
rect 18125 3515 18180 3635
rect 18300 3515 18325 3635
rect 12795 3470 18325 3515
rect 12795 3350 12820 3470
rect 12940 3350 12985 3470
rect 13105 3350 13150 3470
rect 13270 3350 13315 3470
rect 13435 3350 13490 3470
rect 13610 3350 13655 3470
rect 13775 3350 13820 3470
rect 13940 3350 13985 3470
rect 14105 3350 14160 3470
rect 14280 3350 14325 3470
rect 14445 3350 14490 3470
rect 14610 3350 14655 3470
rect 14775 3350 14830 3470
rect 14950 3350 14995 3470
rect 15115 3350 15160 3470
rect 15280 3350 15325 3470
rect 15445 3350 15500 3470
rect 15620 3350 15665 3470
rect 15785 3350 15830 3470
rect 15950 3350 15995 3470
rect 16115 3350 16170 3470
rect 16290 3350 16335 3470
rect 16455 3350 16500 3470
rect 16620 3350 16665 3470
rect 16785 3350 16840 3470
rect 16960 3350 17005 3470
rect 17125 3350 17170 3470
rect 17290 3350 17335 3470
rect 17455 3350 17510 3470
rect 17630 3350 17675 3470
rect 17795 3350 17840 3470
rect 17960 3350 18005 3470
rect 18125 3350 18180 3470
rect 18300 3350 18325 3470
rect 12795 3305 18325 3350
rect 12795 3185 12820 3305
rect 12940 3185 12985 3305
rect 13105 3185 13150 3305
rect 13270 3185 13315 3305
rect 13435 3185 13490 3305
rect 13610 3185 13655 3305
rect 13775 3185 13820 3305
rect 13940 3185 13985 3305
rect 14105 3185 14160 3305
rect 14280 3185 14325 3305
rect 14445 3185 14490 3305
rect 14610 3185 14655 3305
rect 14775 3185 14830 3305
rect 14950 3185 14995 3305
rect 15115 3185 15160 3305
rect 15280 3185 15325 3305
rect 15445 3185 15500 3305
rect 15620 3185 15665 3305
rect 15785 3185 15830 3305
rect 15950 3185 15995 3305
rect 16115 3185 16170 3305
rect 16290 3185 16335 3305
rect 16455 3185 16500 3305
rect 16620 3185 16665 3305
rect 16785 3185 16840 3305
rect 16960 3185 17005 3305
rect 17125 3185 17170 3305
rect 17290 3185 17335 3305
rect 17455 3185 17510 3305
rect 17630 3185 17675 3305
rect 17795 3185 17840 3305
rect 17960 3185 18005 3305
rect 18125 3185 18180 3305
rect 18300 3185 18325 3305
rect 12795 3140 18325 3185
rect 12795 3020 12820 3140
rect 12940 3020 12985 3140
rect 13105 3020 13150 3140
rect 13270 3020 13315 3140
rect 13435 3020 13490 3140
rect 13610 3020 13655 3140
rect 13775 3020 13820 3140
rect 13940 3020 13985 3140
rect 14105 3020 14160 3140
rect 14280 3020 14325 3140
rect 14445 3020 14490 3140
rect 14610 3020 14655 3140
rect 14775 3020 14830 3140
rect 14950 3020 14995 3140
rect 15115 3020 15160 3140
rect 15280 3020 15325 3140
rect 15445 3020 15500 3140
rect 15620 3020 15665 3140
rect 15785 3020 15830 3140
rect 15950 3020 15995 3140
rect 16115 3020 16170 3140
rect 16290 3020 16335 3140
rect 16455 3020 16500 3140
rect 16620 3020 16665 3140
rect 16785 3020 16840 3140
rect 16960 3020 17005 3140
rect 17125 3020 17170 3140
rect 17290 3020 17335 3140
rect 17455 3020 17510 3140
rect 17630 3020 17675 3140
rect 17795 3020 17840 3140
rect 17960 3020 18005 3140
rect 18125 3020 18180 3140
rect 18300 3020 18325 3140
rect 12795 2965 18325 3020
rect 12795 2845 12820 2965
rect 12940 2845 12985 2965
rect 13105 2845 13150 2965
rect 13270 2845 13315 2965
rect 13435 2845 13490 2965
rect 13610 2845 13655 2965
rect 13775 2845 13820 2965
rect 13940 2845 13985 2965
rect 14105 2845 14160 2965
rect 14280 2845 14325 2965
rect 14445 2845 14490 2965
rect 14610 2845 14655 2965
rect 14775 2845 14830 2965
rect 14950 2845 14995 2965
rect 15115 2845 15160 2965
rect 15280 2845 15325 2965
rect 15445 2845 15500 2965
rect 15620 2845 15665 2965
rect 15785 2845 15830 2965
rect 15950 2845 15995 2965
rect 16115 2845 16170 2965
rect 16290 2845 16335 2965
rect 16455 2845 16500 2965
rect 16620 2845 16665 2965
rect 16785 2845 16840 2965
rect 16960 2845 17005 2965
rect 17125 2845 17170 2965
rect 17290 2845 17335 2965
rect 17455 2845 17510 2965
rect 17630 2845 17675 2965
rect 17795 2845 17840 2965
rect 17960 2845 18005 2965
rect 18125 2845 18180 2965
rect 18300 2845 18325 2965
rect 12795 2800 18325 2845
rect 12795 2680 12820 2800
rect 12940 2680 12985 2800
rect 13105 2680 13150 2800
rect 13270 2680 13315 2800
rect 13435 2680 13490 2800
rect 13610 2680 13655 2800
rect 13775 2680 13820 2800
rect 13940 2680 13985 2800
rect 14105 2680 14160 2800
rect 14280 2680 14325 2800
rect 14445 2680 14490 2800
rect 14610 2680 14655 2800
rect 14775 2680 14830 2800
rect 14950 2680 14995 2800
rect 15115 2680 15160 2800
rect 15280 2680 15325 2800
rect 15445 2680 15500 2800
rect 15620 2680 15665 2800
rect 15785 2680 15830 2800
rect 15950 2680 15995 2800
rect 16115 2680 16170 2800
rect 16290 2680 16335 2800
rect 16455 2680 16500 2800
rect 16620 2680 16665 2800
rect 16785 2680 16840 2800
rect 16960 2680 17005 2800
rect 17125 2680 17170 2800
rect 17290 2680 17335 2800
rect 17455 2680 17510 2800
rect 17630 2680 17675 2800
rect 17795 2680 17840 2800
rect 17960 2680 18005 2800
rect 18125 2680 18180 2800
rect 18300 2680 18325 2800
rect 12795 2635 18325 2680
rect 12795 2515 12820 2635
rect 12940 2515 12985 2635
rect 13105 2515 13150 2635
rect 13270 2515 13315 2635
rect 13435 2515 13490 2635
rect 13610 2515 13655 2635
rect 13775 2515 13820 2635
rect 13940 2515 13985 2635
rect 14105 2515 14160 2635
rect 14280 2515 14325 2635
rect 14445 2515 14490 2635
rect 14610 2515 14655 2635
rect 14775 2515 14830 2635
rect 14950 2515 14995 2635
rect 15115 2515 15160 2635
rect 15280 2515 15325 2635
rect 15445 2515 15500 2635
rect 15620 2515 15665 2635
rect 15785 2515 15830 2635
rect 15950 2515 15995 2635
rect 16115 2515 16170 2635
rect 16290 2515 16335 2635
rect 16455 2515 16500 2635
rect 16620 2515 16665 2635
rect 16785 2515 16840 2635
rect 16960 2515 17005 2635
rect 17125 2515 17170 2635
rect 17290 2515 17335 2635
rect 17455 2515 17510 2635
rect 17630 2515 17675 2635
rect 17795 2515 17840 2635
rect 17960 2515 18005 2635
rect 18125 2515 18180 2635
rect 18300 2515 18325 2635
rect 12795 2470 18325 2515
rect 12795 2350 12820 2470
rect 12940 2350 12985 2470
rect 13105 2350 13150 2470
rect 13270 2350 13315 2470
rect 13435 2350 13490 2470
rect 13610 2350 13655 2470
rect 13775 2350 13820 2470
rect 13940 2350 13985 2470
rect 14105 2350 14160 2470
rect 14280 2350 14325 2470
rect 14445 2350 14490 2470
rect 14610 2350 14655 2470
rect 14775 2350 14830 2470
rect 14950 2350 14995 2470
rect 15115 2350 15160 2470
rect 15280 2350 15325 2470
rect 15445 2350 15500 2470
rect 15620 2350 15665 2470
rect 15785 2350 15830 2470
rect 15950 2350 15995 2470
rect 16115 2350 16170 2470
rect 16290 2350 16335 2470
rect 16455 2350 16500 2470
rect 16620 2350 16665 2470
rect 16785 2350 16840 2470
rect 16960 2350 17005 2470
rect 17125 2350 17170 2470
rect 17290 2350 17335 2470
rect 17455 2350 17510 2470
rect 17630 2350 17675 2470
rect 17795 2350 17840 2470
rect 17960 2350 18005 2470
rect 18125 2350 18180 2470
rect 18300 2350 18325 2470
rect 12795 2295 18325 2350
rect 12795 2175 12820 2295
rect 12940 2175 12985 2295
rect 13105 2175 13150 2295
rect 13270 2175 13315 2295
rect 13435 2175 13490 2295
rect 13610 2175 13655 2295
rect 13775 2175 13820 2295
rect 13940 2175 13985 2295
rect 14105 2175 14160 2295
rect 14280 2175 14325 2295
rect 14445 2175 14490 2295
rect 14610 2175 14655 2295
rect 14775 2175 14830 2295
rect 14950 2175 14995 2295
rect 15115 2175 15160 2295
rect 15280 2175 15325 2295
rect 15445 2175 15500 2295
rect 15620 2175 15665 2295
rect 15785 2175 15830 2295
rect 15950 2175 15995 2295
rect 16115 2175 16170 2295
rect 16290 2175 16335 2295
rect 16455 2175 16500 2295
rect 16620 2175 16665 2295
rect 16785 2175 16840 2295
rect 16960 2175 17005 2295
rect 17125 2175 17170 2295
rect 17290 2175 17335 2295
rect 17455 2175 17510 2295
rect 17630 2175 17675 2295
rect 17795 2175 17840 2295
rect 17960 2175 18005 2295
rect 18125 2175 18180 2295
rect 18300 2175 18325 2295
rect 12795 2130 18325 2175
rect 12795 2010 12820 2130
rect 12940 2010 12985 2130
rect 13105 2010 13150 2130
rect 13270 2010 13315 2130
rect 13435 2010 13490 2130
rect 13610 2010 13655 2130
rect 13775 2010 13820 2130
rect 13940 2010 13985 2130
rect 14105 2010 14160 2130
rect 14280 2010 14325 2130
rect 14445 2010 14490 2130
rect 14610 2010 14655 2130
rect 14775 2010 14830 2130
rect 14950 2010 14995 2130
rect 15115 2010 15160 2130
rect 15280 2010 15325 2130
rect 15445 2010 15500 2130
rect 15620 2010 15665 2130
rect 15785 2010 15830 2130
rect 15950 2010 15995 2130
rect 16115 2010 16170 2130
rect 16290 2010 16335 2130
rect 16455 2010 16500 2130
rect 16620 2010 16665 2130
rect 16785 2010 16840 2130
rect 16960 2010 17005 2130
rect 17125 2010 17170 2130
rect 17290 2010 17335 2130
rect 17455 2010 17510 2130
rect 17630 2010 17675 2130
rect 17795 2010 17840 2130
rect 17960 2010 18005 2130
rect 18125 2010 18180 2130
rect 18300 2010 18325 2130
rect 12795 1965 18325 2010
rect 12795 1845 12820 1965
rect 12940 1845 12985 1965
rect 13105 1845 13150 1965
rect 13270 1845 13315 1965
rect 13435 1845 13490 1965
rect 13610 1845 13655 1965
rect 13775 1845 13820 1965
rect 13940 1845 13985 1965
rect 14105 1845 14160 1965
rect 14280 1845 14325 1965
rect 14445 1845 14490 1965
rect 14610 1845 14655 1965
rect 14775 1845 14830 1965
rect 14950 1845 14995 1965
rect 15115 1845 15160 1965
rect 15280 1845 15325 1965
rect 15445 1845 15500 1965
rect 15620 1845 15665 1965
rect 15785 1845 15830 1965
rect 15950 1845 15995 1965
rect 16115 1845 16170 1965
rect 16290 1845 16335 1965
rect 16455 1845 16500 1965
rect 16620 1845 16665 1965
rect 16785 1845 16840 1965
rect 16960 1845 17005 1965
rect 17125 1845 17170 1965
rect 17290 1845 17335 1965
rect 17455 1845 17510 1965
rect 17630 1845 17675 1965
rect 17795 1845 17840 1965
rect 17960 1845 18005 1965
rect 18125 1845 18180 1965
rect 18300 1845 18325 1965
rect 12795 1800 18325 1845
rect 12795 1680 12820 1800
rect 12940 1680 12985 1800
rect 13105 1680 13150 1800
rect 13270 1680 13315 1800
rect 13435 1680 13490 1800
rect 13610 1680 13655 1800
rect 13775 1680 13820 1800
rect 13940 1680 13985 1800
rect 14105 1680 14160 1800
rect 14280 1680 14325 1800
rect 14445 1680 14490 1800
rect 14610 1680 14655 1800
rect 14775 1680 14830 1800
rect 14950 1680 14995 1800
rect 15115 1680 15160 1800
rect 15280 1680 15325 1800
rect 15445 1680 15500 1800
rect 15620 1680 15665 1800
rect 15785 1680 15830 1800
rect 15950 1680 15995 1800
rect 16115 1680 16170 1800
rect 16290 1680 16335 1800
rect 16455 1680 16500 1800
rect 16620 1680 16665 1800
rect 16785 1680 16840 1800
rect 16960 1680 17005 1800
rect 17125 1680 17170 1800
rect 17290 1680 17335 1800
rect 17455 1680 17510 1800
rect 17630 1680 17675 1800
rect 17795 1680 17840 1800
rect 17960 1680 18005 1800
rect 18125 1680 18180 1800
rect 18300 1680 18325 1800
rect 12795 1655 18325 1680
rect 18485 7040 18510 7125
rect 18630 7040 18675 7160
rect 18795 7040 18840 7160
rect 18960 7040 19005 7160
rect 19125 7040 19180 7160
rect 19300 7040 19345 7160
rect 19465 7040 19510 7160
rect 19630 7040 19675 7160
rect 19795 7040 19850 7160
rect 19970 7040 20015 7160
rect 20135 7040 20180 7160
rect 20300 7040 20345 7160
rect 20465 7040 20520 7160
rect 20640 7040 20685 7160
rect 20805 7040 20850 7160
rect 20970 7040 21015 7160
rect 21135 7040 21190 7160
rect 21310 7040 21355 7160
rect 21475 7040 21520 7160
rect 21640 7040 21685 7160
rect 21805 7040 21860 7160
rect 21980 7040 22025 7160
rect 22145 7040 22190 7160
rect 22310 7040 22355 7160
rect 22475 7040 22530 7160
rect 22650 7040 22695 7160
rect 22815 7040 22860 7160
rect 22980 7040 23025 7160
rect 23145 7040 23200 7160
rect 23320 7040 23365 7160
rect 23485 7040 23530 7160
rect 23650 7040 23695 7160
rect 23815 7040 23870 7160
rect 23990 7125 24200 7160
rect 23990 7040 24015 7125
rect 18485 6985 24015 7040
rect 18485 6865 18510 6985
rect 18630 6865 18675 6985
rect 18795 6865 18840 6985
rect 18960 6865 19005 6985
rect 19125 6865 19180 6985
rect 19300 6865 19345 6985
rect 19465 6865 19510 6985
rect 19630 6865 19675 6985
rect 19795 6865 19850 6985
rect 19970 6865 20015 6985
rect 20135 6865 20180 6985
rect 20300 6865 20345 6985
rect 20465 6865 20520 6985
rect 20640 6865 20685 6985
rect 20805 6865 20850 6985
rect 20970 6865 21015 6985
rect 21135 6865 21190 6985
rect 21310 6865 21355 6985
rect 21475 6865 21520 6985
rect 21640 6865 21685 6985
rect 21805 6865 21860 6985
rect 21980 6865 22025 6985
rect 22145 6865 22190 6985
rect 22310 6865 22355 6985
rect 22475 6865 22530 6985
rect 22650 6865 22695 6985
rect 22815 6865 22860 6985
rect 22980 6865 23025 6985
rect 23145 6865 23200 6985
rect 23320 6865 23365 6985
rect 23485 6865 23530 6985
rect 23650 6865 23695 6985
rect 23815 6865 23870 6985
rect 23990 6865 24015 6985
rect 18485 6820 24015 6865
rect 18485 6700 18510 6820
rect 18630 6700 18675 6820
rect 18795 6700 18840 6820
rect 18960 6700 19005 6820
rect 19125 6700 19180 6820
rect 19300 6700 19345 6820
rect 19465 6700 19510 6820
rect 19630 6700 19675 6820
rect 19795 6700 19850 6820
rect 19970 6700 20015 6820
rect 20135 6700 20180 6820
rect 20300 6700 20345 6820
rect 20465 6700 20520 6820
rect 20640 6700 20685 6820
rect 20805 6700 20850 6820
rect 20970 6700 21015 6820
rect 21135 6700 21190 6820
rect 21310 6700 21355 6820
rect 21475 6700 21520 6820
rect 21640 6700 21685 6820
rect 21805 6700 21860 6820
rect 21980 6700 22025 6820
rect 22145 6700 22190 6820
rect 22310 6700 22355 6820
rect 22475 6700 22530 6820
rect 22650 6700 22695 6820
rect 22815 6700 22860 6820
rect 22980 6700 23025 6820
rect 23145 6700 23200 6820
rect 23320 6700 23365 6820
rect 23485 6700 23530 6820
rect 23650 6700 23695 6820
rect 23815 6700 23870 6820
rect 23990 6700 24015 6820
rect 18485 6655 24015 6700
rect 18485 6535 18510 6655
rect 18630 6535 18675 6655
rect 18795 6535 18840 6655
rect 18960 6535 19005 6655
rect 19125 6535 19180 6655
rect 19300 6535 19345 6655
rect 19465 6535 19510 6655
rect 19630 6535 19675 6655
rect 19795 6535 19850 6655
rect 19970 6535 20015 6655
rect 20135 6535 20180 6655
rect 20300 6535 20345 6655
rect 20465 6535 20520 6655
rect 20640 6535 20685 6655
rect 20805 6535 20850 6655
rect 20970 6535 21015 6655
rect 21135 6535 21190 6655
rect 21310 6535 21355 6655
rect 21475 6535 21520 6655
rect 21640 6535 21685 6655
rect 21805 6535 21860 6655
rect 21980 6535 22025 6655
rect 22145 6535 22190 6655
rect 22310 6535 22355 6655
rect 22475 6535 22530 6655
rect 22650 6535 22695 6655
rect 22815 6535 22860 6655
rect 22980 6535 23025 6655
rect 23145 6535 23200 6655
rect 23320 6535 23365 6655
rect 23485 6535 23530 6655
rect 23650 6535 23695 6655
rect 23815 6535 23870 6655
rect 23990 6535 24015 6655
rect 18485 6490 24015 6535
rect 18485 6370 18510 6490
rect 18630 6370 18675 6490
rect 18795 6370 18840 6490
rect 18960 6370 19005 6490
rect 19125 6370 19180 6490
rect 19300 6370 19345 6490
rect 19465 6370 19510 6490
rect 19630 6370 19675 6490
rect 19795 6370 19850 6490
rect 19970 6370 20015 6490
rect 20135 6370 20180 6490
rect 20300 6370 20345 6490
rect 20465 6370 20520 6490
rect 20640 6370 20685 6490
rect 20805 6370 20850 6490
rect 20970 6370 21015 6490
rect 21135 6370 21190 6490
rect 21310 6370 21355 6490
rect 21475 6370 21520 6490
rect 21640 6370 21685 6490
rect 21805 6370 21860 6490
rect 21980 6370 22025 6490
rect 22145 6370 22190 6490
rect 22310 6370 22355 6490
rect 22475 6370 22530 6490
rect 22650 6370 22695 6490
rect 22815 6370 22860 6490
rect 22980 6370 23025 6490
rect 23145 6370 23200 6490
rect 23320 6370 23365 6490
rect 23485 6370 23530 6490
rect 23650 6370 23695 6490
rect 23815 6370 23870 6490
rect 23990 6370 24015 6490
rect 18485 6315 24015 6370
rect 18485 6195 18510 6315
rect 18630 6195 18675 6315
rect 18795 6195 18840 6315
rect 18960 6195 19005 6315
rect 19125 6195 19180 6315
rect 19300 6195 19345 6315
rect 19465 6195 19510 6315
rect 19630 6195 19675 6315
rect 19795 6195 19850 6315
rect 19970 6195 20015 6315
rect 20135 6195 20180 6315
rect 20300 6195 20345 6315
rect 20465 6195 20520 6315
rect 20640 6195 20685 6315
rect 20805 6195 20850 6315
rect 20970 6195 21015 6315
rect 21135 6195 21190 6315
rect 21310 6195 21355 6315
rect 21475 6195 21520 6315
rect 21640 6195 21685 6315
rect 21805 6195 21860 6315
rect 21980 6195 22025 6315
rect 22145 6195 22190 6315
rect 22310 6195 22355 6315
rect 22475 6195 22530 6315
rect 22650 6195 22695 6315
rect 22815 6195 22860 6315
rect 22980 6195 23025 6315
rect 23145 6195 23200 6315
rect 23320 6195 23365 6315
rect 23485 6195 23530 6315
rect 23650 6195 23695 6315
rect 23815 6195 23870 6315
rect 23990 6195 24015 6315
rect 18485 6150 24015 6195
rect 18485 6030 18510 6150
rect 18630 6030 18675 6150
rect 18795 6030 18840 6150
rect 18960 6030 19005 6150
rect 19125 6030 19180 6150
rect 19300 6030 19345 6150
rect 19465 6030 19510 6150
rect 19630 6030 19675 6150
rect 19795 6030 19850 6150
rect 19970 6030 20015 6150
rect 20135 6030 20180 6150
rect 20300 6030 20345 6150
rect 20465 6030 20520 6150
rect 20640 6030 20685 6150
rect 20805 6030 20850 6150
rect 20970 6030 21015 6150
rect 21135 6030 21190 6150
rect 21310 6030 21355 6150
rect 21475 6030 21520 6150
rect 21640 6030 21685 6150
rect 21805 6030 21860 6150
rect 21980 6030 22025 6150
rect 22145 6030 22190 6150
rect 22310 6030 22355 6150
rect 22475 6030 22530 6150
rect 22650 6030 22695 6150
rect 22815 6030 22860 6150
rect 22980 6030 23025 6150
rect 23145 6030 23200 6150
rect 23320 6030 23365 6150
rect 23485 6030 23530 6150
rect 23650 6030 23695 6150
rect 23815 6030 23870 6150
rect 23990 6030 24015 6150
rect 18485 5985 24015 6030
rect 18485 5865 18510 5985
rect 18630 5865 18675 5985
rect 18795 5865 18840 5985
rect 18960 5865 19005 5985
rect 19125 5865 19180 5985
rect 19300 5865 19345 5985
rect 19465 5865 19510 5985
rect 19630 5865 19675 5985
rect 19795 5865 19850 5985
rect 19970 5865 20015 5985
rect 20135 5865 20180 5985
rect 20300 5865 20345 5985
rect 20465 5865 20520 5985
rect 20640 5865 20685 5985
rect 20805 5865 20850 5985
rect 20970 5865 21015 5985
rect 21135 5865 21190 5985
rect 21310 5865 21355 5985
rect 21475 5865 21520 5985
rect 21640 5865 21685 5985
rect 21805 5865 21860 5985
rect 21980 5865 22025 5985
rect 22145 5865 22190 5985
rect 22310 5865 22355 5985
rect 22475 5865 22530 5985
rect 22650 5865 22695 5985
rect 22815 5865 22860 5985
rect 22980 5865 23025 5985
rect 23145 5865 23200 5985
rect 23320 5865 23365 5985
rect 23485 5865 23530 5985
rect 23650 5865 23695 5985
rect 23815 5865 23870 5985
rect 23990 5865 24015 5985
rect 18485 5820 24015 5865
rect 18485 5700 18510 5820
rect 18630 5700 18675 5820
rect 18795 5700 18840 5820
rect 18960 5700 19005 5820
rect 19125 5700 19180 5820
rect 19300 5700 19345 5820
rect 19465 5700 19510 5820
rect 19630 5700 19675 5820
rect 19795 5700 19850 5820
rect 19970 5700 20015 5820
rect 20135 5700 20180 5820
rect 20300 5700 20345 5820
rect 20465 5700 20520 5820
rect 20640 5700 20685 5820
rect 20805 5700 20850 5820
rect 20970 5700 21015 5820
rect 21135 5700 21190 5820
rect 21310 5700 21355 5820
rect 21475 5700 21520 5820
rect 21640 5700 21685 5820
rect 21805 5700 21860 5820
rect 21980 5700 22025 5820
rect 22145 5700 22190 5820
rect 22310 5700 22355 5820
rect 22475 5700 22530 5820
rect 22650 5700 22695 5820
rect 22815 5700 22860 5820
rect 22980 5700 23025 5820
rect 23145 5700 23200 5820
rect 23320 5700 23365 5820
rect 23485 5700 23530 5820
rect 23650 5700 23695 5820
rect 23815 5700 23870 5820
rect 23990 5700 24015 5820
rect 18485 5645 24015 5700
rect 18485 5525 18510 5645
rect 18630 5525 18675 5645
rect 18795 5525 18840 5645
rect 18960 5525 19005 5645
rect 19125 5525 19180 5645
rect 19300 5525 19345 5645
rect 19465 5525 19510 5645
rect 19630 5525 19675 5645
rect 19795 5525 19850 5645
rect 19970 5525 20015 5645
rect 20135 5525 20180 5645
rect 20300 5525 20345 5645
rect 20465 5525 20520 5645
rect 20640 5525 20685 5645
rect 20805 5525 20850 5645
rect 20970 5525 21015 5645
rect 21135 5525 21190 5645
rect 21310 5525 21355 5645
rect 21475 5525 21520 5645
rect 21640 5525 21685 5645
rect 21805 5525 21860 5645
rect 21980 5525 22025 5645
rect 22145 5525 22190 5645
rect 22310 5525 22355 5645
rect 22475 5525 22530 5645
rect 22650 5525 22695 5645
rect 22815 5525 22860 5645
rect 22980 5525 23025 5645
rect 23145 5525 23200 5645
rect 23320 5525 23365 5645
rect 23485 5525 23530 5645
rect 23650 5525 23695 5645
rect 23815 5525 23870 5645
rect 23990 5525 24015 5645
rect 18485 5480 24015 5525
rect 18485 5360 18510 5480
rect 18630 5360 18675 5480
rect 18795 5360 18840 5480
rect 18960 5360 19005 5480
rect 19125 5360 19180 5480
rect 19300 5360 19345 5480
rect 19465 5360 19510 5480
rect 19630 5360 19675 5480
rect 19795 5360 19850 5480
rect 19970 5360 20015 5480
rect 20135 5360 20180 5480
rect 20300 5360 20345 5480
rect 20465 5360 20520 5480
rect 20640 5360 20685 5480
rect 20805 5360 20850 5480
rect 20970 5360 21015 5480
rect 21135 5360 21190 5480
rect 21310 5360 21355 5480
rect 21475 5360 21520 5480
rect 21640 5360 21685 5480
rect 21805 5360 21860 5480
rect 21980 5360 22025 5480
rect 22145 5360 22190 5480
rect 22310 5360 22355 5480
rect 22475 5360 22530 5480
rect 22650 5360 22695 5480
rect 22815 5360 22860 5480
rect 22980 5360 23025 5480
rect 23145 5360 23200 5480
rect 23320 5360 23365 5480
rect 23485 5360 23530 5480
rect 23650 5360 23695 5480
rect 23815 5360 23870 5480
rect 23990 5360 24015 5480
rect 18485 5315 24015 5360
rect 18485 5195 18510 5315
rect 18630 5195 18675 5315
rect 18795 5195 18840 5315
rect 18960 5195 19005 5315
rect 19125 5195 19180 5315
rect 19300 5195 19345 5315
rect 19465 5195 19510 5315
rect 19630 5195 19675 5315
rect 19795 5195 19850 5315
rect 19970 5195 20015 5315
rect 20135 5195 20180 5315
rect 20300 5195 20345 5315
rect 20465 5195 20520 5315
rect 20640 5195 20685 5315
rect 20805 5195 20850 5315
rect 20970 5195 21015 5315
rect 21135 5195 21190 5315
rect 21310 5195 21355 5315
rect 21475 5195 21520 5315
rect 21640 5195 21685 5315
rect 21805 5195 21860 5315
rect 21980 5195 22025 5315
rect 22145 5195 22190 5315
rect 22310 5195 22355 5315
rect 22475 5195 22530 5315
rect 22650 5195 22695 5315
rect 22815 5195 22860 5315
rect 22980 5195 23025 5315
rect 23145 5195 23200 5315
rect 23320 5195 23365 5315
rect 23485 5195 23530 5315
rect 23650 5195 23695 5315
rect 23815 5195 23870 5315
rect 23990 5195 24015 5315
rect 18485 5150 24015 5195
rect 18485 5030 18510 5150
rect 18630 5030 18675 5150
rect 18795 5030 18840 5150
rect 18960 5030 19005 5150
rect 19125 5030 19180 5150
rect 19300 5030 19345 5150
rect 19465 5030 19510 5150
rect 19630 5030 19675 5150
rect 19795 5030 19850 5150
rect 19970 5030 20015 5150
rect 20135 5030 20180 5150
rect 20300 5030 20345 5150
rect 20465 5030 20520 5150
rect 20640 5030 20685 5150
rect 20805 5030 20850 5150
rect 20970 5030 21015 5150
rect 21135 5030 21190 5150
rect 21310 5030 21355 5150
rect 21475 5030 21520 5150
rect 21640 5030 21685 5150
rect 21805 5030 21860 5150
rect 21980 5030 22025 5150
rect 22145 5030 22190 5150
rect 22310 5030 22355 5150
rect 22475 5030 22530 5150
rect 22650 5030 22695 5150
rect 22815 5030 22860 5150
rect 22980 5030 23025 5150
rect 23145 5030 23200 5150
rect 23320 5030 23365 5150
rect 23485 5030 23530 5150
rect 23650 5030 23695 5150
rect 23815 5030 23870 5150
rect 23990 5030 24015 5150
rect 18485 4975 24015 5030
rect 18485 4855 18510 4975
rect 18630 4855 18675 4975
rect 18795 4855 18840 4975
rect 18960 4855 19005 4975
rect 19125 4855 19180 4975
rect 19300 4855 19345 4975
rect 19465 4855 19510 4975
rect 19630 4855 19675 4975
rect 19795 4855 19850 4975
rect 19970 4855 20015 4975
rect 20135 4855 20180 4975
rect 20300 4855 20345 4975
rect 20465 4855 20520 4975
rect 20640 4855 20685 4975
rect 20805 4855 20850 4975
rect 20970 4855 21015 4975
rect 21135 4855 21190 4975
rect 21310 4855 21355 4975
rect 21475 4855 21520 4975
rect 21640 4855 21685 4975
rect 21805 4855 21860 4975
rect 21980 4855 22025 4975
rect 22145 4855 22190 4975
rect 22310 4855 22355 4975
rect 22475 4855 22530 4975
rect 22650 4855 22695 4975
rect 22815 4855 22860 4975
rect 22980 4855 23025 4975
rect 23145 4855 23200 4975
rect 23320 4855 23365 4975
rect 23485 4855 23530 4975
rect 23650 4855 23695 4975
rect 23815 4855 23870 4975
rect 23990 4855 24015 4975
rect 18485 4810 24015 4855
rect 18485 4690 18510 4810
rect 18630 4690 18675 4810
rect 18795 4690 18840 4810
rect 18960 4690 19005 4810
rect 19125 4690 19180 4810
rect 19300 4690 19345 4810
rect 19465 4690 19510 4810
rect 19630 4690 19675 4810
rect 19795 4690 19850 4810
rect 19970 4690 20015 4810
rect 20135 4690 20180 4810
rect 20300 4690 20345 4810
rect 20465 4690 20520 4810
rect 20640 4690 20685 4810
rect 20805 4690 20850 4810
rect 20970 4690 21015 4810
rect 21135 4690 21190 4810
rect 21310 4690 21355 4810
rect 21475 4690 21520 4810
rect 21640 4690 21685 4810
rect 21805 4690 21860 4810
rect 21980 4690 22025 4810
rect 22145 4690 22190 4810
rect 22310 4690 22355 4810
rect 22475 4690 22530 4810
rect 22650 4690 22695 4810
rect 22815 4690 22860 4810
rect 22980 4690 23025 4810
rect 23145 4690 23200 4810
rect 23320 4690 23365 4810
rect 23485 4690 23530 4810
rect 23650 4690 23695 4810
rect 23815 4690 23870 4810
rect 23990 4690 24015 4810
rect 18485 4645 24015 4690
rect 18485 4525 18510 4645
rect 18630 4525 18675 4645
rect 18795 4525 18840 4645
rect 18960 4525 19005 4645
rect 19125 4525 19180 4645
rect 19300 4525 19345 4645
rect 19465 4525 19510 4645
rect 19630 4525 19675 4645
rect 19795 4525 19850 4645
rect 19970 4525 20015 4645
rect 20135 4525 20180 4645
rect 20300 4525 20345 4645
rect 20465 4525 20520 4645
rect 20640 4525 20685 4645
rect 20805 4525 20850 4645
rect 20970 4525 21015 4645
rect 21135 4525 21190 4645
rect 21310 4525 21355 4645
rect 21475 4525 21520 4645
rect 21640 4525 21685 4645
rect 21805 4525 21860 4645
rect 21980 4525 22025 4645
rect 22145 4525 22190 4645
rect 22310 4525 22355 4645
rect 22475 4525 22530 4645
rect 22650 4525 22695 4645
rect 22815 4525 22860 4645
rect 22980 4525 23025 4645
rect 23145 4525 23200 4645
rect 23320 4525 23365 4645
rect 23485 4525 23530 4645
rect 23650 4525 23695 4645
rect 23815 4525 23870 4645
rect 23990 4525 24015 4645
rect 18485 4480 24015 4525
rect 18485 4360 18510 4480
rect 18630 4360 18675 4480
rect 18795 4360 18840 4480
rect 18960 4360 19005 4480
rect 19125 4360 19180 4480
rect 19300 4360 19345 4480
rect 19465 4360 19510 4480
rect 19630 4360 19675 4480
rect 19795 4360 19850 4480
rect 19970 4360 20015 4480
rect 20135 4360 20180 4480
rect 20300 4360 20345 4480
rect 20465 4360 20520 4480
rect 20640 4360 20685 4480
rect 20805 4360 20850 4480
rect 20970 4360 21015 4480
rect 21135 4360 21190 4480
rect 21310 4360 21355 4480
rect 21475 4360 21520 4480
rect 21640 4360 21685 4480
rect 21805 4360 21860 4480
rect 21980 4360 22025 4480
rect 22145 4360 22190 4480
rect 22310 4360 22355 4480
rect 22475 4360 22530 4480
rect 22650 4360 22695 4480
rect 22815 4360 22860 4480
rect 22980 4360 23025 4480
rect 23145 4360 23200 4480
rect 23320 4360 23365 4480
rect 23485 4360 23530 4480
rect 23650 4360 23695 4480
rect 23815 4360 23870 4480
rect 23990 4360 24015 4480
rect 18485 4305 24015 4360
rect 18485 4185 18510 4305
rect 18630 4185 18675 4305
rect 18795 4185 18840 4305
rect 18960 4185 19005 4305
rect 19125 4185 19180 4305
rect 19300 4185 19345 4305
rect 19465 4185 19510 4305
rect 19630 4185 19675 4305
rect 19795 4185 19850 4305
rect 19970 4185 20015 4305
rect 20135 4185 20180 4305
rect 20300 4185 20345 4305
rect 20465 4185 20520 4305
rect 20640 4185 20685 4305
rect 20805 4185 20850 4305
rect 20970 4185 21015 4305
rect 21135 4185 21190 4305
rect 21310 4185 21355 4305
rect 21475 4185 21520 4305
rect 21640 4185 21685 4305
rect 21805 4185 21860 4305
rect 21980 4185 22025 4305
rect 22145 4185 22190 4305
rect 22310 4185 22355 4305
rect 22475 4185 22530 4305
rect 22650 4185 22695 4305
rect 22815 4185 22860 4305
rect 22980 4185 23025 4305
rect 23145 4185 23200 4305
rect 23320 4185 23365 4305
rect 23485 4185 23530 4305
rect 23650 4185 23695 4305
rect 23815 4185 23870 4305
rect 23990 4185 24015 4305
rect 18485 4140 24015 4185
rect 18485 4020 18510 4140
rect 18630 4020 18675 4140
rect 18795 4020 18840 4140
rect 18960 4020 19005 4140
rect 19125 4020 19180 4140
rect 19300 4020 19345 4140
rect 19465 4020 19510 4140
rect 19630 4020 19675 4140
rect 19795 4020 19850 4140
rect 19970 4020 20015 4140
rect 20135 4020 20180 4140
rect 20300 4020 20345 4140
rect 20465 4020 20520 4140
rect 20640 4020 20685 4140
rect 20805 4020 20850 4140
rect 20970 4020 21015 4140
rect 21135 4020 21190 4140
rect 21310 4020 21355 4140
rect 21475 4020 21520 4140
rect 21640 4020 21685 4140
rect 21805 4020 21860 4140
rect 21980 4020 22025 4140
rect 22145 4020 22190 4140
rect 22310 4020 22355 4140
rect 22475 4020 22530 4140
rect 22650 4020 22695 4140
rect 22815 4020 22860 4140
rect 22980 4020 23025 4140
rect 23145 4020 23200 4140
rect 23320 4020 23365 4140
rect 23485 4020 23530 4140
rect 23650 4020 23695 4140
rect 23815 4020 23870 4140
rect 23990 4020 24015 4140
rect 18485 3975 24015 4020
rect 18485 3855 18510 3975
rect 18630 3855 18675 3975
rect 18795 3855 18840 3975
rect 18960 3855 19005 3975
rect 19125 3855 19180 3975
rect 19300 3855 19345 3975
rect 19465 3855 19510 3975
rect 19630 3855 19675 3975
rect 19795 3855 19850 3975
rect 19970 3855 20015 3975
rect 20135 3855 20180 3975
rect 20300 3855 20345 3975
rect 20465 3855 20520 3975
rect 20640 3855 20685 3975
rect 20805 3855 20850 3975
rect 20970 3855 21015 3975
rect 21135 3855 21190 3975
rect 21310 3855 21355 3975
rect 21475 3855 21520 3975
rect 21640 3855 21685 3975
rect 21805 3855 21860 3975
rect 21980 3855 22025 3975
rect 22145 3855 22190 3975
rect 22310 3855 22355 3975
rect 22475 3855 22530 3975
rect 22650 3855 22695 3975
rect 22815 3855 22860 3975
rect 22980 3855 23025 3975
rect 23145 3855 23200 3975
rect 23320 3855 23365 3975
rect 23485 3855 23530 3975
rect 23650 3855 23695 3975
rect 23815 3855 23870 3975
rect 23990 3855 24015 3975
rect 18485 3810 24015 3855
rect 18485 3690 18510 3810
rect 18630 3690 18675 3810
rect 18795 3690 18840 3810
rect 18960 3690 19005 3810
rect 19125 3690 19180 3810
rect 19300 3690 19345 3810
rect 19465 3690 19510 3810
rect 19630 3690 19675 3810
rect 19795 3690 19850 3810
rect 19970 3690 20015 3810
rect 20135 3690 20180 3810
rect 20300 3690 20345 3810
rect 20465 3690 20520 3810
rect 20640 3690 20685 3810
rect 20805 3690 20850 3810
rect 20970 3690 21015 3810
rect 21135 3690 21190 3810
rect 21310 3690 21355 3810
rect 21475 3690 21520 3810
rect 21640 3690 21685 3810
rect 21805 3690 21860 3810
rect 21980 3690 22025 3810
rect 22145 3690 22190 3810
rect 22310 3690 22355 3810
rect 22475 3690 22530 3810
rect 22650 3690 22695 3810
rect 22815 3690 22860 3810
rect 22980 3690 23025 3810
rect 23145 3690 23200 3810
rect 23320 3690 23365 3810
rect 23485 3690 23530 3810
rect 23650 3690 23695 3810
rect 23815 3690 23870 3810
rect 23990 3690 24015 3810
rect 18485 3635 24015 3690
rect 18485 3515 18510 3635
rect 18630 3515 18675 3635
rect 18795 3515 18840 3635
rect 18960 3515 19005 3635
rect 19125 3515 19180 3635
rect 19300 3515 19345 3635
rect 19465 3515 19510 3635
rect 19630 3515 19675 3635
rect 19795 3515 19850 3635
rect 19970 3515 20015 3635
rect 20135 3515 20180 3635
rect 20300 3515 20345 3635
rect 20465 3515 20520 3635
rect 20640 3515 20685 3635
rect 20805 3515 20850 3635
rect 20970 3515 21015 3635
rect 21135 3515 21190 3635
rect 21310 3515 21355 3635
rect 21475 3515 21520 3635
rect 21640 3515 21685 3635
rect 21805 3515 21860 3635
rect 21980 3515 22025 3635
rect 22145 3515 22190 3635
rect 22310 3515 22355 3635
rect 22475 3515 22530 3635
rect 22650 3515 22695 3635
rect 22815 3515 22860 3635
rect 22980 3515 23025 3635
rect 23145 3515 23200 3635
rect 23320 3515 23365 3635
rect 23485 3515 23530 3635
rect 23650 3515 23695 3635
rect 23815 3515 23870 3635
rect 23990 3515 24015 3635
rect 18485 3470 24015 3515
rect 18485 3350 18510 3470
rect 18630 3350 18675 3470
rect 18795 3350 18840 3470
rect 18960 3350 19005 3470
rect 19125 3350 19180 3470
rect 19300 3350 19345 3470
rect 19465 3350 19510 3470
rect 19630 3350 19675 3470
rect 19795 3350 19850 3470
rect 19970 3350 20015 3470
rect 20135 3350 20180 3470
rect 20300 3350 20345 3470
rect 20465 3350 20520 3470
rect 20640 3350 20685 3470
rect 20805 3350 20850 3470
rect 20970 3350 21015 3470
rect 21135 3350 21190 3470
rect 21310 3350 21355 3470
rect 21475 3350 21520 3470
rect 21640 3350 21685 3470
rect 21805 3350 21860 3470
rect 21980 3350 22025 3470
rect 22145 3350 22190 3470
rect 22310 3350 22355 3470
rect 22475 3350 22530 3470
rect 22650 3350 22695 3470
rect 22815 3350 22860 3470
rect 22980 3350 23025 3470
rect 23145 3350 23200 3470
rect 23320 3350 23365 3470
rect 23485 3350 23530 3470
rect 23650 3350 23695 3470
rect 23815 3350 23870 3470
rect 23990 3350 24015 3470
rect 18485 3305 24015 3350
rect 18485 3185 18510 3305
rect 18630 3185 18675 3305
rect 18795 3185 18840 3305
rect 18960 3185 19005 3305
rect 19125 3185 19180 3305
rect 19300 3185 19345 3305
rect 19465 3185 19510 3305
rect 19630 3185 19675 3305
rect 19795 3185 19850 3305
rect 19970 3185 20015 3305
rect 20135 3185 20180 3305
rect 20300 3185 20345 3305
rect 20465 3185 20520 3305
rect 20640 3185 20685 3305
rect 20805 3185 20850 3305
rect 20970 3185 21015 3305
rect 21135 3185 21190 3305
rect 21310 3185 21355 3305
rect 21475 3185 21520 3305
rect 21640 3185 21685 3305
rect 21805 3185 21860 3305
rect 21980 3185 22025 3305
rect 22145 3185 22190 3305
rect 22310 3185 22355 3305
rect 22475 3185 22530 3305
rect 22650 3185 22695 3305
rect 22815 3185 22860 3305
rect 22980 3185 23025 3305
rect 23145 3185 23200 3305
rect 23320 3185 23365 3305
rect 23485 3185 23530 3305
rect 23650 3185 23695 3305
rect 23815 3185 23870 3305
rect 23990 3185 24015 3305
rect 18485 3140 24015 3185
rect 18485 3020 18510 3140
rect 18630 3020 18675 3140
rect 18795 3020 18840 3140
rect 18960 3020 19005 3140
rect 19125 3020 19180 3140
rect 19300 3020 19345 3140
rect 19465 3020 19510 3140
rect 19630 3020 19675 3140
rect 19795 3020 19850 3140
rect 19970 3020 20015 3140
rect 20135 3020 20180 3140
rect 20300 3020 20345 3140
rect 20465 3020 20520 3140
rect 20640 3020 20685 3140
rect 20805 3020 20850 3140
rect 20970 3020 21015 3140
rect 21135 3020 21190 3140
rect 21310 3020 21355 3140
rect 21475 3020 21520 3140
rect 21640 3020 21685 3140
rect 21805 3020 21860 3140
rect 21980 3020 22025 3140
rect 22145 3020 22190 3140
rect 22310 3020 22355 3140
rect 22475 3020 22530 3140
rect 22650 3020 22695 3140
rect 22815 3020 22860 3140
rect 22980 3020 23025 3140
rect 23145 3020 23200 3140
rect 23320 3020 23365 3140
rect 23485 3020 23530 3140
rect 23650 3020 23695 3140
rect 23815 3020 23870 3140
rect 23990 3020 24015 3140
rect 18485 2965 24015 3020
rect 18485 2845 18510 2965
rect 18630 2845 18675 2965
rect 18795 2845 18840 2965
rect 18960 2845 19005 2965
rect 19125 2845 19180 2965
rect 19300 2845 19345 2965
rect 19465 2845 19510 2965
rect 19630 2845 19675 2965
rect 19795 2845 19850 2965
rect 19970 2845 20015 2965
rect 20135 2845 20180 2965
rect 20300 2845 20345 2965
rect 20465 2845 20520 2965
rect 20640 2845 20685 2965
rect 20805 2845 20850 2965
rect 20970 2845 21015 2965
rect 21135 2845 21190 2965
rect 21310 2845 21355 2965
rect 21475 2845 21520 2965
rect 21640 2845 21685 2965
rect 21805 2845 21860 2965
rect 21980 2845 22025 2965
rect 22145 2845 22190 2965
rect 22310 2845 22355 2965
rect 22475 2845 22530 2965
rect 22650 2845 22695 2965
rect 22815 2845 22860 2965
rect 22980 2845 23025 2965
rect 23145 2845 23200 2965
rect 23320 2845 23365 2965
rect 23485 2845 23530 2965
rect 23650 2845 23695 2965
rect 23815 2845 23870 2965
rect 23990 2845 24015 2965
rect 18485 2800 24015 2845
rect 18485 2680 18510 2800
rect 18630 2680 18675 2800
rect 18795 2680 18840 2800
rect 18960 2680 19005 2800
rect 19125 2680 19180 2800
rect 19300 2680 19345 2800
rect 19465 2680 19510 2800
rect 19630 2680 19675 2800
rect 19795 2680 19850 2800
rect 19970 2680 20015 2800
rect 20135 2680 20180 2800
rect 20300 2680 20345 2800
rect 20465 2680 20520 2800
rect 20640 2680 20685 2800
rect 20805 2680 20850 2800
rect 20970 2680 21015 2800
rect 21135 2680 21190 2800
rect 21310 2680 21355 2800
rect 21475 2680 21520 2800
rect 21640 2680 21685 2800
rect 21805 2680 21860 2800
rect 21980 2680 22025 2800
rect 22145 2680 22190 2800
rect 22310 2680 22355 2800
rect 22475 2680 22530 2800
rect 22650 2680 22695 2800
rect 22815 2680 22860 2800
rect 22980 2680 23025 2800
rect 23145 2680 23200 2800
rect 23320 2680 23365 2800
rect 23485 2680 23530 2800
rect 23650 2680 23695 2800
rect 23815 2680 23870 2800
rect 23990 2680 24015 2800
rect 18485 2635 24015 2680
rect 18485 2515 18510 2635
rect 18630 2515 18675 2635
rect 18795 2515 18840 2635
rect 18960 2515 19005 2635
rect 19125 2515 19180 2635
rect 19300 2515 19345 2635
rect 19465 2515 19510 2635
rect 19630 2515 19675 2635
rect 19795 2515 19850 2635
rect 19970 2515 20015 2635
rect 20135 2515 20180 2635
rect 20300 2515 20345 2635
rect 20465 2515 20520 2635
rect 20640 2515 20685 2635
rect 20805 2515 20850 2635
rect 20970 2515 21015 2635
rect 21135 2515 21190 2635
rect 21310 2515 21355 2635
rect 21475 2515 21520 2635
rect 21640 2515 21685 2635
rect 21805 2515 21860 2635
rect 21980 2515 22025 2635
rect 22145 2515 22190 2635
rect 22310 2515 22355 2635
rect 22475 2515 22530 2635
rect 22650 2515 22695 2635
rect 22815 2515 22860 2635
rect 22980 2515 23025 2635
rect 23145 2515 23200 2635
rect 23320 2515 23365 2635
rect 23485 2515 23530 2635
rect 23650 2515 23695 2635
rect 23815 2515 23870 2635
rect 23990 2515 24015 2635
rect 18485 2470 24015 2515
rect 18485 2350 18510 2470
rect 18630 2350 18675 2470
rect 18795 2350 18840 2470
rect 18960 2350 19005 2470
rect 19125 2350 19180 2470
rect 19300 2350 19345 2470
rect 19465 2350 19510 2470
rect 19630 2350 19675 2470
rect 19795 2350 19850 2470
rect 19970 2350 20015 2470
rect 20135 2350 20180 2470
rect 20300 2350 20345 2470
rect 20465 2350 20520 2470
rect 20640 2350 20685 2470
rect 20805 2350 20850 2470
rect 20970 2350 21015 2470
rect 21135 2350 21190 2470
rect 21310 2350 21355 2470
rect 21475 2350 21520 2470
rect 21640 2350 21685 2470
rect 21805 2350 21860 2470
rect 21980 2350 22025 2470
rect 22145 2350 22190 2470
rect 22310 2350 22355 2470
rect 22475 2350 22530 2470
rect 22650 2350 22695 2470
rect 22815 2350 22860 2470
rect 22980 2350 23025 2470
rect 23145 2350 23200 2470
rect 23320 2350 23365 2470
rect 23485 2350 23530 2470
rect 23650 2350 23695 2470
rect 23815 2350 23870 2470
rect 23990 2350 24015 2470
rect 18485 2295 24015 2350
rect 18485 2175 18510 2295
rect 18630 2175 18675 2295
rect 18795 2175 18840 2295
rect 18960 2175 19005 2295
rect 19125 2175 19180 2295
rect 19300 2175 19345 2295
rect 19465 2175 19510 2295
rect 19630 2175 19675 2295
rect 19795 2175 19850 2295
rect 19970 2175 20015 2295
rect 20135 2175 20180 2295
rect 20300 2175 20345 2295
rect 20465 2175 20520 2295
rect 20640 2175 20685 2295
rect 20805 2175 20850 2295
rect 20970 2175 21015 2295
rect 21135 2175 21190 2295
rect 21310 2175 21355 2295
rect 21475 2175 21520 2295
rect 21640 2175 21685 2295
rect 21805 2175 21860 2295
rect 21980 2175 22025 2295
rect 22145 2175 22190 2295
rect 22310 2175 22355 2295
rect 22475 2175 22530 2295
rect 22650 2175 22695 2295
rect 22815 2175 22860 2295
rect 22980 2175 23025 2295
rect 23145 2175 23200 2295
rect 23320 2175 23365 2295
rect 23485 2175 23530 2295
rect 23650 2175 23695 2295
rect 23815 2175 23870 2295
rect 23990 2175 24015 2295
rect 18485 2130 24015 2175
rect 18485 2010 18510 2130
rect 18630 2010 18675 2130
rect 18795 2010 18840 2130
rect 18960 2010 19005 2130
rect 19125 2010 19180 2130
rect 19300 2010 19345 2130
rect 19465 2010 19510 2130
rect 19630 2010 19675 2130
rect 19795 2010 19850 2130
rect 19970 2010 20015 2130
rect 20135 2010 20180 2130
rect 20300 2010 20345 2130
rect 20465 2010 20520 2130
rect 20640 2010 20685 2130
rect 20805 2010 20850 2130
rect 20970 2010 21015 2130
rect 21135 2010 21190 2130
rect 21310 2010 21355 2130
rect 21475 2010 21520 2130
rect 21640 2010 21685 2130
rect 21805 2010 21860 2130
rect 21980 2010 22025 2130
rect 22145 2010 22190 2130
rect 22310 2010 22355 2130
rect 22475 2010 22530 2130
rect 22650 2010 22695 2130
rect 22815 2010 22860 2130
rect 22980 2010 23025 2130
rect 23145 2010 23200 2130
rect 23320 2010 23365 2130
rect 23485 2010 23530 2130
rect 23650 2010 23695 2130
rect 23815 2010 23870 2130
rect 23990 2010 24015 2130
rect 18485 1965 24015 2010
rect 18485 1845 18510 1965
rect 18630 1845 18675 1965
rect 18795 1845 18840 1965
rect 18960 1845 19005 1965
rect 19125 1845 19180 1965
rect 19300 1845 19345 1965
rect 19465 1845 19510 1965
rect 19630 1845 19675 1965
rect 19795 1845 19850 1965
rect 19970 1845 20015 1965
rect 20135 1845 20180 1965
rect 20300 1845 20345 1965
rect 20465 1845 20520 1965
rect 20640 1845 20685 1965
rect 20805 1845 20850 1965
rect 20970 1845 21015 1965
rect 21135 1845 21190 1965
rect 21310 1845 21355 1965
rect 21475 1845 21520 1965
rect 21640 1845 21685 1965
rect 21805 1845 21860 1965
rect 21980 1845 22025 1965
rect 22145 1845 22190 1965
rect 22310 1845 22355 1965
rect 22475 1845 22530 1965
rect 22650 1845 22695 1965
rect 22815 1845 22860 1965
rect 22980 1845 23025 1965
rect 23145 1845 23200 1965
rect 23320 1845 23365 1965
rect 23485 1845 23530 1965
rect 23650 1845 23695 1965
rect 23815 1845 23870 1965
rect 23990 1845 24015 1965
rect 18485 1800 24015 1845
rect 18485 1680 18510 1800
rect 18630 1680 18675 1800
rect 18795 1680 18840 1800
rect 18960 1680 19005 1800
rect 19125 1680 19180 1800
rect 19300 1680 19345 1800
rect 19465 1680 19510 1800
rect 19630 1680 19675 1800
rect 19795 1680 19850 1800
rect 19970 1680 20015 1800
rect 20135 1680 20180 1800
rect 20300 1680 20345 1800
rect 20465 1680 20520 1800
rect 20640 1680 20685 1800
rect 20805 1680 20850 1800
rect 20970 1680 21015 1800
rect 21135 1680 21190 1800
rect 21310 1680 21355 1800
rect 21475 1680 21520 1800
rect 21640 1680 21685 1800
rect 21805 1680 21860 1800
rect 21980 1680 22025 1800
rect 22145 1680 22190 1800
rect 22310 1680 22355 1800
rect 22475 1680 22530 1800
rect 22650 1680 22695 1800
rect 22815 1680 22860 1800
rect 22980 1680 23025 1800
rect 23145 1680 23200 1800
rect 23320 1680 23365 1800
rect 23485 1680 23530 1800
rect 23650 1680 23695 1800
rect 23815 1680 23870 1800
rect 23990 1680 24015 1800
rect 18485 1655 24015 1680
rect 24175 7040 24200 7125
rect 24320 7040 24365 7160
rect 24485 7040 24530 7160
rect 24650 7040 24695 7160
rect 24815 7040 24870 7160
rect 24990 7040 25035 7160
rect 25155 7040 25200 7160
rect 25320 7040 25365 7160
rect 25485 7040 25540 7160
rect 25660 7040 25705 7160
rect 25825 7040 25870 7160
rect 25990 7040 26035 7160
rect 26155 7040 26210 7160
rect 26330 7040 26375 7160
rect 26495 7040 26540 7160
rect 26660 7040 26705 7160
rect 26825 7040 26880 7160
rect 27000 7040 27045 7160
rect 27165 7040 27210 7160
rect 27330 7040 27375 7160
rect 27495 7040 27550 7160
rect 27670 7040 27715 7160
rect 27835 7040 27880 7160
rect 28000 7040 28045 7160
rect 28165 7040 28220 7160
rect 28340 7040 28385 7160
rect 28505 7040 28550 7160
rect 28670 7040 28715 7160
rect 28835 7040 28890 7160
rect 29010 7040 29055 7160
rect 29175 7040 29220 7160
rect 29340 7040 29385 7160
rect 29505 7040 29560 7160
rect 29680 7040 29705 7160
rect 24175 6985 29705 7040
rect 24175 6865 24200 6985
rect 24320 6865 24365 6985
rect 24485 6865 24530 6985
rect 24650 6865 24695 6985
rect 24815 6865 24870 6985
rect 24990 6865 25035 6985
rect 25155 6865 25200 6985
rect 25320 6865 25365 6985
rect 25485 6865 25540 6985
rect 25660 6865 25705 6985
rect 25825 6865 25870 6985
rect 25990 6865 26035 6985
rect 26155 6865 26210 6985
rect 26330 6865 26375 6985
rect 26495 6865 26540 6985
rect 26660 6865 26705 6985
rect 26825 6865 26880 6985
rect 27000 6865 27045 6985
rect 27165 6865 27210 6985
rect 27330 6865 27375 6985
rect 27495 6865 27550 6985
rect 27670 6865 27715 6985
rect 27835 6865 27880 6985
rect 28000 6865 28045 6985
rect 28165 6865 28220 6985
rect 28340 6865 28385 6985
rect 28505 6865 28550 6985
rect 28670 6865 28715 6985
rect 28835 6865 28890 6985
rect 29010 6865 29055 6985
rect 29175 6865 29220 6985
rect 29340 6865 29385 6985
rect 29505 6865 29560 6985
rect 29680 6865 29705 6985
rect 24175 6820 29705 6865
rect 24175 6700 24200 6820
rect 24320 6700 24365 6820
rect 24485 6700 24530 6820
rect 24650 6700 24695 6820
rect 24815 6700 24870 6820
rect 24990 6700 25035 6820
rect 25155 6700 25200 6820
rect 25320 6700 25365 6820
rect 25485 6700 25540 6820
rect 25660 6700 25705 6820
rect 25825 6700 25870 6820
rect 25990 6700 26035 6820
rect 26155 6700 26210 6820
rect 26330 6700 26375 6820
rect 26495 6700 26540 6820
rect 26660 6700 26705 6820
rect 26825 6700 26880 6820
rect 27000 6700 27045 6820
rect 27165 6700 27210 6820
rect 27330 6700 27375 6820
rect 27495 6700 27550 6820
rect 27670 6700 27715 6820
rect 27835 6700 27880 6820
rect 28000 6700 28045 6820
rect 28165 6700 28220 6820
rect 28340 6700 28385 6820
rect 28505 6700 28550 6820
rect 28670 6700 28715 6820
rect 28835 6700 28890 6820
rect 29010 6700 29055 6820
rect 29175 6700 29220 6820
rect 29340 6700 29385 6820
rect 29505 6700 29560 6820
rect 29680 6700 29705 6820
rect 24175 6655 29705 6700
rect 24175 6535 24200 6655
rect 24320 6535 24365 6655
rect 24485 6535 24530 6655
rect 24650 6535 24695 6655
rect 24815 6535 24870 6655
rect 24990 6535 25035 6655
rect 25155 6535 25200 6655
rect 25320 6535 25365 6655
rect 25485 6535 25540 6655
rect 25660 6535 25705 6655
rect 25825 6535 25870 6655
rect 25990 6535 26035 6655
rect 26155 6535 26210 6655
rect 26330 6535 26375 6655
rect 26495 6535 26540 6655
rect 26660 6535 26705 6655
rect 26825 6535 26880 6655
rect 27000 6535 27045 6655
rect 27165 6535 27210 6655
rect 27330 6535 27375 6655
rect 27495 6535 27550 6655
rect 27670 6535 27715 6655
rect 27835 6535 27880 6655
rect 28000 6535 28045 6655
rect 28165 6535 28220 6655
rect 28340 6535 28385 6655
rect 28505 6535 28550 6655
rect 28670 6535 28715 6655
rect 28835 6535 28890 6655
rect 29010 6535 29055 6655
rect 29175 6535 29220 6655
rect 29340 6535 29385 6655
rect 29505 6535 29560 6655
rect 29680 6535 29705 6655
rect 24175 6490 29705 6535
rect 24175 6370 24200 6490
rect 24320 6370 24365 6490
rect 24485 6370 24530 6490
rect 24650 6370 24695 6490
rect 24815 6370 24870 6490
rect 24990 6370 25035 6490
rect 25155 6370 25200 6490
rect 25320 6370 25365 6490
rect 25485 6370 25540 6490
rect 25660 6370 25705 6490
rect 25825 6370 25870 6490
rect 25990 6370 26035 6490
rect 26155 6370 26210 6490
rect 26330 6370 26375 6490
rect 26495 6370 26540 6490
rect 26660 6370 26705 6490
rect 26825 6370 26880 6490
rect 27000 6370 27045 6490
rect 27165 6370 27210 6490
rect 27330 6370 27375 6490
rect 27495 6370 27550 6490
rect 27670 6370 27715 6490
rect 27835 6370 27880 6490
rect 28000 6370 28045 6490
rect 28165 6370 28220 6490
rect 28340 6370 28385 6490
rect 28505 6370 28550 6490
rect 28670 6370 28715 6490
rect 28835 6370 28890 6490
rect 29010 6370 29055 6490
rect 29175 6370 29220 6490
rect 29340 6370 29385 6490
rect 29505 6370 29560 6490
rect 29680 6370 29705 6490
rect 24175 6315 29705 6370
rect 24175 6195 24200 6315
rect 24320 6195 24365 6315
rect 24485 6195 24530 6315
rect 24650 6195 24695 6315
rect 24815 6195 24870 6315
rect 24990 6195 25035 6315
rect 25155 6195 25200 6315
rect 25320 6195 25365 6315
rect 25485 6195 25540 6315
rect 25660 6195 25705 6315
rect 25825 6195 25870 6315
rect 25990 6195 26035 6315
rect 26155 6195 26210 6315
rect 26330 6195 26375 6315
rect 26495 6195 26540 6315
rect 26660 6195 26705 6315
rect 26825 6195 26880 6315
rect 27000 6195 27045 6315
rect 27165 6195 27210 6315
rect 27330 6195 27375 6315
rect 27495 6195 27550 6315
rect 27670 6195 27715 6315
rect 27835 6195 27880 6315
rect 28000 6195 28045 6315
rect 28165 6195 28220 6315
rect 28340 6195 28385 6315
rect 28505 6195 28550 6315
rect 28670 6195 28715 6315
rect 28835 6195 28890 6315
rect 29010 6195 29055 6315
rect 29175 6195 29220 6315
rect 29340 6195 29385 6315
rect 29505 6195 29560 6315
rect 29680 6195 29705 6315
rect 24175 6150 29705 6195
rect 24175 6030 24200 6150
rect 24320 6030 24365 6150
rect 24485 6030 24530 6150
rect 24650 6030 24695 6150
rect 24815 6030 24870 6150
rect 24990 6030 25035 6150
rect 25155 6030 25200 6150
rect 25320 6030 25365 6150
rect 25485 6030 25540 6150
rect 25660 6030 25705 6150
rect 25825 6030 25870 6150
rect 25990 6030 26035 6150
rect 26155 6030 26210 6150
rect 26330 6030 26375 6150
rect 26495 6030 26540 6150
rect 26660 6030 26705 6150
rect 26825 6030 26880 6150
rect 27000 6030 27045 6150
rect 27165 6030 27210 6150
rect 27330 6030 27375 6150
rect 27495 6030 27550 6150
rect 27670 6030 27715 6150
rect 27835 6030 27880 6150
rect 28000 6030 28045 6150
rect 28165 6030 28220 6150
rect 28340 6030 28385 6150
rect 28505 6030 28550 6150
rect 28670 6030 28715 6150
rect 28835 6030 28890 6150
rect 29010 6030 29055 6150
rect 29175 6030 29220 6150
rect 29340 6030 29385 6150
rect 29505 6030 29560 6150
rect 29680 6030 29705 6150
rect 24175 5985 29705 6030
rect 24175 5865 24200 5985
rect 24320 5865 24365 5985
rect 24485 5865 24530 5985
rect 24650 5865 24695 5985
rect 24815 5865 24870 5985
rect 24990 5865 25035 5985
rect 25155 5865 25200 5985
rect 25320 5865 25365 5985
rect 25485 5865 25540 5985
rect 25660 5865 25705 5985
rect 25825 5865 25870 5985
rect 25990 5865 26035 5985
rect 26155 5865 26210 5985
rect 26330 5865 26375 5985
rect 26495 5865 26540 5985
rect 26660 5865 26705 5985
rect 26825 5865 26880 5985
rect 27000 5865 27045 5985
rect 27165 5865 27210 5985
rect 27330 5865 27375 5985
rect 27495 5865 27550 5985
rect 27670 5865 27715 5985
rect 27835 5865 27880 5985
rect 28000 5865 28045 5985
rect 28165 5865 28220 5985
rect 28340 5865 28385 5985
rect 28505 5865 28550 5985
rect 28670 5865 28715 5985
rect 28835 5865 28890 5985
rect 29010 5865 29055 5985
rect 29175 5865 29220 5985
rect 29340 5865 29385 5985
rect 29505 5865 29560 5985
rect 29680 5865 29705 5985
rect 24175 5820 29705 5865
rect 24175 5700 24200 5820
rect 24320 5700 24365 5820
rect 24485 5700 24530 5820
rect 24650 5700 24695 5820
rect 24815 5700 24870 5820
rect 24990 5700 25035 5820
rect 25155 5700 25200 5820
rect 25320 5700 25365 5820
rect 25485 5700 25540 5820
rect 25660 5700 25705 5820
rect 25825 5700 25870 5820
rect 25990 5700 26035 5820
rect 26155 5700 26210 5820
rect 26330 5700 26375 5820
rect 26495 5700 26540 5820
rect 26660 5700 26705 5820
rect 26825 5700 26880 5820
rect 27000 5700 27045 5820
rect 27165 5700 27210 5820
rect 27330 5700 27375 5820
rect 27495 5700 27550 5820
rect 27670 5700 27715 5820
rect 27835 5700 27880 5820
rect 28000 5700 28045 5820
rect 28165 5700 28220 5820
rect 28340 5700 28385 5820
rect 28505 5700 28550 5820
rect 28670 5700 28715 5820
rect 28835 5700 28890 5820
rect 29010 5700 29055 5820
rect 29175 5700 29220 5820
rect 29340 5700 29385 5820
rect 29505 5700 29560 5820
rect 29680 5700 29705 5820
rect 24175 5645 29705 5700
rect 24175 5525 24200 5645
rect 24320 5525 24365 5645
rect 24485 5525 24530 5645
rect 24650 5525 24695 5645
rect 24815 5525 24870 5645
rect 24990 5525 25035 5645
rect 25155 5525 25200 5645
rect 25320 5525 25365 5645
rect 25485 5525 25540 5645
rect 25660 5525 25705 5645
rect 25825 5525 25870 5645
rect 25990 5525 26035 5645
rect 26155 5525 26210 5645
rect 26330 5525 26375 5645
rect 26495 5525 26540 5645
rect 26660 5525 26705 5645
rect 26825 5525 26880 5645
rect 27000 5525 27045 5645
rect 27165 5525 27210 5645
rect 27330 5525 27375 5645
rect 27495 5525 27550 5645
rect 27670 5525 27715 5645
rect 27835 5525 27880 5645
rect 28000 5525 28045 5645
rect 28165 5525 28220 5645
rect 28340 5525 28385 5645
rect 28505 5525 28550 5645
rect 28670 5525 28715 5645
rect 28835 5525 28890 5645
rect 29010 5525 29055 5645
rect 29175 5525 29220 5645
rect 29340 5525 29385 5645
rect 29505 5525 29560 5645
rect 29680 5525 29705 5645
rect 24175 5480 29705 5525
rect 24175 5360 24200 5480
rect 24320 5360 24365 5480
rect 24485 5360 24530 5480
rect 24650 5360 24695 5480
rect 24815 5360 24870 5480
rect 24990 5360 25035 5480
rect 25155 5360 25200 5480
rect 25320 5360 25365 5480
rect 25485 5360 25540 5480
rect 25660 5360 25705 5480
rect 25825 5360 25870 5480
rect 25990 5360 26035 5480
rect 26155 5360 26210 5480
rect 26330 5360 26375 5480
rect 26495 5360 26540 5480
rect 26660 5360 26705 5480
rect 26825 5360 26880 5480
rect 27000 5360 27045 5480
rect 27165 5360 27210 5480
rect 27330 5360 27375 5480
rect 27495 5360 27550 5480
rect 27670 5360 27715 5480
rect 27835 5360 27880 5480
rect 28000 5360 28045 5480
rect 28165 5360 28220 5480
rect 28340 5360 28385 5480
rect 28505 5360 28550 5480
rect 28670 5360 28715 5480
rect 28835 5360 28890 5480
rect 29010 5360 29055 5480
rect 29175 5360 29220 5480
rect 29340 5360 29385 5480
rect 29505 5360 29560 5480
rect 29680 5360 29705 5480
rect 24175 5315 29705 5360
rect 24175 5195 24200 5315
rect 24320 5195 24365 5315
rect 24485 5195 24530 5315
rect 24650 5195 24695 5315
rect 24815 5195 24870 5315
rect 24990 5195 25035 5315
rect 25155 5195 25200 5315
rect 25320 5195 25365 5315
rect 25485 5195 25540 5315
rect 25660 5195 25705 5315
rect 25825 5195 25870 5315
rect 25990 5195 26035 5315
rect 26155 5195 26210 5315
rect 26330 5195 26375 5315
rect 26495 5195 26540 5315
rect 26660 5195 26705 5315
rect 26825 5195 26880 5315
rect 27000 5195 27045 5315
rect 27165 5195 27210 5315
rect 27330 5195 27375 5315
rect 27495 5195 27550 5315
rect 27670 5195 27715 5315
rect 27835 5195 27880 5315
rect 28000 5195 28045 5315
rect 28165 5195 28220 5315
rect 28340 5195 28385 5315
rect 28505 5195 28550 5315
rect 28670 5195 28715 5315
rect 28835 5195 28890 5315
rect 29010 5195 29055 5315
rect 29175 5195 29220 5315
rect 29340 5195 29385 5315
rect 29505 5195 29560 5315
rect 29680 5195 29705 5315
rect 24175 5150 29705 5195
rect 24175 5030 24200 5150
rect 24320 5030 24365 5150
rect 24485 5030 24530 5150
rect 24650 5030 24695 5150
rect 24815 5030 24870 5150
rect 24990 5030 25035 5150
rect 25155 5030 25200 5150
rect 25320 5030 25365 5150
rect 25485 5030 25540 5150
rect 25660 5030 25705 5150
rect 25825 5030 25870 5150
rect 25990 5030 26035 5150
rect 26155 5030 26210 5150
rect 26330 5030 26375 5150
rect 26495 5030 26540 5150
rect 26660 5030 26705 5150
rect 26825 5030 26880 5150
rect 27000 5030 27045 5150
rect 27165 5030 27210 5150
rect 27330 5030 27375 5150
rect 27495 5030 27550 5150
rect 27670 5030 27715 5150
rect 27835 5030 27880 5150
rect 28000 5030 28045 5150
rect 28165 5030 28220 5150
rect 28340 5030 28385 5150
rect 28505 5030 28550 5150
rect 28670 5030 28715 5150
rect 28835 5030 28890 5150
rect 29010 5030 29055 5150
rect 29175 5030 29220 5150
rect 29340 5030 29385 5150
rect 29505 5030 29560 5150
rect 29680 5030 29705 5150
rect 24175 4975 29705 5030
rect 24175 4855 24200 4975
rect 24320 4855 24365 4975
rect 24485 4855 24530 4975
rect 24650 4855 24695 4975
rect 24815 4855 24870 4975
rect 24990 4855 25035 4975
rect 25155 4855 25200 4975
rect 25320 4855 25365 4975
rect 25485 4855 25540 4975
rect 25660 4855 25705 4975
rect 25825 4855 25870 4975
rect 25990 4855 26035 4975
rect 26155 4855 26210 4975
rect 26330 4855 26375 4975
rect 26495 4855 26540 4975
rect 26660 4855 26705 4975
rect 26825 4855 26880 4975
rect 27000 4855 27045 4975
rect 27165 4855 27210 4975
rect 27330 4855 27375 4975
rect 27495 4855 27550 4975
rect 27670 4855 27715 4975
rect 27835 4855 27880 4975
rect 28000 4855 28045 4975
rect 28165 4855 28220 4975
rect 28340 4855 28385 4975
rect 28505 4855 28550 4975
rect 28670 4855 28715 4975
rect 28835 4855 28890 4975
rect 29010 4855 29055 4975
rect 29175 4855 29220 4975
rect 29340 4855 29385 4975
rect 29505 4855 29560 4975
rect 29680 4855 29705 4975
rect 24175 4810 29705 4855
rect 24175 4690 24200 4810
rect 24320 4690 24365 4810
rect 24485 4690 24530 4810
rect 24650 4690 24695 4810
rect 24815 4690 24870 4810
rect 24990 4690 25035 4810
rect 25155 4690 25200 4810
rect 25320 4690 25365 4810
rect 25485 4690 25540 4810
rect 25660 4690 25705 4810
rect 25825 4690 25870 4810
rect 25990 4690 26035 4810
rect 26155 4690 26210 4810
rect 26330 4690 26375 4810
rect 26495 4690 26540 4810
rect 26660 4690 26705 4810
rect 26825 4690 26880 4810
rect 27000 4690 27045 4810
rect 27165 4690 27210 4810
rect 27330 4690 27375 4810
rect 27495 4690 27550 4810
rect 27670 4690 27715 4810
rect 27835 4690 27880 4810
rect 28000 4690 28045 4810
rect 28165 4690 28220 4810
rect 28340 4690 28385 4810
rect 28505 4690 28550 4810
rect 28670 4690 28715 4810
rect 28835 4690 28890 4810
rect 29010 4690 29055 4810
rect 29175 4690 29220 4810
rect 29340 4690 29385 4810
rect 29505 4690 29560 4810
rect 29680 4690 29705 4810
rect 24175 4645 29705 4690
rect 24175 4525 24200 4645
rect 24320 4525 24365 4645
rect 24485 4525 24530 4645
rect 24650 4525 24695 4645
rect 24815 4525 24870 4645
rect 24990 4525 25035 4645
rect 25155 4525 25200 4645
rect 25320 4525 25365 4645
rect 25485 4525 25540 4645
rect 25660 4525 25705 4645
rect 25825 4525 25870 4645
rect 25990 4525 26035 4645
rect 26155 4525 26210 4645
rect 26330 4525 26375 4645
rect 26495 4525 26540 4645
rect 26660 4525 26705 4645
rect 26825 4525 26880 4645
rect 27000 4525 27045 4645
rect 27165 4525 27210 4645
rect 27330 4525 27375 4645
rect 27495 4525 27550 4645
rect 27670 4525 27715 4645
rect 27835 4525 27880 4645
rect 28000 4525 28045 4645
rect 28165 4525 28220 4645
rect 28340 4525 28385 4645
rect 28505 4525 28550 4645
rect 28670 4525 28715 4645
rect 28835 4525 28890 4645
rect 29010 4525 29055 4645
rect 29175 4525 29220 4645
rect 29340 4525 29385 4645
rect 29505 4525 29560 4645
rect 29680 4525 29705 4645
rect 24175 4480 29705 4525
rect 24175 4360 24200 4480
rect 24320 4360 24365 4480
rect 24485 4360 24530 4480
rect 24650 4360 24695 4480
rect 24815 4360 24870 4480
rect 24990 4360 25035 4480
rect 25155 4360 25200 4480
rect 25320 4360 25365 4480
rect 25485 4360 25540 4480
rect 25660 4360 25705 4480
rect 25825 4360 25870 4480
rect 25990 4360 26035 4480
rect 26155 4360 26210 4480
rect 26330 4360 26375 4480
rect 26495 4360 26540 4480
rect 26660 4360 26705 4480
rect 26825 4360 26880 4480
rect 27000 4360 27045 4480
rect 27165 4360 27210 4480
rect 27330 4360 27375 4480
rect 27495 4360 27550 4480
rect 27670 4360 27715 4480
rect 27835 4360 27880 4480
rect 28000 4360 28045 4480
rect 28165 4360 28220 4480
rect 28340 4360 28385 4480
rect 28505 4360 28550 4480
rect 28670 4360 28715 4480
rect 28835 4360 28890 4480
rect 29010 4360 29055 4480
rect 29175 4360 29220 4480
rect 29340 4360 29385 4480
rect 29505 4360 29560 4480
rect 29680 4360 29705 4480
rect 24175 4305 29705 4360
rect 24175 4185 24200 4305
rect 24320 4185 24365 4305
rect 24485 4185 24530 4305
rect 24650 4185 24695 4305
rect 24815 4185 24870 4305
rect 24990 4185 25035 4305
rect 25155 4185 25200 4305
rect 25320 4185 25365 4305
rect 25485 4185 25540 4305
rect 25660 4185 25705 4305
rect 25825 4185 25870 4305
rect 25990 4185 26035 4305
rect 26155 4185 26210 4305
rect 26330 4185 26375 4305
rect 26495 4185 26540 4305
rect 26660 4185 26705 4305
rect 26825 4185 26880 4305
rect 27000 4185 27045 4305
rect 27165 4185 27210 4305
rect 27330 4185 27375 4305
rect 27495 4185 27550 4305
rect 27670 4185 27715 4305
rect 27835 4185 27880 4305
rect 28000 4185 28045 4305
rect 28165 4185 28220 4305
rect 28340 4185 28385 4305
rect 28505 4185 28550 4305
rect 28670 4185 28715 4305
rect 28835 4185 28890 4305
rect 29010 4185 29055 4305
rect 29175 4185 29220 4305
rect 29340 4185 29385 4305
rect 29505 4185 29560 4305
rect 29680 4185 29705 4305
rect 24175 4140 29705 4185
rect 24175 4020 24200 4140
rect 24320 4020 24365 4140
rect 24485 4020 24530 4140
rect 24650 4020 24695 4140
rect 24815 4020 24870 4140
rect 24990 4020 25035 4140
rect 25155 4020 25200 4140
rect 25320 4020 25365 4140
rect 25485 4020 25540 4140
rect 25660 4020 25705 4140
rect 25825 4020 25870 4140
rect 25990 4020 26035 4140
rect 26155 4020 26210 4140
rect 26330 4020 26375 4140
rect 26495 4020 26540 4140
rect 26660 4020 26705 4140
rect 26825 4020 26880 4140
rect 27000 4020 27045 4140
rect 27165 4020 27210 4140
rect 27330 4020 27375 4140
rect 27495 4020 27550 4140
rect 27670 4020 27715 4140
rect 27835 4020 27880 4140
rect 28000 4020 28045 4140
rect 28165 4020 28220 4140
rect 28340 4020 28385 4140
rect 28505 4020 28550 4140
rect 28670 4020 28715 4140
rect 28835 4020 28890 4140
rect 29010 4020 29055 4140
rect 29175 4020 29220 4140
rect 29340 4020 29385 4140
rect 29505 4020 29560 4140
rect 29680 4020 29705 4140
rect 24175 3975 29705 4020
rect 24175 3855 24200 3975
rect 24320 3855 24365 3975
rect 24485 3855 24530 3975
rect 24650 3855 24695 3975
rect 24815 3855 24870 3975
rect 24990 3855 25035 3975
rect 25155 3855 25200 3975
rect 25320 3855 25365 3975
rect 25485 3855 25540 3975
rect 25660 3855 25705 3975
rect 25825 3855 25870 3975
rect 25990 3855 26035 3975
rect 26155 3855 26210 3975
rect 26330 3855 26375 3975
rect 26495 3855 26540 3975
rect 26660 3855 26705 3975
rect 26825 3855 26880 3975
rect 27000 3855 27045 3975
rect 27165 3855 27210 3975
rect 27330 3855 27375 3975
rect 27495 3855 27550 3975
rect 27670 3855 27715 3975
rect 27835 3855 27880 3975
rect 28000 3855 28045 3975
rect 28165 3855 28220 3975
rect 28340 3855 28385 3975
rect 28505 3855 28550 3975
rect 28670 3855 28715 3975
rect 28835 3855 28890 3975
rect 29010 3855 29055 3975
rect 29175 3855 29220 3975
rect 29340 3855 29385 3975
rect 29505 3855 29560 3975
rect 29680 3855 29705 3975
rect 24175 3810 29705 3855
rect 24175 3690 24200 3810
rect 24320 3690 24365 3810
rect 24485 3690 24530 3810
rect 24650 3690 24695 3810
rect 24815 3690 24870 3810
rect 24990 3690 25035 3810
rect 25155 3690 25200 3810
rect 25320 3690 25365 3810
rect 25485 3690 25540 3810
rect 25660 3690 25705 3810
rect 25825 3690 25870 3810
rect 25990 3690 26035 3810
rect 26155 3690 26210 3810
rect 26330 3690 26375 3810
rect 26495 3690 26540 3810
rect 26660 3690 26705 3810
rect 26825 3690 26880 3810
rect 27000 3690 27045 3810
rect 27165 3690 27210 3810
rect 27330 3690 27375 3810
rect 27495 3690 27550 3810
rect 27670 3690 27715 3810
rect 27835 3690 27880 3810
rect 28000 3690 28045 3810
rect 28165 3690 28220 3810
rect 28340 3690 28385 3810
rect 28505 3690 28550 3810
rect 28670 3690 28715 3810
rect 28835 3690 28890 3810
rect 29010 3690 29055 3810
rect 29175 3690 29220 3810
rect 29340 3690 29385 3810
rect 29505 3690 29560 3810
rect 29680 3690 29705 3810
rect 24175 3635 29705 3690
rect 24175 3515 24200 3635
rect 24320 3515 24365 3635
rect 24485 3515 24530 3635
rect 24650 3515 24695 3635
rect 24815 3515 24870 3635
rect 24990 3515 25035 3635
rect 25155 3515 25200 3635
rect 25320 3515 25365 3635
rect 25485 3515 25540 3635
rect 25660 3515 25705 3635
rect 25825 3515 25870 3635
rect 25990 3515 26035 3635
rect 26155 3515 26210 3635
rect 26330 3515 26375 3635
rect 26495 3515 26540 3635
rect 26660 3515 26705 3635
rect 26825 3515 26880 3635
rect 27000 3515 27045 3635
rect 27165 3515 27210 3635
rect 27330 3515 27375 3635
rect 27495 3515 27550 3635
rect 27670 3515 27715 3635
rect 27835 3515 27880 3635
rect 28000 3515 28045 3635
rect 28165 3515 28220 3635
rect 28340 3515 28385 3635
rect 28505 3515 28550 3635
rect 28670 3515 28715 3635
rect 28835 3515 28890 3635
rect 29010 3515 29055 3635
rect 29175 3515 29220 3635
rect 29340 3515 29385 3635
rect 29505 3515 29560 3635
rect 29680 3515 29705 3635
rect 24175 3470 29705 3515
rect 24175 3350 24200 3470
rect 24320 3350 24365 3470
rect 24485 3350 24530 3470
rect 24650 3350 24695 3470
rect 24815 3350 24870 3470
rect 24990 3350 25035 3470
rect 25155 3350 25200 3470
rect 25320 3350 25365 3470
rect 25485 3350 25540 3470
rect 25660 3350 25705 3470
rect 25825 3350 25870 3470
rect 25990 3350 26035 3470
rect 26155 3350 26210 3470
rect 26330 3350 26375 3470
rect 26495 3350 26540 3470
rect 26660 3350 26705 3470
rect 26825 3350 26880 3470
rect 27000 3350 27045 3470
rect 27165 3350 27210 3470
rect 27330 3350 27375 3470
rect 27495 3350 27550 3470
rect 27670 3350 27715 3470
rect 27835 3350 27880 3470
rect 28000 3350 28045 3470
rect 28165 3350 28220 3470
rect 28340 3350 28385 3470
rect 28505 3350 28550 3470
rect 28670 3350 28715 3470
rect 28835 3350 28890 3470
rect 29010 3350 29055 3470
rect 29175 3350 29220 3470
rect 29340 3350 29385 3470
rect 29505 3350 29560 3470
rect 29680 3350 29705 3470
rect 24175 3305 29705 3350
rect 24175 3185 24200 3305
rect 24320 3185 24365 3305
rect 24485 3185 24530 3305
rect 24650 3185 24695 3305
rect 24815 3185 24870 3305
rect 24990 3185 25035 3305
rect 25155 3185 25200 3305
rect 25320 3185 25365 3305
rect 25485 3185 25540 3305
rect 25660 3185 25705 3305
rect 25825 3185 25870 3305
rect 25990 3185 26035 3305
rect 26155 3185 26210 3305
rect 26330 3185 26375 3305
rect 26495 3185 26540 3305
rect 26660 3185 26705 3305
rect 26825 3185 26880 3305
rect 27000 3185 27045 3305
rect 27165 3185 27210 3305
rect 27330 3185 27375 3305
rect 27495 3185 27550 3305
rect 27670 3185 27715 3305
rect 27835 3185 27880 3305
rect 28000 3185 28045 3305
rect 28165 3185 28220 3305
rect 28340 3185 28385 3305
rect 28505 3185 28550 3305
rect 28670 3185 28715 3305
rect 28835 3185 28890 3305
rect 29010 3185 29055 3305
rect 29175 3185 29220 3305
rect 29340 3185 29385 3305
rect 29505 3185 29560 3305
rect 29680 3185 29705 3305
rect 24175 3140 29705 3185
rect 24175 3020 24200 3140
rect 24320 3020 24365 3140
rect 24485 3020 24530 3140
rect 24650 3020 24695 3140
rect 24815 3020 24870 3140
rect 24990 3020 25035 3140
rect 25155 3020 25200 3140
rect 25320 3020 25365 3140
rect 25485 3020 25540 3140
rect 25660 3020 25705 3140
rect 25825 3020 25870 3140
rect 25990 3020 26035 3140
rect 26155 3020 26210 3140
rect 26330 3020 26375 3140
rect 26495 3020 26540 3140
rect 26660 3020 26705 3140
rect 26825 3020 26880 3140
rect 27000 3020 27045 3140
rect 27165 3020 27210 3140
rect 27330 3020 27375 3140
rect 27495 3020 27550 3140
rect 27670 3020 27715 3140
rect 27835 3020 27880 3140
rect 28000 3020 28045 3140
rect 28165 3020 28220 3140
rect 28340 3020 28385 3140
rect 28505 3020 28550 3140
rect 28670 3020 28715 3140
rect 28835 3020 28890 3140
rect 29010 3020 29055 3140
rect 29175 3020 29220 3140
rect 29340 3020 29385 3140
rect 29505 3020 29560 3140
rect 29680 3020 29705 3140
rect 24175 2965 29705 3020
rect 24175 2845 24200 2965
rect 24320 2845 24365 2965
rect 24485 2845 24530 2965
rect 24650 2845 24695 2965
rect 24815 2845 24870 2965
rect 24990 2845 25035 2965
rect 25155 2845 25200 2965
rect 25320 2845 25365 2965
rect 25485 2845 25540 2965
rect 25660 2845 25705 2965
rect 25825 2845 25870 2965
rect 25990 2845 26035 2965
rect 26155 2845 26210 2965
rect 26330 2845 26375 2965
rect 26495 2845 26540 2965
rect 26660 2845 26705 2965
rect 26825 2845 26880 2965
rect 27000 2845 27045 2965
rect 27165 2845 27210 2965
rect 27330 2845 27375 2965
rect 27495 2845 27550 2965
rect 27670 2845 27715 2965
rect 27835 2845 27880 2965
rect 28000 2845 28045 2965
rect 28165 2845 28220 2965
rect 28340 2845 28385 2965
rect 28505 2845 28550 2965
rect 28670 2845 28715 2965
rect 28835 2845 28890 2965
rect 29010 2845 29055 2965
rect 29175 2845 29220 2965
rect 29340 2845 29385 2965
rect 29505 2845 29560 2965
rect 29680 2845 29705 2965
rect 24175 2800 29705 2845
rect 24175 2680 24200 2800
rect 24320 2680 24365 2800
rect 24485 2680 24530 2800
rect 24650 2680 24695 2800
rect 24815 2680 24870 2800
rect 24990 2680 25035 2800
rect 25155 2680 25200 2800
rect 25320 2680 25365 2800
rect 25485 2680 25540 2800
rect 25660 2680 25705 2800
rect 25825 2680 25870 2800
rect 25990 2680 26035 2800
rect 26155 2680 26210 2800
rect 26330 2680 26375 2800
rect 26495 2680 26540 2800
rect 26660 2680 26705 2800
rect 26825 2680 26880 2800
rect 27000 2680 27045 2800
rect 27165 2680 27210 2800
rect 27330 2680 27375 2800
rect 27495 2680 27550 2800
rect 27670 2680 27715 2800
rect 27835 2680 27880 2800
rect 28000 2680 28045 2800
rect 28165 2680 28220 2800
rect 28340 2680 28385 2800
rect 28505 2680 28550 2800
rect 28670 2680 28715 2800
rect 28835 2680 28890 2800
rect 29010 2680 29055 2800
rect 29175 2680 29220 2800
rect 29340 2680 29385 2800
rect 29505 2680 29560 2800
rect 29680 2680 29705 2800
rect 24175 2635 29705 2680
rect 24175 2515 24200 2635
rect 24320 2515 24365 2635
rect 24485 2515 24530 2635
rect 24650 2515 24695 2635
rect 24815 2515 24870 2635
rect 24990 2515 25035 2635
rect 25155 2515 25200 2635
rect 25320 2515 25365 2635
rect 25485 2515 25540 2635
rect 25660 2515 25705 2635
rect 25825 2515 25870 2635
rect 25990 2515 26035 2635
rect 26155 2515 26210 2635
rect 26330 2515 26375 2635
rect 26495 2515 26540 2635
rect 26660 2515 26705 2635
rect 26825 2515 26880 2635
rect 27000 2515 27045 2635
rect 27165 2515 27210 2635
rect 27330 2515 27375 2635
rect 27495 2515 27550 2635
rect 27670 2515 27715 2635
rect 27835 2515 27880 2635
rect 28000 2515 28045 2635
rect 28165 2515 28220 2635
rect 28340 2515 28385 2635
rect 28505 2515 28550 2635
rect 28670 2515 28715 2635
rect 28835 2515 28890 2635
rect 29010 2515 29055 2635
rect 29175 2515 29220 2635
rect 29340 2515 29385 2635
rect 29505 2515 29560 2635
rect 29680 2515 29705 2635
rect 24175 2470 29705 2515
rect 24175 2350 24200 2470
rect 24320 2350 24365 2470
rect 24485 2350 24530 2470
rect 24650 2350 24695 2470
rect 24815 2350 24870 2470
rect 24990 2350 25035 2470
rect 25155 2350 25200 2470
rect 25320 2350 25365 2470
rect 25485 2350 25540 2470
rect 25660 2350 25705 2470
rect 25825 2350 25870 2470
rect 25990 2350 26035 2470
rect 26155 2350 26210 2470
rect 26330 2350 26375 2470
rect 26495 2350 26540 2470
rect 26660 2350 26705 2470
rect 26825 2350 26880 2470
rect 27000 2350 27045 2470
rect 27165 2350 27210 2470
rect 27330 2350 27375 2470
rect 27495 2350 27550 2470
rect 27670 2350 27715 2470
rect 27835 2350 27880 2470
rect 28000 2350 28045 2470
rect 28165 2350 28220 2470
rect 28340 2350 28385 2470
rect 28505 2350 28550 2470
rect 28670 2350 28715 2470
rect 28835 2350 28890 2470
rect 29010 2350 29055 2470
rect 29175 2350 29220 2470
rect 29340 2350 29385 2470
rect 29505 2350 29560 2470
rect 29680 2350 29705 2470
rect 24175 2295 29705 2350
rect 24175 2175 24200 2295
rect 24320 2175 24365 2295
rect 24485 2175 24530 2295
rect 24650 2175 24695 2295
rect 24815 2175 24870 2295
rect 24990 2175 25035 2295
rect 25155 2175 25200 2295
rect 25320 2175 25365 2295
rect 25485 2175 25540 2295
rect 25660 2175 25705 2295
rect 25825 2175 25870 2295
rect 25990 2175 26035 2295
rect 26155 2175 26210 2295
rect 26330 2175 26375 2295
rect 26495 2175 26540 2295
rect 26660 2175 26705 2295
rect 26825 2175 26880 2295
rect 27000 2175 27045 2295
rect 27165 2175 27210 2295
rect 27330 2175 27375 2295
rect 27495 2175 27550 2295
rect 27670 2175 27715 2295
rect 27835 2175 27880 2295
rect 28000 2175 28045 2295
rect 28165 2175 28220 2295
rect 28340 2175 28385 2295
rect 28505 2175 28550 2295
rect 28670 2175 28715 2295
rect 28835 2175 28890 2295
rect 29010 2175 29055 2295
rect 29175 2175 29220 2295
rect 29340 2175 29385 2295
rect 29505 2175 29560 2295
rect 29680 2175 29705 2295
rect 24175 2130 29705 2175
rect 24175 2010 24200 2130
rect 24320 2010 24365 2130
rect 24485 2010 24530 2130
rect 24650 2010 24695 2130
rect 24815 2010 24870 2130
rect 24990 2010 25035 2130
rect 25155 2010 25200 2130
rect 25320 2010 25365 2130
rect 25485 2010 25540 2130
rect 25660 2010 25705 2130
rect 25825 2010 25870 2130
rect 25990 2010 26035 2130
rect 26155 2010 26210 2130
rect 26330 2010 26375 2130
rect 26495 2010 26540 2130
rect 26660 2010 26705 2130
rect 26825 2010 26880 2130
rect 27000 2010 27045 2130
rect 27165 2010 27210 2130
rect 27330 2010 27375 2130
rect 27495 2010 27550 2130
rect 27670 2010 27715 2130
rect 27835 2010 27880 2130
rect 28000 2010 28045 2130
rect 28165 2010 28220 2130
rect 28340 2010 28385 2130
rect 28505 2010 28550 2130
rect 28670 2010 28715 2130
rect 28835 2010 28890 2130
rect 29010 2010 29055 2130
rect 29175 2010 29220 2130
rect 29340 2010 29385 2130
rect 29505 2010 29560 2130
rect 29680 2010 29705 2130
rect 24175 1965 29705 2010
rect 24175 1845 24200 1965
rect 24320 1845 24365 1965
rect 24485 1845 24530 1965
rect 24650 1845 24695 1965
rect 24815 1845 24870 1965
rect 24990 1845 25035 1965
rect 25155 1845 25200 1965
rect 25320 1845 25365 1965
rect 25485 1845 25540 1965
rect 25660 1845 25705 1965
rect 25825 1845 25870 1965
rect 25990 1845 26035 1965
rect 26155 1845 26210 1965
rect 26330 1845 26375 1965
rect 26495 1845 26540 1965
rect 26660 1845 26705 1965
rect 26825 1845 26880 1965
rect 27000 1845 27045 1965
rect 27165 1845 27210 1965
rect 27330 1845 27375 1965
rect 27495 1845 27550 1965
rect 27670 1845 27715 1965
rect 27835 1845 27880 1965
rect 28000 1845 28045 1965
rect 28165 1845 28220 1965
rect 28340 1845 28385 1965
rect 28505 1845 28550 1965
rect 28670 1845 28715 1965
rect 28835 1845 28890 1965
rect 29010 1845 29055 1965
rect 29175 1845 29220 1965
rect 29340 1845 29385 1965
rect 29505 1845 29560 1965
rect 29680 1845 29705 1965
rect 24175 1800 29705 1845
rect 24175 1680 24200 1800
rect 24320 1680 24365 1800
rect 24485 1680 24530 1800
rect 24650 1680 24695 1800
rect 24815 1680 24870 1800
rect 24990 1680 25035 1800
rect 25155 1680 25200 1800
rect 25320 1680 25365 1800
rect 25485 1680 25540 1800
rect 25660 1680 25705 1800
rect 25825 1680 25870 1800
rect 25990 1680 26035 1800
rect 26155 1680 26210 1800
rect 26330 1680 26375 1800
rect 26495 1680 26540 1800
rect 26660 1680 26705 1800
rect 26825 1680 26880 1800
rect 27000 1680 27045 1800
rect 27165 1680 27210 1800
rect 27330 1680 27375 1800
rect 27495 1680 27550 1800
rect 27670 1680 27715 1800
rect 27835 1680 27880 1800
rect 28000 1680 28045 1800
rect 28165 1680 28220 1800
rect 28340 1680 28385 1800
rect 28505 1680 28550 1800
rect 28670 1680 28715 1800
rect 28835 1680 28890 1800
rect 29010 1680 29055 1800
rect 29175 1680 29220 1800
rect 29340 1680 29385 1800
rect 29505 1680 29560 1800
rect 29680 1680 29705 1800
rect 24175 1655 29705 1680
rect 12635 1605 12795 1610
rect 18325 1605 18485 1610
rect 24015 1605 24175 1610
rect 7105 1590 29705 1605
rect 7105 1470 7170 1590
rect 7290 1470 7335 1590
rect 7455 1470 7500 1590
rect 7620 1470 7665 1590
rect 7785 1470 7830 1590
rect 7950 1470 7995 1590
rect 8115 1470 8160 1590
rect 8280 1470 8325 1590
rect 8445 1470 8490 1590
rect 8610 1470 8655 1590
rect 8775 1470 8820 1590
rect 8940 1470 8985 1590
rect 9105 1470 9150 1590
rect 9270 1470 9315 1590
rect 9435 1470 9480 1590
rect 9600 1470 9645 1590
rect 9765 1470 9810 1590
rect 9930 1470 9975 1590
rect 10095 1470 10140 1590
rect 10260 1470 10305 1590
rect 10425 1470 10470 1590
rect 10590 1470 10635 1590
rect 10755 1470 10800 1590
rect 10920 1470 10965 1590
rect 11085 1470 11130 1590
rect 11250 1470 11295 1590
rect 11415 1470 11460 1590
rect 11580 1470 11625 1590
rect 11745 1470 11790 1590
rect 11910 1470 11955 1590
rect 12075 1470 12120 1590
rect 12240 1470 12285 1590
rect 12405 1470 12450 1590
rect 12570 1470 12860 1590
rect 12980 1470 13025 1590
rect 13145 1470 13190 1590
rect 13310 1470 13355 1590
rect 13475 1470 13520 1590
rect 13640 1470 13685 1590
rect 13805 1470 13850 1590
rect 13970 1470 14015 1590
rect 14135 1470 14180 1590
rect 14300 1470 14345 1590
rect 14465 1470 14510 1590
rect 14630 1470 14675 1590
rect 14795 1470 14840 1590
rect 14960 1470 15005 1590
rect 15125 1470 15170 1590
rect 15290 1470 15335 1590
rect 15455 1470 15500 1590
rect 15620 1470 15665 1590
rect 15785 1470 15830 1590
rect 15950 1470 15995 1590
rect 16115 1470 16160 1590
rect 16280 1470 16325 1590
rect 16445 1470 16490 1590
rect 16610 1470 16655 1590
rect 16775 1470 16820 1590
rect 16940 1470 16985 1590
rect 17105 1470 17150 1590
rect 17270 1470 17315 1590
rect 17435 1470 17480 1590
rect 17600 1470 17645 1590
rect 17765 1470 17810 1590
rect 17930 1470 17975 1590
rect 18095 1470 18140 1590
rect 18260 1470 18550 1590
rect 18670 1470 18715 1590
rect 18835 1470 18880 1590
rect 19000 1470 19045 1590
rect 19165 1470 19210 1590
rect 19330 1470 19375 1590
rect 19495 1470 19540 1590
rect 19660 1470 19705 1590
rect 19825 1470 19870 1590
rect 19990 1470 20035 1590
rect 20155 1470 20200 1590
rect 20320 1470 20365 1590
rect 20485 1470 20530 1590
rect 20650 1470 20695 1590
rect 20815 1470 20860 1590
rect 20980 1470 21025 1590
rect 21145 1470 21190 1590
rect 21310 1470 21355 1590
rect 21475 1470 21520 1590
rect 21640 1470 21685 1590
rect 21805 1470 21850 1590
rect 21970 1470 22015 1590
rect 22135 1470 22180 1590
rect 22300 1470 22345 1590
rect 22465 1470 22510 1590
rect 22630 1470 22675 1590
rect 22795 1470 22840 1590
rect 22960 1470 23005 1590
rect 23125 1470 23170 1590
rect 23290 1470 23335 1590
rect 23455 1470 23500 1590
rect 23620 1470 23665 1590
rect 23785 1470 23830 1590
rect 23950 1470 24240 1590
rect 24360 1470 24405 1590
rect 24525 1470 24570 1590
rect 24690 1470 24735 1590
rect 24855 1470 24900 1590
rect 25020 1470 25065 1590
rect 25185 1470 25230 1590
rect 25350 1470 25395 1590
rect 25515 1470 25560 1590
rect 25680 1470 25725 1590
rect 25845 1470 25890 1590
rect 26010 1470 26055 1590
rect 26175 1470 26220 1590
rect 26340 1470 26385 1590
rect 26505 1470 26550 1590
rect 26670 1470 26715 1590
rect 26835 1470 26880 1590
rect 27000 1470 27045 1590
rect 27165 1470 27210 1590
rect 27330 1470 27375 1590
rect 27495 1470 27540 1590
rect 27660 1470 27705 1590
rect 27825 1470 27870 1590
rect 27990 1470 28035 1590
rect 28155 1470 28200 1590
rect 28320 1470 28365 1590
rect 28485 1470 28530 1590
rect 28650 1470 28695 1590
rect 28815 1470 28860 1590
rect 28980 1470 29025 1590
rect 29145 1470 29190 1590
rect 29310 1470 29355 1590
rect 29475 1470 29520 1590
rect 29640 1470 29705 1590
rect 7105 1455 29705 1470
rect 12635 1450 12795 1455
rect 18325 1450 18485 1455
rect 24015 1450 24175 1455
rect 7105 1380 12635 1405
rect 7105 1260 7130 1380
rect 7250 1260 7305 1380
rect 7425 1260 7470 1380
rect 7590 1260 7635 1380
rect 7755 1260 7800 1380
rect 7920 1260 7975 1380
rect 8095 1260 8140 1380
rect 8260 1260 8305 1380
rect 8425 1260 8470 1380
rect 8590 1260 8645 1380
rect 8765 1260 8810 1380
rect 8930 1260 8975 1380
rect 9095 1260 9140 1380
rect 9260 1260 9315 1380
rect 9435 1260 9480 1380
rect 9600 1260 9645 1380
rect 9765 1260 9810 1380
rect 9930 1260 9985 1380
rect 10105 1260 10150 1380
rect 10270 1260 10315 1380
rect 10435 1260 10480 1380
rect 10600 1260 10655 1380
rect 10775 1260 10820 1380
rect 10940 1260 10985 1380
rect 11105 1260 11150 1380
rect 11270 1260 11325 1380
rect 11445 1260 11490 1380
rect 11610 1260 11655 1380
rect 11775 1260 11820 1380
rect 11940 1260 11995 1380
rect 12115 1260 12160 1380
rect 12280 1260 12325 1380
rect 12445 1260 12490 1380
rect 12610 1260 12635 1380
rect 7105 1215 12635 1260
rect 7105 1095 7130 1215
rect 7250 1095 7305 1215
rect 7425 1095 7470 1215
rect 7590 1095 7635 1215
rect 7755 1095 7800 1215
rect 7920 1095 7975 1215
rect 8095 1095 8140 1215
rect 8260 1095 8305 1215
rect 8425 1095 8470 1215
rect 8590 1095 8645 1215
rect 8765 1095 8810 1215
rect 8930 1095 8975 1215
rect 9095 1095 9140 1215
rect 9260 1095 9315 1215
rect 9435 1095 9480 1215
rect 9600 1095 9645 1215
rect 9765 1095 9810 1215
rect 9930 1095 9985 1215
rect 10105 1095 10150 1215
rect 10270 1095 10315 1215
rect 10435 1095 10480 1215
rect 10600 1095 10655 1215
rect 10775 1095 10820 1215
rect 10940 1095 10985 1215
rect 11105 1095 11150 1215
rect 11270 1095 11325 1215
rect 11445 1095 11490 1215
rect 11610 1095 11655 1215
rect 11775 1095 11820 1215
rect 11940 1095 11995 1215
rect 12115 1095 12160 1215
rect 12280 1095 12325 1215
rect 12445 1095 12490 1215
rect 12610 1095 12635 1215
rect 7105 1050 12635 1095
rect 7105 930 7130 1050
rect 7250 930 7305 1050
rect 7425 930 7470 1050
rect 7590 930 7635 1050
rect 7755 930 7800 1050
rect 7920 930 7975 1050
rect 8095 930 8140 1050
rect 8260 930 8305 1050
rect 8425 930 8470 1050
rect 8590 930 8645 1050
rect 8765 930 8810 1050
rect 8930 930 8975 1050
rect 9095 930 9140 1050
rect 9260 930 9315 1050
rect 9435 930 9480 1050
rect 9600 930 9645 1050
rect 9765 930 9810 1050
rect 9930 930 9985 1050
rect 10105 930 10150 1050
rect 10270 930 10315 1050
rect 10435 930 10480 1050
rect 10600 930 10655 1050
rect 10775 930 10820 1050
rect 10940 930 10985 1050
rect 11105 930 11150 1050
rect 11270 930 11325 1050
rect 11445 930 11490 1050
rect 11610 930 11655 1050
rect 11775 930 11820 1050
rect 11940 930 11995 1050
rect 12115 930 12160 1050
rect 12280 930 12325 1050
rect 12445 930 12490 1050
rect 12610 930 12635 1050
rect 7105 885 12635 930
rect 7105 765 7130 885
rect 7250 765 7305 885
rect 7425 765 7470 885
rect 7590 765 7635 885
rect 7755 765 7800 885
rect 7920 765 7975 885
rect 8095 765 8140 885
rect 8260 765 8305 885
rect 8425 765 8470 885
rect 8590 765 8645 885
rect 8765 765 8810 885
rect 8930 765 8975 885
rect 9095 765 9140 885
rect 9260 765 9315 885
rect 9435 765 9480 885
rect 9600 765 9645 885
rect 9765 765 9810 885
rect 9930 765 9985 885
rect 10105 765 10150 885
rect 10270 765 10315 885
rect 10435 765 10480 885
rect 10600 765 10655 885
rect 10775 765 10820 885
rect 10940 765 10985 885
rect 11105 765 11150 885
rect 11270 765 11325 885
rect 11445 765 11490 885
rect 11610 765 11655 885
rect 11775 765 11820 885
rect 11940 765 11995 885
rect 12115 765 12160 885
rect 12280 765 12325 885
rect 12445 765 12490 885
rect 12610 765 12635 885
rect 7105 710 12635 765
rect 7105 590 7130 710
rect 7250 590 7305 710
rect 7425 590 7470 710
rect 7590 590 7635 710
rect 7755 590 7800 710
rect 7920 590 7975 710
rect 8095 590 8140 710
rect 8260 590 8305 710
rect 8425 590 8470 710
rect 8590 590 8645 710
rect 8765 590 8810 710
rect 8930 590 8975 710
rect 9095 590 9140 710
rect 9260 590 9315 710
rect 9435 590 9480 710
rect 9600 590 9645 710
rect 9765 590 9810 710
rect 9930 590 9985 710
rect 10105 590 10150 710
rect 10270 590 10315 710
rect 10435 590 10480 710
rect 10600 590 10655 710
rect 10775 590 10820 710
rect 10940 590 10985 710
rect 11105 590 11150 710
rect 11270 590 11325 710
rect 11445 590 11490 710
rect 11610 590 11655 710
rect 11775 590 11820 710
rect 11940 590 11995 710
rect 12115 590 12160 710
rect 12280 590 12325 710
rect 12445 590 12490 710
rect 12610 590 12635 710
rect 7105 545 12635 590
rect 7105 425 7130 545
rect 7250 425 7305 545
rect 7425 425 7470 545
rect 7590 425 7635 545
rect 7755 425 7800 545
rect 7920 425 7975 545
rect 8095 425 8140 545
rect 8260 425 8305 545
rect 8425 425 8470 545
rect 8590 425 8645 545
rect 8765 425 8810 545
rect 8930 425 8975 545
rect 9095 425 9140 545
rect 9260 425 9315 545
rect 9435 425 9480 545
rect 9600 425 9645 545
rect 9765 425 9810 545
rect 9930 425 9985 545
rect 10105 425 10150 545
rect 10270 425 10315 545
rect 10435 425 10480 545
rect 10600 425 10655 545
rect 10775 425 10820 545
rect 10940 425 10985 545
rect 11105 425 11150 545
rect 11270 425 11325 545
rect 11445 425 11490 545
rect 11610 425 11655 545
rect 11775 425 11820 545
rect 11940 425 11995 545
rect 12115 425 12160 545
rect 12280 425 12325 545
rect 12445 425 12490 545
rect 12610 425 12635 545
rect 7105 380 12635 425
rect 7105 260 7130 380
rect 7250 260 7305 380
rect 7425 260 7470 380
rect 7590 260 7635 380
rect 7755 260 7800 380
rect 7920 260 7975 380
rect 8095 260 8140 380
rect 8260 260 8305 380
rect 8425 260 8470 380
rect 8590 260 8645 380
rect 8765 260 8810 380
rect 8930 260 8975 380
rect 9095 260 9140 380
rect 9260 260 9315 380
rect 9435 260 9480 380
rect 9600 260 9645 380
rect 9765 260 9810 380
rect 9930 260 9985 380
rect 10105 260 10150 380
rect 10270 260 10315 380
rect 10435 260 10480 380
rect 10600 260 10655 380
rect 10775 260 10820 380
rect 10940 260 10985 380
rect 11105 260 11150 380
rect 11270 260 11325 380
rect 11445 260 11490 380
rect 11610 260 11655 380
rect 11775 260 11820 380
rect 11940 260 11995 380
rect 12115 260 12160 380
rect 12280 260 12325 380
rect 12445 260 12490 380
rect 12610 260 12635 380
rect 7105 215 12635 260
rect 7105 95 7130 215
rect 7250 95 7305 215
rect 7425 95 7470 215
rect 7590 95 7635 215
rect 7755 95 7800 215
rect 7920 95 7975 215
rect 8095 95 8140 215
rect 8260 95 8305 215
rect 8425 95 8470 215
rect 8590 95 8645 215
rect 8765 95 8810 215
rect 8930 95 8975 215
rect 9095 95 9140 215
rect 9260 95 9315 215
rect 9435 95 9480 215
rect 9600 95 9645 215
rect 9765 95 9810 215
rect 9930 95 9985 215
rect 10105 95 10150 215
rect 10270 95 10315 215
rect 10435 95 10480 215
rect 10600 95 10655 215
rect 10775 95 10820 215
rect 10940 95 10985 215
rect 11105 95 11150 215
rect 11270 95 11325 215
rect 11445 95 11490 215
rect 11610 95 11655 215
rect 11775 95 11820 215
rect 11940 95 11995 215
rect 12115 95 12160 215
rect 12280 95 12325 215
rect 12445 95 12490 215
rect 12610 95 12635 215
rect 7105 40 12635 95
rect 7105 -80 7130 40
rect 7250 -80 7305 40
rect 7425 -80 7470 40
rect 7590 -80 7635 40
rect 7755 -80 7800 40
rect 7920 -80 7975 40
rect 8095 -80 8140 40
rect 8260 -80 8305 40
rect 8425 -80 8470 40
rect 8590 -80 8645 40
rect 8765 -80 8810 40
rect 8930 -80 8975 40
rect 9095 -80 9140 40
rect 9260 -80 9315 40
rect 9435 -80 9480 40
rect 9600 -80 9645 40
rect 9765 -80 9810 40
rect 9930 -80 9985 40
rect 10105 -80 10150 40
rect 10270 -80 10315 40
rect 10435 -80 10480 40
rect 10600 -80 10655 40
rect 10775 -80 10820 40
rect 10940 -80 10985 40
rect 11105 -80 11150 40
rect 11270 -80 11325 40
rect 11445 -80 11490 40
rect 11610 -80 11655 40
rect 11775 -80 11820 40
rect 11940 -80 11995 40
rect 12115 -80 12160 40
rect 12280 -80 12325 40
rect 12445 -80 12490 40
rect 12610 -80 12635 40
rect 7105 -125 12635 -80
rect 7105 -245 7130 -125
rect 7250 -245 7305 -125
rect 7425 -245 7470 -125
rect 7590 -245 7635 -125
rect 7755 -245 7800 -125
rect 7920 -245 7975 -125
rect 8095 -245 8140 -125
rect 8260 -245 8305 -125
rect 8425 -245 8470 -125
rect 8590 -245 8645 -125
rect 8765 -245 8810 -125
rect 8930 -245 8975 -125
rect 9095 -245 9140 -125
rect 9260 -245 9315 -125
rect 9435 -245 9480 -125
rect 9600 -245 9645 -125
rect 9765 -245 9810 -125
rect 9930 -245 9985 -125
rect 10105 -245 10150 -125
rect 10270 -245 10315 -125
rect 10435 -245 10480 -125
rect 10600 -245 10655 -125
rect 10775 -245 10820 -125
rect 10940 -245 10985 -125
rect 11105 -245 11150 -125
rect 11270 -245 11325 -125
rect 11445 -245 11490 -125
rect 11610 -245 11655 -125
rect 11775 -245 11820 -125
rect 11940 -245 11995 -125
rect 12115 -245 12160 -125
rect 12280 -245 12325 -125
rect 12445 -245 12490 -125
rect 12610 -245 12635 -125
rect 7105 -290 12635 -245
rect 7105 -410 7130 -290
rect 7250 -410 7305 -290
rect 7425 -410 7470 -290
rect 7590 -410 7635 -290
rect 7755 -410 7800 -290
rect 7920 -410 7975 -290
rect 8095 -410 8140 -290
rect 8260 -410 8305 -290
rect 8425 -410 8470 -290
rect 8590 -410 8645 -290
rect 8765 -410 8810 -290
rect 8930 -410 8975 -290
rect 9095 -410 9140 -290
rect 9260 -410 9315 -290
rect 9435 -410 9480 -290
rect 9600 -410 9645 -290
rect 9765 -410 9810 -290
rect 9930 -410 9985 -290
rect 10105 -410 10150 -290
rect 10270 -410 10315 -290
rect 10435 -410 10480 -290
rect 10600 -410 10655 -290
rect 10775 -410 10820 -290
rect 10940 -410 10985 -290
rect 11105 -410 11150 -290
rect 11270 -410 11325 -290
rect 11445 -410 11490 -290
rect 11610 -410 11655 -290
rect 11775 -410 11820 -290
rect 11940 -410 11995 -290
rect 12115 -410 12160 -290
rect 12280 -410 12325 -290
rect 12445 -410 12490 -290
rect 12610 -410 12635 -290
rect 7105 -455 12635 -410
rect 7105 -575 7130 -455
rect 7250 -575 7305 -455
rect 7425 -575 7470 -455
rect 7590 -575 7635 -455
rect 7755 -575 7800 -455
rect 7920 -575 7975 -455
rect 8095 -575 8140 -455
rect 8260 -575 8305 -455
rect 8425 -575 8470 -455
rect 8590 -575 8645 -455
rect 8765 -575 8810 -455
rect 8930 -575 8975 -455
rect 9095 -575 9140 -455
rect 9260 -575 9315 -455
rect 9435 -575 9480 -455
rect 9600 -575 9645 -455
rect 9765 -575 9810 -455
rect 9930 -575 9985 -455
rect 10105 -575 10150 -455
rect 10270 -575 10315 -455
rect 10435 -575 10480 -455
rect 10600 -575 10655 -455
rect 10775 -575 10820 -455
rect 10940 -575 10985 -455
rect 11105 -575 11150 -455
rect 11270 -575 11325 -455
rect 11445 -575 11490 -455
rect 11610 -575 11655 -455
rect 11775 -575 11820 -455
rect 11940 -575 11995 -455
rect 12115 -575 12160 -455
rect 12280 -575 12325 -455
rect 12445 -575 12490 -455
rect 12610 -575 12635 -455
rect 7105 -630 12635 -575
rect 7105 -750 7130 -630
rect 7250 -750 7305 -630
rect 7425 -750 7470 -630
rect 7590 -750 7635 -630
rect 7755 -750 7800 -630
rect 7920 -750 7975 -630
rect 8095 -750 8140 -630
rect 8260 -750 8305 -630
rect 8425 -750 8470 -630
rect 8590 -750 8645 -630
rect 8765 -750 8810 -630
rect 8930 -750 8975 -630
rect 9095 -750 9140 -630
rect 9260 -750 9315 -630
rect 9435 -750 9480 -630
rect 9600 -750 9645 -630
rect 9765 -750 9810 -630
rect 9930 -750 9985 -630
rect 10105 -750 10150 -630
rect 10270 -750 10315 -630
rect 10435 -750 10480 -630
rect 10600 -750 10655 -630
rect 10775 -750 10820 -630
rect 10940 -750 10985 -630
rect 11105 -750 11150 -630
rect 11270 -750 11325 -630
rect 11445 -750 11490 -630
rect 11610 -750 11655 -630
rect 11775 -750 11820 -630
rect 11940 -750 11995 -630
rect 12115 -750 12160 -630
rect 12280 -750 12325 -630
rect 12445 -750 12490 -630
rect 12610 -750 12635 -630
rect 7105 -795 12635 -750
rect 7105 -915 7130 -795
rect 7250 -915 7305 -795
rect 7425 -915 7470 -795
rect 7590 -915 7635 -795
rect 7755 -915 7800 -795
rect 7920 -915 7975 -795
rect 8095 -915 8140 -795
rect 8260 -915 8305 -795
rect 8425 -915 8470 -795
rect 8590 -915 8645 -795
rect 8765 -915 8810 -795
rect 8930 -915 8975 -795
rect 9095 -915 9140 -795
rect 9260 -915 9315 -795
rect 9435 -915 9480 -795
rect 9600 -915 9645 -795
rect 9765 -915 9810 -795
rect 9930 -915 9985 -795
rect 10105 -915 10150 -795
rect 10270 -915 10315 -795
rect 10435 -915 10480 -795
rect 10600 -915 10655 -795
rect 10775 -915 10820 -795
rect 10940 -915 10985 -795
rect 11105 -915 11150 -795
rect 11270 -915 11325 -795
rect 11445 -915 11490 -795
rect 11610 -915 11655 -795
rect 11775 -915 11820 -795
rect 11940 -915 11995 -795
rect 12115 -915 12160 -795
rect 12280 -915 12325 -795
rect 12445 -915 12490 -795
rect 12610 -915 12635 -795
rect 7105 -960 12635 -915
rect 7105 -1080 7130 -960
rect 7250 -1080 7305 -960
rect 7425 -1080 7470 -960
rect 7590 -1080 7635 -960
rect 7755 -1080 7800 -960
rect 7920 -1080 7975 -960
rect 8095 -1080 8140 -960
rect 8260 -1080 8305 -960
rect 8425 -1080 8470 -960
rect 8590 -1080 8645 -960
rect 8765 -1080 8810 -960
rect 8930 -1080 8975 -960
rect 9095 -1080 9140 -960
rect 9260 -1080 9315 -960
rect 9435 -1080 9480 -960
rect 9600 -1080 9645 -960
rect 9765 -1080 9810 -960
rect 9930 -1080 9985 -960
rect 10105 -1080 10150 -960
rect 10270 -1080 10315 -960
rect 10435 -1080 10480 -960
rect 10600 -1080 10655 -960
rect 10775 -1080 10820 -960
rect 10940 -1080 10985 -960
rect 11105 -1080 11150 -960
rect 11270 -1080 11325 -960
rect 11445 -1080 11490 -960
rect 11610 -1080 11655 -960
rect 11775 -1080 11820 -960
rect 11940 -1080 11995 -960
rect 12115 -1080 12160 -960
rect 12280 -1080 12325 -960
rect 12445 -1080 12490 -960
rect 12610 -1080 12635 -960
rect 7105 -1125 12635 -1080
rect 7105 -1245 7130 -1125
rect 7250 -1245 7305 -1125
rect 7425 -1245 7470 -1125
rect 7590 -1245 7635 -1125
rect 7755 -1245 7800 -1125
rect 7920 -1245 7975 -1125
rect 8095 -1245 8140 -1125
rect 8260 -1245 8305 -1125
rect 8425 -1245 8470 -1125
rect 8590 -1245 8645 -1125
rect 8765 -1245 8810 -1125
rect 8930 -1245 8975 -1125
rect 9095 -1245 9140 -1125
rect 9260 -1245 9315 -1125
rect 9435 -1245 9480 -1125
rect 9600 -1245 9645 -1125
rect 9765 -1245 9810 -1125
rect 9930 -1245 9985 -1125
rect 10105 -1245 10150 -1125
rect 10270 -1245 10315 -1125
rect 10435 -1245 10480 -1125
rect 10600 -1245 10655 -1125
rect 10775 -1245 10820 -1125
rect 10940 -1245 10985 -1125
rect 11105 -1245 11150 -1125
rect 11270 -1245 11325 -1125
rect 11445 -1245 11490 -1125
rect 11610 -1245 11655 -1125
rect 11775 -1245 11820 -1125
rect 11940 -1245 11995 -1125
rect 12115 -1245 12160 -1125
rect 12280 -1245 12325 -1125
rect 12445 -1245 12490 -1125
rect 12610 -1245 12635 -1125
rect 7105 -1300 12635 -1245
rect 7105 -1420 7130 -1300
rect 7250 -1420 7305 -1300
rect 7425 -1420 7470 -1300
rect 7590 -1420 7635 -1300
rect 7755 -1420 7800 -1300
rect 7920 -1420 7975 -1300
rect 8095 -1420 8140 -1300
rect 8260 -1420 8305 -1300
rect 8425 -1420 8470 -1300
rect 8590 -1420 8645 -1300
rect 8765 -1420 8810 -1300
rect 8930 -1420 8975 -1300
rect 9095 -1420 9140 -1300
rect 9260 -1420 9315 -1300
rect 9435 -1420 9480 -1300
rect 9600 -1420 9645 -1300
rect 9765 -1420 9810 -1300
rect 9930 -1420 9985 -1300
rect 10105 -1420 10150 -1300
rect 10270 -1420 10315 -1300
rect 10435 -1420 10480 -1300
rect 10600 -1420 10655 -1300
rect 10775 -1420 10820 -1300
rect 10940 -1420 10985 -1300
rect 11105 -1420 11150 -1300
rect 11270 -1420 11325 -1300
rect 11445 -1420 11490 -1300
rect 11610 -1420 11655 -1300
rect 11775 -1420 11820 -1300
rect 11940 -1420 11995 -1300
rect 12115 -1420 12160 -1300
rect 12280 -1420 12325 -1300
rect 12445 -1420 12490 -1300
rect 12610 -1420 12635 -1300
rect 7105 -1465 12635 -1420
rect 7105 -1585 7130 -1465
rect 7250 -1585 7305 -1465
rect 7425 -1585 7470 -1465
rect 7590 -1585 7635 -1465
rect 7755 -1585 7800 -1465
rect 7920 -1585 7975 -1465
rect 8095 -1585 8140 -1465
rect 8260 -1585 8305 -1465
rect 8425 -1585 8470 -1465
rect 8590 -1585 8645 -1465
rect 8765 -1585 8810 -1465
rect 8930 -1585 8975 -1465
rect 9095 -1585 9140 -1465
rect 9260 -1585 9315 -1465
rect 9435 -1585 9480 -1465
rect 9600 -1585 9645 -1465
rect 9765 -1585 9810 -1465
rect 9930 -1585 9985 -1465
rect 10105 -1585 10150 -1465
rect 10270 -1585 10315 -1465
rect 10435 -1585 10480 -1465
rect 10600 -1585 10655 -1465
rect 10775 -1585 10820 -1465
rect 10940 -1585 10985 -1465
rect 11105 -1585 11150 -1465
rect 11270 -1585 11325 -1465
rect 11445 -1585 11490 -1465
rect 11610 -1585 11655 -1465
rect 11775 -1585 11820 -1465
rect 11940 -1585 11995 -1465
rect 12115 -1585 12160 -1465
rect 12280 -1585 12325 -1465
rect 12445 -1585 12490 -1465
rect 12610 -1585 12635 -1465
rect 7105 -1630 12635 -1585
rect 7105 -1750 7130 -1630
rect 7250 -1750 7305 -1630
rect 7425 -1750 7470 -1630
rect 7590 -1750 7635 -1630
rect 7755 -1750 7800 -1630
rect 7920 -1750 7975 -1630
rect 8095 -1750 8140 -1630
rect 8260 -1750 8305 -1630
rect 8425 -1750 8470 -1630
rect 8590 -1750 8645 -1630
rect 8765 -1750 8810 -1630
rect 8930 -1750 8975 -1630
rect 9095 -1750 9140 -1630
rect 9260 -1750 9315 -1630
rect 9435 -1750 9480 -1630
rect 9600 -1750 9645 -1630
rect 9765 -1750 9810 -1630
rect 9930 -1750 9985 -1630
rect 10105 -1750 10150 -1630
rect 10270 -1750 10315 -1630
rect 10435 -1750 10480 -1630
rect 10600 -1750 10655 -1630
rect 10775 -1750 10820 -1630
rect 10940 -1750 10985 -1630
rect 11105 -1750 11150 -1630
rect 11270 -1750 11325 -1630
rect 11445 -1750 11490 -1630
rect 11610 -1750 11655 -1630
rect 11775 -1750 11820 -1630
rect 11940 -1750 11995 -1630
rect 12115 -1750 12160 -1630
rect 12280 -1750 12325 -1630
rect 12445 -1750 12490 -1630
rect 12610 -1750 12635 -1630
rect 7105 -1795 12635 -1750
rect 7105 -1915 7130 -1795
rect 7250 -1915 7305 -1795
rect 7425 -1915 7470 -1795
rect 7590 -1915 7635 -1795
rect 7755 -1915 7800 -1795
rect 7920 -1915 7975 -1795
rect 8095 -1915 8140 -1795
rect 8260 -1915 8305 -1795
rect 8425 -1915 8470 -1795
rect 8590 -1915 8645 -1795
rect 8765 -1915 8810 -1795
rect 8930 -1915 8975 -1795
rect 9095 -1915 9140 -1795
rect 9260 -1915 9315 -1795
rect 9435 -1915 9480 -1795
rect 9600 -1915 9645 -1795
rect 9765 -1915 9810 -1795
rect 9930 -1915 9985 -1795
rect 10105 -1915 10150 -1795
rect 10270 -1915 10315 -1795
rect 10435 -1915 10480 -1795
rect 10600 -1915 10655 -1795
rect 10775 -1915 10820 -1795
rect 10940 -1915 10985 -1795
rect 11105 -1915 11150 -1795
rect 11270 -1915 11325 -1795
rect 11445 -1915 11490 -1795
rect 11610 -1915 11655 -1795
rect 11775 -1915 11820 -1795
rect 11940 -1915 11995 -1795
rect 12115 -1915 12160 -1795
rect 12280 -1915 12325 -1795
rect 12445 -1915 12490 -1795
rect 12610 -1915 12635 -1795
rect 7105 -1970 12635 -1915
rect 7105 -2090 7130 -1970
rect 7250 -2090 7305 -1970
rect 7425 -2090 7470 -1970
rect 7590 -2090 7635 -1970
rect 7755 -2090 7800 -1970
rect 7920 -2090 7975 -1970
rect 8095 -2090 8140 -1970
rect 8260 -2090 8305 -1970
rect 8425 -2090 8470 -1970
rect 8590 -2090 8645 -1970
rect 8765 -2090 8810 -1970
rect 8930 -2090 8975 -1970
rect 9095 -2090 9140 -1970
rect 9260 -2090 9315 -1970
rect 9435 -2090 9480 -1970
rect 9600 -2090 9645 -1970
rect 9765 -2090 9810 -1970
rect 9930 -2090 9985 -1970
rect 10105 -2090 10150 -1970
rect 10270 -2090 10315 -1970
rect 10435 -2090 10480 -1970
rect 10600 -2090 10655 -1970
rect 10775 -2090 10820 -1970
rect 10940 -2090 10985 -1970
rect 11105 -2090 11150 -1970
rect 11270 -2090 11325 -1970
rect 11445 -2090 11490 -1970
rect 11610 -2090 11655 -1970
rect 11775 -2090 11820 -1970
rect 11940 -2090 11995 -1970
rect 12115 -2090 12160 -1970
rect 12280 -2090 12325 -1970
rect 12445 -2090 12490 -1970
rect 12610 -2090 12635 -1970
rect 7105 -2135 12635 -2090
rect 7105 -2255 7130 -2135
rect 7250 -2255 7305 -2135
rect 7425 -2255 7470 -2135
rect 7590 -2255 7635 -2135
rect 7755 -2255 7800 -2135
rect 7920 -2255 7975 -2135
rect 8095 -2255 8140 -2135
rect 8260 -2255 8305 -2135
rect 8425 -2255 8470 -2135
rect 8590 -2255 8645 -2135
rect 8765 -2255 8810 -2135
rect 8930 -2255 8975 -2135
rect 9095 -2255 9140 -2135
rect 9260 -2255 9315 -2135
rect 9435 -2255 9480 -2135
rect 9600 -2255 9645 -2135
rect 9765 -2255 9810 -2135
rect 9930 -2255 9985 -2135
rect 10105 -2255 10150 -2135
rect 10270 -2255 10315 -2135
rect 10435 -2255 10480 -2135
rect 10600 -2255 10655 -2135
rect 10775 -2255 10820 -2135
rect 10940 -2255 10985 -2135
rect 11105 -2255 11150 -2135
rect 11270 -2255 11325 -2135
rect 11445 -2255 11490 -2135
rect 11610 -2255 11655 -2135
rect 11775 -2255 11820 -2135
rect 11940 -2255 11995 -2135
rect 12115 -2255 12160 -2135
rect 12280 -2255 12325 -2135
rect 12445 -2255 12490 -2135
rect 12610 -2255 12635 -2135
rect 7105 -2300 12635 -2255
rect 7105 -2420 7130 -2300
rect 7250 -2420 7305 -2300
rect 7425 -2420 7470 -2300
rect 7590 -2420 7635 -2300
rect 7755 -2420 7800 -2300
rect 7920 -2420 7975 -2300
rect 8095 -2420 8140 -2300
rect 8260 -2420 8305 -2300
rect 8425 -2420 8470 -2300
rect 8590 -2420 8645 -2300
rect 8765 -2420 8810 -2300
rect 8930 -2420 8975 -2300
rect 9095 -2420 9140 -2300
rect 9260 -2420 9315 -2300
rect 9435 -2420 9480 -2300
rect 9600 -2420 9645 -2300
rect 9765 -2420 9810 -2300
rect 9930 -2420 9985 -2300
rect 10105 -2420 10150 -2300
rect 10270 -2420 10315 -2300
rect 10435 -2420 10480 -2300
rect 10600 -2420 10655 -2300
rect 10775 -2420 10820 -2300
rect 10940 -2420 10985 -2300
rect 11105 -2420 11150 -2300
rect 11270 -2420 11325 -2300
rect 11445 -2420 11490 -2300
rect 11610 -2420 11655 -2300
rect 11775 -2420 11820 -2300
rect 11940 -2420 11995 -2300
rect 12115 -2420 12160 -2300
rect 12280 -2420 12325 -2300
rect 12445 -2420 12490 -2300
rect 12610 -2420 12635 -2300
rect 7105 -2465 12635 -2420
rect 7105 -2585 7130 -2465
rect 7250 -2585 7305 -2465
rect 7425 -2585 7470 -2465
rect 7590 -2585 7635 -2465
rect 7755 -2585 7800 -2465
rect 7920 -2585 7975 -2465
rect 8095 -2585 8140 -2465
rect 8260 -2585 8305 -2465
rect 8425 -2585 8470 -2465
rect 8590 -2585 8645 -2465
rect 8765 -2585 8810 -2465
rect 8930 -2585 8975 -2465
rect 9095 -2585 9140 -2465
rect 9260 -2585 9315 -2465
rect 9435 -2585 9480 -2465
rect 9600 -2585 9645 -2465
rect 9765 -2585 9810 -2465
rect 9930 -2585 9985 -2465
rect 10105 -2585 10150 -2465
rect 10270 -2585 10315 -2465
rect 10435 -2585 10480 -2465
rect 10600 -2585 10655 -2465
rect 10775 -2585 10820 -2465
rect 10940 -2585 10985 -2465
rect 11105 -2585 11150 -2465
rect 11270 -2585 11325 -2465
rect 11445 -2585 11490 -2465
rect 11610 -2585 11655 -2465
rect 11775 -2585 11820 -2465
rect 11940 -2585 11995 -2465
rect 12115 -2585 12160 -2465
rect 12280 -2585 12325 -2465
rect 12445 -2585 12490 -2465
rect 12610 -2585 12635 -2465
rect 7105 -2640 12635 -2585
rect 7105 -2760 7130 -2640
rect 7250 -2760 7305 -2640
rect 7425 -2760 7470 -2640
rect 7590 -2760 7635 -2640
rect 7755 -2760 7800 -2640
rect 7920 -2760 7975 -2640
rect 8095 -2760 8140 -2640
rect 8260 -2760 8305 -2640
rect 8425 -2760 8470 -2640
rect 8590 -2760 8645 -2640
rect 8765 -2760 8810 -2640
rect 8930 -2760 8975 -2640
rect 9095 -2760 9140 -2640
rect 9260 -2760 9315 -2640
rect 9435 -2760 9480 -2640
rect 9600 -2760 9645 -2640
rect 9765 -2760 9810 -2640
rect 9930 -2760 9985 -2640
rect 10105 -2760 10150 -2640
rect 10270 -2760 10315 -2640
rect 10435 -2760 10480 -2640
rect 10600 -2760 10655 -2640
rect 10775 -2760 10820 -2640
rect 10940 -2760 10985 -2640
rect 11105 -2760 11150 -2640
rect 11270 -2760 11325 -2640
rect 11445 -2760 11490 -2640
rect 11610 -2760 11655 -2640
rect 11775 -2760 11820 -2640
rect 11940 -2760 11995 -2640
rect 12115 -2760 12160 -2640
rect 12280 -2760 12325 -2640
rect 12445 -2760 12490 -2640
rect 12610 -2760 12635 -2640
rect 7105 -2805 12635 -2760
rect 7105 -2925 7130 -2805
rect 7250 -2925 7305 -2805
rect 7425 -2925 7470 -2805
rect 7590 -2925 7635 -2805
rect 7755 -2925 7800 -2805
rect 7920 -2925 7975 -2805
rect 8095 -2925 8140 -2805
rect 8260 -2925 8305 -2805
rect 8425 -2925 8470 -2805
rect 8590 -2925 8645 -2805
rect 8765 -2925 8810 -2805
rect 8930 -2925 8975 -2805
rect 9095 -2925 9140 -2805
rect 9260 -2925 9315 -2805
rect 9435 -2925 9480 -2805
rect 9600 -2925 9645 -2805
rect 9765 -2925 9810 -2805
rect 9930 -2925 9985 -2805
rect 10105 -2925 10150 -2805
rect 10270 -2925 10315 -2805
rect 10435 -2925 10480 -2805
rect 10600 -2925 10655 -2805
rect 10775 -2925 10820 -2805
rect 10940 -2925 10985 -2805
rect 11105 -2925 11150 -2805
rect 11270 -2925 11325 -2805
rect 11445 -2925 11490 -2805
rect 11610 -2925 11655 -2805
rect 11775 -2925 11820 -2805
rect 11940 -2925 11995 -2805
rect 12115 -2925 12160 -2805
rect 12280 -2925 12325 -2805
rect 12445 -2925 12490 -2805
rect 12610 -2925 12635 -2805
rect 7105 -2970 12635 -2925
rect 7105 -3090 7130 -2970
rect 7250 -3090 7305 -2970
rect 7425 -3090 7470 -2970
rect 7590 -3090 7635 -2970
rect 7755 -3090 7800 -2970
rect 7920 -3090 7975 -2970
rect 8095 -3090 8140 -2970
rect 8260 -3090 8305 -2970
rect 8425 -3090 8470 -2970
rect 8590 -3090 8645 -2970
rect 8765 -3090 8810 -2970
rect 8930 -3090 8975 -2970
rect 9095 -3090 9140 -2970
rect 9260 -3090 9315 -2970
rect 9435 -3090 9480 -2970
rect 9600 -3090 9645 -2970
rect 9765 -3090 9810 -2970
rect 9930 -3090 9985 -2970
rect 10105 -3090 10150 -2970
rect 10270 -3090 10315 -2970
rect 10435 -3090 10480 -2970
rect 10600 -3090 10655 -2970
rect 10775 -3090 10820 -2970
rect 10940 -3090 10985 -2970
rect 11105 -3090 11150 -2970
rect 11270 -3090 11325 -2970
rect 11445 -3090 11490 -2970
rect 11610 -3090 11655 -2970
rect 11775 -3090 11820 -2970
rect 11940 -3090 11995 -2970
rect 12115 -3090 12160 -2970
rect 12280 -3090 12325 -2970
rect 12445 -3090 12490 -2970
rect 12610 -3090 12635 -2970
rect 7105 -3135 12635 -3090
rect 7105 -3255 7130 -3135
rect 7250 -3255 7305 -3135
rect 7425 -3255 7470 -3135
rect 7590 -3255 7635 -3135
rect 7755 -3255 7800 -3135
rect 7920 -3255 7975 -3135
rect 8095 -3255 8140 -3135
rect 8260 -3255 8305 -3135
rect 8425 -3255 8470 -3135
rect 8590 -3255 8645 -3135
rect 8765 -3255 8810 -3135
rect 8930 -3255 8975 -3135
rect 9095 -3255 9140 -3135
rect 9260 -3255 9315 -3135
rect 9435 -3255 9480 -3135
rect 9600 -3255 9645 -3135
rect 9765 -3255 9810 -3135
rect 9930 -3255 9985 -3135
rect 10105 -3255 10150 -3135
rect 10270 -3255 10315 -3135
rect 10435 -3255 10480 -3135
rect 10600 -3255 10655 -3135
rect 10775 -3255 10820 -3135
rect 10940 -3255 10985 -3135
rect 11105 -3255 11150 -3135
rect 11270 -3255 11325 -3135
rect 11445 -3255 11490 -3135
rect 11610 -3255 11655 -3135
rect 11775 -3255 11820 -3135
rect 11940 -3255 11995 -3135
rect 12115 -3255 12160 -3135
rect 12280 -3255 12325 -3135
rect 12445 -3255 12490 -3135
rect 12610 -3255 12635 -3135
rect 7105 -3310 12635 -3255
rect 7105 -3430 7130 -3310
rect 7250 -3430 7305 -3310
rect 7425 -3430 7470 -3310
rect 7590 -3430 7635 -3310
rect 7755 -3430 7800 -3310
rect 7920 -3430 7975 -3310
rect 8095 -3430 8140 -3310
rect 8260 -3430 8305 -3310
rect 8425 -3430 8470 -3310
rect 8590 -3430 8645 -3310
rect 8765 -3430 8810 -3310
rect 8930 -3430 8975 -3310
rect 9095 -3430 9140 -3310
rect 9260 -3430 9315 -3310
rect 9435 -3430 9480 -3310
rect 9600 -3430 9645 -3310
rect 9765 -3430 9810 -3310
rect 9930 -3430 9985 -3310
rect 10105 -3430 10150 -3310
rect 10270 -3430 10315 -3310
rect 10435 -3430 10480 -3310
rect 10600 -3430 10655 -3310
rect 10775 -3430 10820 -3310
rect 10940 -3430 10985 -3310
rect 11105 -3430 11150 -3310
rect 11270 -3430 11325 -3310
rect 11445 -3430 11490 -3310
rect 11610 -3430 11655 -3310
rect 11775 -3430 11820 -3310
rect 11940 -3430 11995 -3310
rect 12115 -3430 12160 -3310
rect 12280 -3430 12325 -3310
rect 12445 -3430 12490 -3310
rect 12610 -3430 12635 -3310
rect 7105 -3475 12635 -3430
rect 7105 -3595 7130 -3475
rect 7250 -3595 7305 -3475
rect 7425 -3595 7470 -3475
rect 7590 -3595 7635 -3475
rect 7755 -3595 7800 -3475
rect 7920 -3595 7975 -3475
rect 8095 -3595 8140 -3475
rect 8260 -3595 8305 -3475
rect 8425 -3595 8470 -3475
rect 8590 -3595 8645 -3475
rect 8765 -3595 8810 -3475
rect 8930 -3595 8975 -3475
rect 9095 -3595 9140 -3475
rect 9260 -3595 9315 -3475
rect 9435 -3595 9480 -3475
rect 9600 -3595 9645 -3475
rect 9765 -3595 9810 -3475
rect 9930 -3595 9985 -3475
rect 10105 -3595 10150 -3475
rect 10270 -3595 10315 -3475
rect 10435 -3595 10480 -3475
rect 10600 -3595 10655 -3475
rect 10775 -3595 10820 -3475
rect 10940 -3595 10985 -3475
rect 11105 -3595 11150 -3475
rect 11270 -3595 11325 -3475
rect 11445 -3595 11490 -3475
rect 11610 -3595 11655 -3475
rect 11775 -3595 11820 -3475
rect 11940 -3595 11995 -3475
rect 12115 -3595 12160 -3475
rect 12280 -3595 12325 -3475
rect 12445 -3595 12490 -3475
rect 12610 -3595 12635 -3475
rect 7105 -3640 12635 -3595
rect 7105 -3760 7130 -3640
rect 7250 -3760 7305 -3640
rect 7425 -3760 7470 -3640
rect 7590 -3760 7635 -3640
rect 7755 -3760 7800 -3640
rect 7920 -3760 7975 -3640
rect 8095 -3760 8140 -3640
rect 8260 -3760 8305 -3640
rect 8425 -3760 8470 -3640
rect 8590 -3760 8645 -3640
rect 8765 -3760 8810 -3640
rect 8930 -3760 8975 -3640
rect 9095 -3760 9140 -3640
rect 9260 -3760 9315 -3640
rect 9435 -3760 9480 -3640
rect 9600 -3760 9645 -3640
rect 9765 -3760 9810 -3640
rect 9930 -3760 9985 -3640
rect 10105 -3760 10150 -3640
rect 10270 -3760 10315 -3640
rect 10435 -3760 10480 -3640
rect 10600 -3760 10655 -3640
rect 10775 -3760 10820 -3640
rect 10940 -3760 10985 -3640
rect 11105 -3760 11150 -3640
rect 11270 -3760 11325 -3640
rect 11445 -3760 11490 -3640
rect 11610 -3760 11655 -3640
rect 11775 -3760 11820 -3640
rect 11940 -3760 11995 -3640
rect 12115 -3760 12160 -3640
rect 12280 -3760 12325 -3640
rect 12445 -3760 12490 -3640
rect 12610 -3760 12635 -3640
rect 7105 -3805 12635 -3760
rect 7105 -3925 7130 -3805
rect 7250 -3925 7305 -3805
rect 7425 -3925 7470 -3805
rect 7590 -3925 7635 -3805
rect 7755 -3925 7800 -3805
rect 7920 -3925 7975 -3805
rect 8095 -3925 8140 -3805
rect 8260 -3925 8305 -3805
rect 8425 -3925 8470 -3805
rect 8590 -3925 8645 -3805
rect 8765 -3925 8810 -3805
rect 8930 -3925 8975 -3805
rect 9095 -3925 9140 -3805
rect 9260 -3925 9315 -3805
rect 9435 -3925 9480 -3805
rect 9600 -3925 9645 -3805
rect 9765 -3925 9810 -3805
rect 9930 -3925 9985 -3805
rect 10105 -3925 10150 -3805
rect 10270 -3925 10315 -3805
rect 10435 -3925 10480 -3805
rect 10600 -3925 10655 -3805
rect 10775 -3925 10820 -3805
rect 10940 -3925 10985 -3805
rect 11105 -3925 11150 -3805
rect 11270 -3925 11325 -3805
rect 11445 -3925 11490 -3805
rect 11610 -3925 11655 -3805
rect 11775 -3925 11820 -3805
rect 11940 -3925 11995 -3805
rect 12115 -3925 12160 -3805
rect 12280 -3925 12325 -3805
rect 12445 -3925 12490 -3805
rect 12610 -3925 12635 -3805
rect 7105 -3980 12635 -3925
rect 7105 -4100 7130 -3980
rect 7250 -4100 7305 -3980
rect 7425 -4100 7470 -3980
rect 7590 -4100 7635 -3980
rect 7755 -4100 7800 -3980
rect 7920 -4100 7975 -3980
rect 8095 -4100 8140 -3980
rect 8260 -4100 8305 -3980
rect 8425 -4100 8470 -3980
rect 8590 -4100 8645 -3980
rect 8765 -4100 8810 -3980
rect 8930 -4100 8975 -3980
rect 9095 -4100 9140 -3980
rect 9260 -4100 9315 -3980
rect 9435 -4100 9480 -3980
rect 9600 -4100 9645 -3980
rect 9765 -4100 9810 -3980
rect 9930 -4100 9985 -3980
rect 10105 -4100 10150 -3980
rect 10270 -4100 10315 -3980
rect 10435 -4100 10480 -3980
rect 10600 -4100 10655 -3980
rect 10775 -4100 10820 -3980
rect 10940 -4100 10985 -3980
rect 11105 -4100 11150 -3980
rect 11270 -4100 11325 -3980
rect 11445 -4100 11490 -3980
rect 11610 -4100 11655 -3980
rect 11775 -4100 11820 -3980
rect 11940 -4100 11995 -3980
rect 12115 -4100 12160 -3980
rect 12280 -4100 12325 -3980
rect 12445 -4100 12490 -3980
rect 12610 -4065 12635 -3980
rect 12795 1380 18325 1405
rect 12795 1260 12820 1380
rect 12940 1260 12995 1380
rect 13115 1260 13160 1380
rect 13280 1260 13325 1380
rect 13445 1260 13490 1380
rect 13610 1260 13665 1380
rect 13785 1260 13830 1380
rect 13950 1260 13995 1380
rect 14115 1260 14160 1380
rect 14280 1260 14335 1380
rect 14455 1260 14500 1380
rect 14620 1260 14665 1380
rect 14785 1260 14830 1380
rect 14950 1260 15005 1380
rect 15125 1260 15170 1380
rect 15290 1260 15335 1380
rect 15455 1260 15500 1380
rect 15620 1260 15675 1380
rect 15795 1260 15840 1380
rect 15960 1260 16005 1380
rect 16125 1260 16170 1380
rect 16290 1260 16345 1380
rect 16465 1260 16510 1380
rect 16630 1260 16675 1380
rect 16795 1260 16840 1380
rect 16960 1260 17015 1380
rect 17135 1260 17180 1380
rect 17300 1260 17345 1380
rect 17465 1260 17510 1380
rect 17630 1260 17685 1380
rect 17805 1260 17850 1380
rect 17970 1260 18015 1380
rect 18135 1260 18180 1380
rect 18300 1260 18325 1380
rect 12795 1215 18325 1260
rect 12795 1095 12820 1215
rect 12940 1095 12995 1215
rect 13115 1095 13160 1215
rect 13280 1095 13325 1215
rect 13445 1095 13490 1215
rect 13610 1095 13665 1215
rect 13785 1095 13830 1215
rect 13950 1095 13995 1215
rect 14115 1095 14160 1215
rect 14280 1095 14335 1215
rect 14455 1095 14500 1215
rect 14620 1095 14665 1215
rect 14785 1095 14830 1215
rect 14950 1095 15005 1215
rect 15125 1095 15170 1215
rect 15290 1095 15335 1215
rect 15455 1095 15500 1215
rect 15620 1095 15675 1215
rect 15795 1095 15840 1215
rect 15960 1095 16005 1215
rect 16125 1095 16170 1215
rect 16290 1095 16345 1215
rect 16465 1095 16510 1215
rect 16630 1095 16675 1215
rect 16795 1095 16840 1215
rect 16960 1095 17015 1215
rect 17135 1095 17180 1215
rect 17300 1095 17345 1215
rect 17465 1095 17510 1215
rect 17630 1095 17685 1215
rect 17805 1095 17850 1215
rect 17970 1095 18015 1215
rect 18135 1095 18180 1215
rect 18300 1095 18325 1215
rect 12795 1050 18325 1095
rect 12795 930 12820 1050
rect 12940 930 12995 1050
rect 13115 930 13160 1050
rect 13280 930 13325 1050
rect 13445 930 13490 1050
rect 13610 930 13665 1050
rect 13785 930 13830 1050
rect 13950 930 13995 1050
rect 14115 930 14160 1050
rect 14280 930 14335 1050
rect 14455 930 14500 1050
rect 14620 930 14665 1050
rect 14785 930 14830 1050
rect 14950 930 15005 1050
rect 15125 930 15170 1050
rect 15290 930 15335 1050
rect 15455 930 15500 1050
rect 15620 930 15675 1050
rect 15795 930 15840 1050
rect 15960 930 16005 1050
rect 16125 930 16170 1050
rect 16290 930 16345 1050
rect 16465 930 16510 1050
rect 16630 930 16675 1050
rect 16795 930 16840 1050
rect 16960 930 17015 1050
rect 17135 930 17180 1050
rect 17300 930 17345 1050
rect 17465 930 17510 1050
rect 17630 930 17685 1050
rect 17805 930 17850 1050
rect 17970 930 18015 1050
rect 18135 930 18180 1050
rect 18300 930 18325 1050
rect 12795 885 18325 930
rect 12795 765 12820 885
rect 12940 765 12995 885
rect 13115 765 13160 885
rect 13280 765 13325 885
rect 13445 765 13490 885
rect 13610 765 13665 885
rect 13785 765 13830 885
rect 13950 765 13995 885
rect 14115 765 14160 885
rect 14280 765 14335 885
rect 14455 765 14500 885
rect 14620 765 14665 885
rect 14785 765 14830 885
rect 14950 765 15005 885
rect 15125 765 15170 885
rect 15290 765 15335 885
rect 15455 765 15500 885
rect 15620 765 15675 885
rect 15795 765 15840 885
rect 15960 765 16005 885
rect 16125 765 16170 885
rect 16290 765 16345 885
rect 16465 765 16510 885
rect 16630 765 16675 885
rect 16795 765 16840 885
rect 16960 765 17015 885
rect 17135 765 17180 885
rect 17300 765 17345 885
rect 17465 765 17510 885
rect 17630 765 17685 885
rect 17805 765 17850 885
rect 17970 765 18015 885
rect 18135 765 18180 885
rect 18300 765 18325 885
rect 12795 710 18325 765
rect 12795 590 12820 710
rect 12940 590 12995 710
rect 13115 590 13160 710
rect 13280 590 13325 710
rect 13445 590 13490 710
rect 13610 590 13665 710
rect 13785 590 13830 710
rect 13950 590 13995 710
rect 14115 590 14160 710
rect 14280 590 14335 710
rect 14455 590 14500 710
rect 14620 590 14665 710
rect 14785 590 14830 710
rect 14950 590 15005 710
rect 15125 590 15170 710
rect 15290 590 15335 710
rect 15455 590 15500 710
rect 15620 590 15675 710
rect 15795 590 15840 710
rect 15960 590 16005 710
rect 16125 590 16170 710
rect 16290 590 16345 710
rect 16465 590 16510 710
rect 16630 590 16675 710
rect 16795 590 16840 710
rect 16960 590 17015 710
rect 17135 590 17180 710
rect 17300 590 17345 710
rect 17465 590 17510 710
rect 17630 590 17685 710
rect 17805 590 17850 710
rect 17970 590 18015 710
rect 18135 590 18180 710
rect 18300 590 18325 710
rect 12795 545 18325 590
rect 12795 425 12820 545
rect 12940 425 12995 545
rect 13115 425 13160 545
rect 13280 425 13325 545
rect 13445 425 13490 545
rect 13610 425 13665 545
rect 13785 425 13830 545
rect 13950 425 13995 545
rect 14115 425 14160 545
rect 14280 425 14335 545
rect 14455 425 14500 545
rect 14620 425 14665 545
rect 14785 425 14830 545
rect 14950 425 15005 545
rect 15125 425 15170 545
rect 15290 425 15335 545
rect 15455 425 15500 545
rect 15620 425 15675 545
rect 15795 425 15840 545
rect 15960 425 16005 545
rect 16125 425 16170 545
rect 16290 425 16345 545
rect 16465 425 16510 545
rect 16630 425 16675 545
rect 16795 425 16840 545
rect 16960 425 17015 545
rect 17135 425 17180 545
rect 17300 425 17345 545
rect 17465 425 17510 545
rect 17630 425 17685 545
rect 17805 425 17850 545
rect 17970 425 18015 545
rect 18135 425 18180 545
rect 18300 425 18325 545
rect 12795 380 18325 425
rect 12795 260 12820 380
rect 12940 260 12995 380
rect 13115 260 13160 380
rect 13280 260 13325 380
rect 13445 260 13490 380
rect 13610 260 13665 380
rect 13785 260 13830 380
rect 13950 260 13995 380
rect 14115 260 14160 380
rect 14280 260 14335 380
rect 14455 260 14500 380
rect 14620 260 14665 380
rect 14785 260 14830 380
rect 14950 260 15005 380
rect 15125 260 15170 380
rect 15290 260 15335 380
rect 15455 260 15500 380
rect 15620 260 15675 380
rect 15795 260 15840 380
rect 15960 260 16005 380
rect 16125 260 16170 380
rect 16290 260 16345 380
rect 16465 260 16510 380
rect 16630 260 16675 380
rect 16795 260 16840 380
rect 16960 260 17015 380
rect 17135 260 17180 380
rect 17300 260 17345 380
rect 17465 260 17510 380
rect 17630 260 17685 380
rect 17805 260 17850 380
rect 17970 260 18015 380
rect 18135 260 18180 380
rect 18300 260 18325 380
rect 12795 215 18325 260
rect 12795 95 12820 215
rect 12940 95 12995 215
rect 13115 95 13160 215
rect 13280 95 13325 215
rect 13445 95 13490 215
rect 13610 95 13665 215
rect 13785 95 13830 215
rect 13950 95 13995 215
rect 14115 95 14160 215
rect 14280 95 14335 215
rect 14455 95 14500 215
rect 14620 95 14665 215
rect 14785 95 14830 215
rect 14950 95 15005 215
rect 15125 95 15170 215
rect 15290 95 15335 215
rect 15455 95 15500 215
rect 15620 95 15675 215
rect 15795 95 15840 215
rect 15960 95 16005 215
rect 16125 95 16170 215
rect 16290 95 16345 215
rect 16465 95 16510 215
rect 16630 95 16675 215
rect 16795 95 16840 215
rect 16960 95 17015 215
rect 17135 95 17180 215
rect 17300 95 17345 215
rect 17465 95 17510 215
rect 17630 95 17685 215
rect 17805 95 17850 215
rect 17970 95 18015 215
rect 18135 95 18180 215
rect 18300 95 18325 215
rect 12795 40 18325 95
rect 12795 -80 12820 40
rect 12940 -80 12995 40
rect 13115 -80 13160 40
rect 13280 -80 13325 40
rect 13445 -80 13490 40
rect 13610 -80 13665 40
rect 13785 -80 13830 40
rect 13950 -80 13995 40
rect 14115 -80 14160 40
rect 14280 -80 14335 40
rect 14455 -80 14500 40
rect 14620 -80 14665 40
rect 14785 -80 14830 40
rect 14950 -80 15005 40
rect 15125 -80 15170 40
rect 15290 -80 15335 40
rect 15455 -80 15500 40
rect 15620 -80 15675 40
rect 15795 -80 15840 40
rect 15960 -80 16005 40
rect 16125 -80 16170 40
rect 16290 -80 16345 40
rect 16465 -80 16510 40
rect 16630 -80 16675 40
rect 16795 -80 16840 40
rect 16960 -80 17015 40
rect 17135 -80 17180 40
rect 17300 -80 17345 40
rect 17465 -80 17510 40
rect 17630 -80 17685 40
rect 17805 -80 17850 40
rect 17970 -80 18015 40
rect 18135 -80 18180 40
rect 18300 -80 18325 40
rect 12795 -125 18325 -80
rect 12795 -245 12820 -125
rect 12940 -245 12995 -125
rect 13115 -245 13160 -125
rect 13280 -245 13325 -125
rect 13445 -245 13490 -125
rect 13610 -245 13665 -125
rect 13785 -245 13830 -125
rect 13950 -245 13995 -125
rect 14115 -245 14160 -125
rect 14280 -245 14335 -125
rect 14455 -245 14500 -125
rect 14620 -245 14665 -125
rect 14785 -245 14830 -125
rect 14950 -245 15005 -125
rect 15125 -245 15170 -125
rect 15290 -245 15335 -125
rect 15455 -245 15500 -125
rect 15620 -245 15675 -125
rect 15795 -245 15840 -125
rect 15960 -245 16005 -125
rect 16125 -245 16170 -125
rect 16290 -245 16345 -125
rect 16465 -245 16510 -125
rect 16630 -245 16675 -125
rect 16795 -245 16840 -125
rect 16960 -245 17015 -125
rect 17135 -245 17180 -125
rect 17300 -245 17345 -125
rect 17465 -245 17510 -125
rect 17630 -245 17685 -125
rect 17805 -245 17850 -125
rect 17970 -245 18015 -125
rect 18135 -245 18180 -125
rect 18300 -245 18325 -125
rect 12795 -290 18325 -245
rect 12795 -410 12820 -290
rect 12940 -410 12995 -290
rect 13115 -410 13160 -290
rect 13280 -410 13325 -290
rect 13445 -410 13490 -290
rect 13610 -410 13665 -290
rect 13785 -410 13830 -290
rect 13950 -410 13995 -290
rect 14115 -410 14160 -290
rect 14280 -410 14335 -290
rect 14455 -410 14500 -290
rect 14620 -410 14665 -290
rect 14785 -410 14830 -290
rect 14950 -410 15005 -290
rect 15125 -410 15170 -290
rect 15290 -410 15335 -290
rect 15455 -410 15500 -290
rect 15620 -410 15675 -290
rect 15795 -410 15840 -290
rect 15960 -410 16005 -290
rect 16125 -410 16170 -290
rect 16290 -410 16345 -290
rect 16465 -410 16510 -290
rect 16630 -410 16675 -290
rect 16795 -410 16840 -290
rect 16960 -410 17015 -290
rect 17135 -410 17180 -290
rect 17300 -410 17345 -290
rect 17465 -410 17510 -290
rect 17630 -410 17685 -290
rect 17805 -410 17850 -290
rect 17970 -410 18015 -290
rect 18135 -410 18180 -290
rect 18300 -410 18325 -290
rect 12795 -455 18325 -410
rect 12795 -575 12820 -455
rect 12940 -575 12995 -455
rect 13115 -575 13160 -455
rect 13280 -575 13325 -455
rect 13445 -575 13490 -455
rect 13610 -575 13665 -455
rect 13785 -575 13830 -455
rect 13950 -575 13995 -455
rect 14115 -575 14160 -455
rect 14280 -575 14335 -455
rect 14455 -575 14500 -455
rect 14620 -575 14665 -455
rect 14785 -575 14830 -455
rect 14950 -575 15005 -455
rect 15125 -575 15170 -455
rect 15290 -575 15335 -455
rect 15455 -575 15500 -455
rect 15620 -575 15675 -455
rect 15795 -575 15840 -455
rect 15960 -575 16005 -455
rect 16125 -575 16170 -455
rect 16290 -575 16345 -455
rect 16465 -575 16510 -455
rect 16630 -575 16675 -455
rect 16795 -575 16840 -455
rect 16960 -575 17015 -455
rect 17135 -575 17180 -455
rect 17300 -575 17345 -455
rect 17465 -575 17510 -455
rect 17630 -575 17685 -455
rect 17805 -575 17850 -455
rect 17970 -575 18015 -455
rect 18135 -575 18180 -455
rect 18300 -575 18325 -455
rect 12795 -630 18325 -575
rect 12795 -750 12820 -630
rect 12940 -750 12995 -630
rect 13115 -750 13160 -630
rect 13280 -750 13325 -630
rect 13445 -750 13490 -630
rect 13610 -750 13665 -630
rect 13785 -750 13830 -630
rect 13950 -750 13995 -630
rect 14115 -750 14160 -630
rect 14280 -750 14335 -630
rect 14455 -750 14500 -630
rect 14620 -750 14665 -630
rect 14785 -750 14830 -630
rect 14950 -750 15005 -630
rect 15125 -750 15170 -630
rect 15290 -750 15335 -630
rect 15455 -750 15500 -630
rect 15620 -750 15675 -630
rect 15795 -750 15840 -630
rect 15960 -750 16005 -630
rect 16125 -750 16170 -630
rect 16290 -750 16345 -630
rect 16465 -750 16510 -630
rect 16630 -750 16675 -630
rect 16795 -750 16840 -630
rect 16960 -750 17015 -630
rect 17135 -750 17180 -630
rect 17300 -750 17345 -630
rect 17465 -750 17510 -630
rect 17630 -750 17685 -630
rect 17805 -750 17850 -630
rect 17970 -750 18015 -630
rect 18135 -750 18180 -630
rect 18300 -750 18325 -630
rect 12795 -795 18325 -750
rect 12795 -915 12820 -795
rect 12940 -915 12995 -795
rect 13115 -915 13160 -795
rect 13280 -915 13325 -795
rect 13445 -915 13490 -795
rect 13610 -915 13665 -795
rect 13785 -915 13830 -795
rect 13950 -915 13995 -795
rect 14115 -915 14160 -795
rect 14280 -915 14335 -795
rect 14455 -915 14500 -795
rect 14620 -915 14665 -795
rect 14785 -915 14830 -795
rect 14950 -915 15005 -795
rect 15125 -915 15170 -795
rect 15290 -915 15335 -795
rect 15455 -915 15500 -795
rect 15620 -915 15675 -795
rect 15795 -915 15840 -795
rect 15960 -915 16005 -795
rect 16125 -915 16170 -795
rect 16290 -915 16345 -795
rect 16465 -915 16510 -795
rect 16630 -915 16675 -795
rect 16795 -915 16840 -795
rect 16960 -915 17015 -795
rect 17135 -915 17180 -795
rect 17300 -915 17345 -795
rect 17465 -915 17510 -795
rect 17630 -915 17685 -795
rect 17805 -915 17850 -795
rect 17970 -915 18015 -795
rect 18135 -915 18180 -795
rect 18300 -915 18325 -795
rect 12795 -960 18325 -915
rect 12795 -1080 12820 -960
rect 12940 -1080 12995 -960
rect 13115 -1080 13160 -960
rect 13280 -1080 13325 -960
rect 13445 -1080 13490 -960
rect 13610 -1080 13665 -960
rect 13785 -1080 13830 -960
rect 13950 -1080 13995 -960
rect 14115 -1080 14160 -960
rect 14280 -1080 14335 -960
rect 14455 -1080 14500 -960
rect 14620 -1080 14665 -960
rect 14785 -1080 14830 -960
rect 14950 -1080 15005 -960
rect 15125 -1080 15170 -960
rect 15290 -1080 15335 -960
rect 15455 -1080 15500 -960
rect 15620 -1080 15675 -960
rect 15795 -1080 15840 -960
rect 15960 -1080 16005 -960
rect 16125 -1080 16170 -960
rect 16290 -1080 16345 -960
rect 16465 -1080 16510 -960
rect 16630 -1080 16675 -960
rect 16795 -1080 16840 -960
rect 16960 -1080 17015 -960
rect 17135 -1080 17180 -960
rect 17300 -1080 17345 -960
rect 17465 -1080 17510 -960
rect 17630 -1080 17685 -960
rect 17805 -1080 17850 -960
rect 17970 -1080 18015 -960
rect 18135 -1080 18180 -960
rect 18300 -1080 18325 -960
rect 12795 -1125 18325 -1080
rect 12795 -1245 12820 -1125
rect 12940 -1245 12995 -1125
rect 13115 -1245 13160 -1125
rect 13280 -1245 13325 -1125
rect 13445 -1245 13490 -1125
rect 13610 -1245 13665 -1125
rect 13785 -1245 13830 -1125
rect 13950 -1245 13995 -1125
rect 14115 -1245 14160 -1125
rect 14280 -1245 14335 -1125
rect 14455 -1245 14500 -1125
rect 14620 -1245 14665 -1125
rect 14785 -1245 14830 -1125
rect 14950 -1245 15005 -1125
rect 15125 -1245 15170 -1125
rect 15290 -1245 15335 -1125
rect 15455 -1245 15500 -1125
rect 15620 -1245 15675 -1125
rect 15795 -1245 15840 -1125
rect 15960 -1245 16005 -1125
rect 16125 -1245 16170 -1125
rect 16290 -1245 16345 -1125
rect 16465 -1245 16510 -1125
rect 16630 -1245 16675 -1125
rect 16795 -1245 16840 -1125
rect 16960 -1245 17015 -1125
rect 17135 -1245 17180 -1125
rect 17300 -1245 17345 -1125
rect 17465 -1245 17510 -1125
rect 17630 -1245 17685 -1125
rect 17805 -1245 17850 -1125
rect 17970 -1245 18015 -1125
rect 18135 -1245 18180 -1125
rect 18300 -1245 18325 -1125
rect 12795 -1300 18325 -1245
rect 12795 -1420 12820 -1300
rect 12940 -1420 12995 -1300
rect 13115 -1420 13160 -1300
rect 13280 -1420 13325 -1300
rect 13445 -1420 13490 -1300
rect 13610 -1420 13665 -1300
rect 13785 -1420 13830 -1300
rect 13950 -1420 13995 -1300
rect 14115 -1420 14160 -1300
rect 14280 -1420 14335 -1300
rect 14455 -1420 14500 -1300
rect 14620 -1420 14665 -1300
rect 14785 -1420 14830 -1300
rect 14950 -1420 15005 -1300
rect 15125 -1420 15170 -1300
rect 15290 -1420 15335 -1300
rect 15455 -1420 15500 -1300
rect 15620 -1420 15675 -1300
rect 15795 -1420 15840 -1300
rect 15960 -1420 16005 -1300
rect 16125 -1420 16170 -1300
rect 16290 -1420 16345 -1300
rect 16465 -1420 16510 -1300
rect 16630 -1420 16675 -1300
rect 16795 -1420 16840 -1300
rect 16960 -1420 17015 -1300
rect 17135 -1420 17180 -1300
rect 17300 -1420 17345 -1300
rect 17465 -1420 17510 -1300
rect 17630 -1420 17685 -1300
rect 17805 -1420 17850 -1300
rect 17970 -1420 18015 -1300
rect 18135 -1420 18180 -1300
rect 18300 -1420 18325 -1300
rect 12795 -1465 18325 -1420
rect 12795 -1585 12820 -1465
rect 12940 -1585 12995 -1465
rect 13115 -1585 13160 -1465
rect 13280 -1585 13325 -1465
rect 13445 -1585 13490 -1465
rect 13610 -1585 13665 -1465
rect 13785 -1585 13830 -1465
rect 13950 -1585 13995 -1465
rect 14115 -1585 14160 -1465
rect 14280 -1585 14335 -1465
rect 14455 -1585 14500 -1465
rect 14620 -1585 14665 -1465
rect 14785 -1585 14830 -1465
rect 14950 -1585 15005 -1465
rect 15125 -1585 15170 -1465
rect 15290 -1585 15335 -1465
rect 15455 -1585 15500 -1465
rect 15620 -1585 15675 -1465
rect 15795 -1585 15840 -1465
rect 15960 -1585 16005 -1465
rect 16125 -1585 16170 -1465
rect 16290 -1585 16345 -1465
rect 16465 -1585 16510 -1465
rect 16630 -1585 16675 -1465
rect 16795 -1585 16840 -1465
rect 16960 -1585 17015 -1465
rect 17135 -1585 17180 -1465
rect 17300 -1585 17345 -1465
rect 17465 -1585 17510 -1465
rect 17630 -1585 17685 -1465
rect 17805 -1585 17850 -1465
rect 17970 -1585 18015 -1465
rect 18135 -1585 18180 -1465
rect 18300 -1585 18325 -1465
rect 12795 -1630 18325 -1585
rect 12795 -1750 12820 -1630
rect 12940 -1750 12995 -1630
rect 13115 -1750 13160 -1630
rect 13280 -1750 13325 -1630
rect 13445 -1750 13490 -1630
rect 13610 -1750 13665 -1630
rect 13785 -1750 13830 -1630
rect 13950 -1750 13995 -1630
rect 14115 -1750 14160 -1630
rect 14280 -1750 14335 -1630
rect 14455 -1750 14500 -1630
rect 14620 -1750 14665 -1630
rect 14785 -1750 14830 -1630
rect 14950 -1750 15005 -1630
rect 15125 -1750 15170 -1630
rect 15290 -1750 15335 -1630
rect 15455 -1750 15500 -1630
rect 15620 -1750 15675 -1630
rect 15795 -1750 15840 -1630
rect 15960 -1750 16005 -1630
rect 16125 -1750 16170 -1630
rect 16290 -1750 16345 -1630
rect 16465 -1750 16510 -1630
rect 16630 -1750 16675 -1630
rect 16795 -1750 16840 -1630
rect 16960 -1750 17015 -1630
rect 17135 -1750 17180 -1630
rect 17300 -1750 17345 -1630
rect 17465 -1750 17510 -1630
rect 17630 -1750 17685 -1630
rect 17805 -1750 17850 -1630
rect 17970 -1750 18015 -1630
rect 18135 -1750 18180 -1630
rect 18300 -1750 18325 -1630
rect 12795 -1795 18325 -1750
rect 12795 -1915 12820 -1795
rect 12940 -1915 12995 -1795
rect 13115 -1915 13160 -1795
rect 13280 -1915 13325 -1795
rect 13445 -1915 13490 -1795
rect 13610 -1915 13665 -1795
rect 13785 -1915 13830 -1795
rect 13950 -1915 13995 -1795
rect 14115 -1915 14160 -1795
rect 14280 -1915 14335 -1795
rect 14455 -1915 14500 -1795
rect 14620 -1915 14665 -1795
rect 14785 -1915 14830 -1795
rect 14950 -1915 15005 -1795
rect 15125 -1915 15170 -1795
rect 15290 -1915 15335 -1795
rect 15455 -1915 15500 -1795
rect 15620 -1915 15675 -1795
rect 15795 -1915 15840 -1795
rect 15960 -1915 16005 -1795
rect 16125 -1915 16170 -1795
rect 16290 -1915 16345 -1795
rect 16465 -1915 16510 -1795
rect 16630 -1915 16675 -1795
rect 16795 -1915 16840 -1795
rect 16960 -1915 17015 -1795
rect 17135 -1915 17180 -1795
rect 17300 -1915 17345 -1795
rect 17465 -1915 17510 -1795
rect 17630 -1915 17685 -1795
rect 17805 -1915 17850 -1795
rect 17970 -1915 18015 -1795
rect 18135 -1915 18180 -1795
rect 18300 -1915 18325 -1795
rect 12795 -1970 18325 -1915
rect 12795 -2090 12820 -1970
rect 12940 -2090 12995 -1970
rect 13115 -2090 13160 -1970
rect 13280 -2090 13325 -1970
rect 13445 -2090 13490 -1970
rect 13610 -2090 13665 -1970
rect 13785 -2090 13830 -1970
rect 13950 -2090 13995 -1970
rect 14115 -2090 14160 -1970
rect 14280 -2090 14335 -1970
rect 14455 -2090 14500 -1970
rect 14620 -2090 14665 -1970
rect 14785 -2090 14830 -1970
rect 14950 -2090 15005 -1970
rect 15125 -2090 15170 -1970
rect 15290 -2090 15335 -1970
rect 15455 -2090 15500 -1970
rect 15620 -2090 15675 -1970
rect 15795 -2090 15840 -1970
rect 15960 -2090 16005 -1970
rect 16125 -2090 16170 -1970
rect 16290 -2090 16345 -1970
rect 16465 -2090 16510 -1970
rect 16630 -2090 16675 -1970
rect 16795 -2090 16840 -1970
rect 16960 -2090 17015 -1970
rect 17135 -2090 17180 -1970
rect 17300 -2090 17345 -1970
rect 17465 -2090 17510 -1970
rect 17630 -2090 17685 -1970
rect 17805 -2090 17850 -1970
rect 17970 -2090 18015 -1970
rect 18135 -2090 18180 -1970
rect 18300 -2090 18325 -1970
rect 12795 -2135 18325 -2090
rect 12795 -2255 12820 -2135
rect 12940 -2255 12995 -2135
rect 13115 -2255 13160 -2135
rect 13280 -2255 13325 -2135
rect 13445 -2255 13490 -2135
rect 13610 -2255 13665 -2135
rect 13785 -2255 13830 -2135
rect 13950 -2255 13995 -2135
rect 14115 -2255 14160 -2135
rect 14280 -2255 14335 -2135
rect 14455 -2255 14500 -2135
rect 14620 -2255 14665 -2135
rect 14785 -2255 14830 -2135
rect 14950 -2255 15005 -2135
rect 15125 -2255 15170 -2135
rect 15290 -2255 15335 -2135
rect 15455 -2255 15500 -2135
rect 15620 -2255 15675 -2135
rect 15795 -2255 15840 -2135
rect 15960 -2255 16005 -2135
rect 16125 -2255 16170 -2135
rect 16290 -2255 16345 -2135
rect 16465 -2255 16510 -2135
rect 16630 -2255 16675 -2135
rect 16795 -2255 16840 -2135
rect 16960 -2255 17015 -2135
rect 17135 -2255 17180 -2135
rect 17300 -2255 17345 -2135
rect 17465 -2255 17510 -2135
rect 17630 -2255 17685 -2135
rect 17805 -2255 17850 -2135
rect 17970 -2255 18015 -2135
rect 18135 -2255 18180 -2135
rect 18300 -2255 18325 -2135
rect 12795 -2300 18325 -2255
rect 12795 -2420 12820 -2300
rect 12940 -2420 12995 -2300
rect 13115 -2420 13160 -2300
rect 13280 -2420 13325 -2300
rect 13445 -2420 13490 -2300
rect 13610 -2420 13665 -2300
rect 13785 -2420 13830 -2300
rect 13950 -2420 13995 -2300
rect 14115 -2420 14160 -2300
rect 14280 -2420 14335 -2300
rect 14455 -2420 14500 -2300
rect 14620 -2420 14665 -2300
rect 14785 -2420 14830 -2300
rect 14950 -2420 15005 -2300
rect 15125 -2420 15170 -2300
rect 15290 -2420 15335 -2300
rect 15455 -2420 15500 -2300
rect 15620 -2420 15675 -2300
rect 15795 -2420 15840 -2300
rect 15960 -2420 16005 -2300
rect 16125 -2420 16170 -2300
rect 16290 -2420 16345 -2300
rect 16465 -2420 16510 -2300
rect 16630 -2420 16675 -2300
rect 16795 -2420 16840 -2300
rect 16960 -2420 17015 -2300
rect 17135 -2420 17180 -2300
rect 17300 -2420 17345 -2300
rect 17465 -2420 17510 -2300
rect 17630 -2420 17685 -2300
rect 17805 -2420 17850 -2300
rect 17970 -2420 18015 -2300
rect 18135 -2420 18180 -2300
rect 18300 -2420 18325 -2300
rect 12795 -2465 18325 -2420
rect 12795 -2585 12820 -2465
rect 12940 -2585 12995 -2465
rect 13115 -2585 13160 -2465
rect 13280 -2585 13325 -2465
rect 13445 -2585 13490 -2465
rect 13610 -2585 13665 -2465
rect 13785 -2585 13830 -2465
rect 13950 -2585 13995 -2465
rect 14115 -2585 14160 -2465
rect 14280 -2585 14335 -2465
rect 14455 -2585 14500 -2465
rect 14620 -2585 14665 -2465
rect 14785 -2585 14830 -2465
rect 14950 -2585 15005 -2465
rect 15125 -2585 15170 -2465
rect 15290 -2585 15335 -2465
rect 15455 -2585 15500 -2465
rect 15620 -2585 15675 -2465
rect 15795 -2585 15840 -2465
rect 15960 -2585 16005 -2465
rect 16125 -2585 16170 -2465
rect 16290 -2585 16345 -2465
rect 16465 -2585 16510 -2465
rect 16630 -2585 16675 -2465
rect 16795 -2585 16840 -2465
rect 16960 -2585 17015 -2465
rect 17135 -2585 17180 -2465
rect 17300 -2585 17345 -2465
rect 17465 -2585 17510 -2465
rect 17630 -2585 17685 -2465
rect 17805 -2585 17850 -2465
rect 17970 -2585 18015 -2465
rect 18135 -2585 18180 -2465
rect 18300 -2585 18325 -2465
rect 12795 -2640 18325 -2585
rect 12795 -2760 12820 -2640
rect 12940 -2760 12995 -2640
rect 13115 -2760 13160 -2640
rect 13280 -2760 13325 -2640
rect 13445 -2760 13490 -2640
rect 13610 -2760 13665 -2640
rect 13785 -2760 13830 -2640
rect 13950 -2760 13995 -2640
rect 14115 -2760 14160 -2640
rect 14280 -2760 14335 -2640
rect 14455 -2760 14500 -2640
rect 14620 -2760 14665 -2640
rect 14785 -2760 14830 -2640
rect 14950 -2760 15005 -2640
rect 15125 -2760 15170 -2640
rect 15290 -2760 15335 -2640
rect 15455 -2760 15500 -2640
rect 15620 -2760 15675 -2640
rect 15795 -2760 15840 -2640
rect 15960 -2760 16005 -2640
rect 16125 -2760 16170 -2640
rect 16290 -2760 16345 -2640
rect 16465 -2760 16510 -2640
rect 16630 -2760 16675 -2640
rect 16795 -2760 16840 -2640
rect 16960 -2760 17015 -2640
rect 17135 -2760 17180 -2640
rect 17300 -2760 17345 -2640
rect 17465 -2760 17510 -2640
rect 17630 -2760 17685 -2640
rect 17805 -2760 17850 -2640
rect 17970 -2760 18015 -2640
rect 18135 -2760 18180 -2640
rect 18300 -2760 18325 -2640
rect 12795 -2805 18325 -2760
rect 12795 -2925 12820 -2805
rect 12940 -2925 12995 -2805
rect 13115 -2925 13160 -2805
rect 13280 -2925 13325 -2805
rect 13445 -2925 13490 -2805
rect 13610 -2925 13665 -2805
rect 13785 -2925 13830 -2805
rect 13950 -2925 13995 -2805
rect 14115 -2925 14160 -2805
rect 14280 -2925 14335 -2805
rect 14455 -2925 14500 -2805
rect 14620 -2925 14665 -2805
rect 14785 -2925 14830 -2805
rect 14950 -2925 15005 -2805
rect 15125 -2925 15170 -2805
rect 15290 -2925 15335 -2805
rect 15455 -2925 15500 -2805
rect 15620 -2925 15675 -2805
rect 15795 -2925 15840 -2805
rect 15960 -2925 16005 -2805
rect 16125 -2925 16170 -2805
rect 16290 -2925 16345 -2805
rect 16465 -2925 16510 -2805
rect 16630 -2925 16675 -2805
rect 16795 -2925 16840 -2805
rect 16960 -2925 17015 -2805
rect 17135 -2925 17180 -2805
rect 17300 -2925 17345 -2805
rect 17465 -2925 17510 -2805
rect 17630 -2925 17685 -2805
rect 17805 -2925 17850 -2805
rect 17970 -2925 18015 -2805
rect 18135 -2925 18180 -2805
rect 18300 -2925 18325 -2805
rect 12795 -2970 18325 -2925
rect 12795 -3090 12820 -2970
rect 12940 -3090 12995 -2970
rect 13115 -3090 13160 -2970
rect 13280 -3090 13325 -2970
rect 13445 -3090 13490 -2970
rect 13610 -3090 13665 -2970
rect 13785 -3090 13830 -2970
rect 13950 -3090 13995 -2970
rect 14115 -3090 14160 -2970
rect 14280 -3090 14335 -2970
rect 14455 -3090 14500 -2970
rect 14620 -3090 14665 -2970
rect 14785 -3090 14830 -2970
rect 14950 -3090 15005 -2970
rect 15125 -3090 15170 -2970
rect 15290 -3090 15335 -2970
rect 15455 -3090 15500 -2970
rect 15620 -3090 15675 -2970
rect 15795 -3090 15840 -2970
rect 15960 -3090 16005 -2970
rect 16125 -3090 16170 -2970
rect 16290 -3090 16345 -2970
rect 16465 -3090 16510 -2970
rect 16630 -3090 16675 -2970
rect 16795 -3090 16840 -2970
rect 16960 -3090 17015 -2970
rect 17135 -3090 17180 -2970
rect 17300 -3090 17345 -2970
rect 17465 -3090 17510 -2970
rect 17630 -3090 17685 -2970
rect 17805 -3090 17850 -2970
rect 17970 -3090 18015 -2970
rect 18135 -3090 18180 -2970
rect 18300 -3090 18325 -2970
rect 12795 -3135 18325 -3090
rect 12795 -3255 12820 -3135
rect 12940 -3255 12995 -3135
rect 13115 -3255 13160 -3135
rect 13280 -3255 13325 -3135
rect 13445 -3255 13490 -3135
rect 13610 -3255 13665 -3135
rect 13785 -3255 13830 -3135
rect 13950 -3255 13995 -3135
rect 14115 -3255 14160 -3135
rect 14280 -3255 14335 -3135
rect 14455 -3255 14500 -3135
rect 14620 -3255 14665 -3135
rect 14785 -3255 14830 -3135
rect 14950 -3255 15005 -3135
rect 15125 -3255 15170 -3135
rect 15290 -3255 15335 -3135
rect 15455 -3255 15500 -3135
rect 15620 -3255 15675 -3135
rect 15795 -3255 15840 -3135
rect 15960 -3255 16005 -3135
rect 16125 -3255 16170 -3135
rect 16290 -3255 16345 -3135
rect 16465 -3255 16510 -3135
rect 16630 -3255 16675 -3135
rect 16795 -3255 16840 -3135
rect 16960 -3255 17015 -3135
rect 17135 -3255 17180 -3135
rect 17300 -3255 17345 -3135
rect 17465 -3255 17510 -3135
rect 17630 -3255 17685 -3135
rect 17805 -3255 17850 -3135
rect 17970 -3255 18015 -3135
rect 18135 -3255 18180 -3135
rect 18300 -3255 18325 -3135
rect 12795 -3310 18325 -3255
rect 12795 -3430 12820 -3310
rect 12940 -3430 12995 -3310
rect 13115 -3430 13160 -3310
rect 13280 -3430 13325 -3310
rect 13445 -3430 13490 -3310
rect 13610 -3430 13665 -3310
rect 13785 -3430 13830 -3310
rect 13950 -3430 13995 -3310
rect 14115 -3430 14160 -3310
rect 14280 -3430 14335 -3310
rect 14455 -3430 14500 -3310
rect 14620 -3430 14665 -3310
rect 14785 -3430 14830 -3310
rect 14950 -3430 15005 -3310
rect 15125 -3430 15170 -3310
rect 15290 -3430 15335 -3310
rect 15455 -3430 15500 -3310
rect 15620 -3430 15675 -3310
rect 15795 -3430 15840 -3310
rect 15960 -3430 16005 -3310
rect 16125 -3430 16170 -3310
rect 16290 -3430 16345 -3310
rect 16465 -3430 16510 -3310
rect 16630 -3430 16675 -3310
rect 16795 -3430 16840 -3310
rect 16960 -3430 17015 -3310
rect 17135 -3430 17180 -3310
rect 17300 -3430 17345 -3310
rect 17465 -3430 17510 -3310
rect 17630 -3430 17685 -3310
rect 17805 -3430 17850 -3310
rect 17970 -3430 18015 -3310
rect 18135 -3430 18180 -3310
rect 18300 -3430 18325 -3310
rect 12795 -3475 18325 -3430
rect 12795 -3595 12820 -3475
rect 12940 -3595 12995 -3475
rect 13115 -3595 13160 -3475
rect 13280 -3595 13325 -3475
rect 13445 -3595 13490 -3475
rect 13610 -3595 13665 -3475
rect 13785 -3595 13830 -3475
rect 13950 -3595 13995 -3475
rect 14115 -3595 14160 -3475
rect 14280 -3595 14335 -3475
rect 14455 -3595 14500 -3475
rect 14620 -3595 14665 -3475
rect 14785 -3595 14830 -3475
rect 14950 -3595 15005 -3475
rect 15125 -3595 15170 -3475
rect 15290 -3595 15335 -3475
rect 15455 -3595 15500 -3475
rect 15620 -3595 15675 -3475
rect 15795 -3595 15840 -3475
rect 15960 -3595 16005 -3475
rect 16125 -3595 16170 -3475
rect 16290 -3595 16345 -3475
rect 16465 -3595 16510 -3475
rect 16630 -3595 16675 -3475
rect 16795 -3595 16840 -3475
rect 16960 -3595 17015 -3475
rect 17135 -3595 17180 -3475
rect 17300 -3595 17345 -3475
rect 17465 -3595 17510 -3475
rect 17630 -3595 17685 -3475
rect 17805 -3595 17850 -3475
rect 17970 -3595 18015 -3475
rect 18135 -3595 18180 -3475
rect 18300 -3595 18325 -3475
rect 12795 -3640 18325 -3595
rect 12795 -3760 12820 -3640
rect 12940 -3760 12995 -3640
rect 13115 -3760 13160 -3640
rect 13280 -3760 13325 -3640
rect 13445 -3760 13490 -3640
rect 13610 -3760 13665 -3640
rect 13785 -3760 13830 -3640
rect 13950 -3760 13995 -3640
rect 14115 -3760 14160 -3640
rect 14280 -3760 14335 -3640
rect 14455 -3760 14500 -3640
rect 14620 -3760 14665 -3640
rect 14785 -3760 14830 -3640
rect 14950 -3760 15005 -3640
rect 15125 -3760 15170 -3640
rect 15290 -3760 15335 -3640
rect 15455 -3760 15500 -3640
rect 15620 -3760 15675 -3640
rect 15795 -3760 15840 -3640
rect 15960 -3760 16005 -3640
rect 16125 -3760 16170 -3640
rect 16290 -3760 16345 -3640
rect 16465 -3760 16510 -3640
rect 16630 -3760 16675 -3640
rect 16795 -3760 16840 -3640
rect 16960 -3760 17015 -3640
rect 17135 -3760 17180 -3640
rect 17300 -3760 17345 -3640
rect 17465 -3760 17510 -3640
rect 17630 -3760 17685 -3640
rect 17805 -3760 17850 -3640
rect 17970 -3760 18015 -3640
rect 18135 -3760 18180 -3640
rect 18300 -3760 18325 -3640
rect 12795 -3805 18325 -3760
rect 12795 -3925 12820 -3805
rect 12940 -3925 12995 -3805
rect 13115 -3925 13160 -3805
rect 13280 -3925 13325 -3805
rect 13445 -3925 13490 -3805
rect 13610 -3925 13665 -3805
rect 13785 -3925 13830 -3805
rect 13950 -3925 13995 -3805
rect 14115 -3925 14160 -3805
rect 14280 -3925 14335 -3805
rect 14455 -3925 14500 -3805
rect 14620 -3925 14665 -3805
rect 14785 -3925 14830 -3805
rect 14950 -3925 15005 -3805
rect 15125 -3925 15170 -3805
rect 15290 -3925 15335 -3805
rect 15455 -3925 15500 -3805
rect 15620 -3925 15675 -3805
rect 15795 -3925 15840 -3805
rect 15960 -3925 16005 -3805
rect 16125 -3925 16170 -3805
rect 16290 -3925 16345 -3805
rect 16465 -3925 16510 -3805
rect 16630 -3925 16675 -3805
rect 16795 -3925 16840 -3805
rect 16960 -3925 17015 -3805
rect 17135 -3925 17180 -3805
rect 17300 -3925 17345 -3805
rect 17465 -3925 17510 -3805
rect 17630 -3925 17685 -3805
rect 17805 -3925 17850 -3805
rect 17970 -3925 18015 -3805
rect 18135 -3925 18180 -3805
rect 18300 -3925 18325 -3805
rect 12795 -3980 18325 -3925
rect 12795 -4065 12820 -3980
rect 12610 -4100 12820 -4065
rect 12940 -4100 12995 -3980
rect 13115 -4100 13160 -3980
rect 13280 -4100 13325 -3980
rect 13445 -4100 13490 -3980
rect 13610 -4100 13665 -3980
rect 13785 -4100 13830 -3980
rect 13950 -4100 13995 -3980
rect 14115 -4100 14160 -3980
rect 14280 -4100 14335 -3980
rect 14455 -4100 14500 -3980
rect 14620 -4100 14665 -3980
rect 14785 -4100 14830 -3980
rect 14950 -4100 15005 -3980
rect 15125 -4100 15170 -3980
rect 15290 -4100 15335 -3980
rect 15455 -4100 15500 -3980
rect 15620 -4100 15675 -3980
rect 15795 -4100 15840 -3980
rect 15960 -4100 16005 -3980
rect 16125 -4100 16170 -3980
rect 16290 -4100 16345 -3980
rect 16465 -4100 16510 -3980
rect 16630 -4100 16675 -3980
rect 16795 -4100 16840 -3980
rect 16960 -4100 17015 -3980
rect 17135 -4100 17180 -3980
rect 17300 -4100 17345 -3980
rect 17465 -4100 17510 -3980
rect 17630 -4100 17685 -3980
rect 17805 -4100 17850 -3980
rect 17970 -4100 18015 -3980
rect 18135 -4100 18180 -3980
rect 18300 -4065 18325 -3980
rect 18485 1380 24015 1405
rect 18485 1260 18510 1380
rect 18630 1260 18685 1380
rect 18805 1260 18850 1380
rect 18970 1260 19015 1380
rect 19135 1260 19180 1380
rect 19300 1260 19355 1380
rect 19475 1260 19520 1380
rect 19640 1260 19685 1380
rect 19805 1260 19850 1380
rect 19970 1260 20025 1380
rect 20145 1260 20190 1380
rect 20310 1260 20355 1380
rect 20475 1260 20520 1380
rect 20640 1260 20695 1380
rect 20815 1260 20860 1380
rect 20980 1260 21025 1380
rect 21145 1260 21190 1380
rect 21310 1260 21365 1380
rect 21485 1260 21530 1380
rect 21650 1260 21695 1380
rect 21815 1260 21860 1380
rect 21980 1260 22035 1380
rect 22155 1260 22200 1380
rect 22320 1260 22365 1380
rect 22485 1260 22530 1380
rect 22650 1260 22705 1380
rect 22825 1260 22870 1380
rect 22990 1260 23035 1380
rect 23155 1260 23200 1380
rect 23320 1260 23375 1380
rect 23495 1260 23540 1380
rect 23660 1260 23705 1380
rect 23825 1260 23870 1380
rect 23990 1260 24015 1380
rect 18485 1215 24015 1260
rect 18485 1095 18510 1215
rect 18630 1095 18685 1215
rect 18805 1095 18850 1215
rect 18970 1095 19015 1215
rect 19135 1095 19180 1215
rect 19300 1095 19355 1215
rect 19475 1095 19520 1215
rect 19640 1095 19685 1215
rect 19805 1095 19850 1215
rect 19970 1095 20025 1215
rect 20145 1095 20190 1215
rect 20310 1095 20355 1215
rect 20475 1095 20520 1215
rect 20640 1095 20695 1215
rect 20815 1095 20860 1215
rect 20980 1095 21025 1215
rect 21145 1095 21190 1215
rect 21310 1095 21365 1215
rect 21485 1095 21530 1215
rect 21650 1095 21695 1215
rect 21815 1095 21860 1215
rect 21980 1095 22035 1215
rect 22155 1095 22200 1215
rect 22320 1095 22365 1215
rect 22485 1095 22530 1215
rect 22650 1095 22705 1215
rect 22825 1095 22870 1215
rect 22990 1095 23035 1215
rect 23155 1095 23200 1215
rect 23320 1095 23375 1215
rect 23495 1095 23540 1215
rect 23660 1095 23705 1215
rect 23825 1095 23870 1215
rect 23990 1095 24015 1215
rect 18485 1050 24015 1095
rect 18485 930 18510 1050
rect 18630 930 18685 1050
rect 18805 930 18850 1050
rect 18970 930 19015 1050
rect 19135 930 19180 1050
rect 19300 930 19355 1050
rect 19475 930 19520 1050
rect 19640 930 19685 1050
rect 19805 930 19850 1050
rect 19970 930 20025 1050
rect 20145 930 20190 1050
rect 20310 930 20355 1050
rect 20475 930 20520 1050
rect 20640 930 20695 1050
rect 20815 930 20860 1050
rect 20980 930 21025 1050
rect 21145 930 21190 1050
rect 21310 930 21365 1050
rect 21485 930 21530 1050
rect 21650 930 21695 1050
rect 21815 930 21860 1050
rect 21980 930 22035 1050
rect 22155 930 22200 1050
rect 22320 930 22365 1050
rect 22485 930 22530 1050
rect 22650 930 22705 1050
rect 22825 930 22870 1050
rect 22990 930 23035 1050
rect 23155 930 23200 1050
rect 23320 930 23375 1050
rect 23495 930 23540 1050
rect 23660 930 23705 1050
rect 23825 930 23870 1050
rect 23990 930 24015 1050
rect 18485 885 24015 930
rect 18485 765 18510 885
rect 18630 765 18685 885
rect 18805 765 18850 885
rect 18970 765 19015 885
rect 19135 765 19180 885
rect 19300 765 19355 885
rect 19475 765 19520 885
rect 19640 765 19685 885
rect 19805 765 19850 885
rect 19970 765 20025 885
rect 20145 765 20190 885
rect 20310 765 20355 885
rect 20475 765 20520 885
rect 20640 765 20695 885
rect 20815 765 20860 885
rect 20980 765 21025 885
rect 21145 765 21190 885
rect 21310 765 21365 885
rect 21485 765 21530 885
rect 21650 765 21695 885
rect 21815 765 21860 885
rect 21980 765 22035 885
rect 22155 765 22200 885
rect 22320 765 22365 885
rect 22485 765 22530 885
rect 22650 765 22705 885
rect 22825 765 22870 885
rect 22990 765 23035 885
rect 23155 765 23200 885
rect 23320 765 23375 885
rect 23495 765 23540 885
rect 23660 765 23705 885
rect 23825 765 23870 885
rect 23990 765 24015 885
rect 18485 710 24015 765
rect 18485 590 18510 710
rect 18630 590 18685 710
rect 18805 590 18850 710
rect 18970 590 19015 710
rect 19135 590 19180 710
rect 19300 590 19355 710
rect 19475 590 19520 710
rect 19640 590 19685 710
rect 19805 590 19850 710
rect 19970 590 20025 710
rect 20145 590 20190 710
rect 20310 590 20355 710
rect 20475 590 20520 710
rect 20640 590 20695 710
rect 20815 590 20860 710
rect 20980 590 21025 710
rect 21145 590 21190 710
rect 21310 590 21365 710
rect 21485 590 21530 710
rect 21650 590 21695 710
rect 21815 590 21860 710
rect 21980 590 22035 710
rect 22155 590 22200 710
rect 22320 590 22365 710
rect 22485 590 22530 710
rect 22650 590 22705 710
rect 22825 590 22870 710
rect 22990 590 23035 710
rect 23155 590 23200 710
rect 23320 590 23375 710
rect 23495 590 23540 710
rect 23660 590 23705 710
rect 23825 590 23870 710
rect 23990 590 24015 710
rect 18485 545 24015 590
rect 18485 425 18510 545
rect 18630 425 18685 545
rect 18805 425 18850 545
rect 18970 425 19015 545
rect 19135 425 19180 545
rect 19300 425 19355 545
rect 19475 425 19520 545
rect 19640 425 19685 545
rect 19805 425 19850 545
rect 19970 425 20025 545
rect 20145 425 20190 545
rect 20310 425 20355 545
rect 20475 425 20520 545
rect 20640 425 20695 545
rect 20815 425 20860 545
rect 20980 425 21025 545
rect 21145 425 21190 545
rect 21310 425 21365 545
rect 21485 425 21530 545
rect 21650 425 21695 545
rect 21815 425 21860 545
rect 21980 425 22035 545
rect 22155 425 22200 545
rect 22320 425 22365 545
rect 22485 425 22530 545
rect 22650 425 22705 545
rect 22825 425 22870 545
rect 22990 425 23035 545
rect 23155 425 23200 545
rect 23320 425 23375 545
rect 23495 425 23540 545
rect 23660 425 23705 545
rect 23825 425 23870 545
rect 23990 425 24015 545
rect 18485 380 24015 425
rect 18485 260 18510 380
rect 18630 260 18685 380
rect 18805 260 18850 380
rect 18970 260 19015 380
rect 19135 260 19180 380
rect 19300 260 19355 380
rect 19475 260 19520 380
rect 19640 260 19685 380
rect 19805 260 19850 380
rect 19970 260 20025 380
rect 20145 260 20190 380
rect 20310 260 20355 380
rect 20475 260 20520 380
rect 20640 260 20695 380
rect 20815 260 20860 380
rect 20980 260 21025 380
rect 21145 260 21190 380
rect 21310 260 21365 380
rect 21485 260 21530 380
rect 21650 260 21695 380
rect 21815 260 21860 380
rect 21980 260 22035 380
rect 22155 260 22200 380
rect 22320 260 22365 380
rect 22485 260 22530 380
rect 22650 260 22705 380
rect 22825 260 22870 380
rect 22990 260 23035 380
rect 23155 260 23200 380
rect 23320 260 23375 380
rect 23495 260 23540 380
rect 23660 260 23705 380
rect 23825 260 23870 380
rect 23990 260 24015 380
rect 18485 215 24015 260
rect 18485 95 18510 215
rect 18630 95 18685 215
rect 18805 95 18850 215
rect 18970 95 19015 215
rect 19135 95 19180 215
rect 19300 95 19355 215
rect 19475 95 19520 215
rect 19640 95 19685 215
rect 19805 95 19850 215
rect 19970 95 20025 215
rect 20145 95 20190 215
rect 20310 95 20355 215
rect 20475 95 20520 215
rect 20640 95 20695 215
rect 20815 95 20860 215
rect 20980 95 21025 215
rect 21145 95 21190 215
rect 21310 95 21365 215
rect 21485 95 21530 215
rect 21650 95 21695 215
rect 21815 95 21860 215
rect 21980 95 22035 215
rect 22155 95 22200 215
rect 22320 95 22365 215
rect 22485 95 22530 215
rect 22650 95 22705 215
rect 22825 95 22870 215
rect 22990 95 23035 215
rect 23155 95 23200 215
rect 23320 95 23375 215
rect 23495 95 23540 215
rect 23660 95 23705 215
rect 23825 95 23870 215
rect 23990 95 24015 215
rect 18485 40 24015 95
rect 18485 -80 18510 40
rect 18630 -80 18685 40
rect 18805 -80 18850 40
rect 18970 -80 19015 40
rect 19135 -80 19180 40
rect 19300 -80 19355 40
rect 19475 -80 19520 40
rect 19640 -80 19685 40
rect 19805 -80 19850 40
rect 19970 -80 20025 40
rect 20145 -80 20190 40
rect 20310 -80 20355 40
rect 20475 -80 20520 40
rect 20640 -80 20695 40
rect 20815 -80 20860 40
rect 20980 -80 21025 40
rect 21145 -80 21190 40
rect 21310 -80 21365 40
rect 21485 -80 21530 40
rect 21650 -80 21695 40
rect 21815 -80 21860 40
rect 21980 -80 22035 40
rect 22155 -80 22200 40
rect 22320 -80 22365 40
rect 22485 -80 22530 40
rect 22650 -80 22705 40
rect 22825 -80 22870 40
rect 22990 -80 23035 40
rect 23155 -80 23200 40
rect 23320 -80 23375 40
rect 23495 -80 23540 40
rect 23660 -80 23705 40
rect 23825 -80 23870 40
rect 23990 -80 24015 40
rect 18485 -125 24015 -80
rect 18485 -245 18510 -125
rect 18630 -245 18685 -125
rect 18805 -245 18850 -125
rect 18970 -245 19015 -125
rect 19135 -245 19180 -125
rect 19300 -245 19355 -125
rect 19475 -245 19520 -125
rect 19640 -245 19685 -125
rect 19805 -245 19850 -125
rect 19970 -245 20025 -125
rect 20145 -245 20190 -125
rect 20310 -245 20355 -125
rect 20475 -245 20520 -125
rect 20640 -245 20695 -125
rect 20815 -245 20860 -125
rect 20980 -245 21025 -125
rect 21145 -245 21190 -125
rect 21310 -245 21365 -125
rect 21485 -245 21530 -125
rect 21650 -245 21695 -125
rect 21815 -245 21860 -125
rect 21980 -245 22035 -125
rect 22155 -245 22200 -125
rect 22320 -245 22365 -125
rect 22485 -245 22530 -125
rect 22650 -245 22705 -125
rect 22825 -245 22870 -125
rect 22990 -245 23035 -125
rect 23155 -245 23200 -125
rect 23320 -245 23375 -125
rect 23495 -245 23540 -125
rect 23660 -245 23705 -125
rect 23825 -245 23870 -125
rect 23990 -245 24015 -125
rect 18485 -290 24015 -245
rect 18485 -410 18510 -290
rect 18630 -410 18685 -290
rect 18805 -410 18850 -290
rect 18970 -410 19015 -290
rect 19135 -410 19180 -290
rect 19300 -410 19355 -290
rect 19475 -410 19520 -290
rect 19640 -410 19685 -290
rect 19805 -410 19850 -290
rect 19970 -410 20025 -290
rect 20145 -410 20190 -290
rect 20310 -410 20355 -290
rect 20475 -410 20520 -290
rect 20640 -410 20695 -290
rect 20815 -410 20860 -290
rect 20980 -410 21025 -290
rect 21145 -410 21190 -290
rect 21310 -410 21365 -290
rect 21485 -410 21530 -290
rect 21650 -410 21695 -290
rect 21815 -410 21860 -290
rect 21980 -410 22035 -290
rect 22155 -410 22200 -290
rect 22320 -410 22365 -290
rect 22485 -410 22530 -290
rect 22650 -410 22705 -290
rect 22825 -410 22870 -290
rect 22990 -410 23035 -290
rect 23155 -410 23200 -290
rect 23320 -410 23375 -290
rect 23495 -410 23540 -290
rect 23660 -410 23705 -290
rect 23825 -410 23870 -290
rect 23990 -410 24015 -290
rect 18485 -455 24015 -410
rect 18485 -575 18510 -455
rect 18630 -575 18685 -455
rect 18805 -575 18850 -455
rect 18970 -575 19015 -455
rect 19135 -575 19180 -455
rect 19300 -575 19355 -455
rect 19475 -575 19520 -455
rect 19640 -575 19685 -455
rect 19805 -575 19850 -455
rect 19970 -575 20025 -455
rect 20145 -575 20190 -455
rect 20310 -575 20355 -455
rect 20475 -575 20520 -455
rect 20640 -575 20695 -455
rect 20815 -575 20860 -455
rect 20980 -575 21025 -455
rect 21145 -575 21190 -455
rect 21310 -575 21365 -455
rect 21485 -575 21530 -455
rect 21650 -575 21695 -455
rect 21815 -575 21860 -455
rect 21980 -575 22035 -455
rect 22155 -575 22200 -455
rect 22320 -575 22365 -455
rect 22485 -575 22530 -455
rect 22650 -575 22705 -455
rect 22825 -575 22870 -455
rect 22990 -575 23035 -455
rect 23155 -575 23200 -455
rect 23320 -575 23375 -455
rect 23495 -575 23540 -455
rect 23660 -575 23705 -455
rect 23825 -575 23870 -455
rect 23990 -575 24015 -455
rect 18485 -630 24015 -575
rect 18485 -750 18510 -630
rect 18630 -750 18685 -630
rect 18805 -750 18850 -630
rect 18970 -750 19015 -630
rect 19135 -750 19180 -630
rect 19300 -750 19355 -630
rect 19475 -750 19520 -630
rect 19640 -750 19685 -630
rect 19805 -750 19850 -630
rect 19970 -750 20025 -630
rect 20145 -750 20190 -630
rect 20310 -750 20355 -630
rect 20475 -750 20520 -630
rect 20640 -750 20695 -630
rect 20815 -750 20860 -630
rect 20980 -750 21025 -630
rect 21145 -750 21190 -630
rect 21310 -750 21365 -630
rect 21485 -750 21530 -630
rect 21650 -750 21695 -630
rect 21815 -750 21860 -630
rect 21980 -750 22035 -630
rect 22155 -750 22200 -630
rect 22320 -750 22365 -630
rect 22485 -750 22530 -630
rect 22650 -750 22705 -630
rect 22825 -750 22870 -630
rect 22990 -750 23035 -630
rect 23155 -750 23200 -630
rect 23320 -750 23375 -630
rect 23495 -750 23540 -630
rect 23660 -750 23705 -630
rect 23825 -750 23870 -630
rect 23990 -750 24015 -630
rect 18485 -795 24015 -750
rect 18485 -915 18510 -795
rect 18630 -915 18685 -795
rect 18805 -915 18850 -795
rect 18970 -915 19015 -795
rect 19135 -915 19180 -795
rect 19300 -915 19355 -795
rect 19475 -915 19520 -795
rect 19640 -915 19685 -795
rect 19805 -915 19850 -795
rect 19970 -915 20025 -795
rect 20145 -915 20190 -795
rect 20310 -915 20355 -795
rect 20475 -915 20520 -795
rect 20640 -915 20695 -795
rect 20815 -915 20860 -795
rect 20980 -915 21025 -795
rect 21145 -915 21190 -795
rect 21310 -915 21365 -795
rect 21485 -915 21530 -795
rect 21650 -915 21695 -795
rect 21815 -915 21860 -795
rect 21980 -915 22035 -795
rect 22155 -915 22200 -795
rect 22320 -915 22365 -795
rect 22485 -915 22530 -795
rect 22650 -915 22705 -795
rect 22825 -915 22870 -795
rect 22990 -915 23035 -795
rect 23155 -915 23200 -795
rect 23320 -915 23375 -795
rect 23495 -915 23540 -795
rect 23660 -915 23705 -795
rect 23825 -915 23870 -795
rect 23990 -915 24015 -795
rect 18485 -960 24015 -915
rect 18485 -1080 18510 -960
rect 18630 -1080 18685 -960
rect 18805 -1080 18850 -960
rect 18970 -1080 19015 -960
rect 19135 -1080 19180 -960
rect 19300 -1080 19355 -960
rect 19475 -1080 19520 -960
rect 19640 -1080 19685 -960
rect 19805 -1080 19850 -960
rect 19970 -1080 20025 -960
rect 20145 -1080 20190 -960
rect 20310 -1080 20355 -960
rect 20475 -1080 20520 -960
rect 20640 -1080 20695 -960
rect 20815 -1080 20860 -960
rect 20980 -1080 21025 -960
rect 21145 -1080 21190 -960
rect 21310 -1080 21365 -960
rect 21485 -1080 21530 -960
rect 21650 -1080 21695 -960
rect 21815 -1080 21860 -960
rect 21980 -1080 22035 -960
rect 22155 -1080 22200 -960
rect 22320 -1080 22365 -960
rect 22485 -1080 22530 -960
rect 22650 -1080 22705 -960
rect 22825 -1080 22870 -960
rect 22990 -1080 23035 -960
rect 23155 -1080 23200 -960
rect 23320 -1080 23375 -960
rect 23495 -1080 23540 -960
rect 23660 -1080 23705 -960
rect 23825 -1080 23870 -960
rect 23990 -1080 24015 -960
rect 18485 -1125 24015 -1080
rect 18485 -1245 18510 -1125
rect 18630 -1245 18685 -1125
rect 18805 -1245 18850 -1125
rect 18970 -1245 19015 -1125
rect 19135 -1245 19180 -1125
rect 19300 -1245 19355 -1125
rect 19475 -1245 19520 -1125
rect 19640 -1245 19685 -1125
rect 19805 -1245 19850 -1125
rect 19970 -1245 20025 -1125
rect 20145 -1245 20190 -1125
rect 20310 -1245 20355 -1125
rect 20475 -1245 20520 -1125
rect 20640 -1245 20695 -1125
rect 20815 -1245 20860 -1125
rect 20980 -1245 21025 -1125
rect 21145 -1245 21190 -1125
rect 21310 -1245 21365 -1125
rect 21485 -1245 21530 -1125
rect 21650 -1245 21695 -1125
rect 21815 -1245 21860 -1125
rect 21980 -1245 22035 -1125
rect 22155 -1245 22200 -1125
rect 22320 -1245 22365 -1125
rect 22485 -1245 22530 -1125
rect 22650 -1245 22705 -1125
rect 22825 -1245 22870 -1125
rect 22990 -1245 23035 -1125
rect 23155 -1245 23200 -1125
rect 23320 -1245 23375 -1125
rect 23495 -1245 23540 -1125
rect 23660 -1245 23705 -1125
rect 23825 -1245 23870 -1125
rect 23990 -1245 24015 -1125
rect 18485 -1300 24015 -1245
rect 18485 -1420 18510 -1300
rect 18630 -1420 18685 -1300
rect 18805 -1420 18850 -1300
rect 18970 -1420 19015 -1300
rect 19135 -1420 19180 -1300
rect 19300 -1420 19355 -1300
rect 19475 -1420 19520 -1300
rect 19640 -1420 19685 -1300
rect 19805 -1420 19850 -1300
rect 19970 -1420 20025 -1300
rect 20145 -1420 20190 -1300
rect 20310 -1420 20355 -1300
rect 20475 -1420 20520 -1300
rect 20640 -1420 20695 -1300
rect 20815 -1420 20860 -1300
rect 20980 -1420 21025 -1300
rect 21145 -1420 21190 -1300
rect 21310 -1420 21365 -1300
rect 21485 -1420 21530 -1300
rect 21650 -1420 21695 -1300
rect 21815 -1420 21860 -1300
rect 21980 -1420 22035 -1300
rect 22155 -1420 22200 -1300
rect 22320 -1420 22365 -1300
rect 22485 -1420 22530 -1300
rect 22650 -1420 22705 -1300
rect 22825 -1420 22870 -1300
rect 22990 -1420 23035 -1300
rect 23155 -1420 23200 -1300
rect 23320 -1420 23375 -1300
rect 23495 -1420 23540 -1300
rect 23660 -1420 23705 -1300
rect 23825 -1420 23870 -1300
rect 23990 -1420 24015 -1300
rect 18485 -1465 24015 -1420
rect 18485 -1585 18510 -1465
rect 18630 -1585 18685 -1465
rect 18805 -1585 18850 -1465
rect 18970 -1585 19015 -1465
rect 19135 -1585 19180 -1465
rect 19300 -1585 19355 -1465
rect 19475 -1585 19520 -1465
rect 19640 -1585 19685 -1465
rect 19805 -1585 19850 -1465
rect 19970 -1585 20025 -1465
rect 20145 -1585 20190 -1465
rect 20310 -1585 20355 -1465
rect 20475 -1585 20520 -1465
rect 20640 -1585 20695 -1465
rect 20815 -1585 20860 -1465
rect 20980 -1585 21025 -1465
rect 21145 -1585 21190 -1465
rect 21310 -1585 21365 -1465
rect 21485 -1585 21530 -1465
rect 21650 -1585 21695 -1465
rect 21815 -1585 21860 -1465
rect 21980 -1585 22035 -1465
rect 22155 -1585 22200 -1465
rect 22320 -1585 22365 -1465
rect 22485 -1585 22530 -1465
rect 22650 -1585 22705 -1465
rect 22825 -1585 22870 -1465
rect 22990 -1585 23035 -1465
rect 23155 -1585 23200 -1465
rect 23320 -1585 23375 -1465
rect 23495 -1585 23540 -1465
rect 23660 -1585 23705 -1465
rect 23825 -1585 23870 -1465
rect 23990 -1585 24015 -1465
rect 18485 -1630 24015 -1585
rect 18485 -1750 18510 -1630
rect 18630 -1750 18685 -1630
rect 18805 -1750 18850 -1630
rect 18970 -1750 19015 -1630
rect 19135 -1750 19180 -1630
rect 19300 -1750 19355 -1630
rect 19475 -1750 19520 -1630
rect 19640 -1750 19685 -1630
rect 19805 -1750 19850 -1630
rect 19970 -1750 20025 -1630
rect 20145 -1750 20190 -1630
rect 20310 -1750 20355 -1630
rect 20475 -1750 20520 -1630
rect 20640 -1750 20695 -1630
rect 20815 -1750 20860 -1630
rect 20980 -1750 21025 -1630
rect 21145 -1750 21190 -1630
rect 21310 -1750 21365 -1630
rect 21485 -1750 21530 -1630
rect 21650 -1750 21695 -1630
rect 21815 -1750 21860 -1630
rect 21980 -1750 22035 -1630
rect 22155 -1750 22200 -1630
rect 22320 -1750 22365 -1630
rect 22485 -1750 22530 -1630
rect 22650 -1750 22705 -1630
rect 22825 -1750 22870 -1630
rect 22990 -1750 23035 -1630
rect 23155 -1750 23200 -1630
rect 23320 -1750 23375 -1630
rect 23495 -1750 23540 -1630
rect 23660 -1750 23705 -1630
rect 23825 -1750 23870 -1630
rect 23990 -1750 24015 -1630
rect 18485 -1795 24015 -1750
rect 18485 -1915 18510 -1795
rect 18630 -1915 18685 -1795
rect 18805 -1915 18850 -1795
rect 18970 -1915 19015 -1795
rect 19135 -1915 19180 -1795
rect 19300 -1915 19355 -1795
rect 19475 -1915 19520 -1795
rect 19640 -1915 19685 -1795
rect 19805 -1915 19850 -1795
rect 19970 -1915 20025 -1795
rect 20145 -1915 20190 -1795
rect 20310 -1915 20355 -1795
rect 20475 -1915 20520 -1795
rect 20640 -1915 20695 -1795
rect 20815 -1915 20860 -1795
rect 20980 -1915 21025 -1795
rect 21145 -1915 21190 -1795
rect 21310 -1915 21365 -1795
rect 21485 -1915 21530 -1795
rect 21650 -1915 21695 -1795
rect 21815 -1915 21860 -1795
rect 21980 -1915 22035 -1795
rect 22155 -1915 22200 -1795
rect 22320 -1915 22365 -1795
rect 22485 -1915 22530 -1795
rect 22650 -1915 22705 -1795
rect 22825 -1915 22870 -1795
rect 22990 -1915 23035 -1795
rect 23155 -1915 23200 -1795
rect 23320 -1915 23375 -1795
rect 23495 -1915 23540 -1795
rect 23660 -1915 23705 -1795
rect 23825 -1915 23870 -1795
rect 23990 -1915 24015 -1795
rect 18485 -1970 24015 -1915
rect 18485 -2090 18510 -1970
rect 18630 -2090 18685 -1970
rect 18805 -2090 18850 -1970
rect 18970 -2090 19015 -1970
rect 19135 -2090 19180 -1970
rect 19300 -2090 19355 -1970
rect 19475 -2090 19520 -1970
rect 19640 -2090 19685 -1970
rect 19805 -2090 19850 -1970
rect 19970 -2090 20025 -1970
rect 20145 -2090 20190 -1970
rect 20310 -2090 20355 -1970
rect 20475 -2090 20520 -1970
rect 20640 -2090 20695 -1970
rect 20815 -2090 20860 -1970
rect 20980 -2090 21025 -1970
rect 21145 -2090 21190 -1970
rect 21310 -2090 21365 -1970
rect 21485 -2090 21530 -1970
rect 21650 -2090 21695 -1970
rect 21815 -2090 21860 -1970
rect 21980 -2090 22035 -1970
rect 22155 -2090 22200 -1970
rect 22320 -2090 22365 -1970
rect 22485 -2090 22530 -1970
rect 22650 -2090 22705 -1970
rect 22825 -2090 22870 -1970
rect 22990 -2090 23035 -1970
rect 23155 -2090 23200 -1970
rect 23320 -2090 23375 -1970
rect 23495 -2090 23540 -1970
rect 23660 -2090 23705 -1970
rect 23825 -2090 23870 -1970
rect 23990 -2090 24015 -1970
rect 18485 -2135 24015 -2090
rect 18485 -2255 18510 -2135
rect 18630 -2255 18685 -2135
rect 18805 -2255 18850 -2135
rect 18970 -2255 19015 -2135
rect 19135 -2255 19180 -2135
rect 19300 -2255 19355 -2135
rect 19475 -2255 19520 -2135
rect 19640 -2255 19685 -2135
rect 19805 -2255 19850 -2135
rect 19970 -2255 20025 -2135
rect 20145 -2255 20190 -2135
rect 20310 -2255 20355 -2135
rect 20475 -2255 20520 -2135
rect 20640 -2255 20695 -2135
rect 20815 -2255 20860 -2135
rect 20980 -2255 21025 -2135
rect 21145 -2255 21190 -2135
rect 21310 -2255 21365 -2135
rect 21485 -2255 21530 -2135
rect 21650 -2255 21695 -2135
rect 21815 -2255 21860 -2135
rect 21980 -2255 22035 -2135
rect 22155 -2255 22200 -2135
rect 22320 -2255 22365 -2135
rect 22485 -2255 22530 -2135
rect 22650 -2255 22705 -2135
rect 22825 -2255 22870 -2135
rect 22990 -2255 23035 -2135
rect 23155 -2255 23200 -2135
rect 23320 -2255 23375 -2135
rect 23495 -2255 23540 -2135
rect 23660 -2255 23705 -2135
rect 23825 -2255 23870 -2135
rect 23990 -2255 24015 -2135
rect 18485 -2300 24015 -2255
rect 18485 -2420 18510 -2300
rect 18630 -2420 18685 -2300
rect 18805 -2420 18850 -2300
rect 18970 -2420 19015 -2300
rect 19135 -2420 19180 -2300
rect 19300 -2420 19355 -2300
rect 19475 -2420 19520 -2300
rect 19640 -2420 19685 -2300
rect 19805 -2420 19850 -2300
rect 19970 -2420 20025 -2300
rect 20145 -2420 20190 -2300
rect 20310 -2420 20355 -2300
rect 20475 -2420 20520 -2300
rect 20640 -2420 20695 -2300
rect 20815 -2420 20860 -2300
rect 20980 -2420 21025 -2300
rect 21145 -2420 21190 -2300
rect 21310 -2420 21365 -2300
rect 21485 -2420 21530 -2300
rect 21650 -2420 21695 -2300
rect 21815 -2420 21860 -2300
rect 21980 -2420 22035 -2300
rect 22155 -2420 22200 -2300
rect 22320 -2420 22365 -2300
rect 22485 -2420 22530 -2300
rect 22650 -2420 22705 -2300
rect 22825 -2420 22870 -2300
rect 22990 -2420 23035 -2300
rect 23155 -2420 23200 -2300
rect 23320 -2420 23375 -2300
rect 23495 -2420 23540 -2300
rect 23660 -2420 23705 -2300
rect 23825 -2420 23870 -2300
rect 23990 -2420 24015 -2300
rect 18485 -2465 24015 -2420
rect 18485 -2585 18510 -2465
rect 18630 -2585 18685 -2465
rect 18805 -2585 18850 -2465
rect 18970 -2585 19015 -2465
rect 19135 -2585 19180 -2465
rect 19300 -2585 19355 -2465
rect 19475 -2585 19520 -2465
rect 19640 -2585 19685 -2465
rect 19805 -2585 19850 -2465
rect 19970 -2585 20025 -2465
rect 20145 -2585 20190 -2465
rect 20310 -2585 20355 -2465
rect 20475 -2585 20520 -2465
rect 20640 -2585 20695 -2465
rect 20815 -2585 20860 -2465
rect 20980 -2585 21025 -2465
rect 21145 -2585 21190 -2465
rect 21310 -2585 21365 -2465
rect 21485 -2585 21530 -2465
rect 21650 -2585 21695 -2465
rect 21815 -2585 21860 -2465
rect 21980 -2585 22035 -2465
rect 22155 -2585 22200 -2465
rect 22320 -2585 22365 -2465
rect 22485 -2585 22530 -2465
rect 22650 -2585 22705 -2465
rect 22825 -2585 22870 -2465
rect 22990 -2585 23035 -2465
rect 23155 -2585 23200 -2465
rect 23320 -2585 23375 -2465
rect 23495 -2585 23540 -2465
rect 23660 -2585 23705 -2465
rect 23825 -2585 23870 -2465
rect 23990 -2585 24015 -2465
rect 18485 -2640 24015 -2585
rect 18485 -2760 18510 -2640
rect 18630 -2760 18685 -2640
rect 18805 -2760 18850 -2640
rect 18970 -2760 19015 -2640
rect 19135 -2760 19180 -2640
rect 19300 -2760 19355 -2640
rect 19475 -2760 19520 -2640
rect 19640 -2760 19685 -2640
rect 19805 -2760 19850 -2640
rect 19970 -2760 20025 -2640
rect 20145 -2760 20190 -2640
rect 20310 -2760 20355 -2640
rect 20475 -2760 20520 -2640
rect 20640 -2760 20695 -2640
rect 20815 -2760 20860 -2640
rect 20980 -2760 21025 -2640
rect 21145 -2760 21190 -2640
rect 21310 -2760 21365 -2640
rect 21485 -2760 21530 -2640
rect 21650 -2760 21695 -2640
rect 21815 -2760 21860 -2640
rect 21980 -2760 22035 -2640
rect 22155 -2760 22200 -2640
rect 22320 -2760 22365 -2640
rect 22485 -2760 22530 -2640
rect 22650 -2760 22705 -2640
rect 22825 -2760 22870 -2640
rect 22990 -2760 23035 -2640
rect 23155 -2760 23200 -2640
rect 23320 -2760 23375 -2640
rect 23495 -2760 23540 -2640
rect 23660 -2760 23705 -2640
rect 23825 -2760 23870 -2640
rect 23990 -2760 24015 -2640
rect 18485 -2805 24015 -2760
rect 18485 -2925 18510 -2805
rect 18630 -2925 18685 -2805
rect 18805 -2925 18850 -2805
rect 18970 -2925 19015 -2805
rect 19135 -2925 19180 -2805
rect 19300 -2925 19355 -2805
rect 19475 -2925 19520 -2805
rect 19640 -2925 19685 -2805
rect 19805 -2925 19850 -2805
rect 19970 -2925 20025 -2805
rect 20145 -2925 20190 -2805
rect 20310 -2925 20355 -2805
rect 20475 -2925 20520 -2805
rect 20640 -2925 20695 -2805
rect 20815 -2925 20860 -2805
rect 20980 -2925 21025 -2805
rect 21145 -2925 21190 -2805
rect 21310 -2925 21365 -2805
rect 21485 -2925 21530 -2805
rect 21650 -2925 21695 -2805
rect 21815 -2925 21860 -2805
rect 21980 -2925 22035 -2805
rect 22155 -2925 22200 -2805
rect 22320 -2925 22365 -2805
rect 22485 -2925 22530 -2805
rect 22650 -2925 22705 -2805
rect 22825 -2925 22870 -2805
rect 22990 -2925 23035 -2805
rect 23155 -2925 23200 -2805
rect 23320 -2925 23375 -2805
rect 23495 -2925 23540 -2805
rect 23660 -2925 23705 -2805
rect 23825 -2925 23870 -2805
rect 23990 -2925 24015 -2805
rect 18485 -2970 24015 -2925
rect 18485 -3090 18510 -2970
rect 18630 -3090 18685 -2970
rect 18805 -3090 18850 -2970
rect 18970 -3090 19015 -2970
rect 19135 -3090 19180 -2970
rect 19300 -3090 19355 -2970
rect 19475 -3090 19520 -2970
rect 19640 -3090 19685 -2970
rect 19805 -3090 19850 -2970
rect 19970 -3090 20025 -2970
rect 20145 -3090 20190 -2970
rect 20310 -3090 20355 -2970
rect 20475 -3090 20520 -2970
rect 20640 -3090 20695 -2970
rect 20815 -3090 20860 -2970
rect 20980 -3090 21025 -2970
rect 21145 -3090 21190 -2970
rect 21310 -3090 21365 -2970
rect 21485 -3090 21530 -2970
rect 21650 -3090 21695 -2970
rect 21815 -3090 21860 -2970
rect 21980 -3090 22035 -2970
rect 22155 -3090 22200 -2970
rect 22320 -3090 22365 -2970
rect 22485 -3090 22530 -2970
rect 22650 -3090 22705 -2970
rect 22825 -3090 22870 -2970
rect 22990 -3090 23035 -2970
rect 23155 -3090 23200 -2970
rect 23320 -3090 23375 -2970
rect 23495 -3090 23540 -2970
rect 23660 -3090 23705 -2970
rect 23825 -3090 23870 -2970
rect 23990 -3090 24015 -2970
rect 18485 -3135 24015 -3090
rect 18485 -3255 18510 -3135
rect 18630 -3255 18685 -3135
rect 18805 -3255 18850 -3135
rect 18970 -3255 19015 -3135
rect 19135 -3255 19180 -3135
rect 19300 -3255 19355 -3135
rect 19475 -3255 19520 -3135
rect 19640 -3255 19685 -3135
rect 19805 -3255 19850 -3135
rect 19970 -3255 20025 -3135
rect 20145 -3255 20190 -3135
rect 20310 -3255 20355 -3135
rect 20475 -3255 20520 -3135
rect 20640 -3255 20695 -3135
rect 20815 -3255 20860 -3135
rect 20980 -3255 21025 -3135
rect 21145 -3255 21190 -3135
rect 21310 -3255 21365 -3135
rect 21485 -3255 21530 -3135
rect 21650 -3255 21695 -3135
rect 21815 -3255 21860 -3135
rect 21980 -3255 22035 -3135
rect 22155 -3255 22200 -3135
rect 22320 -3255 22365 -3135
rect 22485 -3255 22530 -3135
rect 22650 -3255 22705 -3135
rect 22825 -3255 22870 -3135
rect 22990 -3255 23035 -3135
rect 23155 -3255 23200 -3135
rect 23320 -3255 23375 -3135
rect 23495 -3255 23540 -3135
rect 23660 -3255 23705 -3135
rect 23825 -3255 23870 -3135
rect 23990 -3255 24015 -3135
rect 18485 -3310 24015 -3255
rect 18485 -3430 18510 -3310
rect 18630 -3430 18685 -3310
rect 18805 -3430 18850 -3310
rect 18970 -3430 19015 -3310
rect 19135 -3430 19180 -3310
rect 19300 -3430 19355 -3310
rect 19475 -3430 19520 -3310
rect 19640 -3430 19685 -3310
rect 19805 -3430 19850 -3310
rect 19970 -3430 20025 -3310
rect 20145 -3430 20190 -3310
rect 20310 -3430 20355 -3310
rect 20475 -3430 20520 -3310
rect 20640 -3430 20695 -3310
rect 20815 -3430 20860 -3310
rect 20980 -3430 21025 -3310
rect 21145 -3430 21190 -3310
rect 21310 -3430 21365 -3310
rect 21485 -3430 21530 -3310
rect 21650 -3430 21695 -3310
rect 21815 -3430 21860 -3310
rect 21980 -3430 22035 -3310
rect 22155 -3430 22200 -3310
rect 22320 -3430 22365 -3310
rect 22485 -3430 22530 -3310
rect 22650 -3430 22705 -3310
rect 22825 -3430 22870 -3310
rect 22990 -3430 23035 -3310
rect 23155 -3430 23200 -3310
rect 23320 -3430 23375 -3310
rect 23495 -3430 23540 -3310
rect 23660 -3430 23705 -3310
rect 23825 -3430 23870 -3310
rect 23990 -3430 24015 -3310
rect 18485 -3475 24015 -3430
rect 18485 -3595 18510 -3475
rect 18630 -3595 18685 -3475
rect 18805 -3595 18850 -3475
rect 18970 -3595 19015 -3475
rect 19135 -3595 19180 -3475
rect 19300 -3595 19355 -3475
rect 19475 -3595 19520 -3475
rect 19640 -3595 19685 -3475
rect 19805 -3595 19850 -3475
rect 19970 -3595 20025 -3475
rect 20145 -3595 20190 -3475
rect 20310 -3595 20355 -3475
rect 20475 -3595 20520 -3475
rect 20640 -3595 20695 -3475
rect 20815 -3595 20860 -3475
rect 20980 -3595 21025 -3475
rect 21145 -3595 21190 -3475
rect 21310 -3595 21365 -3475
rect 21485 -3595 21530 -3475
rect 21650 -3595 21695 -3475
rect 21815 -3595 21860 -3475
rect 21980 -3595 22035 -3475
rect 22155 -3595 22200 -3475
rect 22320 -3595 22365 -3475
rect 22485 -3595 22530 -3475
rect 22650 -3595 22705 -3475
rect 22825 -3595 22870 -3475
rect 22990 -3595 23035 -3475
rect 23155 -3595 23200 -3475
rect 23320 -3595 23375 -3475
rect 23495 -3595 23540 -3475
rect 23660 -3595 23705 -3475
rect 23825 -3595 23870 -3475
rect 23990 -3595 24015 -3475
rect 18485 -3640 24015 -3595
rect 18485 -3760 18510 -3640
rect 18630 -3760 18685 -3640
rect 18805 -3760 18850 -3640
rect 18970 -3760 19015 -3640
rect 19135 -3760 19180 -3640
rect 19300 -3760 19355 -3640
rect 19475 -3760 19520 -3640
rect 19640 -3760 19685 -3640
rect 19805 -3760 19850 -3640
rect 19970 -3760 20025 -3640
rect 20145 -3760 20190 -3640
rect 20310 -3760 20355 -3640
rect 20475 -3760 20520 -3640
rect 20640 -3760 20695 -3640
rect 20815 -3760 20860 -3640
rect 20980 -3760 21025 -3640
rect 21145 -3760 21190 -3640
rect 21310 -3760 21365 -3640
rect 21485 -3760 21530 -3640
rect 21650 -3760 21695 -3640
rect 21815 -3760 21860 -3640
rect 21980 -3760 22035 -3640
rect 22155 -3760 22200 -3640
rect 22320 -3760 22365 -3640
rect 22485 -3760 22530 -3640
rect 22650 -3760 22705 -3640
rect 22825 -3760 22870 -3640
rect 22990 -3760 23035 -3640
rect 23155 -3760 23200 -3640
rect 23320 -3760 23375 -3640
rect 23495 -3760 23540 -3640
rect 23660 -3760 23705 -3640
rect 23825 -3760 23870 -3640
rect 23990 -3760 24015 -3640
rect 18485 -3805 24015 -3760
rect 18485 -3925 18510 -3805
rect 18630 -3925 18685 -3805
rect 18805 -3925 18850 -3805
rect 18970 -3925 19015 -3805
rect 19135 -3925 19180 -3805
rect 19300 -3925 19355 -3805
rect 19475 -3925 19520 -3805
rect 19640 -3925 19685 -3805
rect 19805 -3925 19850 -3805
rect 19970 -3925 20025 -3805
rect 20145 -3925 20190 -3805
rect 20310 -3925 20355 -3805
rect 20475 -3925 20520 -3805
rect 20640 -3925 20695 -3805
rect 20815 -3925 20860 -3805
rect 20980 -3925 21025 -3805
rect 21145 -3925 21190 -3805
rect 21310 -3925 21365 -3805
rect 21485 -3925 21530 -3805
rect 21650 -3925 21695 -3805
rect 21815 -3925 21860 -3805
rect 21980 -3925 22035 -3805
rect 22155 -3925 22200 -3805
rect 22320 -3925 22365 -3805
rect 22485 -3925 22530 -3805
rect 22650 -3925 22705 -3805
rect 22825 -3925 22870 -3805
rect 22990 -3925 23035 -3805
rect 23155 -3925 23200 -3805
rect 23320 -3925 23375 -3805
rect 23495 -3925 23540 -3805
rect 23660 -3925 23705 -3805
rect 23825 -3925 23870 -3805
rect 23990 -3925 24015 -3805
rect 18485 -3980 24015 -3925
rect 18485 -4065 18510 -3980
rect 18300 -4100 18510 -4065
rect 18630 -4100 18685 -3980
rect 18805 -4100 18850 -3980
rect 18970 -4100 19015 -3980
rect 19135 -4100 19180 -3980
rect 19300 -4100 19355 -3980
rect 19475 -4100 19520 -3980
rect 19640 -4100 19685 -3980
rect 19805 -4100 19850 -3980
rect 19970 -4100 20025 -3980
rect 20145 -4100 20190 -3980
rect 20310 -4100 20355 -3980
rect 20475 -4100 20520 -3980
rect 20640 -4100 20695 -3980
rect 20815 -4100 20860 -3980
rect 20980 -4100 21025 -3980
rect 21145 -4100 21190 -3980
rect 21310 -4100 21365 -3980
rect 21485 -4100 21530 -3980
rect 21650 -4100 21695 -3980
rect 21815 -4100 21860 -3980
rect 21980 -4100 22035 -3980
rect 22155 -4100 22200 -3980
rect 22320 -4100 22365 -3980
rect 22485 -4100 22530 -3980
rect 22650 -4100 22705 -3980
rect 22825 -4100 22870 -3980
rect 22990 -4100 23035 -3980
rect 23155 -4100 23200 -3980
rect 23320 -4100 23375 -3980
rect 23495 -4100 23540 -3980
rect 23660 -4100 23705 -3980
rect 23825 -4100 23870 -3980
rect 23990 -4065 24015 -3980
rect 24175 1380 29705 1405
rect 24175 1260 24200 1380
rect 24320 1260 24375 1380
rect 24495 1260 24540 1380
rect 24660 1260 24705 1380
rect 24825 1260 24870 1380
rect 24990 1260 25045 1380
rect 25165 1260 25210 1380
rect 25330 1260 25375 1380
rect 25495 1260 25540 1380
rect 25660 1260 25715 1380
rect 25835 1260 25880 1380
rect 26000 1260 26045 1380
rect 26165 1260 26210 1380
rect 26330 1260 26385 1380
rect 26505 1260 26550 1380
rect 26670 1260 26715 1380
rect 26835 1260 26880 1380
rect 27000 1260 27055 1380
rect 27175 1260 27220 1380
rect 27340 1260 27385 1380
rect 27505 1260 27550 1380
rect 27670 1260 27725 1380
rect 27845 1260 27890 1380
rect 28010 1260 28055 1380
rect 28175 1260 28220 1380
rect 28340 1260 28395 1380
rect 28515 1260 28560 1380
rect 28680 1260 28725 1380
rect 28845 1260 28890 1380
rect 29010 1260 29065 1380
rect 29185 1260 29230 1380
rect 29350 1260 29395 1380
rect 29515 1260 29560 1380
rect 29680 1260 29705 1380
rect 24175 1215 29705 1260
rect 24175 1095 24200 1215
rect 24320 1095 24375 1215
rect 24495 1095 24540 1215
rect 24660 1095 24705 1215
rect 24825 1095 24870 1215
rect 24990 1095 25045 1215
rect 25165 1095 25210 1215
rect 25330 1095 25375 1215
rect 25495 1095 25540 1215
rect 25660 1095 25715 1215
rect 25835 1095 25880 1215
rect 26000 1095 26045 1215
rect 26165 1095 26210 1215
rect 26330 1095 26385 1215
rect 26505 1095 26550 1215
rect 26670 1095 26715 1215
rect 26835 1095 26880 1215
rect 27000 1095 27055 1215
rect 27175 1095 27220 1215
rect 27340 1095 27385 1215
rect 27505 1095 27550 1215
rect 27670 1095 27725 1215
rect 27845 1095 27890 1215
rect 28010 1095 28055 1215
rect 28175 1095 28220 1215
rect 28340 1095 28395 1215
rect 28515 1095 28560 1215
rect 28680 1095 28725 1215
rect 28845 1095 28890 1215
rect 29010 1095 29065 1215
rect 29185 1095 29230 1215
rect 29350 1095 29395 1215
rect 29515 1095 29560 1215
rect 29680 1095 29705 1215
rect 24175 1050 29705 1095
rect 24175 930 24200 1050
rect 24320 930 24375 1050
rect 24495 930 24540 1050
rect 24660 930 24705 1050
rect 24825 930 24870 1050
rect 24990 930 25045 1050
rect 25165 930 25210 1050
rect 25330 930 25375 1050
rect 25495 930 25540 1050
rect 25660 930 25715 1050
rect 25835 930 25880 1050
rect 26000 930 26045 1050
rect 26165 930 26210 1050
rect 26330 930 26385 1050
rect 26505 930 26550 1050
rect 26670 930 26715 1050
rect 26835 930 26880 1050
rect 27000 930 27055 1050
rect 27175 930 27220 1050
rect 27340 930 27385 1050
rect 27505 930 27550 1050
rect 27670 930 27725 1050
rect 27845 930 27890 1050
rect 28010 930 28055 1050
rect 28175 930 28220 1050
rect 28340 930 28395 1050
rect 28515 930 28560 1050
rect 28680 930 28725 1050
rect 28845 930 28890 1050
rect 29010 930 29065 1050
rect 29185 930 29230 1050
rect 29350 930 29395 1050
rect 29515 930 29560 1050
rect 29680 930 29705 1050
rect 24175 885 29705 930
rect 24175 765 24200 885
rect 24320 765 24375 885
rect 24495 765 24540 885
rect 24660 765 24705 885
rect 24825 765 24870 885
rect 24990 765 25045 885
rect 25165 765 25210 885
rect 25330 765 25375 885
rect 25495 765 25540 885
rect 25660 765 25715 885
rect 25835 765 25880 885
rect 26000 765 26045 885
rect 26165 765 26210 885
rect 26330 765 26385 885
rect 26505 765 26550 885
rect 26670 765 26715 885
rect 26835 765 26880 885
rect 27000 765 27055 885
rect 27175 765 27220 885
rect 27340 765 27385 885
rect 27505 765 27550 885
rect 27670 765 27725 885
rect 27845 765 27890 885
rect 28010 765 28055 885
rect 28175 765 28220 885
rect 28340 765 28395 885
rect 28515 765 28560 885
rect 28680 765 28725 885
rect 28845 765 28890 885
rect 29010 765 29065 885
rect 29185 765 29230 885
rect 29350 765 29395 885
rect 29515 765 29560 885
rect 29680 765 29705 885
rect 24175 710 29705 765
rect 24175 590 24200 710
rect 24320 590 24375 710
rect 24495 590 24540 710
rect 24660 590 24705 710
rect 24825 590 24870 710
rect 24990 590 25045 710
rect 25165 590 25210 710
rect 25330 590 25375 710
rect 25495 590 25540 710
rect 25660 590 25715 710
rect 25835 590 25880 710
rect 26000 590 26045 710
rect 26165 590 26210 710
rect 26330 590 26385 710
rect 26505 590 26550 710
rect 26670 590 26715 710
rect 26835 590 26880 710
rect 27000 590 27055 710
rect 27175 590 27220 710
rect 27340 590 27385 710
rect 27505 590 27550 710
rect 27670 590 27725 710
rect 27845 590 27890 710
rect 28010 590 28055 710
rect 28175 590 28220 710
rect 28340 590 28395 710
rect 28515 590 28560 710
rect 28680 590 28725 710
rect 28845 590 28890 710
rect 29010 590 29065 710
rect 29185 590 29230 710
rect 29350 590 29395 710
rect 29515 590 29560 710
rect 29680 590 29705 710
rect 24175 545 29705 590
rect 24175 425 24200 545
rect 24320 425 24375 545
rect 24495 425 24540 545
rect 24660 425 24705 545
rect 24825 425 24870 545
rect 24990 425 25045 545
rect 25165 425 25210 545
rect 25330 425 25375 545
rect 25495 425 25540 545
rect 25660 425 25715 545
rect 25835 425 25880 545
rect 26000 425 26045 545
rect 26165 425 26210 545
rect 26330 425 26385 545
rect 26505 425 26550 545
rect 26670 425 26715 545
rect 26835 425 26880 545
rect 27000 425 27055 545
rect 27175 425 27220 545
rect 27340 425 27385 545
rect 27505 425 27550 545
rect 27670 425 27725 545
rect 27845 425 27890 545
rect 28010 425 28055 545
rect 28175 425 28220 545
rect 28340 425 28395 545
rect 28515 425 28560 545
rect 28680 425 28725 545
rect 28845 425 28890 545
rect 29010 425 29065 545
rect 29185 425 29230 545
rect 29350 425 29395 545
rect 29515 425 29560 545
rect 29680 425 29705 545
rect 24175 380 29705 425
rect 24175 260 24200 380
rect 24320 260 24375 380
rect 24495 260 24540 380
rect 24660 260 24705 380
rect 24825 260 24870 380
rect 24990 260 25045 380
rect 25165 260 25210 380
rect 25330 260 25375 380
rect 25495 260 25540 380
rect 25660 260 25715 380
rect 25835 260 25880 380
rect 26000 260 26045 380
rect 26165 260 26210 380
rect 26330 260 26385 380
rect 26505 260 26550 380
rect 26670 260 26715 380
rect 26835 260 26880 380
rect 27000 260 27055 380
rect 27175 260 27220 380
rect 27340 260 27385 380
rect 27505 260 27550 380
rect 27670 260 27725 380
rect 27845 260 27890 380
rect 28010 260 28055 380
rect 28175 260 28220 380
rect 28340 260 28395 380
rect 28515 260 28560 380
rect 28680 260 28725 380
rect 28845 260 28890 380
rect 29010 260 29065 380
rect 29185 260 29230 380
rect 29350 260 29395 380
rect 29515 260 29560 380
rect 29680 260 29705 380
rect 24175 215 29705 260
rect 24175 95 24200 215
rect 24320 95 24375 215
rect 24495 95 24540 215
rect 24660 95 24705 215
rect 24825 95 24870 215
rect 24990 95 25045 215
rect 25165 95 25210 215
rect 25330 95 25375 215
rect 25495 95 25540 215
rect 25660 95 25715 215
rect 25835 95 25880 215
rect 26000 95 26045 215
rect 26165 95 26210 215
rect 26330 95 26385 215
rect 26505 95 26550 215
rect 26670 95 26715 215
rect 26835 95 26880 215
rect 27000 95 27055 215
rect 27175 95 27220 215
rect 27340 95 27385 215
rect 27505 95 27550 215
rect 27670 95 27725 215
rect 27845 95 27890 215
rect 28010 95 28055 215
rect 28175 95 28220 215
rect 28340 95 28395 215
rect 28515 95 28560 215
rect 28680 95 28725 215
rect 28845 95 28890 215
rect 29010 95 29065 215
rect 29185 95 29230 215
rect 29350 95 29395 215
rect 29515 95 29560 215
rect 29680 95 29705 215
rect 24175 40 29705 95
rect 24175 -80 24200 40
rect 24320 -80 24375 40
rect 24495 -80 24540 40
rect 24660 -80 24705 40
rect 24825 -80 24870 40
rect 24990 -80 25045 40
rect 25165 -80 25210 40
rect 25330 -80 25375 40
rect 25495 -80 25540 40
rect 25660 -80 25715 40
rect 25835 -80 25880 40
rect 26000 -80 26045 40
rect 26165 -80 26210 40
rect 26330 -80 26385 40
rect 26505 -80 26550 40
rect 26670 -80 26715 40
rect 26835 -80 26880 40
rect 27000 -80 27055 40
rect 27175 -80 27220 40
rect 27340 -80 27385 40
rect 27505 -80 27550 40
rect 27670 -80 27725 40
rect 27845 -80 27890 40
rect 28010 -80 28055 40
rect 28175 -80 28220 40
rect 28340 -80 28395 40
rect 28515 -80 28560 40
rect 28680 -80 28725 40
rect 28845 -80 28890 40
rect 29010 -80 29065 40
rect 29185 -80 29230 40
rect 29350 -80 29395 40
rect 29515 -80 29560 40
rect 29680 -80 29705 40
rect 24175 -125 29705 -80
rect 24175 -245 24200 -125
rect 24320 -245 24375 -125
rect 24495 -245 24540 -125
rect 24660 -245 24705 -125
rect 24825 -245 24870 -125
rect 24990 -245 25045 -125
rect 25165 -245 25210 -125
rect 25330 -245 25375 -125
rect 25495 -245 25540 -125
rect 25660 -245 25715 -125
rect 25835 -245 25880 -125
rect 26000 -245 26045 -125
rect 26165 -245 26210 -125
rect 26330 -245 26385 -125
rect 26505 -245 26550 -125
rect 26670 -245 26715 -125
rect 26835 -245 26880 -125
rect 27000 -245 27055 -125
rect 27175 -245 27220 -125
rect 27340 -245 27385 -125
rect 27505 -245 27550 -125
rect 27670 -245 27725 -125
rect 27845 -245 27890 -125
rect 28010 -245 28055 -125
rect 28175 -245 28220 -125
rect 28340 -245 28395 -125
rect 28515 -245 28560 -125
rect 28680 -245 28725 -125
rect 28845 -245 28890 -125
rect 29010 -245 29065 -125
rect 29185 -245 29230 -125
rect 29350 -245 29395 -125
rect 29515 -245 29560 -125
rect 29680 -245 29705 -125
rect 24175 -290 29705 -245
rect 24175 -410 24200 -290
rect 24320 -410 24375 -290
rect 24495 -410 24540 -290
rect 24660 -410 24705 -290
rect 24825 -410 24870 -290
rect 24990 -410 25045 -290
rect 25165 -410 25210 -290
rect 25330 -410 25375 -290
rect 25495 -410 25540 -290
rect 25660 -410 25715 -290
rect 25835 -410 25880 -290
rect 26000 -410 26045 -290
rect 26165 -410 26210 -290
rect 26330 -410 26385 -290
rect 26505 -410 26550 -290
rect 26670 -410 26715 -290
rect 26835 -410 26880 -290
rect 27000 -410 27055 -290
rect 27175 -410 27220 -290
rect 27340 -410 27385 -290
rect 27505 -410 27550 -290
rect 27670 -410 27725 -290
rect 27845 -410 27890 -290
rect 28010 -410 28055 -290
rect 28175 -410 28220 -290
rect 28340 -410 28395 -290
rect 28515 -410 28560 -290
rect 28680 -410 28725 -290
rect 28845 -410 28890 -290
rect 29010 -410 29065 -290
rect 29185 -410 29230 -290
rect 29350 -410 29395 -290
rect 29515 -410 29560 -290
rect 29680 -410 29705 -290
rect 24175 -455 29705 -410
rect 24175 -575 24200 -455
rect 24320 -575 24375 -455
rect 24495 -575 24540 -455
rect 24660 -575 24705 -455
rect 24825 -575 24870 -455
rect 24990 -575 25045 -455
rect 25165 -575 25210 -455
rect 25330 -575 25375 -455
rect 25495 -575 25540 -455
rect 25660 -575 25715 -455
rect 25835 -575 25880 -455
rect 26000 -575 26045 -455
rect 26165 -575 26210 -455
rect 26330 -575 26385 -455
rect 26505 -575 26550 -455
rect 26670 -575 26715 -455
rect 26835 -575 26880 -455
rect 27000 -575 27055 -455
rect 27175 -575 27220 -455
rect 27340 -575 27385 -455
rect 27505 -575 27550 -455
rect 27670 -575 27725 -455
rect 27845 -575 27890 -455
rect 28010 -575 28055 -455
rect 28175 -575 28220 -455
rect 28340 -575 28395 -455
rect 28515 -575 28560 -455
rect 28680 -575 28725 -455
rect 28845 -575 28890 -455
rect 29010 -575 29065 -455
rect 29185 -575 29230 -455
rect 29350 -575 29395 -455
rect 29515 -575 29560 -455
rect 29680 -575 29705 -455
rect 24175 -630 29705 -575
rect 24175 -750 24200 -630
rect 24320 -750 24375 -630
rect 24495 -750 24540 -630
rect 24660 -750 24705 -630
rect 24825 -750 24870 -630
rect 24990 -750 25045 -630
rect 25165 -750 25210 -630
rect 25330 -750 25375 -630
rect 25495 -750 25540 -630
rect 25660 -750 25715 -630
rect 25835 -750 25880 -630
rect 26000 -750 26045 -630
rect 26165 -750 26210 -630
rect 26330 -750 26385 -630
rect 26505 -750 26550 -630
rect 26670 -750 26715 -630
rect 26835 -750 26880 -630
rect 27000 -750 27055 -630
rect 27175 -750 27220 -630
rect 27340 -750 27385 -630
rect 27505 -750 27550 -630
rect 27670 -750 27725 -630
rect 27845 -750 27890 -630
rect 28010 -750 28055 -630
rect 28175 -750 28220 -630
rect 28340 -750 28395 -630
rect 28515 -750 28560 -630
rect 28680 -750 28725 -630
rect 28845 -750 28890 -630
rect 29010 -750 29065 -630
rect 29185 -750 29230 -630
rect 29350 -750 29395 -630
rect 29515 -750 29560 -630
rect 29680 -750 29705 -630
rect 24175 -795 29705 -750
rect 24175 -915 24200 -795
rect 24320 -915 24375 -795
rect 24495 -915 24540 -795
rect 24660 -915 24705 -795
rect 24825 -915 24870 -795
rect 24990 -915 25045 -795
rect 25165 -915 25210 -795
rect 25330 -915 25375 -795
rect 25495 -915 25540 -795
rect 25660 -915 25715 -795
rect 25835 -915 25880 -795
rect 26000 -915 26045 -795
rect 26165 -915 26210 -795
rect 26330 -915 26385 -795
rect 26505 -915 26550 -795
rect 26670 -915 26715 -795
rect 26835 -915 26880 -795
rect 27000 -915 27055 -795
rect 27175 -915 27220 -795
rect 27340 -915 27385 -795
rect 27505 -915 27550 -795
rect 27670 -915 27725 -795
rect 27845 -915 27890 -795
rect 28010 -915 28055 -795
rect 28175 -915 28220 -795
rect 28340 -915 28395 -795
rect 28515 -915 28560 -795
rect 28680 -915 28725 -795
rect 28845 -915 28890 -795
rect 29010 -915 29065 -795
rect 29185 -915 29230 -795
rect 29350 -915 29395 -795
rect 29515 -915 29560 -795
rect 29680 -915 29705 -795
rect 24175 -960 29705 -915
rect 24175 -1080 24200 -960
rect 24320 -1080 24375 -960
rect 24495 -1080 24540 -960
rect 24660 -1080 24705 -960
rect 24825 -1080 24870 -960
rect 24990 -1080 25045 -960
rect 25165 -1080 25210 -960
rect 25330 -1080 25375 -960
rect 25495 -1080 25540 -960
rect 25660 -1080 25715 -960
rect 25835 -1080 25880 -960
rect 26000 -1080 26045 -960
rect 26165 -1080 26210 -960
rect 26330 -1080 26385 -960
rect 26505 -1080 26550 -960
rect 26670 -1080 26715 -960
rect 26835 -1080 26880 -960
rect 27000 -1080 27055 -960
rect 27175 -1080 27220 -960
rect 27340 -1080 27385 -960
rect 27505 -1080 27550 -960
rect 27670 -1080 27725 -960
rect 27845 -1080 27890 -960
rect 28010 -1080 28055 -960
rect 28175 -1080 28220 -960
rect 28340 -1080 28395 -960
rect 28515 -1080 28560 -960
rect 28680 -1080 28725 -960
rect 28845 -1080 28890 -960
rect 29010 -1080 29065 -960
rect 29185 -1080 29230 -960
rect 29350 -1080 29395 -960
rect 29515 -1080 29560 -960
rect 29680 -1080 29705 -960
rect 24175 -1125 29705 -1080
rect 24175 -1245 24200 -1125
rect 24320 -1245 24375 -1125
rect 24495 -1245 24540 -1125
rect 24660 -1245 24705 -1125
rect 24825 -1245 24870 -1125
rect 24990 -1245 25045 -1125
rect 25165 -1245 25210 -1125
rect 25330 -1245 25375 -1125
rect 25495 -1245 25540 -1125
rect 25660 -1245 25715 -1125
rect 25835 -1245 25880 -1125
rect 26000 -1245 26045 -1125
rect 26165 -1245 26210 -1125
rect 26330 -1245 26385 -1125
rect 26505 -1245 26550 -1125
rect 26670 -1245 26715 -1125
rect 26835 -1245 26880 -1125
rect 27000 -1245 27055 -1125
rect 27175 -1245 27220 -1125
rect 27340 -1245 27385 -1125
rect 27505 -1245 27550 -1125
rect 27670 -1245 27725 -1125
rect 27845 -1245 27890 -1125
rect 28010 -1245 28055 -1125
rect 28175 -1245 28220 -1125
rect 28340 -1245 28395 -1125
rect 28515 -1245 28560 -1125
rect 28680 -1245 28725 -1125
rect 28845 -1245 28890 -1125
rect 29010 -1245 29065 -1125
rect 29185 -1245 29230 -1125
rect 29350 -1245 29395 -1125
rect 29515 -1245 29560 -1125
rect 29680 -1245 29705 -1125
rect 24175 -1300 29705 -1245
rect 24175 -1420 24200 -1300
rect 24320 -1420 24375 -1300
rect 24495 -1420 24540 -1300
rect 24660 -1420 24705 -1300
rect 24825 -1420 24870 -1300
rect 24990 -1420 25045 -1300
rect 25165 -1420 25210 -1300
rect 25330 -1420 25375 -1300
rect 25495 -1420 25540 -1300
rect 25660 -1420 25715 -1300
rect 25835 -1420 25880 -1300
rect 26000 -1420 26045 -1300
rect 26165 -1420 26210 -1300
rect 26330 -1420 26385 -1300
rect 26505 -1420 26550 -1300
rect 26670 -1420 26715 -1300
rect 26835 -1420 26880 -1300
rect 27000 -1420 27055 -1300
rect 27175 -1420 27220 -1300
rect 27340 -1420 27385 -1300
rect 27505 -1420 27550 -1300
rect 27670 -1420 27725 -1300
rect 27845 -1420 27890 -1300
rect 28010 -1420 28055 -1300
rect 28175 -1420 28220 -1300
rect 28340 -1420 28395 -1300
rect 28515 -1420 28560 -1300
rect 28680 -1420 28725 -1300
rect 28845 -1420 28890 -1300
rect 29010 -1420 29065 -1300
rect 29185 -1420 29230 -1300
rect 29350 -1420 29395 -1300
rect 29515 -1420 29560 -1300
rect 29680 -1420 29705 -1300
rect 24175 -1465 29705 -1420
rect 24175 -1585 24200 -1465
rect 24320 -1585 24375 -1465
rect 24495 -1585 24540 -1465
rect 24660 -1585 24705 -1465
rect 24825 -1585 24870 -1465
rect 24990 -1585 25045 -1465
rect 25165 -1585 25210 -1465
rect 25330 -1585 25375 -1465
rect 25495 -1585 25540 -1465
rect 25660 -1585 25715 -1465
rect 25835 -1585 25880 -1465
rect 26000 -1585 26045 -1465
rect 26165 -1585 26210 -1465
rect 26330 -1585 26385 -1465
rect 26505 -1585 26550 -1465
rect 26670 -1585 26715 -1465
rect 26835 -1585 26880 -1465
rect 27000 -1585 27055 -1465
rect 27175 -1585 27220 -1465
rect 27340 -1585 27385 -1465
rect 27505 -1585 27550 -1465
rect 27670 -1585 27725 -1465
rect 27845 -1585 27890 -1465
rect 28010 -1585 28055 -1465
rect 28175 -1585 28220 -1465
rect 28340 -1585 28395 -1465
rect 28515 -1585 28560 -1465
rect 28680 -1585 28725 -1465
rect 28845 -1585 28890 -1465
rect 29010 -1585 29065 -1465
rect 29185 -1585 29230 -1465
rect 29350 -1585 29395 -1465
rect 29515 -1585 29560 -1465
rect 29680 -1585 29705 -1465
rect 24175 -1630 29705 -1585
rect 24175 -1750 24200 -1630
rect 24320 -1750 24375 -1630
rect 24495 -1750 24540 -1630
rect 24660 -1750 24705 -1630
rect 24825 -1750 24870 -1630
rect 24990 -1750 25045 -1630
rect 25165 -1750 25210 -1630
rect 25330 -1750 25375 -1630
rect 25495 -1750 25540 -1630
rect 25660 -1750 25715 -1630
rect 25835 -1750 25880 -1630
rect 26000 -1750 26045 -1630
rect 26165 -1750 26210 -1630
rect 26330 -1750 26385 -1630
rect 26505 -1750 26550 -1630
rect 26670 -1750 26715 -1630
rect 26835 -1750 26880 -1630
rect 27000 -1750 27055 -1630
rect 27175 -1750 27220 -1630
rect 27340 -1750 27385 -1630
rect 27505 -1750 27550 -1630
rect 27670 -1750 27725 -1630
rect 27845 -1750 27890 -1630
rect 28010 -1750 28055 -1630
rect 28175 -1750 28220 -1630
rect 28340 -1750 28395 -1630
rect 28515 -1750 28560 -1630
rect 28680 -1750 28725 -1630
rect 28845 -1750 28890 -1630
rect 29010 -1750 29065 -1630
rect 29185 -1750 29230 -1630
rect 29350 -1750 29395 -1630
rect 29515 -1750 29560 -1630
rect 29680 -1750 29705 -1630
rect 24175 -1795 29705 -1750
rect 24175 -1915 24200 -1795
rect 24320 -1915 24375 -1795
rect 24495 -1915 24540 -1795
rect 24660 -1915 24705 -1795
rect 24825 -1915 24870 -1795
rect 24990 -1915 25045 -1795
rect 25165 -1915 25210 -1795
rect 25330 -1915 25375 -1795
rect 25495 -1915 25540 -1795
rect 25660 -1915 25715 -1795
rect 25835 -1915 25880 -1795
rect 26000 -1915 26045 -1795
rect 26165 -1915 26210 -1795
rect 26330 -1915 26385 -1795
rect 26505 -1915 26550 -1795
rect 26670 -1915 26715 -1795
rect 26835 -1915 26880 -1795
rect 27000 -1915 27055 -1795
rect 27175 -1915 27220 -1795
rect 27340 -1915 27385 -1795
rect 27505 -1915 27550 -1795
rect 27670 -1915 27725 -1795
rect 27845 -1915 27890 -1795
rect 28010 -1915 28055 -1795
rect 28175 -1915 28220 -1795
rect 28340 -1915 28395 -1795
rect 28515 -1915 28560 -1795
rect 28680 -1915 28725 -1795
rect 28845 -1915 28890 -1795
rect 29010 -1915 29065 -1795
rect 29185 -1915 29230 -1795
rect 29350 -1915 29395 -1795
rect 29515 -1915 29560 -1795
rect 29680 -1915 29705 -1795
rect 24175 -1970 29705 -1915
rect 24175 -2090 24200 -1970
rect 24320 -2090 24375 -1970
rect 24495 -2090 24540 -1970
rect 24660 -2090 24705 -1970
rect 24825 -2090 24870 -1970
rect 24990 -2090 25045 -1970
rect 25165 -2090 25210 -1970
rect 25330 -2090 25375 -1970
rect 25495 -2090 25540 -1970
rect 25660 -2090 25715 -1970
rect 25835 -2090 25880 -1970
rect 26000 -2090 26045 -1970
rect 26165 -2090 26210 -1970
rect 26330 -2090 26385 -1970
rect 26505 -2090 26550 -1970
rect 26670 -2090 26715 -1970
rect 26835 -2090 26880 -1970
rect 27000 -2090 27055 -1970
rect 27175 -2090 27220 -1970
rect 27340 -2090 27385 -1970
rect 27505 -2090 27550 -1970
rect 27670 -2090 27725 -1970
rect 27845 -2090 27890 -1970
rect 28010 -2090 28055 -1970
rect 28175 -2090 28220 -1970
rect 28340 -2090 28395 -1970
rect 28515 -2090 28560 -1970
rect 28680 -2090 28725 -1970
rect 28845 -2090 28890 -1970
rect 29010 -2090 29065 -1970
rect 29185 -2090 29230 -1970
rect 29350 -2090 29395 -1970
rect 29515 -2090 29560 -1970
rect 29680 -2090 29705 -1970
rect 24175 -2135 29705 -2090
rect 24175 -2255 24200 -2135
rect 24320 -2255 24375 -2135
rect 24495 -2255 24540 -2135
rect 24660 -2255 24705 -2135
rect 24825 -2255 24870 -2135
rect 24990 -2255 25045 -2135
rect 25165 -2255 25210 -2135
rect 25330 -2255 25375 -2135
rect 25495 -2255 25540 -2135
rect 25660 -2255 25715 -2135
rect 25835 -2255 25880 -2135
rect 26000 -2255 26045 -2135
rect 26165 -2255 26210 -2135
rect 26330 -2255 26385 -2135
rect 26505 -2255 26550 -2135
rect 26670 -2255 26715 -2135
rect 26835 -2255 26880 -2135
rect 27000 -2255 27055 -2135
rect 27175 -2255 27220 -2135
rect 27340 -2255 27385 -2135
rect 27505 -2255 27550 -2135
rect 27670 -2255 27725 -2135
rect 27845 -2255 27890 -2135
rect 28010 -2255 28055 -2135
rect 28175 -2255 28220 -2135
rect 28340 -2255 28395 -2135
rect 28515 -2255 28560 -2135
rect 28680 -2255 28725 -2135
rect 28845 -2255 28890 -2135
rect 29010 -2255 29065 -2135
rect 29185 -2255 29230 -2135
rect 29350 -2255 29395 -2135
rect 29515 -2255 29560 -2135
rect 29680 -2255 29705 -2135
rect 24175 -2300 29705 -2255
rect 24175 -2420 24200 -2300
rect 24320 -2420 24375 -2300
rect 24495 -2420 24540 -2300
rect 24660 -2420 24705 -2300
rect 24825 -2420 24870 -2300
rect 24990 -2420 25045 -2300
rect 25165 -2420 25210 -2300
rect 25330 -2420 25375 -2300
rect 25495 -2420 25540 -2300
rect 25660 -2420 25715 -2300
rect 25835 -2420 25880 -2300
rect 26000 -2420 26045 -2300
rect 26165 -2420 26210 -2300
rect 26330 -2420 26385 -2300
rect 26505 -2420 26550 -2300
rect 26670 -2420 26715 -2300
rect 26835 -2420 26880 -2300
rect 27000 -2420 27055 -2300
rect 27175 -2420 27220 -2300
rect 27340 -2420 27385 -2300
rect 27505 -2420 27550 -2300
rect 27670 -2420 27725 -2300
rect 27845 -2420 27890 -2300
rect 28010 -2420 28055 -2300
rect 28175 -2420 28220 -2300
rect 28340 -2420 28395 -2300
rect 28515 -2420 28560 -2300
rect 28680 -2420 28725 -2300
rect 28845 -2420 28890 -2300
rect 29010 -2420 29065 -2300
rect 29185 -2420 29230 -2300
rect 29350 -2420 29395 -2300
rect 29515 -2420 29560 -2300
rect 29680 -2420 29705 -2300
rect 24175 -2465 29705 -2420
rect 24175 -2585 24200 -2465
rect 24320 -2585 24375 -2465
rect 24495 -2585 24540 -2465
rect 24660 -2585 24705 -2465
rect 24825 -2585 24870 -2465
rect 24990 -2585 25045 -2465
rect 25165 -2585 25210 -2465
rect 25330 -2585 25375 -2465
rect 25495 -2585 25540 -2465
rect 25660 -2585 25715 -2465
rect 25835 -2585 25880 -2465
rect 26000 -2585 26045 -2465
rect 26165 -2585 26210 -2465
rect 26330 -2585 26385 -2465
rect 26505 -2585 26550 -2465
rect 26670 -2585 26715 -2465
rect 26835 -2585 26880 -2465
rect 27000 -2585 27055 -2465
rect 27175 -2585 27220 -2465
rect 27340 -2585 27385 -2465
rect 27505 -2585 27550 -2465
rect 27670 -2585 27725 -2465
rect 27845 -2585 27890 -2465
rect 28010 -2585 28055 -2465
rect 28175 -2585 28220 -2465
rect 28340 -2585 28395 -2465
rect 28515 -2585 28560 -2465
rect 28680 -2585 28725 -2465
rect 28845 -2585 28890 -2465
rect 29010 -2585 29065 -2465
rect 29185 -2585 29230 -2465
rect 29350 -2585 29395 -2465
rect 29515 -2585 29560 -2465
rect 29680 -2585 29705 -2465
rect 24175 -2640 29705 -2585
rect 24175 -2760 24200 -2640
rect 24320 -2760 24375 -2640
rect 24495 -2760 24540 -2640
rect 24660 -2760 24705 -2640
rect 24825 -2760 24870 -2640
rect 24990 -2760 25045 -2640
rect 25165 -2760 25210 -2640
rect 25330 -2760 25375 -2640
rect 25495 -2760 25540 -2640
rect 25660 -2760 25715 -2640
rect 25835 -2760 25880 -2640
rect 26000 -2760 26045 -2640
rect 26165 -2760 26210 -2640
rect 26330 -2760 26385 -2640
rect 26505 -2760 26550 -2640
rect 26670 -2760 26715 -2640
rect 26835 -2760 26880 -2640
rect 27000 -2760 27055 -2640
rect 27175 -2760 27220 -2640
rect 27340 -2760 27385 -2640
rect 27505 -2760 27550 -2640
rect 27670 -2760 27725 -2640
rect 27845 -2760 27890 -2640
rect 28010 -2760 28055 -2640
rect 28175 -2760 28220 -2640
rect 28340 -2760 28395 -2640
rect 28515 -2760 28560 -2640
rect 28680 -2760 28725 -2640
rect 28845 -2760 28890 -2640
rect 29010 -2760 29065 -2640
rect 29185 -2760 29230 -2640
rect 29350 -2760 29395 -2640
rect 29515 -2760 29560 -2640
rect 29680 -2760 29705 -2640
rect 24175 -2805 29705 -2760
rect 24175 -2925 24200 -2805
rect 24320 -2925 24375 -2805
rect 24495 -2925 24540 -2805
rect 24660 -2925 24705 -2805
rect 24825 -2925 24870 -2805
rect 24990 -2925 25045 -2805
rect 25165 -2925 25210 -2805
rect 25330 -2925 25375 -2805
rect 25495 -2925 25540 -2805
rect 25660 -2925 25715 -2805
rect 25835 -2925 25880 -2805
rect 26000 -2925 26045 -2805
rect 26165 -2925 26210 -2805
rect 26330 -2925 26385 -2805
rect 26505 -2925 26550 -2805
rect 26670 -2925 26715 -2805
rect 26835 -2925 26880 -2805
rect 27000 -2925 27055 -2805
rect 27175 -2925 27220 -2805
rect 27340 -2925 27385 -2805
rect 27505 -2925 27550 -2805
rect 27670 -2925 27725 -2805
rect 27845 -2925 27890 -2805
rect 28010 -2925 28055 -2805
rect 28175 -2925 28220 -2805
rect 28340 -2925 28395 -2805
rect 28515 -2925 28560 -2805
rect 28680 -2925 28725 -2805
rect 28845 -2925 28890 -2805
rect 29010 -2925 29065 -2805
rect 29185 -2925 29230 -2805
rect 29350 -2925 29395 -2805
rect 29515 -2925 29560 -2805
rect 29680 -2925 29705 -2805
rect 24175 -2970 29705 -2925
rect 24175 -3090 24200 -2970
rect 24320 -3090 24375 -2970
rect 24495 -3090 24540 -2970
rect 24660 -3090 24705 -2970
rect 24825 -3090 24870 -2970
rect 24990 -3090 25045 -2970
rect 25165 -3090 25210 -2970
rect 25330 -3090 25375 -2970
rect 25495 -3090 25540 -2970
rect 25660 -3090 25715 -2970
rect 25835 -3090 25880 -2970
rect 26000 -3090 26045 -2970
rect 26165 -3090 26210 -2970
rect 26330 -3090 26385 -2970
rect 26505 -3090 26550 -2970
rect 26670 -3090 26715 -2970
rect 26835 -3090 26880 -2970
rect 27000 -3090 27055 -2970
rect 27175 -3090 27220 -2970
rect 27340 -3090 27385 -2970
rect 27505 -3090 27550 -2970
rect 27670 -3090 27725 -2970
rect 27845 -3090 27890 -2970
rect 28010 -3090 28055 -2970
rect 28175 -3090 28220 -2970
rect 28340 -3090 28395 -2970
rect 28515 -3090 28560 -2970
rect 28680 -3090 28725 -2970
rect 28845 -3090 28890 -2970
rect 29010 -3090 29065 -2970
rect 29185 -3090 29230 -2970
rect 29350 -3090 29395 -2970
rect 29515 -3090 29560 -2970
rect 29680 -3090 29705 -2970
rect 24175 -3135 29705 -3090
rect 24175 -3255 24200 -3135
rect 24320 -3255 24375 -3135
rect 24495 -3255 24540 -3135
rect 24660 -3255 24705 -3135
rect 24825 -3255 24870 -3135
rect 24990 -3255 25045 -3135
rect 25165 -3255 25210 -3135
rect 25330 -3255 25375 -3135
rect 25495 -3255 25540 -3135
rect 25660 -3255 25715 -3135
rect 25835 -3255 25880 -3135
rect 26000 -3255 26045 -3135
rect 26165 -3255 26210 -3135
rect 26330 -3255 26385 -3135
rect 26505 -3255 26550 -3135
rect 26670 -3255 26715 -3135
rect 26835 -3255 26880 -3135
rect 27000 -3255 27055 -3135
rect 27175 -3255 27220 -3135
rect 27340 -3255 27385 -3135
rect 27505 -3255 27550 -3135
rect 27670 -3255 27725 -3135
rect 27845 -3255 27890 -3135
rect 28010 -3255 28055 -3135
rect 28175 -3255 28220 -3135
rect 28340 -3255 28395 -3135
rect 28515 -3255 28560 -3135
rect 28680 -3255 28725 -3135
rect 28845 -3255 28890 -3135
rect 29010 -3255 29065 -3135
rect 29185 -3255 29230 -3135
rect 29350 -3255 29395 -3135
rect 29515 -3255 29560 -3135
rect 29680 -3255 29705 -3135
rect 24175 -3310 29705 -3255
rect 24175 -3430 24200 -3310
rect 24320 -3430 24375 -3310
rect 24495 -3430 24540 -3310
rect 24660 -3430 24705 -3310
rect 24825 -3430 24870 -3310
rect 24990 -3430 25045 -3310
rect 25165 -3430 25210 -3310
rect 25330 -3430 25375 -3310
rect 25495 -3430 25540 -3310
rect 25660 -3430 25715 -3310
rect 25835 -3430 25880 -3310
rect 26000 -3430 26045 -3310
rect 26165 -3430 26210 -3310
rect 26330 -3430 26385 -3310
rect 26505 -3430 26550 -3310
rect 26670 -3430 26715 -3310
rect 26835 -3430 26880 -3310
rect 27000 -3430 27055 -3310
rect 27175 -3430 27220 -3310
rect 27340 -3430 27385 -3310
rect 27505 -3430 27550 -3310
rect 27670 -3430 27725 -3310
rect 27845 -3430 27890 -3310
rect 28010 -3430 28055 -3310
rect 28175 -3430 28220 -3310
rect 28340 -3430 28395 -3310
rect 28515 -3430 28560 -3310
rect 28680 -3430 28725 -3310
rect 28845 -3430 28890 -3310
rect 29010 -3430 29065 -3310
rect 29185 -3430 29230 -3310
rect 29350 -3430 29395 -3310
rect 29515 -3430 29560 -3310
rect 29680 -3430 29705 -3310
rect 24175 -3475 29705 -3430
rect 24175 -3595 24200 -3475
rect 24320 -3595 24375 -3475
rect 24495 -3595 24540 -3475
rect 24660 -3595 24705 -3475
rect 24825 -3595 24870 -3475
rect 24990 -3595 25045 -3475
rect 25165 -3595 25210 -3475
rect 25330 -3595 25375 -3475
rect 25495 -3595 25540 -3475
rect 25660 -3595 25715 -3475
rect 25835 -3595 25880 -3475
rect 26000 -3595 26045 -3475
rect 26165 -3595 26210 -3475
rect 26330 -3595 26385 -3475
rect 26505 -3595 26550 -3475
rect 26670 -3595 26715 -3475
rect 26835 -3595 26880 -3475
rect 27000 -3595 27055 -3475
rect 27175 -3595 27220 -3475
rect 27340 -3595 27385 -3475
rect 27505 -3595 27550 -3475
rect 27670 -3595 27725 -3475
rect 27845 -3595 27890 -3475
rect 28010 -3595 28055 -3475
rect 28175 -3595 28220 -3475
rect 28340 -3595 28395 -3475
rect 28515 -3595 28560 -3475
rect 28680 -3595 28725 -3475
rect 28845 -3595 28890 -3475
rect 29010 -3595 29065 -3475
rect 29185 -3595 29230 -3475
rect 29350 -3595 29395 -3475
rect 29515 -3595 29560 -3475
rect 29680 -3595 29705 -3475
rect 24175 -3640 29705 -3595
rect 24175 -3760 24200 -3640
rect 24320 -3760 24375 -3640
rect 24495 -3760 24540 -3640
rect 24660 -3760 24705 -3640
rect 24825 -3760 24870 -3640
rect 24990 -3760 25045 -3640
rect 25165 -3760 25210 -3640
rect 25330 -3760 25375 -3640
rect 25495 -3760 25540 -3640
rect 25660 -3760 25715 -3640
rect 25835 -3760 25880 -3640
rect 26000 -3760 26045 -3640
rect 26165 -3760 26210 -3640
rect 26330 -3760 26385 -3640
rect 26505 -3760 26550 -3640
rect 26670 -3760 26715 -3640
rect 26835 -3760 26880 -3640
rect 27000 -3760 27055 -3640
rect 27175 -3760 27220 -3640
rect 27340 -3760 27385 -3640
rect 27505 -3760 27550 -3640
rect 27670 -3760 27725 -3640
rect 27845 -3760 27890 -3640
rect 28010 -3760 28055 -3640
rect 28175 -3760 28220 -3640
rect 28340 -3760 28395 -3640
rect 28515 -3760 28560 -3640
rect 28680 -3760 28725 -3640
rect 28845 -3760 28890 -3640
rect 29010 -3760 29065 -3640
rect 29185 -3760 29230 -3640
rect 29350 -3760 29395 -3640
rect 29515 -3760 29560 -3640
rect 29680 -3760 29705 -3640
rect 24175 -3805 29705 -3760
rect 24175 -3925 24200 -3805
rect 24320 -3925 24375 -3805
rect 24495 -3925 24540 -3805
rect 24660 -3925 24705 -3805
rect 24825 -3925 24870 -3805
rect 24990 -3925 25045 -3805
rect 25165 -3925 25210 -3805
rect 25330 -3925 25375 -3805
rect 25495 -3925 25540 -3805
rect 25660 -3925 25715 -3805
rect 25835 -3925 25880 -3805
rect 26000 -3925 26045 -3805
rect 26165 -3925 26210 -3805
rect 26330 -3925 26385 -3805
rect 26505 -3925 26550 -3805
rect 26670 -3925 26715 -3805
rect 26835 -3925 26880 -3805
rect 27000 -3925 27055 -3805
rect 27175 -3925 27220 -3805
rect 27340 -3925 27385 -3805
rect 27505 -3925 27550 -3805
rect 27670 -3925 27725 -3805
rect 27845 -3925 27890 -3805
rect 28010 -3925 28055 -3805
rect 28175 -3925 28220 -3805
rect 28340 -3925 28395 -3805
rect 28515 -3925 28560 -3805
rect 28680 -3925 28725 -3805
rect 28845 -3925 28890 -3805
rect 29010 -3925 29065 -3805
rect 29185 -3925 29230 -3805
rect 29350 -3925 29395 -3805
rect 29515 -3925 29560 -3805
rect 29680 -3925 29705 -3805
rect 24175 -3980 29705 -3925
rect 24175 -4065 24200 -3980
rect 23990 -4100 24200 -4065
rect 24320 -4100 24375 -3980
rect 24495 -4100 24540 -3980
rect 24660 -4100 24705 -3980
rect 24825 -4100 24870 -3980
rect 24990 -4100 25045 -3980
rect 25165 -4100 25210 -3980
rect 25330 -4100 25375 -3980
rect 25495 -4100 25540 -3980
rect 25660 -4100 25715 -3980
rect 25835 -4100 25880 -3980
rect 26000 -4100 26045 -3980
rect 26165 -4100 26210 -3980
rect 26330 -4100 26385 -3980
rect 26505 -4100 26550 -3980
rect 26670 -4100 26715 -3980
rect 26835 -4100 26880 -3980
rect 27000 -4100 27055 -3980
rect 27175 -4100 27220 -3980
rect 27340 -4100 27385 -3980
rect 27505 -4100 27550 -3980
rect 27670 -4100 27725 -3980
rect 27845 -4100 27890 -3980
rect 28010 -4100 28055 -3980
rect 28175 -4100 28220 -3980
rect 28340 -4100 28395 -3980
rect 28515 -4100 28560 -3980
rect 28680 -4100 28725 -3980
rect 28845 -4100 28890 -3980
rect 29010 -4100 29065 -3980
rect 29185 -4100 29230 -3980
rect 29350 -4100 29395 -3980
rect 29515 -4100 29560 -3980
rect 29680 -4100 29705 -3980
rect 7105 -4310 29705 -4100
rect 7105 -4430 7130 -4310
rect 7250 -4430 7295 -4310
rect 7415 -4430 7460 -4310
rect 7580 -4430 7625 -4310
rect 7745 -4430 7800 -4310
rect 7920 -4430 7965 -4310
rect 8085 -4430 8130 -4310
rect 8250 -4430 8295 -4310
rect 8415 -4430 8470 -4310
rect 8590 -4430 8635 -4310
rect 8755 -4430 8800 -4310
rect 8920 -4430 8965 -4310
rect 9085 -4430 9140 -4310
rect 9260 -4430 9305 -4310
rect 9425 -4430 9470 -4310
rect 9590 -4430 9635 -4310
rect 9755 -4430 9810 -4310
rect 9930 -4430 9975 -4310
rect 10095 -4430 10140 -4310
rect 10260 -4430 10305 -4310
rect 10425 -4430 10480 -4310
rect 10600 -4430 10645 -4310
rect 10765 -4430 10810 -4310
rect 10930 -4430 10975 -4310
rect 11095 -4430 11150 -4310
rect 11270 -4430 11315 -4310
rect 11435 -4430 11480 -4310
rect 11600 -4430 11645 -4310
rect 11765 -4430 11820 -4310
rect 11940 -4430 11985 -4310
rect 12105 -4430 12150 -4310
rect 12270 -4430 12315 -4310
rect 12435 -4430 12490 -4310
rect 12610 -4345 12820 -4310
rect 12610 -4430 12635 -4345
rect 7105 -4485 12635 -4430
rect 7105 -4605 7130 -4485
rect 7250 -4605 7295 -4485
rect 7415 -4605 7460 -4485
rect 7580 -4605 7625 -4485
rect 7745 -4605 7800 -4485
rect 7920 -4605 7965 -4485
rect 8085 -4605 8130 -4485
rect 8250 -4605 8295 -4485
rect 8415 -4605 8470 -4485
rect 8590 -4605 8635 -4485
rect 8755 -4605 8800 -4485
rect 8920 -4605 8965 -4485
rect 9085 -4605 9140 -4485
rect 9260 -4605 9305 -4485
rect 9425 -4605 9470 -4485
rect 9590 -4605 9635 -4485
rect 9755 -4605 9810 -4485
rect 9930 -4605 9975 -4485
rect 10095 -4605 10140 -4485
rect 10260 -4605 10305 -4485
rect 10425 -4605 10480 -4485
rect 10600 -4605 10645 -4485
rect 10765 -4605 10810 -4485
rect 10930 -4605 10975 -4485
rect 11095 -4605 11150 -4485
rect 11270 -4605 11315 -4485
rect 11435 -4605 11480 -4485
rect 11600 -4605 11645 -4485
rect 11765 -4605 11820 -4485
rect 11940 -4605 11985 -4485
rect 12105 -4605 12150 -4485
rect 12270 -4605 12315 -4485
rect 12435 -4605 12490 -4485
rect 12610 -4605 12635 -4485
rect 7105 -4650 12635 -4605
rect 7105 -4770 7130 -4650
rect 7250 -4770 7295 -4650
rect 7415 -4770 7460 -4650
rect 7580 -4770 7625 -4650
rect 7745 -4770 7800 -4650
rect 7920 -4770 7965 -4650
rect 8085 -4770 8130 -4650
rect 8250 -4770 8295 -4650
rect 8415 -4770 8470 -4650
rect 8590 -4770 8635 -4650
rect 8755 -4770 8800 -4650
rect 8920 -4770 8965 -4650
rect 9085 -4770 9140 -4650
rect 9260 -4770 9305 -4650
rect 9425 -4770 9470 -4650
rect 9590 -4770 9635 -4650
rect 9755 -4770 9810 -4650
rect 9930 -4770 9975 -4650
rect 10095 -4770 10140 -4650
rect 10260 -4770 10305 -4650
rect 10425 -4770 10480 -4650
rect 10600 -4770 10645 -4650
rect 10765 -4770 10810 -4650
rect 10930 -4770 10975 -4650
rect 11095 -4770 11150 -4650
rect 11270 -4770 11315 -4650
rect 11435 -4770 11480 -4650
rect 11600 -4770 11645 -4650
rect 11765 -4770 11820 -4650
rect 11940 -4770 11985 -4650
rect 12105 -4770 12150 -4650
rect 12270 -4770 12315 -4650
rect 12435 -4770 12490 -4650
rect 12610 -4770 12635 -4650
rect 7105 -4815 12635 -4770
rect 7105 -4935 7130 -4815
rect 7250 -4935 7295 -4815
rect 7415 -4935 7460 -4815
rect 7580 -4935 7625 -4815
rect 7745 -4935 7800 -4815
rect 7920 -4935 7965 -4815
rect 8085 -4935 8130 -4815
rect 8250 -4935 8295 -4815
rect 8415 -4935 8470 -4815
rect 8590 -4935 8635 -4815
rect 8755 -4935 8800 -4815
rect 8920 -4935 8965 -4815
rect 9085 -4935 9140 -4815
rect 9260 -4935 9305 -4815
rect 9425 -4935 9470 -4815
rect 9590 -4935 9635 -4815
rect 9755 -4935 9810 -4815
rect 9930 -4935 9975 -4815
rect 10095 -4935 10140 -4815
rect 10260 -4935 10305 -4815
rect 10425 -4935 10480 -4815
rect 10600 -4935 10645 -4815
rect 10765 -4935 10810 -4815
rect 10930 -4935 10975 -4815
rect 11095 -4935 11150 -4815
rect 11270 -4935 11315 -4815
rect 11435 -4935 11480 -4815
rect 11600 -4935 11645 -4815
rect 11765 -4935 11820 -4815
rect 11940 -4935 11985 -4815
rect 12105 -4935 12150 -4815
rect 12270 -4935 12315 -4815
rect 12435 -4935 12490 -4815
rect 12610 -4935 12635 -4815
rect 7105 -4980 12635 -4935
rect 7105 -5100 7130 -4980
rect 7250 -5100 7295 -4980
rect 7415 -5100 7460 -4980
rect 7580 -5100 7625 -4980
rect 7745 -5100 7800 -4980
rect 7920 -5100 7965 -4980
rect 8085 -5100 8130 -4980
rect 8250 -5100 8295 -4980
rect 8415 -5100 8470 -4980
rect 8590 -5100 8635 -4980
rect 8755 -5100 8800 -4980
rect 8920 -5100 8965 -4980
rect 9085 -5100 9140 -4980
rect 9260 -5100 9305 -4980
rect 9425 -5100 9470 -4980
rect 9590 -5100 9635 -4980
rect 9755 -5100 9810 -4980
rect 9930 -5100 9975 -4980
rect 10095 -5100 10140 -4980
rect 10260 -5100 10305 -4980
rect 10425 -5100 10480 -4980
rect 10600 -5100 10645 -4980
rect 10765 -5100 10810 -4980
rect 10930 -5100 10975 -4980
rect 11095 -5100 11150 -4980
rect 11270 -5100 11315 -4980
rect 11435 -5100 11480 -4980
rect 11600 -5100 11645 -4980
rect 11765 -5100 11820 -4980
rect 11940 -5100 11985 -4980
rect 12105 -5100 12150 -4980
rect 12270 -5100 12315 -4980
rect 12435 -5100 12490 -4980
rect 12610 -5100 12635 -4980
rect 7105 -5155 12635 -5100
rect 7105 -5275 7130 -5155
rect 7250 -5275 7295 -5155
rect 7415 -5275 7460 -5155
rect 7580 -5275 7625 -5155
rect 7745 -5275 7800 -5155
rect 7920 -5275 7965 -5155
rect 8085 -5275 8130 -5155
rect 8250 -5275 8295 -5155
rect 8415 -5275 8470 -5155
rect 8590 -5275 8635 -5155
rect 8755 -5275 8800 -5155
rect 8920 -5275 8965 -5155
rect 9085 -5275 9140 -5155
rect 9260 -5275 9305 -5155
rect 9425 -5275 9470 -5155
rect 9590 -5275 9635 -5155
rect 9755 -5275 9810 -5155
rect 9930 -5275 9975 -5155
rect 10095 -5275 10140 -5155
rect 10260 -5275 10305 -5155
rect 10425 -5275 10480 -5155
rect 10600 -5275 10645 -5155
rect 10765 -5275 10810 -5155
rect 10930 -5275 10975 -5155
rect 11095 -5275 11150 -5155
rect 11270 -5275 11315 -5155
rect 11435 -5275 11480 -5155
rect 11600 -5275 11645 -5155
rect 11765 -5275 11820 -5155
rect 11940 -5275 11985 -5155
rect 12105 -5275 12150 -5155
rect 12270 -5275 12315 -5155
rect 12435 -5275 12490 -5155
rect 12610 -5275 12635 -5155
rect 7105 -5320 12635 -5275
rect 7105 -5440 7130 -5320
rect 7250 -5440 7295 -5320
rect 7415 -5440 7460 -5320
rect 7580 -5440 7625 -5320
rect 7745 -5440 7800 -5320
rect 7920 -5440 7965 -5320
rect 8085 -5440 8130 -5320
rect 8250 -5440 8295 -5320
rect 8415 -5440 8470 -5320
rect 8590 -5440 8635 -5320
rect 8755 -5440 8800 -5320
rect 8920 -5440 8965 -5320
rect 9085 -5440 9140 -5320
rect 9260 -5440 9305 -5320
rect 9425 -5440 9470 -5320
rect 9590 -5440 9635 -5320
rect 9755 -5440 9810 -5320
rect 9930 -5440 9975 -5320
rect 10095 -5440 10140 -5320
rect 10260 -5440 10305 -5320
rect 10425 -5440 10480 -5320
rect 10600 -5440 10645 -5320
rect 10765 -5440 10810 -5320
rect 10930 -5440 10975 -5320
rect 11095 -5440 11150 -5320
rect 11270 -5440 11315 -5320
rect 11435 -5440 11480 -5320
rect 11600 -5440 11645 -5320
rect 11765 -5440 11820 -5320
rect 11940 -5440 11985 -5320
rect 12105 -5440 12150 -5320
rect 12270 -5440 12315 -5320
rect 12435 -5440 12490 -5320
rect 12610 -5440 12635 -5320
rect 7105 -5485 12635 -5440
rect 7105 -5605 7130 -5485
rect 7250 -5605 7295 -5485
rect 7415 -5605 7460 -5485
rect 7580 -5605 7625 -5485
rect 7745 -5605 7800 -5485
rect 7920 -5605 7965 -5485
rect 8085 -5605 8130 -5485
rect 8250 -5605 8295 -5485
rect 8415 -5605 8470 -5485
rect 8590 -5605 8635 -5485
rect 8755 -5605 8800 -5485
rect 8920 -5605 8965 -5485
rect 9085 -5605 9140 -5485
rect 9260 -5605 9305 -5485
rect 9425 -5605 9470 -5485
rect 9590 -5605 9635 -5485
rect 9755 -5605 9810 -5485
rect 9930 -5605 9975 -5485
rect 10095 -5605 10140 -5485
rect 10260 -5605 10305 -5485
rect 10425 -5605 10480 -5485
rect 10600 -5605 10645 -5485
rect 10765 -5605 10810 -5485
rect 10930 -5605 10975 -5485
rect 11095 -5605 11150 -5485
rect 11270 -5605 11315 -5485
rect 11435 -5605 11480 -5485
rect 11600 -5605 11645 -5485
rect 11765 -5605 11820 -5485
rect 11940 -5605 11985 -5485
rect 12105 -5605 12150 -5485
rect 12270 -5605 12315 -5485
rect 12435 -5605 12490 -5485
rect 12610 -5605 12635 -5485
rect 7105 -5650 12635 -5605
rect 7105 -5770 7130 -5650
rect 7250 -5770 7295 -5650
rect 7415 -5770 7460 -5650
rect 7580 -5770 7625 -5650
rect 7745 -5770 7800 -5650
rect 7920 -5770 7965 -5650
rect 8085 -5770 8130 -5650
rect 8250 -5770 8295 -5650
rect 8415 -5770 8470 -5650
rect 8590 -5770 8635 -5650
rect 8755 -5770 8800 -5650
rect 8920 -5770 8965 -5650
rect 9085 -5770 9140 -5650
rect 9260 -5770 9305 -5650
rect 9425 -5770 9470 -5650
rect 9590 -5770 9635 -5650
rect 9755 -5770 9810 -5650
rect 9930 -5770 9975 -5650
rect 10095 -5770 10140 -5650
rect 10260 -5770 10305 -5650
rect 10425 -5770 10480 -5650
rect 10600 -5770 10645 -5650
rect 10765 -5770 10810 -5650
rect 10930 -5770 10975 -5650
rect 11095 -5770 11150 -5650
rect 11270 -5770 11315 -5650
rect 11435 -5770 11480 -5650
rect 11600 -5770 11645 -5650
rect 11765 -5770 11820 -5650
rect 11940 -5770 11985 -5650
rect 12105 -5770 12150 -5650
rect 12270 -5770 12315 -5650
rect 12435 -5770 12490 -5650
rect 12610 -5770 12635 -5650
rect 7105 -5825 12635 -5770
rect 7105 -5945 7130 -5825
rect 7250 -5945 7295 -5825
rect 7415 -5945 7460 -5825
rect 7580 -5945 7625 -5825
rect 7745 -5945 7800 -5825
rect 7920 -5945 7965 -5825
rect 8085 -5945 8130 -5825
rect 8250 -5945 8295 -5825
rect 8415 -5945 8470 -5825
rect 8590 -5945 8635 -5825
rect 8755 -5945 8800 -5825
rect 8920 -5945 8965 -5825
rect 9085 -5945 9140 -5825
rect 9260 -5945 9305 -5825
rect 9425 -5945 9470 -5825
rect 9590 -5945 9635 -5825
rect 9755 -5945 9810 -5825
rect 9930 -5945 9975 -5825
rect 10095 -5945 10140 -5825
rect 10260 -5945 10305 -5825
rect 10425 -5945 10480 -5825
rect 10600 -5945 10645 -5825
rect 10765 -5945 10810 -5825
rect 10930 -5945 10975 -5825
rect 11095 -5945 11150 -5825
rect 11270 -5945 11315 -5825
rect 11435 -5945 11480 -5825
rect 11600 -5945 11645 -5825
rect 11765 -5945 11820 -5825
rect 11940 -5945 11985 -5825
rect 12105 -5945 12150 -5825
rect 12270 -5945 12315 -5825
rect 12435 -5945 12490 -5825
rect 12610 -5945 12635 -5825
rect 7105 -5990 12635 -5945
rect 7105 -6110 7130 -5990
rect 7250 -6110 7295 -5990
rect 7415 -6110 7460 -5990
rect 7580 -6110 7625 -5990
rect 7745 -6110 7800 -5990
rect 7920 -6110 7965 -5990
rect 8085 -6110 8130 -5990
rect 8250 -6110 8295 -5990
rect 8415 -6110 8470 -5990
rect 8590 -6110 8635 -5990
rect 8755 -6110 8800 -5990
rect 8920 -6110 8965 -5990
rect 9085 -6110 9140 -5990
rect 9260 -6110 9305 -5990
rect 9425 -6110 9470 -5990
rect 9590 -6110 9635 -5990
rect 9755 -6110 9810 -5990
rect 9930 -6110 9975 -5990
rect 10095 -6110 10140 -5990
rect 10260 -6110 10305 -5990
rect 10425 -6110 10480 -5990
rect 10600 -6110 10645 -5990
rect 10765 -6110 10810 -5990
rect 10930 -6110 10975 -5990
rect 11095 -6110 11150 -5990
rect 11270 -6110 11315 -5990
rect 11435 -6110 11480 -5990
rect 11600 -6110 11645 -5990
rect 11765 -6110 11820 -5990
rect 11940 -6110 11985 -5990
rect 12105 -6110 12150 -5990
rect 12270 -6110 12315 -5990
rect 12435 -6110 12490 -5990
rect 12610 -6110 12635 -5990
rect 7105 -6155 12635 -6110
rect 7105 -6275 7130 -6155
rect 7250 -6275 7295 -6155
rect 7415 -6275 7460 -6155
rect 7580 -6275 7625 -6155
rect 7745 -6275 7800 -6155
rect 7920 -6275 7965 -6155
rect 8085 -6275 8130 -6155
rect 8250 -6275 8295 -6155
rect 8415 -6275 8470 -6155
rect 8590 -6275 8635 -6155
rect 8755 -6275 8800 -6155
rect 8920 -6275 8965 -6155
rect 9085 -6275 9140 -6155
rect 9260 -6275 9305 -6155
rect 9425 -6275 9470 -6155
rect 9590 -6275 9635 -6155
rect 9755 -6275 9810 -6155
rect 9930 -6275 9975 -6155
rect 10095 -6275 10140 -6155
rect 10260 -6275 10305 -6155
rect 10425 -6275 10480 -6155
rect 10600 -6275 10645 -6155
rect 10765 -6275 10810 -6155
rect 10930 -6275 10975 -6155
rect 11095 -6275 11150 -6155
rect 11270 -6275 11315 -6155
rect 11435 -6275 11480 -6155
rect 11600 -6275 11645 -6155
rect 11765 -6275 11820 -6155
rect 11940 -6275 11985 -6155
rect 12105 -6275 12150 -6155
rect 12270 -6275 12315 -6155
rect 12435 -6275 12490 -6155
rect 12610 -6275 12635 -6155
rect 7105 -6320 12635 -6275
rect 7105 -6440 7130 -6320
rect 7250 -6440 7295 -6320
rect 7415 -6440 7460 -6320
rect 7580 -6440 7625 -6320
rect 7745 -6440 7800 -6320
rect 7920 -6440 7965 -6320
rect 8085 -6440 8130 -6320
rect 8250 -6440 8295 -6320
rect 8415 -6440 8470 -6320
rect 8590 -6440 8635 -6320
rect 8755 -6440 8800 -6320
rect 8920 -6440 8965 -6320
rect 9085 -6440 9140 -6320
rect 9260 -6440 9305 -6320
rect 9425 -6440 9470 -6320
rect 9590 -6440 9635 -6320
rect 9755 -6440 9810 -6320
rect 9930 -6440 9975 -6320
rect 10095 -6440 10140 -6320
rect 10260 -6440 10305 -6320
rect 10425 -6440 10480 -6320
rect 10600 -6440 10645 -6320
rect 10765 -6440 10810 -6320
rect 10930 -6440 10975 -6320
rect 11095 -6440 11150 -6320
rect 11270 -6440 11315 -6320
rect 11435 -6440 11480 -6320
rect 11600 -6440 11645 -6320
rect 11765 -6440 11820 -6320
rect 11940 -6440 11985 -6320
rect 12105 -6440 12150 -6320
rect 12270 -6440 12315 -6320
rect 12435 -6440 12490 -6320
rect 12610 -6440 12635 -6320
rect 7105 -6495 12635 -6440
rect 7105 -6615 7130 -6495
rect 7250 -6615 7295 -6495
rect 7415 -6615 7460 -6495
rect 7580 -6615 7625 -6495
rect 7745 -6615 7800 -6495
rect 7920 -6615 7965 -6495
rect 8085 -6615 8130 -6495
rect 8250 -6615 8295 -6495
rect 8415 -6615 8470 -6495
rect 8590 -6615 8635 -6495
rect 8755 -6615 8800 -6495
rect 8920 -6615 8965 -6495
rect 9085 -6615 9140 -6495
rect 9260 -6615 9305 -6495
rect 9425 -6615 9470 -6495
rect 9590 -6615 9635 -6495
rect 9755 -6615 9810 -6495
rect 9930 -6615 9975 -6495
rect 10095 -6615 10140 -6495
rect 10260 -6615 10305 -6495
rect 10425 -6615 10480 -6495
rect 10600 -6615 10645 -6495
rect 10765 -6615 10810 -6495
rect 10930 -6615 10975 -6495
rect 11095 -6615 11150 -6495
rect 11270 -6615 11315 -6495
rect 11435 -6615 11480 -6495
rect 11600 -6615 11645 -6495
rect 11765 -6615 11820 -6495
rect 11940 -6615 11985 -6495
rect 12105 -6615 12150 -6495
rect 12270 -6615 12315 -6495
rect 12435 -6615 12490 -6495
rect 12610 -6615 12635 -6495
rect 7105 -6660 12635 -6615
rect 7105 -6780 7130 -6660
rect 7250 -6780 7295 -6660
rect 7415 -6780 7460 -6660
rect 7580 -6780 7625 -6660
rect 7745 -6780 7800 -6660
rect 7920 -6780 7965 -6660
rect 8085 -6780 8130 -6660
rect 8250 -6780 8295 -6660
rect 8415 -6780 8470 -6660
rect 8590 -6780 8635 -6660
rect 8755 -6780 8800 -6660
rect 8920 -6780 8965 -6660
rect 9085 -6780 9140 -6660
rect 9260 -6780 9305 -6660
rect 9425 -6780 9470 -6660
rect 9590 -6780 9635 -6660
rect 9755 -6780 9810 -6660
rect 9930 -6780 9975 -6660
rect 10095 -6780 10140 -6660
rect 10260 -6780 10305 -6660
rect 10425 -6780 10480 -6660
rect 10600 -6780 10645 -6660
rect 10765 -6780 10810 -6660
rect 10930 -6780 10975 -6660
rect 11095 -6780 11150 -6660
rect 11270 -6780 11315 -6660
rect 11435 -6780 11480 -6660
rect 11600 -6780 11645 -6660
rect 11765 -6780 11820 -6660
rect 11940 -6780 11985 -6660
rect 12105 -6780 12150 -6660
rect 12270 -6780 12315 -6660
rect 12435 -6780 12490 -6660
rect 12610 -6780 12635 -6660
rect 7105 -6825 12635 -6780
rect 7105 -6945 7130 -6825
rect 7250 -6945 7295 -6825
rect 7415 -6945 7460 -6825
rect 7580 -6945 7625 -6825
rect 7745 -6945 7800 -6825
rect 7920 -6945 7965 -6825
rect 8085 -6945 8130 -6825
rect 8250 -6945 8295 -6825
rect 8415 -6945 8470 -6825
rect 8590 -6945 8635 -6825
rect 8755 -6945 8800 -6825
rect 8920 -6945 8965 -6825
rect 9085 -6945 9140 -6825
rect 9260 -6945 9305 -6825
rect 9425 -6945 9470 -6825
rect 9590 -6945 9635 -6825
rect 9755 -6945 9810 -6825
rect 9930 -6945 9975 -6825
rect 10095 -6945 10140 -6825
rect 10260 -6945 10305 -6825
rect 10425 -6945 10480 -6825
rect 10600 -6945 10645 -6825
rect 10765 -6945 10810 -6825
rect 10930 -6945 10975 -6825
rect 11095 -6945 11150 -6825
rect 11270 -6945 11315 -6825
rect 11435 -6945 11480 -6825
rect 11600 -6945 11645 -6825
rect 11765 -6945 11820 -6825
rect 11940 -6945 11985 -6825
rect 12105 -6945 12150 -6825
rect 12270 -6945 12315 -6825
rect 12435 -6945 12490 -6825
rect 12610 -6945 12635 -6825
rect 7105 -6990 12635 -6945
rect 7105 -7110 7130 -6990
rect 7250 -7110 7295 -6990
rect 7415 -7110 7460 -6990
rect 7580 -7110 7625 -6990
rect 7745 -7110 7800 -6990
rect 7920 -7110 7965 -6990
rect 8085 -7110 8130 -6990
rect 8250 -7110 8295 -6990
rect 8415 -7110 8470 -6990
rect 8590 -7110 8635 -6990
rect 8755 -7110 8800 -6990
rect 8920 -7110 8965 -6990
rect 9085 -7110 9140 -6990
rect 9260 -7110 9305 -6990
rect 9425 -7110 9470 -6990
rect 9590 -7110 9635 -6990
rect 9755 -7110 9810 -6990
rect 9930 -7110 9975 -6990
rect 10095 -7110 10140 -6990
rect 10260 -7110 10305 -6990
rect 10425 -7110 10480 -6990
rect 10600 -7110 10645 -6990
rect 10765 -7110 10810 -6990
rect 10930 -7110 10975 -6990
rect 11095 -7110 11150 -6990
rect 11270 -7110 11315 -6990
rect 11435 -7110 11480 -6990
rect 11600 -7110 11645 -6990
rect 11765 -7110 11820 -6990
rect 11940 -7110 11985 -6990
rect 12105 -7110 12150 -6990
rect 12270 -7110 12315 -6990
rect 12435 -7110 12490 -6990
rect 12610 -7110 12635 -6990
rect 7105 -7165 12635 -7110
rect 7105 -7285 7130 -7165
rect 7250 -7285 7295 -7165
rect 7415 -7285 7460 -7165
rect 7580 -7285 7625 -7165
rect 7745 -7285 7800 -7165
rect 7920 -7285 7965 -7165
rect 8085 -7285 8130 -7165
rect 8250 -7285 8295 -7165
rect 8415 -7285 8470 -7165
rect 8590 -7285 8635 -7165
rect 8755 -7285 8800 -7165
rect 8920 -7285 8965 -7165
rect 9085 -7285 9140 -7165
rect 9260 -7285 9305 -7165
rect 9425 -7285 9470 -7165
rect 9590 -7285 9635 -7165
rect 9755 -7285 9810 -7165
rect 9930 -7285 9975 -7165
rect 10095 -7285 10140 -7165
rect 10260 -7285 10305 -7165
rect 10425 -7285 10480 -7165
rect 10600 -7285 10645 -7165
rect 10765 -7285 10810 -7165
rect 10930 -7285 10975 -7165
rect 11095 -7285 11150 -7165
rect 11270 -7285 11315 -7165
rect 11435 -7285 11480 -7165
rect 11600 -7285 11645 -7165
rect 11765 -7285 11820 -7165
rect 11940 -7285 11985 -7165
rect 12105 -7285 12150 -7165
rect 12270 -7285 12315 -7165
rect 12435 -7285 12490 -7165
rect 12610 -7285 12635 -7165
rect 7105 -7330 12635 -7285
rect 7105 -7450 7130 -7330
rect 7250 -7450 7295 -7330
rect 7415 -7450 7460 -7330
rect 7580 -7450 7625 -7330
rect 7745 -7450 7800 -7330
rect 7920 -7450 7965 -7330
rect 8085 -7450 8130 -7330
rect 8250 -7450 8295 -7330
rect 8415 -7450 8470 -7330
rect 8590 -7450 8635 -7330
rect 8755 -7450 8800 -7330
rect 8920 -7450 8965 -7330
rect 9085 -7450 9140 -7330
rect 9260 -7450 9305 -7330
rect 9425 -7450 9470 -7330
rect 9590 -7450 9635 -7330
rect 9755 -7450 9810 -7330
rect 9930 -7450 9975 -7330
rect 10095 -7450 10140 -7330
rect 10260 -7450 10305 -7330
rect 10425 -7450 10480 -7330
rect 10600 -7450 10645 -7330
rect 10765 -7450 10810 -7330
rect 10930 -7450 10975 -7330
rect 11095 -7450 11150 -7330
rect 11270 -7450 11315 -7330
rect 11435 -7450 11480 -7330
rect 11600 -7450 11645 -7330
rect 11765 -7450 11820 -7330
rect 11940 -7450 11985 -7330
rect 12105 -7450 12150 -7330
rect 12270 -7450 12315 -7330
rect 12435 -7450 12490 -7330
rect 12610 -7450 12635 -7330
rect 7105 -7495 12635 -7450
rect 7105 -7615 7130 -7495
rect 7250 -7615 7295 -7495
rect 7415 -7615 7460 -7495
rect 7580 -7615 7625 -7495
rect 7745 -7615 7800 -7495
rect 7920 -7615 7965 -7495
rect 8085 -7615 8130 -7495
rect 8250 -7615 8295 -7495
rect 8415 -7615 8470 -7495
rect 8590 -7615 8635 -7495
rect 8755 -7615 8800 -7495
rect 8920 -7615 8965 -7495
rect 9085 -7615 9140 -7495
rect 9260 -7615 9305 -7495
rect 9425 -7615 9470 -7495
rect 9590 -7615 9635 -7495
rect 9755 -7615 9810 -7495
rect 9930 -7615 9975 -7495
rect 10095 -7615 10140 -7495
rect 10260 -7615 10305 -7495
rect 10425 -7615 10480 -7495
rect 10600 -7615 10645 -7495
rect 10765 -7615 10810 -7495
rect 10930 -7615 10975 -7495
rect 11095 -7615 11150 -7495
rect 11270 -7615 11315 -7495
rect 11435 -7615 11480 -7495
rect 11600 -7615 11645 -7495
rect 11765 -7615 11820 -7495
rect 11940 -7615 11985 -7495
rect 12105 -7615 12150 -7495
rect 12270 -7615 12315 -7495
rect 12435 -7615 12490 -7495
rect 12610 -7615 12635 -7495
rect 7105 -7660 12635 -7615
rect 7105 -7780 7130 -7660
rect 7250 -7780 7295 -7660
rect 7415 -7780 7460 -7660
rect 7580 -7780 7625 -7660
rect 7745 -7780 7800 -7660
rect 7920 -7780 7965 -7660
rect 8085 -7780 8130 -7660
rect 8250 -7780 8295 -7660
rect 8415 -7780 8470 -7660
rect 8590 -7780 8635 -7660
rect 8755 -7780 8800 -7660
rect 8920 -7780 8965 -7660
rect 9085 -7780 9140 -7660
rect 9260 -7780 9305 -7660
rect 9425 -7780 9470 -7660
rect 9590 -7780 9635 -7660
rect 9755 -7780 9810 -7660
rect 9930 -7780 9975 -7660
rect 10095 -7780 10140 -7660
rect 10260 -7780 10305 -7660
rect 10425 -7780 10480 -7660
rect 10600 -7780 10645 -7660
rect 10765 -7780 10810 -7660
rect 10930 -7780 10975 -7660
rect 11095 -7780 11150 -7660
rect 11270 -7780 11315 -7660
rect 11435 -7780 11480 -7660
rect 11600 -7780 11645 -7660
rect 11765 -7780 11820 -7660
rect 11940 -7780 11985 -7660
rect 12105 -7780 12150 -7660
rect 12270 -7780 12315 -7660
rect 12435 -7780 12490 -7660
rect 12610 -7780 12635 -7660
rect 7105 -7835 12635 -7780
rect 7105 -7955 7130 -7835
rect 7250 -7955 7295 -7835
rect 7415 -7955 7460 -7835
rect 7580 -7955 7625 -7835
rect 7745 -7955 7800 -7835
rect 7920 -7955 7965 -7835
rect 8085 -7955 8130 -7835
rect 8250 -7955 8295 -7835
rect 8415 -7955 8470 -7835
rect 8590 -7955 8635 -7835
rect 8755 -7955 8800 -7835
rect 8920 -7955 8965 -7835
rect 9085 -7955 9140 -7835
rect 9260 -7955 9305 -7835
rect 9425 -7955 9470 -7835
rect 9590 -7955 9635 -7835
rect 9755 -7955 9810 -7835
rect 9930 -7955 9975 -7835
rect 10095 -7955 10140 -7835
rect 10260 -7955 10305 -7835
rect 10425 -7955 10480 -7835
rect 10600 -7955 10645 -7835
rect 10765 -7955 10810 -7835
rect 10930 -7955 10975 -7835
rect 11095 -7955 11150 -7835
rect 11270 -7955 11315 -7835
rect 11435 -7955 11480 -7835
rect 11600 -7955 11645 -7835
rect 11765 -7955 11820 -7835
rect 11940 -7955 11985 -7835
rect 12105 -7955 12150 -7835
rect 12270 -7955 12315 -7835
rect 12435 -7955 12490 -7835
rect 12610 -7955 12635 -7835
rect 7105 -8000 12635 -7955
rect 7105 -8120 7130 -8000
rect 7250 -8120 7295 -8000
rect 7415 -8120 7460 -8000
rect 7580 -8120 7625 -8000
rect 7745 -8120 7800 -8000
rect 7920 -8120 7965 -8000
rect 8085 -8120 8130 -8000
rect 8250 -8120 8295 -8000
rect 8415 -8120 8470 -8000
rect 8590 -8120 8635 -8000
rect 8755 -8120 8800 -8000
rect 8920 -8120 8965 -8000
rect 9085 -8120 9140 -8000
rect 9260 -8120 9305 -8000
rect 9425 -8120 9470 -8000
rect 9590 -8120 9635 -8000
rect 9755 -8120 9810 -8000
rect 9930 -8120 9975 -8000
rect 10095 -8120 10140 -8000
rect 10260 -8120 10305 -8000
rect 10425 -8120 10480 -8000
rect 10600 -8120 10645 -8000
rect 10765 -8120 10810 -8000
rect 10930 -8120 10975 -8000
rect 11095 -8120 11150 -8000
rect 11270 -8120 11315 -8000
rect 11435 -8120 11480 -8000
rect 11600 -8120 11645 -8000
rect 11765 -8120 11820 -8000
rect 11940 -8120 11985 -8000
rect 12105 -8120 12150 -8000
rect 12270 -8120 12315 -8000
rect 12435 -8120 12490 -8000
rect 12610 -8120 12635 -8000
rect 7105 -8165 12635 -8120
rect 7105 -8285 7130 -8165
rect 7250 -8285 7295 -8165
rect 7415 -8285 7460 -8165
rect 7580 -8285 7625 -8165
rect 7745 -8285 7800 -8165
rect 7920 -8285 7965 -8165
rect 8085 -8285 8130 -8165
rect 8250 -8285 8295 -8165
rect 8415 -8285 8470 -8165
rect 8590 -8285 8635 -8165
rect 8755 -8285 8800 -8165
rect 8920 -8285 8965 -8165
rect 9085 -8285 9140 -8165
rect 9260 -8285 9305 -8165
rect 9425 -8285 9470 -8165
rect 9590 -8285 9635 -8165
rect 9755 -8285 9810 -8165
rect 9930 -8285 9975 -8165
rect 10095 -8285 10140 -8165
rect 10260 -8285 10305 -8165
rect 10425 -8285 10480 -8165
rect 10600 -8285 10645 -8165
rect 10765 -8285 10810 -8165
rect 10930 -8285 10975 -8165
rect 11095 -8285 11150 -8165
rect 11270 -8285 11315 -8165
rect 11435 -8285 11480 -8165
rect 11600 -8285 11645 -8165
rect 11765 -8285 11820 -8165
rect 11940 -8285 11985 -8165
rect 12105 -8285 12150 -8165
rect 12270 -8285 12315 -8165
rect 12435 -8285 12490 -8165
rect 12610 -8285 12635 -8165
rect 7105 -8330 12635 -8285
rect 7105 -8450 7130 -8330
rect 7250 -8450 7295 -8330
rect 7415 -8450 7460 -8330
rect 7580 -8450 7625 -8330
rect 7745 -8450 7800 -8330
rect 7920 -8450 7965 -8330
rect 8085 -8450 8130 -8330
rect 8250 -8450 8295 -8330
rect 8415 -8450 8470 -8330
rect 8590 -8450 8635 -8330
rect 8755 -8450 8800 -8330
rect 8920 -8450 8965 -8330
rect 9085 -8450 9140 -8330
rect 9260 -8450 9305 -8330
rect 9425 -8450 9470 -8330
rect 9590 -8450 9635 -8330
rect 9755 -8450 9810 -8330
rect 9930 -8450 9975 -8330
rect 10095 -8450 10140 -8330
rect 10260 -8450 10305 -8330
rect 10425 -8450 10480 -8330
rect 10600 -8450 10645 -8330
rect 10765 -8450 10810 -8330
rect 10930 -8450 10975 -8330
rect 11095 -8450 11150 -8330
rect 11270 -8450 11315 -8330
rect 11435 -8450 11480 -8330
rect 11600 -8450 11645 -8330
rect 11765 -8450 11820 -8330
rect 11940 -8450 11985 -8330
rect 12105 -8450 12150 -8330
rect 12270 -8450 12315 -8330
rect 12435 -8450 12490 -8330
rect 12610 -8450 12635 -8330
rect 7105 -8505 12635 -8450
rect 7105 -8625 7130 -8505
rect 7250 -8625 7295 -8505
rect 7415 -8625 7460 -8505
rect 7580 -8625 7625 -8505
rect 7745 -8625 7800 -8505
rect 7920 -8625 7965 -8505
rect 8085 -8625 8130 -8505
rect 8250 -8625 8295 -8505
rect 8415 -8625 8470 -8505
rect 8590 -8625 8635 -8505
rect 8755 -8625 8800 -8505
rect 8920 -8625 8965 -8505
rect 9085 -8625 9140 -8505
rect 9260 -8625 9305 -8505
rect 9425 -8625 9470 -8505
rect 9590 -8625 9635 -8505
rect 9755 -8625 9810 -8505
rect 9930 -8625 9975 -8505
rect 10095 -8625 10140 -8505
rect 10260 -8625 10305 -8505
rect 10425 -8625 10480 -8505
rect 10600 -8625 10645 -8505
rect 10765 -8625 10810 -8505
rect 10930 -8625 10975 -8505
rect 11095 -8625 11150 -8505
rect 11270 -8625 11315 -8505
rect 11435 -8625 11480 -8505
rect 11600 -8625 11645 -8505
rect 11765 -8625 11820 -8505
rect 11940 -8625 11985 -8505
rect 12105 -8625 12150 -8505
rect 12270 -8625 12315 -8505
rect 12435 -8625 12490 -8505
rect 12610 -8625 12635 -8505
rect 7105 -8670 12635 -8625
rect 7105 -8790 7130 -8670
rect 7250 -8790 7295 -8670
rect 7415 -8790 7460 -8670
rect 7580 -8790 7625 -8670
rect 7745 -8790 7800 -8670
rect 7920 -8790 7965 -8670
rect 8085 -8790 8130 -8670
rect 8250 -8790 8295 -8670
rect 8415 -8790 8470 -8670
rect 8590 -8790 8635 -8670
rect 8755 -8790 8800 -8670
rect 8920 -8790 8965 -8670
rect 9085 -8790 9140 -8670
rect 9260 -8790 9305 -8670
rect 9425 -8790 9470 -8670
rect 9590 -8790 9635 -8670
rect 9755 -8790 9810 -8670
rect 9930 -8790 9975 -8670
rect 10095 -8790 10140 -8670
rect 10260 -8790 10305 -8670
rect 10425 -8790 10480 -8670
rect 10600 -8790 10645 -8670
rect 10765 -8790 10810 -8670
rect 10930 -8790 10975 -8670
rect 11095 -8790 11150 -8670
rect 11270 -8790 11315 -8670
rect 11435 -8790 11480 -8670
rect 11600 -8790 11645 -8670
rect 11765 -8790 11820 -8670
rect 11940 -8790 11985 -8670
rect 12105 -8790 12150 -8670
rect 12270 -8790 12315 -8670
rect 12435 -8790 12490 -8670
rect 12610 -8790 12635 -8670
rect 7105 -8835 12635 -8790
rect 7105 -8955 7130 -8835
rect 7250 -8955 7295 -8835
rect 7415 -8955 7460 -8835
rect 7580 -8955 7625 -8835
rect 7745 -8955 7800 -8835
rect 7920 -8955 7965 -8835
rect 8085 -8955 8130 -8835
rect 8250 -8955 8295 -8835
rect 8415 -8955 8470 -8835
rect 8590 -8955 8635 -8835
rect 8755 -8955 8800 -8835
rect 8920 -8955 8965 -8835
rect 9085 -8955 9140 -8835
rect 9260 -8955 9305 -8835
rect 9425 -8955 9470 -8835
rect 9590 -8955 9635 -8835
rect 9755 -8955 9810 -8835
rect 9930 -8955 9975 -8835
rect 10095 -8955 10140 -8835
rect 10260 -8955 10305 -8835
rect 10425 -8955 10480 -8835
rect 10600 -8955 10645 -8835
rect 10765 -8955 10810 -8835
rect 10930 -8955 10975 -8835
rect 11095 -8955 11150 -8835
rect 11270 -8955 11315 -8835
rect 11435 -8955 11480 -8835
rect 11600 -8955 11645 -8835
rect 11765 -8955 11820 -8835
rect 11940 -8955 11985 -8835
rect 12105 -8955 12150 -8835
rect 12270 -8955 12315 -8835
rect 12435 -8955 12490 -8835
rect 12610 -8955 12635 -8835
rect 7105 -9000 12635 -8955
rect 7105 -9120 7130 -9000
rect 7250 -9120 7295 -9000
rect 7415 -9120 7460 -9000
rect 7580 -9120 7625 -9000
rect 7745 -9120 7800 -9000
rect 7920 -9120 7965 -9000
rect 8085 -9120 8130 -9000
rect 8250 -9120 8295 -9000
rect 8415 -9120 8470 -9000
rect 8590 -9120 8635 -9000
rect 8755 -9120 8800 -9000
rect 8920 -9120 8965 -9000
rect 9085 -9120 9140 -9000
rect 9260 -9120 9305 -9000
rect 9425 -9120 9470 -9000
rect 9590 -9120 9635 -9000
rect 9755 -9120 9810 -9000
rect 9930 -9120 9975 -9000
rect 10095 -9120 10140 -9000
rect 10260 -9120 10305 -9000
rect 10425 -9120 10480 -9000
rect 10600 -9120 10645 -9000
rect 10765 -9120 10810 -9000
rect 10930 -9120 10975 -9000
rect 11095 -9120 11150 -9000
rect 11270 -9120 11315 -9000
rect 11435 -9120 11480 -9000
rect 11600 -9120 11645 -9000
rect 11765 -9120 11820 -9000
rect 11940 -9120 11985 -9000
rect 12105 -9120 12150 -9000
rect 12270 -9120 12315 -9000
rect 12435 -9120 12490 -9000
rect 12610 -9120 12635 -9000
rect 7105 -9175 12635 -9120
rect 7105 -9295 7130 -9175
rect 7250 -9295 7295 -9175
rect 7415 -9295 7460 -9175
rect 7580 -9295 7625 -9175
rect 7745 -9295 7800 -9175
rect 7920 -9295 7965 -9175
rect 8085 -9295 8130 -9175
rect 8250 -9295 8295 -9175
rect 8415 -9295 8470 -9175
rect 8590 -9295 8635 -9175
rect 8755 -9295 8800 -9175
rect 8920 -9295 8965 -9175
rect 9085 -9295 9140 -9175
rect 9260 -9295 9305 -9175
rect 9425 -9295 9470 -9175
rect 9590 -9295 9635 -9175
rect 9755 -9295 9810 -9175
rect 9930 -9295 9975 -9175
rect 10095 -9295 10140 -9175
rect 10260 -9295 10305 -9175
rect 10425 -9295 10480 -9175
rect 10600 -9295 10645 -9175
rect 10765 -9295 10810 -9175
rect 10930 -9295 10975 -9175
rect 11095 -9295 11150 -9175
rect 11270 -9295 11315 -9175
rect 11435 -9295 11480 -9175
rect 11600 -9295 11645 -9175
rect 11765 -9295 11820 -9175
rect 11940 -9295 11985 -9175
rect 12105 -9295 12150 -9175
rect 12270 -9295 12315 -9175
rect 12435 -9295 12490 -9175
rect 12610 -9295 12635 -9175
rect 7105 -9340 12635 -9295
rect 7105 -9460 7130 -9340
rect 7250 -9460 7295 -9340
rect 7415 -9460 7460 -9340
rect 7580 -9460 7625 -9340
rect 7745 -9460 7800 -9340
rect 7920 -9460 7965 -9340
rect 8085 -9460 8130 -9340
rect 8250 -9460 8295 -9340
rect 8415 -9460 8470 -9340
rect 8590 -9460 8635 -9340
rect 8755 -9460 8800 -9340
rect 8920 -9460 8965 -9340
rect 9085 -9460 9140 -9340
rect 9260 -9460 9305 -9340
rect 9425 -9460 9470 -9340
rect 9590 -9460 9635 -9340
rect 9755 -9460 9810 -9340
rect 9930 -9460 9975 -9340
rect 10095 -9460 10140 -9340
rect 10260 -9460 10305 -9340
rect 10425 -9460 10480 -9340
rect 10600 -9460 10645 -9340
rect 10765 -9460 10810 -9340
rect 10930 -9460 10975 -9340
rect 11095 -9460 11150 -9340
rect 11270 -9460 11315 -9340
rect 11435 -9460 11480 -9340
rect 11600 -9460 11645 -9340
rect 11765 -9460 11820 -9340
rect 11940 -9460 11985 -9340
rect 12105 -9460 12150 -9340
rect 12270 -9460 12315 -9340
rect 12435 -9460 12490 -9340
rect 12610 -9460 12635 -9340
rect 7105 -9505 12635 -9460
rect 7105 -9625 7130 -9505
rect 7250 -9625 7295 -9505
rect 7415 -9625 7460 -9505
rect 7580 -9625 7625 -9505
rect 7745 -9625 7800 -9505
rect 7920 -9625 7965 -9505
rect 8085 -9625 8130 -9505
rect 8250 -9625 8295 -9505
rect 8415 -9625 8470 -9505
rect 8590 -9625 8635 -9505
rect 8755 -9625 8800 -9505
rect 8920 -9625 8965 -9505
rect 9085 -9625 9140 -9505
rect 9260 -9625 9305 -9505
rect 9425 -9625 9470 -9505
rect 9590 -9625 9635 -9505
rect 9755 -9625 9810 -9505
rect 9930 -9625 9975 -9505
rect 10095 -9625 10140 -9505
rect 10260 -9625 10305 -9505
rect 10425 -9625 10480 -9505
rect 10600 -9625 10645 -9505
rect 10765 -9625 10810 -9505
rect 10930 -9625 10975 -9505
rect 11095 -9625 11150 -9505
rect 11270 -9625 11315 -9505
rect 11435 -9625 11480 -9505
rect 11600 -9625 11645 -9505
rect 11765 -9625 11820 -9505
rect 11940 -9625 11985 -9505
rect 12105 -9625 12150 -9505
rect 12270 -9625 12315 -9505
rect 12435 -9625 12490 -9505
rect 12610 -9625 12635 -9505
rect 7105 -9670 12635 -9625
rect 7105 -9790 7130 -9670
rect 7250 -9790 7295 -9670
rect 7415 -9790 7460 -9670
rect 7580 -9790 7625 -9670
rect 7745 -9790 7800 -9670
rect 7920 -9790 7965 -9670
rect 8085 -9790 8130 -9670
rect 8250 -9790 8295 -9670
rect 8415 -9790 8470 -9670
rect 8590 -9790 8635 -9670
rect 8755 -9790 8800 -9670
rect 8920 -9790 8965 -9670
rect 9085 -9790 9140 -9670
rect 9260 -9790 9305 -9670
rect 9425 -9790 9470 -9670
rect 9590 -9790 9635 -9670
rect 9755 -9790 9810 -9670
rect 9930 -9790 9975 -9670
rect 10095 -9790 10140 -9670
rect 10260 -9790 10305 -9670
rect 10425 -9790 10480 -9670
rect 10600 -9790 10645 -9670
rect 10765 -9790 10810 -9670
rect 10930 -9790 10975 -9670
rect 11095 -9790 11150 -9670
rect 11270 -9790 11315 -9670
rect 11435 -9790 11480 -9670
rect 11600 -9790 11645 -9670
rect 11765 -9790 11820 -9670
rect 11940 -9790 11985 -9670
rect 12105 -9790 12150 -9670
rect 12270 -9790 12315 -9670
rect 12435 -9790 12490 -9670
rect 12610 -9790 12635 -9670
rect 7105 -9815 12635 -9790
rect 12795 -4430 12820 -4345
rect 12940 -4430 12985 -4310
rect 13105 -4430 13150 -4310
rect 13270 -4430 13315 -4310
rect 13435 -4430 13490 -4310
rect 13610 -4430 13655 -4310
rect 13775 -4430 13820 -4310
rect 13940 -4430 13985 -4310
rect 14105 -4430 14160 -4310
rect 14280 -4430 14325 -4310
rect 14445 -4430 14490 -4310
rect 14610 -4430 14655 -4310
rect 14775 -4430 14830 -4310
rect 14950 -4430 14995 -4310
rect 15115 -4430 15160 -4310
rect 15280 -4430 15325 -4310
rect 15445 -4430 15500 -4310
rect 15620 -4430 15665 -4310
rect 15785 -4430 15830 -4310
rect 15950 -4430 15995 -4310
rect 16115 -4430 16170 -4310
rect 16290 -4430 16335 -4310
rect 16455 -4430 16500 -4310
rect 16620 -4430 16665 -4310
rect 16785 -4430 16840 -4310
rect 16960 -4430 17005 -4310
rect 17125 -4430 17170 -4310
rect 17290 -4430 17335 -4310
rect 17455 -4430 17510 -4310
rect 17630 -4430 17675 -4310
rect 17795 -4430 17840 -4310
rect 17960 -4430 18005 -4310
rect 18125 -4430 18180 -4310
rect 18300 -4345 18510 -4310
rect 18300 -4430 18325 -4345
rect 12795 -4485 18325 -4430
rect 12795 -4605 12820 -4485
rect 12940 -4605 12985 -4485
rect 13105 -4605 13150 -4485
rect 13270 -4605 13315 -4485
rect 13435 -4605 13490 -4485
rect 13610 -4605 13655 -4485
rect 13775 -4605 13820 -4485
rect 13940 -4605 13985 -4485
rect 14105 -4605 14160 -4485
rect 14280 -4605 14325 -4485
rect 14445 -4605 14490 -4485
rect 14610 -4605 14655 -4485
rect 14775 -4605 14830 -4485
rect 14950 -4605 14995 -4485
rect 15115 -4605 15160 -4485
rect 15280 -4605 15325 -4485
rect 15445 -4605 15500 -4485
rect 15620 -4605 15665 -4485
rect 15785 -4605 15830 -4485
rect 15950 -4605 15995 -4485
rect 16115 -4605 16170 -4485
rect 16290 -4605 16335 -4485
rect 16455 -4605 16500 -4485
rect 16620 -4605 16665 -4485
rect 16785 -4605 16840 -4485
rect 16960 -4605 17005 -4485
rect 17125 -4605 17170 -4485
rect 17290 -4605 17335 -4485
rect 17455 -4605 17510 -4485
rect 17630 -4605 17675 -4485
rect 17795 -4605 17840 -4485
rect 17960 -4605 18005 -4485
rect 18125 -4605 18180 -4485
rect 18300 -4605 18325 -4485
rect 12795 -4650 18325 -4605
rect 12795 -4770 12820 -4650
rect 12940 -4770 12985 -4650
rect 13105 -4770 13150 -4650
rect 13270 -4770 13315 -4650
rect 13435 -4770 13490 -4650
rect 13610 -4770 13655 -4650
rect 13775 -4770 13820 -4650
rect 13940 -4770 13985 -4650
rect 14105 -4770 14160 -4650
rect 14280 -4770 14325 -4650
rect 14445 -4770 14490 -4650
rect 14610 -4770 14655 -4650
rect 14775 -4770 14830 -4650
rect 14950 -4770 14995 -4650
rect 15115 -4770 15160 -4650
rect 15280 -4770 15325 -4650
rect 15445 -4770 15500 -4650
rect 15620 -4770 15665 -4650
rect 15785 -4770 15830 -4650
rect 15950 -4770 15995 -4650
rect 16115 -4770 16170 -4650
rect 16290 -4770 16335 -4650
rect 16455 -4770 16500 -4650
rect 16620 -4770 16665 -4650
rect 16785 -4770 16840 -4650
rect 16960 -4770 17005 -4650
rect 17125 -4770 17170 -4650
rect 17290 -4770 17335 -4650
rect 17455 -4770 17510 -4650
rect 17630 -4770 17675 -4650
rect 17795 -4770 17840 -4650
rect 17960 -4770 18005 -4650
rect 18125 -4770 18180 -4650
rect 18300 -4770 18325 -4650
rect 12795 -4815 18325 -4770
rect 12795 -4935 12820 -4815
rect 12940 -4935 12985 -4815
rect 13105 -4935 13150 -4815
rect 13270 -4935 13315 -4815
rect 13435 -4935 13490 -4815
rect 13610 -4935 13655 -4815
rect 13775 -4935 13820 -4815
rect 13940 -4935 13985 -4815
rect 14105 -4935 14160 -4815
rect 14280 -4935 14325 -4815
rect 14445 -4935 14490 -4815
rect 14610 -4935 14655 -4815
rect 14775 -4935 14830 -4815
rect 14950 -4935 14995 -4815
rect 15115 -4935 15160 -4815
rect 15280 -4935 15325 -4815
rect 15445 -4935 15500 -4815
rect 15620 -4935 15665 -4815
rect 15785 -4935 15830 -4815
rect 15950 -4935 15995 -4815
rect 16115 -4935 16170 -4815
rect 16290 -4935 16335 -4815
rect 16455 -4935 16500 -4815
rect 16620 -4935 16665 -4815
rect 16785 -4935 16840 -4815
rect 16960 -4935 17005 -4815
rect 17125 -4935 17170 -4815
rect 17290 -4935 17335 -4815
rect 17455 -4935 17510 -4815
rect 17630 -4935 17675 -4815
rect 17795 -4935 17840 -4815
rect 17960 -4935 18005 -4815
rect 18125 -4935 18180 -4815
rect 18300 -4935 18325 -4815
rect 12795 -4980 18325 -4935
rect 12795 -5100 12820 -4980
rect 12940 -5100 12985 -4980
rect 13105 -5100 13150 -4980
rect 13270 -5100 13315 -4980
rect 13435 -5100 13490 -4980
rect 13610 -5100 13655 -4980
rect 13775 -5100 13820 -4980
rect 13940 -5100 13985 -4980
rect 14105 -5100 14160 -4980
rect 14280 -5100 14325 -4980
rect 14445 -5100 14490 -4980
rect 14610 -5100 14655 -4980
rect 14775 -5100 14830 -4980
rect 14950 -5100 14995 -4980
rect 15115 -5100 15160 -4980
rect 15280 -5100 15325 -4980
rect 15445 -5100 15500 -4980
rect 15620 -5100 15665 -4980
rect 15785 -5100 15830 -4980
rect 15950 -5100 15995 -4980
rect 16115 -5100 16170 -4980
rect 16290 -5100 16335 -4980
rect 16455 -5100 16500 -4980
rect 16620 -5100 16665 -4980
rect 16785 -5100 16840 -4980
rect 16960 -5100 17005 -4980
rect 17125 -5100 17170 -4980
rect 17290 -5100 17335 -4980
rect 17455 -5100 17510 -4980
rect 17630 -5100 17675 -4980
rect 17795 -5100 17840 -4980
rect 17960 -5100 18005 -4980
rect 18125 -5100 18180 -4980
rect 18300 -5100 18325 -4980
rect 12795 -5155 18325 -5100
rect 12795 -5275 12820 -5155
rect 12940 -5275 12985 -5155
rect 13105 -5275 13150 -5155
rect 13270 -5275 13315 -5155
rect 13435 -5275 13490 -5155
rect 13610 -5275 13655 -5155
rect 13775 -5275 13820 -5155
rect 13940 -5275 13985 -5155
rect 14105 -5275 14160 -5155
rect 14280 -5275 14325 -5155
rect 14445 -5275 14490 -5155
rect 14610 -5275 14655 -5155
rect 14775 -5275 14830 -5155
rect 14950 -5275 14995 -5155
rect 15115 -5275 15160 -5155
rect 15280 -5275 15325 -5155
rect 15445 -5275 15500 -5155
rect 15620 -5275 15665 -5155
rect 15785 -5275 15830 -5155
rect 15950 -5275 15995 -5155
rect 16115 -5275 16170 -5155
rect 16290 -5275 16335 -5155
rect 16455 -5275 16500 -5155
rect 16620 -5275 16665 -5155
rect 16785 -5275 16840 -5155
rect 16960 -5275 17005 -5155
rect 17125 -5275 17170 -5155
rect 17290 -5275 17335 -5155
rect 17455 -5275 17510 -5155
rect 17630 -5275 17675 -5155
rect 17795 -5275 17840 -5155
rect 17960 -5275 18005 -5155
rect 18125 -5275 18180 -5155
rect 18300 -5275 18325 -5155
rect 12795 -5320 18325 -5275
rect 12795 -5440 12820 -5320
rect 12940 -5440 12985 -5320
rect 13105 -5440 13150 -5320
rect 13270 -5440 13315 -5320
rect 13435 -5440 13490 -5320
rect 13610 -5440 13655 -5320
rect 13775 -5440 13820 -5320
rect 13940 -5440 13985 -5320
rect 14105 -5440 14160 -5320
rect 14280 -5440 14325 -5320
rect 14445 -5440 14490 -5320
rect 14610 -5440 14655 -5320
rect 14775 -5440 14830 -5320
rect 14950 -5440 14995 -5320
rect 15115 -5440 15160 -5320
rect 15280 -5440 15325 -5320
rect 15445 -5440 15500 -5320
rect 15620 -5440 15665 -5320
rect 15785 -5440 15830 -5320
rect 15950 -5440 15995 -5320
rect 16115 -5440 16170 -5320
rect 16290 -5440 16335 -5320
rect 16455 -5440 16500 -5320
rect 16620 -5440 16665 -5320
rect 16785 -5440 16840 -5320
rect 16960 -5440 17005 -5320
rect 17125 -5440 17170 -5320
rect 17290 -5440 17335 -5320
rect 17455 -5440 17510 -5320
rect 17630 -5440 17675 -5320
rect 17795 -5440 17840 -5320
rect 17960 -5440 18005 -5320
rect 18125 -5440 18180 -5320
rect 18300 -5440 18325 -5320
rect 12795 -5485 18325 -5440
rect 12795 -5605 12820 -5485
rect 12940 -5605 12985 -5485
rect 13105 -5605 13150 -5485
rect 13270 -5605 13315 -5485
rect 13435 -5605 13490 -5485
rect 13610 -5605 13655 -5485
rect 13775 -5605 13820 -5485
rect 13940 -5605 13985 -5485
rect 14105 -5605 14160 -5485
rect 14280 -5605 14325 -5485
rect 14445 -5605 14490 -5485
rect 14610 -5605 14655 -5485
rect 14775 -5605 14830 -5485
rect 14950 -5605 14995 -5485
rect 15115 -5605 15160 -5485
rect 15280 -5605 15325 -5485
rect 15445 -5605 15500 -5485
rect 15620 -5605 15665 -5485
rect 15785 -5605 15830 -5485
rect 15950 -5605 15995 -5485
rect 16115 -5605 16170 -5485
rect 16290 -5605 16335 -5485
rect 16455 -5605 16500 -5485
rect 16620 -5605 16665 -5485
rect 16785 -5605 16840 -5485
rect 16960 -5605 17005 -5485
rect 17125 -5605 17170 -5485
rect 17290 -5605 17335 -5485
rect 17455 -5605 17510 -5485
rect 17630 -5605 17675 -5485
rect 17795 -5605 17840 -5485
rect 17960 -5605 18005 -5485
rect 18125 -5605 18180 -5485
rect 18300 -5605 18325 -5485
rect 12795 -5650 18325 -5605
rect 12795 -5770 12820 -5650
rect 12940 -5770 12985 -5650
rect 13105 -5770 13150 -5650
rect 13270 -5770 13315 -5650
rect 13435 -5770 13490 -5650
rect 13610 -5770 13655 -5650
rect 13775 -5770 13820 -5650
rect 13940 -5770 13985 -5650
rect 14105 -5770 14160 -5650
rect 14280 -5770 14325 -5650
rect 14445 -5770 14490 -5650
rect 14610 -5770 14655 -5650
rect 14775 -5770 14830 -5650
rect 14950 -5770 14995 -5650
rect 15115 -5770 15160 -5650
rect 15280 -5770 15325 -5650
rect 15445 -5770 15500 -5650
rect 15620 -5770 15665 -5650
rect 15785 -5770 15830 -5650
rect 15950 -5770 15995 -5650
rect 16115 -5770 16170 -5650
rect 16290 -5770 16335 -5650
rect 16455 -5770 16500 -5650
rect 16620 -5770 16665 -5650
rect 16785 -5770 16840 -5650
rect 16960 -5770 17005 -5650
rect 17125 -5770 17170 -5650
rect 17290 -5770 17335 -5650
rect 17455 -5770 17510 -5650
rect 17630 -5770 17675 -5650
rect 17795 -5770 17840 -5650
rect 17960 -5770 18005 -5650
rect 18125 -5770 18180 -5650
rect 18300 -5770 18325 -5650
rect 12795 -5825 18325 -5770
rect 12795 -5945 12820 -5825
rect 12940 -5945 12985 -5825
rect 13105 -5945 13150 -5825
rect 13270 -5945 13315 -5825
rect 13435 -5945 13490 -5825
rect 13610 -5945 13655 -5825
rect 13775 -5945 13820 -5825
rect 13940 -5945 13985 -5825
rect 14105 -5945 14160 -5825
rect 14280 -5945 14325 -5825
rect 14445 -5945 14490 -5825
rect 14610 -5945 14655 -5825
rect 14775 -5945 14830 -5825
rect 14950 -5945 14995 -5825
rect 15115 -5945 15160 -5825
rect 15280 -5945 15325 -5825
rect 15445 -5945 15500 -5825
rect 15620 -5945 15665 -5825
rect 15785 -5945 15830 -5825
rect 15950 -5945 15995 -5825
rect 16115 -5945 16170 -5825
rect 16290 -5945 16335 -5825
rect 16455 -5945 16500 -5825
rect 16620 -5945 16665 -5825
rect 16785 -5945 16840 -5825
rect 16960 -5945 17005 -5825
rect 17125 -5945 17170 -5825
rect 17290 -5945 17335 -5825
rect 17455 -5945 17510 -5825
rect 17630 -5945 17675 -5825
rect 17795 -5945 17840 -5825
rect 17960 -5945 18005 -5825
rect 18125 -5945 18180 -5825
rect 18300 -5945 18325 -5825
rect 12795 -5990 18325 -5945
rect 12795 -6110 12820 -5990
rect 12940 -6110 12985 -5990
rect 13105 -6110 13150 -5990
rect 13270 -6110 13315 -5990
rect 13435 -6110 13490 -5990
rect 13610 -6110 13655 -5990
rect 13775 -6110 13820 -5990
rect 13940 -6110 13985 -5990
rect 14105 -6110 14160 -5990
rect 14280 -6110 14325 -5990
rect 14445 -6110 14490 -5990
rect 14610 -6110 14655 -5990
rect 14775 -6110 14830 -5990
rect 14950 -6110 14995 -5990
rect 15115 -6110 15160 -5990
rect 15280 -6110 15325 -5990
rect 15445 -6110 15500 -5990
rect 15620 -6110 15665 -5990
rect 15785 -6110 15830 -5990
rect 15950 -6110 15995 -5990
rect 16115 -6110 16170 -5990
rect 16290 -6110 16335 -5990
rect 16455 -6110 16500 -5990
rect 16620 -6110 16665 -5990
rect 16785 -6110 16840 -5990
rect 16960 -6110 17005 -5990
rect 17125 -6110 17170 -5990
rect 17290 -6110 17335 -5990
rect 17455 -6110 17510 -5990
rect 17630 -6110 17675 -5990
rect 17795 -6110 17840 -5990
rect 17960 -6110 18005 -5990
rect 18125 -6110 18180 -5990
rect 18300 -6110 18325 -5990
rect 12795 -6155 18325 -6110
rect 12795 -6275 12820 -6155
rect 12940 -6275 12985 -6155
rect 13105 -6275 13150 -6155
rect 13270 -6275 13315 -6155
rect 13435 -6275 13490 -6155
rect 13610 -6275 13655 -6155
rect 13775 -6275 13820 -6155
rect 13940 -6275 13985 -6155
rect 14105 -6275 14160 -6155
rect 14280 -6275 14325 -6155
rect 14445 -6275 14490 -6155
rect 14610 -6275 14655 -6155
rect 14775 -6275 14830 -6155
rect 14950 -6275 14995 -6155
rect 15115 -6275 15160 -6155
rect 15280 -6275 15325 -6155
rect 15445 -6275 15500 -6155
rect 15620 -6275 15665 -6155
rect 15785 -6275 15830 -6155
rect 15950 -6275 15995 -6155
rect 16115 -6275 16170 -6155
rect 16290 -6275 16335 -6155
rect 16455 -6275 16500 -6155
rect 16620 -6275 16665 -6155
rect 16785 -6275 16840 -6155
rect 16960 -6275 17005 -6155
rect 17125 -6275 17170 -6155
rect 17290 -6275 17335 -6155
rect 17455 -6275 17510 -6155
rect 17630 -6275 17675 -6155
rect 17795 -6275 17840 -6155
rect 17960 -6275 18005 -6155
rect 18125 -6275 18180 -6155
rect 18300 -6275 18325 -6155
rect 12795 -6320 18325 -6275
rect 12795 -6440 12820 -6320
rect 12940 -6440 12985 -6320
rect 13105 -6440 13150 -6320
rect 13270 -6440 13315 -6320
rect 13435 -6440 13490 -6320
rect 13610 -6440 13655 -6320
rect 13775 -6440 13820 -6320
rect 13940 -6440 13985 -6320
rect 14105 -6440 14160 -6320
rect 14280 -6440 14325 -6320
rect 14445 -6440 14490 -6320
rect 14610 -6440 14655 -6320
rect 14775 -6440 14830 -6320
rect 14950 -6440 14995 -6320
rect 15115 -6440 15160 -6320
rect 15280 -6440 15325 -6320
rect 15445 -6440 15500 -6320
rect 15620 -6440 15665 -6320
rect 15785 -6440 15830 -6320
rect 15950 -6440 15995 -6320
rect 16115 -6440 16170 -6320
rect 16290 -6440 16335 -6320
rect 16455 -6440 16500 -6320
rect 16620 -6440 16665 -6320
rect 16785 -6440 16840 -6320
rect 16960 -6440 17005 -6320
rect 17125 -6440 17170 -6320
rect 17290 -6440 17335 -6320
rect 17455 -6440 17510 -6320
rect 17630 -6440 17675 -6320
rect 17795 -6440 17840 -6320
rect 17960 -6440 18005 -6320
rect 18125 -6440 18180 -6320
rect 18300 -6440 18325 -6320
rect 12795 -6495 18325 -6440
rect 12795 -6615 12820 -6495
rect 12940 -6615 12985 -6495
rect 13105 -6615 13150 -6495
rect 13270 -6615 13315 -6495
rect 13435 -6615 13490 -6495
rect 13610 -6615 13655 -6495
rect 13775 -6615 13820 -6495
rect 13940 -6615 13985 -6495
rect 14105 -6615 14160 -6495
rect 14280 -6615 14325 -6495
rect 14445 -6615 14490 -6495
rect 14610 -6615 14655 -6495
rect 14775 -6615 14830 -6495
rect 14950 -6615 14995 -6495
rect 15115 -6615 15160 -6495
rect 15280 -6615 15325 -6495
rect 15445 -6615 15500 -6495
rect 15620 -6615 15665 -6495
rect 15785 -6615 15830 -6495
rect 15950 -6615 15995 -6495
rect 16115 -6615 16170 -6495
rect 16290 -6615 16335 -6495
rect 16455 -6615 16500 -6495
rect 16620 -6615 16665 -6495
rect 16785 -6615 16840 -6495
rect 16960 -6615 17005 -6495
rect 17125 -6615 17170 -6495
rect 17290 -6615 17335 -6495
rect 17455 -6615 17510 -6495
rect 17630 -6615 17675 -6495
rect 17795 -6615 17840 -6495
rect 17960 -6615 18005 -6495
rect 18125 -6615 18180 -6495
rect 18300 -6615 18325 -6495
rect 12795 -6660 18325 -6615
rect 12795 -6780 12820 -6660
rect 12940 -6780 12985 -6660
rect 13105 -6780 13150 -6660
rect 13270 -6780 13315 -6660
rect 13435 -6780 13490 -6660
rect 13610 -6780 13655 -6660
rect 13775 -6780 13820 -6660
rect 13940 -6780 13985 -6660
rect 14105 -6780 14160 -6660
rect 14280 -6780 14325 -6660
rect 14445 -6780 14490 -6660
rect 14610 -6780 14655 -6660
rect 14775 -6780 14830 -6660
rect 14950 -6780 14995 -6660
rect 15115 -6780 15160 -6660
rect 15280 -6780 15325 -6660
rect 15445 -6780 15500 -6660
rect 15620 -6780 15665 -6660
rect 15785 -6780 15830 -6660
rect 15950 -6780 15995 -6660
rect 16115 -6780 16170 -6660
rect 16290 -6780 16335 -6660
rect 16455 -6780 16500 -6660
rect 16620 -6780 16665 -6660
rect 16785 -6780 16840 -6660
rect 16960 -6780 17005 -6660
rect 17125 -6780 17170 -6660
rect 17290 -6780 17335 -6660
rect 17455 -6780 17510 -6660
rect 17630 -6780 17675 -6660
rect 17795 -6780 17840 -6660
rect 17960 -6780 18005 -6660
rect 18125 -6780 18180 -6660
rect 18300 -6780 18325 -6660
rect 12795 -6825 18325 -6780
rect 12795 -6945 12820 -6825
rect 12940 -6945 12985 -6825
rect 13105 -6945 13150 -6825
rect 13270 -6945 13315 -6825
rect 13435 -6945 13490 -6825
rect 13610 -6945 13655 -6825
rect 13775 -6945 13820 -6825
rect 13940 -6945 13985 -6825
rect 14105 -6945 14160 -6825
rect 14280 -6945 14325 -6825
rect 14445 -6945 14490 -6825
rect 14610 -6945 14655 -6825
rect 14775 -6945 14830 -6825
rect 14950 -6945 14995 -6825
rect 15115 -6945 15160 -6825
rect 15280 -6945 15325 -6825
rect 15445 -6945 15500 -6825
rect 15620 -6945 15665 -6825
rect 15785 -6945 15830 -6825
rect 15950 -6945 15995 -6825
rect 16115 -6945 16170 -6825
rect 16290 -6945 16335 -6825
rect 16455 -6945 16500 -6825
rect 16620 -6945 16665 -6825
rect 16785 -6945 16840 -6825
rect 16960 -6945 17005 -6825
rect 17125 -6945 17170 -6825
rect 17290 -6945 17335 -6825
rect 17455 -6945 17510 -6825
rect 17630 -6945 17675 -6825
rect 17795 -6945 17840 -6825
rect 17960 -6945 18005 -6825
rect 18125 -6945 18180 -6825
rect 18300 -6945 18325 -6825
rect 12795 -6990 18325 -6945
rect 12795 -7110 12820 -6990
rect 12940 -7110 12985 -6990
rect 13105 -7110 13150 -6990
rect 13270 -7110 13315 -6990
rect 13435 -7110 13490 -6990
rect 13610 -7110 13655 -6990
rect 13775 -7110 13820 -6990
rect 13940 -7110 13985 -6990
rect 14105 -7110 14160 -6990
rect 14280 -7110 14325 -6990
rect 14445 -7110 14490 -6990
rect 14610 -7110 14655 -6990
rect 14775 -7110 14830 -6990
rect 14950 -7110 14995 -6990
rect 15115 -7110 15160 -6990
rect 15280 -7110 15325 -6990
rect 15445 -7110 15500 -6990
rect 15620 -7110 15665 -6990
rect 15785 -7110 15830 -6990
rect 15950 -7110 15995 -6990
rect 16115 -7110 16170 -6990
rect 16290 -7110 16335 -6990
rect 16455 -7110 16500 -6990
rect 16620 -7110 16665 -6990
rect 16785 -7110 16840 -6990
rect 16960 -7110 17005 -6990
rect 17125 -7110 17170 -6990
rect 17290 -7110 17335 -6990
rect 17455 -7110 17510 -6990
rect 17630 -7110 17675 -6990
rect 17795 -7110 17840 -6990
rect 17960 -7110 18005 -6990
rect 18125 -7110 18180 -6990
rect 18300 -7110 18325 -6990
rect 12795 -7165 18325 -7110
rect 12795 -7285 12820 -7165
rect 12940 -7285 12985 -7165
rect 13105 -7285 13150 -7165
rect 13270 -7285 13315 -7165
rect 13435 -7285 13490 -7165
rect 13610 -7285 13655 -7165
rect 13775 -7285 13820 -7165
rect 13940 -7285 13985 -7165
rect 14105 -7285 14160 -7165
rect 14280 -7285 14325 -7165
rect 14445 -7285 14490 -7165
rect 14610 -7285 14655 -7165
rect 14775 -7285 14830 -7165
rect 14950 -7285 14995 -7165
rect 15115 -7285 15160 -7165
rect 15280 -7285 15325 -7165
rect 15445 -7285 15500 -7165
rect 15620 -7285 15665 -7165
rect 15785 -7285 15830 -7165
rect 15950 -7285 15995 -7165
rect 16115 -7285 16170 -7165
rect 16290 -7285 16335 -7165
rect 16455 -7285 16500 -7165
rect 16620 -7285 16665 -7165
rect 16785 -7285 16840 -7165
rect 16960 -7285 17005 -7165
rect 17125 -7285 17170 -7165
rect 17290 -7285 17335 -7165
rect 17455 -7285 17510 -7165
rect 17630 -7285 17675 -7165
rect 17795 -7285 17840 -7165
rect 17960 -7285 18005 -7165
rect 18125 -7285 18180 -7165
rect 18300 -7285 18325 -7165
rect 12795 -7330 18325 -7285
rect 12795 -7450 12820 -7330
rect 12940 -7450 12985 -7330
rect 13105 -7450 13150 -7330
rect 13270 -7450 13315 -7330
rect 13435 -7450 13490 -7330
rect 13610 -7450 13655 -7330
rect 13775 -7450 13820 -7330
rect 13940 -7450 13985 -7330
rect 14105 -7450 14160 -7330
rect 14280 -7450 14325 -7330
rect 14445 -7450 14490 -7330
rect 14610 -7450 14655 -7330
rect 14775 -7450 14830 -7330
rect 14950 -7450 14995 -7330
rect 15115 -7450 15160 -7330
rect 15280 -7450 15325 -7330
rect 15445 -7450 15500 -7330
rect 15620 -7450 15665 -7330
rect 15785 -7450 15830 -7330
rect 15950 -7450 15995 -7330
rect 16115 -7450 16170 -7330
rect 16290 -7450 16335 -7330
rect 16455 -7450 16500 -7330
rect 16620 -7450 16665 -7330
rect 16785 -7450 16840 -7330
rect 16960 -7450 17005 -7330
rect 17125 -7450 17170 -7330
rect 17290 -7450 17335 -7330
rect 17455 -7450 17510 -7330
rect 17630 -7450 17675 -7330
rect 17795 -7450 17840 -7330
rect 17960 -7450 18005 -7330
rect 18125 -7450 18180 -7330
rect 18300 -7450 18325 -7330
rect 12795 -7495 18325 -7450
rect 12795 -7615 12820 -7495
rect 12940 -7615 12985 -7495
rect 13105 -7615 13150 -7495
rect 13270 -7615 13315 -7495
rect 13435 -7615 13490 -7495
rect 13610 -7615 13655 -7495
rect 13775 -7615 13820 -7495
rect 13940 -7615 13985 -7495
rect 14105 -7615 14160 -7495
rect 14280 -7615 14325 -7495
rect 14445 -7615 14490 -7495
rect 14610 -7615 14655 -7495
rect 14775 -7615 14830 -7495
rect 14950 -7615 14995 -7495
rect 15115 -7615 15160 -7495
rect 15280 -7615 15325 -7495
rect 15445 -7615 15500 -7495
rect 15620 -7615 15665 -7495
rect 15785 -7615 15830 -7495
rect 15950 -7615 15995 -7495
rect 16115 -7615 16170 -7495
rect 16290 -7615 16335 -7495
rect 16455 -7615 16500 -7495
rect 16620 -7615 16665 -7495
rect 16785 -7615 16840 -7495
rect 16960 -7615 17005 -7495
rect 17125 -7615 17170 -7495
rect 17290 -7615 17335 -7495
rect 17455 -7615 17510 -7495
rect 17630 -7615 17675 -7495
rect 17795 -7615 17840 -7495
rect 17960 -7615 18005 -7495
rect 18125 -7615 18180 -7495
rect 18300 -7615 18325 -7495
rect 12795 -7660 18325 -7615
rect 12795 -7780 12820 -7660
rect 12940 -7780 12985 -7660
rect 13105 -7780 13150 -7660
rect 13270 -7780 13315 -7660
rect 13435 -7780 13490 -7660
rect 13610 -7780 13655 -7660
rect 13775 -7780 13820 -7660
rect 13940 -7780 13985 -7660
rect 14105 -7780 14160 -7660
rect 14280 -7780 14325 -7660
rect 14445 -7780 14490 -7660
rect 14610 -7780 14655 -7660
rect 14775 -7780 14830 -7660
rect 14950 -7780 14995 -7660
rect 15115 -7780 15160 -7660
rect 15280 -7780 15325 -7660
rect 15445 -7780 15500 -7660
rect 15620 -7780 15665 -7660
rect 15785 -7780 15830 -7660
rect 15950 -7780 15995 -7660
rect 16115 -7780 16170 -7660
rect 16290 -7780 16335 -7660
rect 16455 -7780 16500 -7660
rect 16620 -7780 16665 -7660
rect 16785 -7780 16840 -7660
rect 16960 -7780 17005 -7660
rect 17125 -7780 17170 -7660
rect 17290 -7780 17335 -7660
rect 17455 -7780 17510 -7660
rect 17630 -7780 17675 -7660
rect 17795 -7780 17840 -7660
rect 17960 -7780 18005 -7660
rect 18125 -7780 18180 -7660
rect 18300 -7780 18325 -7660
rect 12795 -7835 18325 -7780
rect 12795 -7955 12820 -7835
rect 12940 -7955 12985 -7835
rect 13105 -7955 13150 -7835
rect 13270 -7955 13315 -7835
rect 13435 -7955 13490 -7835
rect 13610 -7955 13655 -7835
rect 13775 -7955 13820 -7835
rect 13940 -7955 13985 -7835
rect 14105 -7955 14160 -7835
rect 14280 -7955 14325 -7835
rect 14445 -7955 14490 -7835
rect 14610 -7955 14655 -7835
rect 14775 -7955 14830 -7835
rect 14950 -7955 14995 -7835
rect 15115 -7955 15160 -7835
rect 15280 -7955 15325 -7835
rect 15445 -7955 15500 -7835
rect 15620 -7955 15665 -7835
rect 15785 -7955 15830 -7835
rect 15950 -7955 15995 -7835
rect 16115 -7955 16170 -7835
rect 16290 -7955 16335 -7835
rect 16455 -7955 16500 -7835
rect 16620 -7955 16665 -7835
rect 16785 -7955 16840 -7835
rect 16960 -7955 17005 -7835
rect 17125 -7955 17170 -7835
rect 17290 -7955 17335 -7835
rect 17455 -7955 17510 -7835
rect 17630 -7955 17675 -7835
rect 17795 -7955 17840 -7835
rect 17960 -7955 18005 -7835
rect 18125 -7955 18180 -7835
rect 18300 -7955 18325 -7835
rect 12795 -8000 18325 -7955
rect 12795 -8120 12820 -8000
rect 12940 -8120 12985 -8000
rect 13105 -8120 13150 -8000
rect 13270 -8120 13315 -8000
rect 13435 -8120 13490 -8000
rect 13610 -8120 13655 -8000
rect 13775 -8120 13820 -8000
rect 13940 -8120 13985 -8000
rect 14105 -8120 14160 -8000
rect 14280 -8120 14325 -8000
rect 14445 -8120 14490 -8000
rect 14610 -8120 14655 -8000
rect 14775 -8120 14830 -8000
rect 14950 -8120 14995 -8000
rect 15115 -8120 15160 -8000
rect 15280 -8120 15325 -8000
rect 15445 -8120 15500 -8000
rect 15620 -8120 15665 -8000
rect 15785 -8120 15830 -8000
rect 15950 -8120 15995 -8000
rect 16115 -8120 16170 -8000
rect 16290 -8120 16335 -8000
rect 16455 -8120 16500 -8000
rect 16620 -8120 16665 -8000
rect 16785 -8120 16840 -8000
rect 16960 -8120 17005 -8000
rect 17125 -8120 17170 -8000
rect 17290 -8120 17335 -8000
rect 17455 -8120 17510 -8000
rect 17630 -8120 17675 -8000
rect 17795 -8120 17840 -8000
rect 17960 -8120 18005 -8000
rect 18125 -8120 18180 -8000
rect 18300 -8120 18325 -8000
rect 12795 -8165 18325 -8120
rect 12795 -8285 12820 -8165
rect 12940 -8285 12985 -8165
rect 13105 -8285 13150 -8165
rect 13270 -8285 13315 -8165
rect 13435 -8285 13490 -8165
rect 13610 -8285 13655 -8165
rect 13775 -8285 13820 -8165
rect 13940 -8285 13985 -8165
rect 14105 -8285 14160 -8165
rect 14280 -8285 14325 -8165
rect 14445 -8285 14490 -8165
rect 14610 -8285 14655 -8165
rect 14775 -8285 14830 -8165
rect 14950 -8285 14995 -8165
rect 15115 -8285 15160 -8165
rect 15280 -8285 15325 -8165
rect 15445 -8285 15500 -8165
rect 15620 -8285 15665 -8165
rect 15785 -8285 15830 -8165
rect 15950 -8285 15995 -8165
rect 16115 -8285 16170 -8165
rect 16290 -8285 16335 -8165
rect 16455 -8285 16500 -8165
rect 16620 -8285 16665 -8165
rect 16785 -8285 16840 -8165
rect 16960 -8285 17005 -8165
rect 17125 -8285 17170 -8165
rect 17290 -8285 17335 -8165
rect 17455 -8285 17510 -8165
rect 17630 -8285 17675 -8165
rect 17795 -8285 17840 -8165
rect 17960 -8285 18005 -8165
rect 18125 -8285 18180 -8165
rect 18300 -8285 18325 -8165
rect 12795 -8330 18325 -8285
rect 12795 -8450 12820 -8330
rect 12940 -8450 12985 -8330
rect 13105 -8450 13150 -8330
rect 13270 -8450 13315 -8330
rect 13435 -8450 13490 -8330
rect 13610 -8450 13655 -8330
rect 13775 -8450 13820 -8330
rect 13940 -8450 13985 -8330
rect 14105 -8450 14160 -8330
rect 14280 -8450 14325 -8330
rect 14445 -8450 14490 -8330
rect 14610 -8450 14655 -8330
rect 14775 -8450 14830 -8330
rect 14950 -8450 14995 -8330
rect 15115 -8450 15160 -8330
rect 15280 -8450 15325 -8330
rect 15445 -8450 15500 -8330
rect 15620 -8450 15665 -8330
rect 15785 -8450 15830 -8330
rect 15950 -8450 15995 -8330
rect 16115 -8450 16170 -8330
rect 16290 -8450 16335 -8330
rect 16455 -8450 16500 -8330
rect 16620 -8450 16665 -8330
rect 16785 -8450 16840 -8330
rect 16960 -8450 17005 -8330
rect 17125 -8450 17170 -8330
rect 17290 -8450 17335 -8330
rect 17455 -8450 17510 -8330
rect 17630 -8450 17675 -8330
rect 17795 -8450 17840 -8330
rect 17960 -8450 18005 -8330
rect 18125 -8450 18180 -8330
rect 18300 -8450 18325 -8330
rect 12795 -8505 18325 -8450
rect 12795 -8625 12820 -8505
rect 12940 -8625 12985 -8505
rect 13105 -8625 13150 -8505
rect 13270 -8625 13315 -8505
rect 13435 -8625 13490 -8505
rect 13610 -8625 13655 -8505
rect 13775 -8625 13820 -8505
rect 13940 -8625 13985 -8505
rect 14105 -8625 14160 -8505
rect 14280 -8625 14325 -8505
rect 14445 -8625 14490 -8505
rect 14610 -8625 14655 -8505
rect 14775 -8625 14830 -8505
rect 14950 -8625 14995 -8505
rect 15115 -8625 15160 -8505
rect 15280 -8625 15325 -8505
rect 15445 -8625 15500 -8505
rect 15620 -8625 15665 -8505
rect 15785 -8625 15830 -8505
rect 15950 -8625 15995 -8505
rect 16115 -8625 16170 -8505
rect 16290 -8625 16335 -8505
rect 16455 -8625 16500 -8505
rect 16620 -8625 16665 -8505
rect 16785 -8625 16840 -8505
rect 16960 -8625 17005 -8505
rect 17125 -8625 17170 -8505
rect 17290 -8625 17335 -8505
rect 17455 -8625 17510 -8505
rect 17630 -8625 17675 -8505
rect 17795 -8625 17840 -8505
rect 17960 -8625 18005 -8505
rect 18125 -8625 18180 -8505
rect 18300 -8625 18325 -8505
rect 12795 -8670 18325 -8625
rect 12795 -8790 12820 -8670
rect 12940 -8790 12985 -8670
rect 13105 -8790 13150 -8670
rect 13270 -8790 13315 -8670
rect 13435 -8790 13490 -8670
rect 13610 -8790 13655 -8670
rect 13775 -8790 13820 -8670
rect 13940 -8790 13985 -8670
rect 14105 -8790 14160 -8670
rect 14280 -8790 14325 -8670
rect 14445 -8790 14490 -8670
rect 14610 -8790 14655 -8670
rect 14775 -8790 14830 -8670
rect 14950 -8790 14995 -8670
rect 15115 -8790 15160 -8670
rect 15280 -8790 15325 -8670
rect 15445 -8790 15500 -8670
rect 15620 -8790 15665 -8670
rect 15785 -8790 15830 -8670
rect 15950 -8790 15995 -8670
rect 16115 -8790 16170 -8670
rect 16290 -8790 16335 -8670
rect 16455 -8790 16500 -8670
rect 16620 -8790 16665 -8670
rect 16785 -8790 16840 -8670
rect 16960 -8790 17005 -8670
rect 17125 -8790 17170 -8670
rect 17290 -8790 17335 -8670
rect 17455 -8790 17510 -8670
rect 17630 -8790 17675 -8670
rect 17795 -8790 17840 -8670
rect 17960 -8790 18005 -8670
rect 18125 -8790 18180 -8670
rect 18300 -8790 18325 -8670
rect 12795 -8835 18325 -8790
rect 12795 -8955 12820 -8835
rect 12940 -8955 12985 -8835
rect 13105 -8955 13150 -8835
rect 13270 -8955 13315 -8835
rect 13435 -8955 13490 -8835
rect 13610 -8955 13655 -8835
rect 13775 -8955 13820 -8835
rect 13940 -8955 13985 -8835
rect 14105 -8955 14160 -8835
rect 14280 -8955 14325 -8835
rect 14445 -8955 14490 -8835
rect 14610 -8955 14655 -8835
rect 14775 -8955 14830 -8835
rect 14950 -8955 14995 -8835
rect 15115 -8955 15160 -8835
rect 15280 -8955 15325 -8835
rect 15445 -8955 15500 -8835
rect 15620 -8955 15665 -8835
rect 15785 -8955 15830 -8835
rect 15950 -8955 15995 -8835
rect 16115 -8955 16170 -8835
rect 16290 -8955 16335 -8835
rect 16455 -8955 16500 -8835
rect 16620 -8955 16665 -8835
rect 16785 -8955 16840 -8835
rect 16960 -8955 17005 -8835
rect 17125 -8955 17170 -8835
rect 17290 -8955 17335 -8835
rect 17455 -8955 17510 -8835
rect 17630 -8955 17675 -8835
rect 17795 -8955 17840 -8835
rect 17960 -8955 18005 -8835
rect 18125 -8955 18180 -8835
rect 18300 -8955 18325 -8835
rect 12795 -9000 18325 -8955
rect 12795 -9120 12820 -9000
rect 12940 -9120 12985 -9000
rect 13105 -9120 13150 -9000
rect 13270 -9120 13315 -9000
rect 13435 -9120 13490 -9000
rect 13610 -9120 13655 -9000
rect 13775 -9120 13820 -9000
rect 13940 -9120 13985 -9000
rect 14105 -9120 14160 -9000
rect 14280 -9120 14325 -9000
rect 14445 -9120 14490 -9000
rect 14610 -9120 14655 -9000
rect 14775 -9120 14830 -9000
rect 14950 -9120 14995 -9000
rect 15115 -9120 15160 -9000
rect 15280 -9120 15325 -9000
rect 15445 -9120 15500 -9000
rect 15620 -9120 15665 -9000
rect 15785 -9120 15830 -9000
rect 15950 -9120 15995 -9000
rect 16115 -9120 16170 -9000
rect 16290 -9120 16335 -9000
rect 16455 -9120 16500 -9000
rect 16620 -9120 16665 -9000
rect 16785 -9120 16840 -9000
rect 16960 -9120 17005 -9000
rect 17125 -9120 17170 -9000
rect 17290 -9120 17335 -9000
rect 17455 -9120 17510 -9000
rect 17630 -9120 17675 -9000
rect 17795 -9120 17840 -9000
rect 17960 -9120 18005 -9000
rect 18125 -9120 18180 -9000
rect 18300 -9120 18325 -9000
rect 12795 -9175 18325 -9120
rect 12795 -9295 12820 -9175
rect 12940 -9295 12985 -9175
rect 13105 -9295 13150 -9175
rect 13270 -9295 13315 -9175
rect 13435 -9295 13490 -9175
rect 13610 -9295 13655 -9175
rect 13775 -9295 13820 -9175
rect 13940 -9295 13985 -9175
rect 14105 -9295 14160 -9175
rect 14280 -9295 14325 -9175
rect 14445 -9295 14490 -9175
rect 14610 -9295 14655 -9175
rect 14775 -9295 14830 -9175
rect 14950 -9295 14995 -9175
rect 15115 -9295 15160 -9175
rect 15280 -9295 15325 -9175
rect 15445 -9295 15500 -9175
rect 15620 -9295 15665 -9175
rect 15785 -9295 15830 -9175
rect 15950 -9295 15995 -9175
rect 16115 -9295 16170 -9175
rect 16290 -9295 16335 -9175
rect 16455 -9295 16500 -9175
rect 16620 -9295 16665 -9175
rect 16785 -9295 16840 -9175
rect 16960 -9295 17005 -9175
rect 17125 -9295 17170 -9175
rect 17290 -9295 17335 -9175
rect 17455 -9295 17510 -9175
rect 17630 -9295 17675 -9175
rect 17795 -9295 17840 -9175
rect 17960 -9295 18005 -9175
rect 18125 -9295 18180 -9175
rect 18300 -9295 18325 -9175
rect 12795 -9340 18325 -9295
rect 12795 -9460 12820 -9340
rect 12940 -9460 12985 -9340
rect 13105 -9460 13150 -9340
rect 13270 -9460 13315 -9340
rect 13435 -9460 13490 -9340
rect 13610 -9460 13655 -9340
rect 13775 -9460 13820 -9340
rect 13940 -9460 13985 -9340
rect 14105 -9460 14160 -9340
rect 14280 -9460 14325 -9340
rect 14445 -9460 14490 -9340
rect 14610 -9460 14655 -9340
rect 14775 -9460 14830 -9340
rect 14950 -9460 14995 -9340
rect 15115 -9460 15160 -9340
rect 15280 -9460 15325 -9340
rect 15445 -9460 15500 -9340
rect 15620 -9460 15665 -9340
rect 15785 -9460 15830 -9340
rect 15950 -9460 15995 -9340
rect 16115 -9460 16170 -9340
rect 16290 -9460 16335 -9340
rect 16455 -9460 16500 -9340
rect 16620 -9460 16665 -9340
rect 16785 -9460 16840 -9340
rect 16960 -9460 17005 -9340
rect 17125 -9460 17170 -9340
rect 17290 -9460 17335 -9340
rect 17455 -9460 17510 -9340
rect 17630 -9460 17675 -9340
rect 17795 -9460 17840 -9340
rect 17960 -9460 18005 -9340
rect 18125 -9460 18180 -9340
rect 18300 -9460 18325 -9340
rect 12795 -9505 18325 -9460
rect 12795 -9625 12820 -9505
rect 12940 -9625 12985 -9505
rect 13105 -9625 13150 -9505
rect 13270 -9625 13315 -9505
rect 13435 -9625 13490 -9505
rect 13610 -9625 13655 -9505
rect 13775 -9625 13820 -9505
rect 13940 -9625 13985 -9505
rect 14105 -9625 14160 -9505
rect 14280 -9625 14325 -9505
rect 14445 -9625 14490 -9505
rect 14610 -9625 14655 -9505
rect 14775 -9625 14830 -9505
rect 14950 -9625 14995 -9505
rect 15115 -9625 15160 -9505
rect 15280 -9625 15325 -9505
rect 15445 -9625 15500 -9505
rect 15620 -9625 15665 -9505
rect 15785 -9625 15830 -9505
rect 15950 -9625 15995 -9505
rect 16115 -9625 16170 -9505
rect 16290 -9625 16335 -9505
rect 16455 -9625 16500 -9505
rect 16620 -9625 16665 -9505
rect 16785 -9625 16840 -9505
rect 16960 -9625 17005 -9505
rect 17125 -9625 17170 -9505
rect 17290 -9625 17335 -9505
rect 17455 -9625 17510 -9505
rect 17630 -9625 17675 -9505
rect 17795 -9625 17840 -9505
rect 17960 -9625 18005 -9505
rect 18125 -9625 18180 -9505
rect 18300 -9625 18325 -9505
rect 12795 -9670 18325 -9625
rect 12795 -9790 12820 -9670
rect 12940 -9790 12985 -9670
rect 13105 -9790 13150 -9670
rect 13270 -9790 13315 -9670
rect 13435 -9790 13490 -9670
rect 13610 -9790 13655 -9670
rect 13775 -9790 13820 -9670
rect 13940 -9790 13985 -9670
rect 14105 -9790 14160 -9670
rect 14280 -9790 14325 -9670
rect 14445 -9790 14490 -9670
rect 14610 -9790 14655 -9670
rect 14775 -9790 14830 -9670
rect 14950 -9790 14995 -9670
rect 15115 -9790 15160 -9670
rect 15280 -9790 15325 -9670
rect 15445 -9790 15500 -9670
rect 15620 -9790 15665 -9670
rect 15785 -9790 15830 -9670
rect 15950 -9790 15995 -9670
rect 16115 -9790 16170 -9670
rect 16290 -9790 16335 -9670
rect 16455 -9790 16500 -9670
rect 16620 -9790 16665 -9670
rect 16785 -9790 16840 -9670
rect 16960 -9790 17005 -9670
rect 17125 -9790 17170 -9670
rect 17290 -9790 17335 -9670
rect 17455 -9790 17510 -9670
rect 17630 -9790 17675 -9670
rect 17795 -9790 17840 -9670
rect 17960 -9790 18005 -9670
rect 18125 -9790 18180 -9670
rect 18300 -9790 18325 -9670
rect 12795 -9815 18325 -9790
rect 18485 -4430 18510 -4345
rect 18630 -4430 18675 -4310
rect 18795 -4430 18840 -4310
rect 18960 -4430 19005 -4310
rect 19125 -4430 19180 -4310
rect 19300 -4430 19345 -4310
rect 19465 -4430 19510 -4310
rect 19630 -4430 19675 -4310
rect 19795 -4430 19850 -4310
rect 19970 -4430 20015 -4310
rect 20135 -4430 20180 -4310
rect 20300 -4430 20345 -4310
rect 20465 -4430 20520 -4310
rect 20640 -4430 20685 -4310
rect 20805 -4430 20850 -4310
rect 20970 -4430 21015 -4310
rect 21135 -4430 21190 -4310
rect 21310 -4430 21355 -4310
rect 21475 -4430 21520 -4310
rect 21640 -4430 21685 -4310
rect 21805 -4430 21860 -4310
rect 21980 -4430 22025 -4310
rect 22145 -4430 22190 -4310
rect 22310 -4430 22355 -4310
rect 22475 -4430 22530 -4310
rect 22650 -4430 22695 -4310
rect 22815 -4430 22860 -4310
rect 22980 -4430 23025 -4310
rect 23145 -4430 23200 -4310
rect 23320 -4430 23365 -4310
rect 23485 -4430 23530 -4310
rect 23650 -4430 23695 -4310
rect 23815 -4430 23870 -4310
rect 23990 -4345 24200 -4310
rect 23990 -4430 24015 -4345
rect 18485 -4485 24015 -4430
rect 18485 -4605 18510 -4485
rect 18630 -4605 18675 -4485
rect 18795 -4605 18840 -4485
rect 18960 -4605 19005 -4485
rect 19125 -4605 19180 -4485
rect 19300 -4605 19345 -4485
rect 19465 -4605 19510 -4485
rect 19630 -4605 19675 -4485
rect 19795 -4605 19850 -4485
rect 19970 -4605 20015 -4485
rect 20135 -4605 20180 -4485
rect 20300 -4605 20345 -4485
rect 20465 -4605 20520 -4485
rect 20640 -4605 20685 -4485
rect 20805 -4605 20850 -4485
rect 20970 -4605 21015 -4485
rect 21135 -4605 21190 -4485
rect 21310 -4605 21355 -4485
rect 21475 -4605 21520 -4485
rect 21640 -4605 21685 -4485
rect 21805 -4605 21860 -4485
rect 21980 -4605 22025 -4485
rect 22145 -4605 22190 -4485
rect 22310 -4605 22355 -4485
rect 22475 -4605 22530 -4485
rect 22650 -4605 22695 -4485
rect 22815 -4605 22860 -4485
rect 22980 -4605 23025 -4485
rect 23145 -4605 23200 -4485
rect 23320 -4605 23365 -4485
rect 23485 -4605 23530 -4485
rect 23650 -4605 23695 -4485
rect 23815 -4605 23870 -4485
rect 23990 -4605 24015 -4485
rect 18485 -4650 24015 -4605
rect 18485 -4770 18510 -4650
rect 18630 -4770 18675 -4650
rect 18795 -4770 18840 -4650
rect 18960 -4770 19005 -4650
rect 19125 -4770 19180 -4650
rect 19300 -4770 19345 -4650
rect 19465 -4770 19510 -4650
rect 19630 -4770 19675 -4650
rect 19795 -4770 19850 -4650
rect 19970 -4770 20015 -4650
rect 20135 -4770 20180 -4650
rect 20300 -4770 20345 -4650
rect 20465 -4770 20520 -4650
rect 20640 -4770 20685 -4650
rect 20805 -4770 20850 -4650
rect 20970 -4770 21015 -4650
rect 21135 -4770 21190 -4650
rect 21310 -4770 21355 -4650
rect 21475 -4770 21520 -4650
rect 21640 -4770 21685 -4650
rect 21805 -4770 21860 -4650
rect 21980 -4770 22025 -4650
rect 22145 -4770 22190 -4650
rect 22310 -4770 22355 -4650
rect 22475 -4770 22530 -4650
rect 22650 -4770 22695 -4650
rect 22815 -4770 22860 -4650
rect 22980 -4770 23025 -4650
rect 23145 -4770 23200 -4650
rect 23320 -4770 23365 -4650
rect 23485 -4770 23530 -4650
rect 23650 -4770 23695 -4650
rect 23815 -4770 23870 -4650
rect 23990 -4770 24015 -4650
rect 18485 -4815 24015 -4770
rect 18485 -4935 18510 -4815
rect 18630 -4935 18675 -4815
rect 18795 -4935 18840 -4815
rect 18960 -4935 19005 -4815
rect 19125 -4935 19180 -4815
rect 19300 -4935 19345 -4815
rect 19465 -4935 19510 -4815
rect 19630 -4935 19675 -4815
rect 19795 -4935 19850 -4815
rect 19970 -4935 20015 -4815
rect 20135 -4935 20180 -4815
rect 20300 -4935 20345 -4815
rect 20465 -4935 20520 -4815
rect 20640 -4935 20685 -4815
rect 20805 -4935 20850 -4815
rect 20970 -4935 21015 -4815
rect 21135 -4935 21190 -4815
rect 21310 -4935 21355 -4815
rect 21475 -4935 21520 -4815
rect 21640 -4935 21685 -4815
rect 21805 -4935 21860 -4815
rect 21980 -4935 22025 -4815
rect 22145 -4935 22190 -4815
rect 22310 -4935 22355 -4815
rect 22475 -4935 22530 -4815
rect 22650 -4935 22695 -4815
rect 22815 -4935 22860 -4815
rect 22980 -4935 23025 -4815
rect 23145 -4935 23200 -4815
rect 23320 -4935 23365 -4815
rect 23485 -4935 23530 -4815
rect 23650 -4935 23695 -4815
rect 23815 -4935 23870 -4815
rect 23990 -4935 24015 -4815
rect 18485 -4980 24015 -4935
rect 18485 -5100 18510 -4980
rect 18630 -5100 18675 -4980
rect 18795 -5100 18840 -4980
rect 18960 -5100 19005 -4980
rect 19125 -5100 19180 -4980
rect 19300 -5100 19345 -4980
rect 19465 -5100 19510 -4980
rect 19630 -5100 19675 -4980
rect 19795 -5100 19850 -4980
rect 19970 -5100 20015 -4980
rect 20135 -5100 20180 -4980
rect 20300 -5100 20345 -4980
rect 20465 -5100 20520 -4980
rect 20640 -5100 20685 -4980
rect 20805 -5100 20850 -4980
rect 20970 -5100 21015 -4980
rect 21135 -5100 21190 -4980
rect 21310 -5100 21355 -4980
rect 21475 -5100 21520 -4980
rect 21640 -5100 21685 -4980
rect 21805 -5100 21860 -4980
rect 21980 -5100 22025 -4980
rect 22145 -5100 22190 -4980
rect 22310 -5100 22355 -4980
rect 22475 -5100 22530 -4980
rect 22650 -5100 22695 -4980
rect 22815 -5100 22860 -4980
rect 22980 -5100 23025 -4980
rect 23145 -5100 23200 -4980
rect 23320 -5100 23365 -4980
rect 23485 -5100 23530 -4980
rect 23650 -5100 23695 -4980
rect 23815 -5100 23870 -4980
rect 23990 -5100 24015 -4980
rect 18485 -5155 24015 -5100
rect 18485 -5275 18510 -5155
rect 18630 -5275 18675 -5155
rect 18795 -5275 18840 -5155
rect 18960 -5275 19005 -5155
rect 19125 -5275 19180 -5155
rect 19300 -5275 19345 -5155
rect 19465 -5275 19510 -5155
rect 19630 -5275 19675 -5155
rect 19795 -5275 19850 -5155
rect 19970 -5275 20015 -5155
rect 20135 -5275 20180 -5155
rect 20300 -5275 20345 -5155
rect 20465 -5275 20520 -5155
rect 20640 -5275 20685 -5155
rect 20805 -5275 20850 -5155
rect 20970 -5275 21015 -5155
rect 21135 -5275 21190 -5155
rect 21310 -5275 21355 -5155
rect 21475 -5275 21520 -5155
rect 21640 -5275 21685 -5155
rect 21805 -5275 21860 -5155
rect 21980 -5275 22025 -5155
rect 22145 -5275 22190 -5155
rect 22310 -5275 22355 -5155
rect 22475 -5275 22530 -5155
rect 22650 -5275 22695 -5155
rect 22815 -5275 22860 -5155
rect 22980 -5275 23025 -5155
rect 23145 -5275 23200 -5155
rect 23320 -5275 23365 -5155
rect 23485 -5275 23530 -5155
rect 23650 -5275 23695 -5155
rect 23815 -5275 23870 -5155
rect 23990 -5275 24015 -5155
rect 18485 -5320 24015 -5275
rect 18485 -5440 18510 -5320
rect 18630 -5440 18675 -5320
rect 18795 -5440 18840 -5320
rect 18960 -5440 19005 -5320
rect 19125 -5440 19180 -5320
rect 19300 -5440 19345 -5320
rect 19465 -5440 19510 -5320
rect 19630 -5440 19675 -5320
rect 19795 -5440 19850 -5320
rect 19970 -5440 20015 -5320
rect 20135 -5440 20180 -5320
rect 20300 -5440 20345 -5320
rect 20465 -5440 20520 -5320
rect 20640 -5440 20685 -5320
rect 20805 -5440 20850 -5320
rect 20970 -5440 21015 -5320
rect 21135 -5440 21190 -5320
rect 21310 -5440 21355 -5320
rect 21475 -5440 21520 -5320
rect 21640 -5440 21685 -5320
rect 21805 -5440 21860 -5320
rect 21980 -5440 22025 -5320
rect 22145 -5440 22190 -5320
rect 22310 -5440 22355 -5320
rect 22475 -5440 22530 -5320
rect 22650 -5440 22695 -5320
rect 22815 -5440 22860 -5320
rect 22980 -5440 23025 -5320
rect 23145 -5440 23200 -5320
rect 23320 -5440 23365 -5320
rect 23485 -5440 23530 -5320
rect 23650 -5440 23695 -5320
rect 23815 -5440 23870 -5320
rect 23990 -5440 24015 -5320
rect 18485 -5485 24015 -5440
rect 18485 -5605 18510 -5485
rect 18630 -5605 18675 -5485
rect 18795 -5605 18840 -5485
rect 18960 -5605 19005 -5485
rect 19125 -5605 19180 -5485
rect 19300 -5605 19345 -5485
rect 19465 -5605 19510 -5485
rect 19630 -5605 19675 -5485
rect 19795 -5605 19850 -5485
rect 19970 -5605 20015 -5485
rect 20135 -5605 20180 -5485
rect 20300 -5605 20345 -5485
rect 20465 -5605 20520 -5485
rect 20640 -5605 20685 -5485
rect 20805 -5605 20850 -5485
rect 20970 -5605 21015 -5485
rect 21135 -5605 21190 -5485
rect 21310 -5605 21355 -5485
rect 21475 -5605 21520 -5485
rect 21640 -5605 21685 -5485
rect 21805 -5605 21860 -5485
rect 21980 -5605 22025 -5485
rect 22145 -5605 22190 -5485
rect 22310 -5605 22355 -5485
rect 22475 -5605 22530 -5485
rect 22650 -5605 22695 -5485
rect 22815 -5605 22860 -5485
rect 22980 -5605 23025 -5485
rect 23145 -5605 23200 -5485
rect 23320 -5605 23365 -5485
rect 23485 -5605 23530 -5485
rect 23650 -5605 23695 -5485
rect 23815 -5605 23870 -5485
rect 23990 -5605 24015 -5485
rect 18485 -5650 24015 -5605
rect 18485 -5770 18510 -5650
rect 18630 -5770 18675 -5650
rect 18795 -5770 18840 -5650
rect 18960 -5770 19005 -5650
rect 19125 -5770 19180 -5650
rect 19300 -5770 19345 -5650
rect 19465 -5770 19510 -5650
rect 19630 -5770 19675 -5650
rect 19795 -5770 19850 -5650
rect 19970 -5770 20015 -5650
rect 20135 -5770 20180 -5650
rect 20300 -5770 20345 -5650
rect 20465 -5770 20520 -5650
rect 20640 -5770 20685 -5650
rect 20805 -5770 20850 -5650
rect 20970 -5770 21015 -5650
rect 21135 -5770 21190 -5650
rect 21310 -5770 21355 -5650
rect 21475 -5770 21520 -5650
rect 21640 -5770 21685 -5650
rect 21805 -5770 21860 -5650
rect 21980 -5770 22025 -5650
rect 22145 -5770 22190 -5650
rect 22310 -5770 22355 -5650
rect 22475 -5770 22530 -5650
rect 22650 -5770 22695 -5650
rect 22815 -5770 22860 -5650
rect 22980 -5770 23025 -5650
rect 23145 -5770 23200 -5650
rect 23320 -5770 23365 -5650
rect 23485 -5770 23530 -5650
rect 23650 -5770 23695 -5650
rect 23815 -5770 23870 -5650
rect 23990 -5770 24015 -5650
rect 18485 -5825 24015 -5770
rect 18485 -5945 18510 -5825
rect 18630 -5945 18675 -5825
rect 18795 -5945 18840 -5825
rect 18960 -5945 19005 -5825
rect 19125 -5945 19180 -5825
rect 19300 -5945 19345 -5825
rect 19465 -5945 19510 -5825
rect 19630 -5945 19675 -5825
rect 19795 -5945 19850 -5825
rect 19970 -5945 20015 -5825
rect 20135 -5945 20180 -5825
rect 20300 -5945 20345 -5825
rect 20465 -5945 20520 -5825
rect 20640 -5945 20685 -5825
rect 20805 -5945 20850 -5825
rect 20970 -5945 21015 -5825
rect 21135 -5945 21190 -5825
rect 21310 -5945 21355 -5825
rect 21475 -5945 21520 -5825
rect 21640 -5945 21685 -5825
rect 21805 -5945 21860 -5825
rect 21980 -5945 22025 -5825
rect 22145 -5945 22190 -5825
rect 22310 -5945 22355 -5825
rect 22475 -5945 22530 -5825
rect 22650 -5945 22695 -5825
rect 22815 -5945 22860 -5825
rect 22980 -5945 23025 -5825
rect 23145 -5945 23200 -5825
rect 23320 -5945 23365 -5825
rect 23485 -5945 23530 -5825
rect 23650 -5945 23695 -5825
rect 23815 -5945 23870 -5825
rect 23990 -5945 24015 -5825
rect 18485 -5990 24015 -5945
rect 18485 -6110 18510 -5990
rect 18630 -6110 18675 -5990
rect 18795 -6110 18840 -5990
rect 18960 -6110 19005 -5990
rect 19125 -6110 19180 -5990
rect 19300 -6110 19345 -5990
rect 19465 -6110 19510 -5990
rect 19630 -6110 19675 -5990
rect 19795 -6110 19850 -5990
rect 19970 -6110 20015 -5990
rect 20135 -6110 20180 -5990
rect 20300 -6110 20345 -5990
rect 20465 -6110 20520 -5990
rect 20640 -6110 20685 -5990
rect 20805 -6110 20850 -5990
rect 20970 -6110 21015 -5990
rect 21135 -6110 21190 -5990
rect 21310 -6110 21355 -5990
rect 21475 -6110 21520 -5990
rect 21640 -6110 21685 -5990
rect 21805 -6110 21860 -5990
rect 21980 -6110 22025 -5990
rect 22145 -6110 22190 -5990
rect 22310 -6110 22355 -5990
rect 22475 -6110 22530 -5990
rect 22650 -6110 22695 -5990
rect 22815 -6110 22860 -5990
rect 22980 -6110 23025 -5990
rect 23145 -6110 23200 -5990
rect 23320 -6110 23365 -5990
rect 23485 -6110 23530 -5990
rect 23650 -6110 23695 -5990
rect 23815 -6110 23870 -5990
rect 23990 -6110 24015 -5990
rect 18485 -6155 24015 -6110
rect 18485 -6275 18510 -6155
rect 18630 -6275 18675 -6155
rect 18795 -6275 18840 -6155
rect 18960 -6275 19005 -6155
rect 19125 -6275 19180 -6155
rect 19300 -6275 19345 -6155
rect 19465 -6275 19510 -6155
rect 19630 -6275 19675 -6155
rect 19795 -6275 19850 -6155
rect 19970 -6275 20015 -6155
rect 20135 -6275 20180 -6155
rect 20300 -6275 20345 -6155
rect 20465 -6275 20520 -6155
rect 20640 -6275 20685 -6155
rect 20805 -6275 20850 -6155
rect 20970 -6275 21015 -6155
rect 21135 -6275 21190 -6155
rect 21310 -6275 21355 -6155
rect 21475 -6275 21520 -6155
rect 21640 -6275 21685 -6155
rect 21805 -6275 21860 -6155
rect 21980 -6275 22025 -6155
rect 22145 -6275 22190 -6155
rect 22310 -6275 22355 -6155
rect 22475 -6275 22530 -6155
rect 22650 -6275 22695 -6155
rect 22815 -6275 22860 -6155
rect 22980 -6275 23025 -6155
rect 23145 -6275 23200 -6155
rect 23320 -6275 23365 -6155
rect 23485 -6275 23530 -6155
rect 23650 -6275 23695 -6155
rect 23815 -6275 23870 -6155
rect 23990 -6275 24015 -6155
rect 18485 -6320 24015 -6275
rect 18485 -6440 18510 -6320
rect 18630 -6440 18675 -6320
rect 18795 -6440 18840 -6320
rect 18960 -6440 19005 -6320
rect 19125 -6440 19180 -6320
rect 19300 -6440 19345 -6320
rect 19465 -6440 19510 -6320
rect 19630 -6440 19675 -6320
rect 19795 -6440 19850 -6320
rect 19970 -6440 20015 -6320
rect 20135 -6440 20180 -6320
rect 20300 -6440 20345 -6320
rect 20465 -6440 20520 -6320
rect 20640 -6440 20685 -6320
rect 20805 -6440 20850 -6320
rect 20970 -6440 21015 -6320
rect 21135 -6440 21190 -6320
rect 21310 -6440 21355 -6320
rect 21475 -6440 21520 -6320
rect 21640 -6440 21685 -6320
rect 21805 -6440 21860 -6320
rect 21980 -6440 22025 -6320
rect 22145 -6440 22190 -6320
rect 22310 -6440 22355 -6320
rect 22475 -6440 22530 -6320
rect 22650 -6440 22695 -6320
rect 22815 -6440 22860 -6320
rect 22980 -6440 23025 -6320
rect 23145 -6440 23200 -6320
rect 23320 -6440 23365 -6320
rect 23485 -6440 23530 -6320
rect 23650 -6440 23695 -6320
rect 23815 -6440 23870 -6320
rect 23990 -6440 24015 -6320
rect 18485 -6495 24015 -6440
rect 18485 -6615 18510 -6495
rect 18630 -6615 18675 -6495
rect 18795 -6615 18840 -6495
rect 18960 -6615 19005 -6495
rect 19125 -6615 19180 -6495
rect 19300 -6615 19345 -6495
rect 19465 -6615 19510 -6495
rect 19630 -6615 19675 -6495
rect 19795 -6615 19850 -6495
rect 19970 -6615 20015 -6495
rect 20135 -6615 20180 -6495
rect 20300 -6615 20345 -6495
rect 20465 -6615 20520 -6495
rect 20640 -6615 20685 -6495
rect 20805 -6615 20850 -6495
rect 20970 -6615 21015 -6495
rect 21135 -6615 21190 -6495
rect 21310 -6615 21355 -6495
rect 21475 -6615 21520 -6495
rect 21640 -6615 21685 -6495
rect 21805 -6615 21860 -6495
rect 21980 -6615 22025 -6495
rect 22145 -6615 22190 -6495
rect 22310 -6615 22355 -6495
rect 22475 -6615 22530 -6495
rect 22650 -6615 22695 -6495
rect 22815 -6615 22860 -6495
rect 22980 -6615 23025 -6495
rect 23145 -6615 23200 -6495
rect 23320 -6615 23365 -6495
rect 23485 -6615 23530 -6495
rect 23650 -6615 23695 -6495
rect 23815 -6615 23870 -6495
rect 23990 -6615 24015 -6495
rect 18485 -6660 24015 -6615
rect 18485 -6780 18510 -6660
rect 18630 -6780 18675 -6660
rect 18795 -6780 18840 -6660
rect 18960 -6780 19005 -6660
rect 19125 -6780 19180 -6660
rect 19300 -6780 19345 -6660
rect 19465 -6780 19510 -6660
rect 19630 -6780 19675 -6660
rect 19795 -6780 19850 -6660
rect 19970 -6780 20015 -6660
rect 20135 -6780 20180 -6660
rect 20300 -6780 20345 -6660
rect 20465 -6780 20520 -6660
rect 20640 -6780 20685 -6660
rect 20805 -6780 20850 -6660
rect 20970 -6780 21015 -6660
rect 21135 -6780 21190 -6660
rect 21310 -6780 21355 -6660
rect 21475 -6780 21520 -6660
rect 21640 -6780 21685 -6660
rect 21805 -6780 21860 -6660
rect 21980 -6780 22025 -6660
rect 22145 -6780 22190 -6660
rect 22310 -6780 22355 -6660
rect 22475 -6780 22530 -6660
rect 22650 -6780 22695 -6660
rect 22815 -6780 22860 -6660
rect 22980 -6780 23025 -6660
rect 23145 -6780 23200 -6660
rect 23320 -6780 23365 -6660
rect 23485 -6780 23530 -6660
rect 23650 -6780 23695 -6660
rect 23815 -6780 23870 -6660
rect 23990 -6780 24015 -6660
rect 18485 -6825 24015 -6780
rect 18485 -6945 18510 -6825
rect 18630 -6945 18675 -6825
rect 18795 -6945 18840 -6825
rect 18960 -6945 19005 -6825
rect 19125 -6945 19180 -6825
rect 19300 -6945 19345 -6825
rect 19465 -6945 19510 -6825
rect 19630 -6945 19675 -6825
rect 19795 -6945 19850 -6825
rect 19970 -6945 20015 -6825
rect 20135 -6945 20180 -6825
rect 20300 -6945 20345 -6825
rect 20465 -6945 20520 -6825
rect 20640 -6945 20685 -6825
rect 20805 -6945 20850 -6825
rect 20970 -6945 21015 -6825
rect 21135 -6945 21190 -6825
rect 21310 -6945 21355 -6825
rect 21475 -6945 21520 -6825
rect 21640 -6945 21685 -6825
rect 21805 -6945 21860 -6825
rect 21980 -6945 22025 -6825
rect 22145 -6945 22190 -6825
rect 22310 -6945 22355 -6825
rect 22475 -6945 22530 -6825
rect 22650 -6945 22695 -6825
rect 22815 -6945 22860 -6825
rect 22980 -6945 23025 -6825
rect 23145 -6945 23200 -6825
rect 23320 -6945 23365 -6825
rect 23485 -6945 23530 -6825
rect 23650 -6945 23695 -6825
rect 23815 -6945 23870 -6825
rect 23990 -6945 24015 -6825
rect 18485 -6990 24015 -6945
rect 18485 -7110 18510 -6990
rect 18630 -7110 18675 -6990
rect 18795 -7110 18840 -6990
rect 18960 -7110 19005 -6990
rect 19125 -7110 19180 -6990
rect 19300 -7110 19345 -6990
rect 19465 -7110 19510 -6990
rect 19630 -7110 19675 -6990
rect 19795 -7110 19850 -6990
rect 19970 -7110 20015 -6990
rect 20135 -7110 20180 -6990
rect 20300 -7110 20345 -6990
rect 20465 -7110 20520 -6990
rect 20640 -7110 20685 -6990
rect 20805 -7110 20850 -6990
rect 20970 -7110 21015 -6990
rect 21135 -7110 21190 -6990
rect 21310 -7110 21355 -6990
rect 21475 -7110 21520 -6990
rect 21640 -7110 21685 -6990
rect 21805 -7110 21860 -6990
rect 21980 -7110 22025 -6990
rect 22145 -7110 22190 -6990
rect 22310 -7110 22355 -6990
rect 22475 -7110 22530 -6990
rect 22650 -7110 22695 -6990
rect 22815 -7110 22860 -6990
rect 22980 -7110 23025 -6990
rect 23145 -7110 23200 -6990
rect 23320 -7110 23365 -6990
rect 23485 -7110 23530 -6990
rect 23650 -7110 23695 -6990
rect 23815 -7110 23870 -6990
rect 23990 -7110 24015 -6990
rect 18485 -7165 24015 -7110
rect 18485 -7285 18510 -7165
rect 18630 -7285 18675 -7165
rect 18795 -7285 18840 -7165
rect 18960 -7285 19005 -7165
rect 19125 -7285 19180 -7165
rect 19300 -7285 19345 -7165
rect 19465 -7285 19510 -7165
rect 19630 -7285 19675 -7165
rect 19795 -7285 19850 -7165
rect 19970 -7285 20015 -7165
rect 20135 -7285 20180 -7165
rect 20300 -7285 20345 -7165
rect 20465 -7285 20520 -7165
rect 20640 -7285 20685 -7165
rect 20805 -7285 20850 -7165
rect 20970 -7285 21015 -7165
rect 21135 -7285 21190 -7165
rect 21310 -7285 21355 -7165
rect 21475 -7285 21520 -7165
rect 21640 -7285 21685 -7165
rect 21805 -7285 21860 -7165
rect 21980 -7285 22025 -7165
rect 22145 -7285 22190 -7165
rect 22310 -7285 22355 -7165
rect 22475 -7285 22530 -7165
rect 22650 -7285 22695 -7165
rect 22815 -7285 22860 -7165
rect 22980 -7285 23025 -7165
rect 23145 -7285 23200 -7165
rect 23320 -7285 23365 -7165
rect 23485 -7285 23530 -7165
rect 23650 -7285 23695 -7165
rect 23815 -7285 23870 -7165
rect 23990 -7285 24015 -7165
rect 18485 -7330 24015 -7285
rect 18485 -7450 18510 -7330
rect 18630 -7450 18675 -7330
rect 18795 -7450 18840 -7330
rect 18960 -7450 19005 -7330
rect 19125 -7450 19180 -7330
rect 19300 -7450 19345 -7330
rect 19465 -7450 19510 -7330
rect 19630 -7450 19675 -7330
rect 19795 -7450 19850 -7330
rect 19970 -7450 20015 -7330
rect 20135 -7450 20180 -7330
rect 20300 -7450 20345 -7330
rect 20465 -7450 20520 -7330
rect 20640 -7450 20685 -7330
rect 20805 -7450 20850 -7330
rect 20970 -7450 21015 -7330
rect 21135 -7450 21190 -7330
rect 21310 -7450 21355 -7330
rect 21475 -7450 21520 -7330
rect 21640 -7450 21685 -7330
rect 21805 -7450 21860 -7330
rect 21980 -7450 22025 -7330
rect 22145 -7450 22190 -7330
rect 22310 -7450 22355 -7330
rect 22475 -7450 22530 -7330
rect 22650 -7450 22695 -7330
rect 22815 -7450 22860 -7330
rect 22980 -7450 23025 -7330
rect 23145 -7450 23200 -7330
rect 23320 -7450 23365 -7330
rect 23485 -7450 23530 -7330
rect 23650 -7450 23695 -7330
rect 23815 -7450 23870 -7330
rect 23990 -7450 24015 -7330
rect 18485 -7495 24015 -7450
rect 18485 -7615 18510 -7495
rect 18630 -7615 18675 -7495
rect 18795 -7615 18840 -7495
rect 18960 -7615 19005 -7495
rect 19125 -7615 19180 -7495
rect 19300 -7615 19345 -7495
rect 19465 -7615 19510 -7495
rect 19630 -7615 19675 -7495
rect 19795 -7615 19850 -7495
rect 19970 -7615 20015 -7495
rect 20135 -7615 20180 -7495
rect 20300 -7615 20345 -7495
rect 20465 -7615 20520 -7495
rect 20640 -7615 20685 -7495
rect 20805 -7615 20850 -7495
rect 20970 -7615 21015 -7495
rect 21135 -7615 21190 -7495
rect 21310 -7615 21355 -7495
rect 21475 -7615 21520 -7495
rect 21640 -7615 21685 -7495
rect 21805 -7615 21860 -7495
rect 21980 -7615 22025 -7495
rect 22145 -7615 22190 -7495
rect 22310 -7615 22355 -7495
rect 22475 -7615 22530 -7495
rect 22650 -7615 22695 -7495
rect 22815 -7615 22860 -7495
rect 22980 -7615 23025 -7495
rect 23145 -7615 23200 -7495
rect 23320 -7615 23365 -7495
rect 23485 -7615 23530 -7495
rect 23650 -7615 23695 -7495
rect 23815 -7615 23870 -7495
rect 23990 -7615 24015 -7495
rect 18485 -7660 24015 -7615
rect 18485 -7780 18510 -7660
rect 18630 -7780 18675 -7660
rect 18795 -7780 18840 -7660
rect 18960 -7780 19005 -7660
rect 19125 -7780 19180 -7660
rect 19300 -7780 19345 -7660
rect 19465 -7780 19510 -7660
rect 19630 -7780 19675 -7660
rect 19795 -7780 19850 -7660
rect 19970 -7780 20015 -7660
rect 20135 -7780 20180 -7660
rect 20300 -7780 20345 -7660
rect 20465 -7780 20520 -7660
rect 20640 -7780 20685 -7660
rect 20805 -7780 20850 -7660
rect 20970 -7780 21015 -7660
rect 21135 -7780 21190 -7660
rect 21310 -7780 21355 -7660
rect 21475 -7780 21520 -7660
rect 21640 -7780 21685 -7660
rect 21805 -7780 21860 -7660
rect 21980 -7780 22025 -7660
rect 22145 -7780 22190 -7660
rect 22310 -7780 22355 -7660
rect 22475 -7780 22530 -7660
rect 22650 -7780 22695 -7660
rect 22815 -7780 22860 -7660
rect 22980 -7780 23025 -7660
rect 23145 -7780 23200 -7660
rect 23320 -7780 23365 -7660
rect 23485 -7780 23530 -7660
rect 23650 -7780 23695 -7660
rect 23815 -7780 23870 -7660
rect 23990 -7780 24015 -7660
rect 18485 -7835 24015 -7780
rect 18485 -7955 18510 -7835
rect 18630 -7955 18675 -7835
rect 18795 -7955 18840 -7835
rect 18960 -7955 19005 -7835
rect 19125 -7955 19180 -7835
rect 19300 -7955 19345 -7835
rect 19465 -7955 19510 -7835
rect 19630 -7955 19675 -7835
rect 19795 -7955 19850 -7835
rect 19970 -7955 20015 -7835
rect 20135 -7955 20180 -7835
rect 20300 -7955 20345 -7835
rect 20465 -7955 20520 -7835
rect 20640 -7955 20685 -7835
rect 20805 -7955 20850 -7835
rect 20970 -7955 21015 -7835
rect 21135 -7955 21190 -7835
rect 21310 -7955 21355 -7835
rect 21475 -7955 21520 -7835
rect 21640 -7955 21685 -7835
rect 21805 -7955 21860 -7835
rect 21980 -7955 22025 -7835
rect 22145 -7955 22190 -7835
rect 22310 -7955 22355 -7835
rect 22475 -7955 22530 -7835
rect 22650 -7955 22695 -7835
rect 22815 -7955 22860 -7835
rect 22980 -7955 23025 -7835
rect 23145 -7955 23200 -7835
rect 23320 -7955 23365 -7835
rect 23485 -7955 23530 -7835
rect 23650 -7955 23695 -7835
rect 23815 -7955 23870 -7835
rect 23990 -7955 24015 -7835
rect 18485 -8000 24015 -7955
rect 18485 -8120 18510 -8000
rect 18630 -8120 18675 -8000
rect 18795 -8120 18840 -8000
rect 18960 -8120 19005 -8000
rect 19125 -8120 19180 -8000
rect 19300 -8120 19345 -8000
rect 19465 -8120 19510 -8000
rect 19630 -8120 19675 -8000
rect 19795 -8120 19850 -8000
rect 19970 -8120 20015 -8000
rect 20135 -8120 20180 -8000
rect 20300 -8120 20345 -8000
rect 20465 -8120 20520 -8000
rect 20640 -8120 20685 -8000
rect 20805 -8120 20850 -8000
rect 20970 -8120 21015 -8000
rect 21135 -8120 21190 -8000
rect 21310 -8120 21355 -8000
rect 21475 -8120 21520 -8000
rect 21640 -8120 21685 -8000
rect 21805 -8120 21860 -8000
rect 21980 -8120 22025 -8000
rect 22145 -8120 22190 -8000
rect 22310 -8120 22355 -8000
rect 22475 -8120 22530 -8000
rect 22650 -8120 22695 -8000
rect 22815 -8120 22860 -8000
rect 22980 -8120 23025 -8000
rect 23145 -8120 23200 -8000
rect 23320 -8120 23365 -8000
rect 23485 -8120 23530 -8000
rect 23650 -8120 23695 -8000
rect 23815 -8120 23870 -8000
rect 23990 -8120 24015 -8000
rect 18485 -8165 24015 -8120
rect 18485 -8285 18510 -8165
rect 18630 -8285 18675 -8165
rect 18795 -8285 18840 -8165
rect 18960 -8285 19005 -8165
rect 19125 -8285 19180 -8165
rect 19300 -8285 19345 -8165
rect 19465 -8285 19510 -8165
rect 19630 -8285 19675 -8165
rect 19795 -8285 19850 -8165
rect 19970 -8285 20015 -8165
rect 20135 -8285 20180 -8165
rect 20300 -8285 20345 -8165
rect 20465 -8285 20520 -8165
rect 20640 -8285 20685 -8165
rect 20805 -8285 20850 -8165
rect 20970 -8285 21015 -8165
rect 21135 -8285 21190 -8165
rect 21310 -8285 21355 -8165
rect 21475 -8285 21520 -8165
rect 21640 -8285 21685 -8165
rect 21805 -8285 21860 -8165
rect 21980 -8285 22025 -8165
rect 22145 -8285 22190 -8165
rect 22310 -8285 22355 -8165
rect 22475 -8285 22530 -8165
rect 22650 -8285 22695 -8165
rect 22815 -8285 22860 -8165
rect 22980 -8285 23025 -8165
rect 23145 -8285 23200 -8165
rect 23320 -8285 23365 -8165
rect 23485 -8285 23530 -8165
rect 23650 -8285 23695 -8165
rect 23815 -8285 23870 -8165
rect 23990 -8285 24015 -8165
rect 18485 -8330 24015 -8285
rect 18485 -8450 18510 -8330
rect 18630 -8450 18675 -8330
rect 18795 -8450 18840 -8330
rect 18960 -8450 19005 -8330
rect 19125 -8450 19180 -8330
rect 19300 -8450 19345 -8330
rect 19465 -8450 19510 -8330
rect 19630 -8450 19675 -8330
rect 19795 -8450 19850 -8330
rect 19970 -8450 20015 -8330
rect 20135 -8450 20180 -8330
rect 20300 -8450 20345 -8330
rect 20465 -8450 20520 -8330
rect 20640 -8450 20685 -8330
rect 20805 -8450 20850 -8330
rect 20970 -8450 21015 -8330
rect 21135 -8450 21190 -8330
rect 21310 -8450 21355 -8330
rect 21475 -8450 21520 -8330
rect 21640 -8450 21685 -8330
rect 21805 -8450 21860 -8330
rect 21980 -8450 22025 -8330
rect 22145 -8450 22190 -8330
rect 22310 -8450 22355 -8330
rect 22475 -8450 22530 -8330
rect 22650 -8450 22695 -8330
rect 22815 -8450 22860 -8330
rect 22980 -8450 23025 -8330
rect 23145 -8450 23200 -8330
rect 23320 -8450 23365 -8330
rect 23485 -8450 23530 -8330
rect 23650 -8450 23695 -8330
rect 23815 -8450 23870 -8330
rect 23990 -8450 24015 -8330
rect 18485 -8505 24015 -8450
rect 18485 -8625 18510 -8505
rect 18630 -8625 18675 -8505
rect 18795 -8625 18840 -8505
rect 18960 -8625 19005 -8505
rect 19125 -8625 19180 -8505
rect 19300 -8625 19345 -8505
rect 19465 -8625 19510 -8505
rect 19630 -8625 19675 -8505
rect 19795 -8625 19850 -8505
rect 19970 -8625 20015 -8505
rect 20135 -8625 20180 -8505
rect 20300 -8625 20345 -8505
rect 20465 -8625 20520 -8505
rect 20640 -8625 20685 -8505
rect 20805 -8625 20850 -8505
rect 20970 -8625 21015 -8505
rect 21135 -8625 21190 -8505
rect 21310 -8625 21355 -8505
rect 21475 -8625 21520 -8505
rect 21640 -8625 21685 -8505
rect 21805 -8625 21860 -8505
rect 21980 -8625 22025 -8505
rect 22145 -8625 22190 -8505
rect 22310 -8625 22355 -8505
rect 22475 -8625 22530 -8505
rect 22650 -8625 22695 -8505
rect 22815 -8625 22860 -8505
rect 22980 -8625 23025 -8505
rect 23145 -8625 23200 -8505
rect 23320 -8625 23365 -8505
rect 23485 -8625 23530 -8505
rect 23650 -8625 23695 -8505
rect 23815 -8625 23870 -8505
rect 23990 -8625 24015 -8505
rect 18485 -8670 24015 -8625
rect 18485 -8790 18510 -8670
rect 18630 -8790 18675 -8670
rect 18795 -8790 18840 -8670
rect 18960 -8790 19005 -8670
rect 19125 -8790 19180 -8670
rect 19300 -8790 19345 -8670
rect 19465 -8790 19510 -8670
rect 19630 -8790 19675 -8670
rect 19795 -8790 19850 -8670
rect 19970 -8790 20015 -8670
rect 20135 -8790 20180 -8670
rect 20300 -8790 20345 -8670
rect 20465 -8790 20520 -8670
rect 20640 -8790 20685 -8670
rect 20805 -8790 20850 -8670
rect 20970 -8790 21015 -8670
rect 21135 -8790 21190 -8670
rect 21310 -8790 21355 -8670
rect 21475 -8790 21520 -8670
rect 21640 -8790 21685 -8670
rect 21805 -8790 21860 -8670
rect 21980 -8790 22025 -8670
rect 22145 -8790 22190 -8670
rect 22310 -8790 22355 -8670
rect 22475 -8790 22530 -8670
rect 22650 -8790 22695 -8670
rect 22815 -8790 22860 -8670
rect 22980 -8790 23025 -8670
rect 23145 -8790 23200 -8670
rect 23320 -8790 23365 -8670
rect 23485 -8790 23530 -8670
rect 23650 -8790 23695 -8670
rect 23815 -8790 23870 -8670
rect 23990 -8790 24015 -8670
rect 18485 -8835 24015 -8790
rect 18485 -8955 18510 -8835
rect 18630 -8955 18675 -8835
rect 18795 -8955 18840 -8835
rect 18960 -8955 19005 -8835
rect 19125 -8955 19180 -8835
rect 19300 -8955 19345 -8835
rect 19465 -8955 19510 -8835
rect 19630 -8955 19675 -8835
rect 19795 -8955 19850 -8835
rect 19970 -8955 20015 -8835
rect 20135 -8955 20180 -8835
rect 20300 -8955 20345 -8835
rect 20465 -8955 20520 -8835
rect 20640 -8955 20685 -8835
rect 20805 -8955 20850 -8835
rect 20970 -8955 21015 -8835
rect 21135 -8955 21190 -8835
rect 21310 -8955 21355 -8835
rect 21475 -8955 21520 -8835
rect 21640 -8955 21685 -8835
rect 21805 -8955 21860 -8835
rect 21980 -8955 22025 -8835
rect 22145 -8955 22190 -8835
rect 22310 -8955 22355 -8835
rect 22475 -8955 22530 -8835
rect 22650 -8955 22695 -8835
rect 22815 -8955 22860 -8835
rect 22980 -8955 23025 -8835
rect 23145 -8955 23200 -8835
rect 23320 -8955 23365 -8835
rect 23485 -8955 23530 -8835
rect 23650 -8955 23695 -8835
rect 23815 -8955 23870 -8835
rect 23990 -8955 24015 -8835
rect 18485 -9000 24015 -8955
rect 18485 -9120 18510 -9000
rect 18630 -9120 18675 -9000
rect 18795 -9120 18840 -9000
rect 18960 -9120 19005 -9000
rect 19125 -9120 19180 -9000
rect 19300 -9120 19345 -9000
rect 19465 -9120 19510 -9000
rect 19630 -9120 19675 -9000
rect 19795 -9120 19850 -9000
rect 19970 -9120 20015 -9000
rect 20135 -9120 20180 -9000
rect 20300 -9120 20345 -9000
rect 20465 -9120 20520 -9000
rect 20640 -9120 20685 -9000
rect 20805 -9120 20850 -9000
rect 20970 -9120 21015 -9000
rect 21135 -9120 21190 -9000
rect 21310 -9120 21355 -9000
rect 21475 -9120 21520 -9000
rect 21640 -9120 21685 -9000
rect 21805 -9120 21860 -9000
rect 21980 -9120 22025 -9000
rect 22145 -9120 22190 -9000
rect 22310 -9120 22355 -9000
rect 22475 -9120 22530 -9000
rect 22650 -9120 22695 -9000
rect 22815 -9120 22860 -9000
rect 22980 -9120 23025 -9000
rect 23145 -9120 23200 -9000
rect 23320 -9120 23365 -9000
rect 23485 -9120 23530 -9000
rect 23650 -9120 23695 -9000
rect 23815 -9120 23870 -9000
rect 23990 -9120 24015 -9000
rect 18485 -9175 24015 -9120
rect 18485 -9295 18510 -9175
rect 18630 -9295 18675 -9175
rect 18795 -9295 18840 -9175
rect 18960 -9295 19005 -9175
rect 19125 -9295 19180 -9175
rect 19300 -9295 19345 -9175
rect 19465 -9295 19510 -9175
rect 19630 -9295 19675 -9175
rect 19795 -9295 19850 -9175
rect 19970 -9295 20015 -9175
rect 20135 -9295 20180 -9175
rect 20300 -9295 20345 -9175
rect 20465 -9295 20520 -9175
rect 20640 -9295 20685 -9175
rect 20805 -9295 20850 -9175
rect 20970 -9295 21015 -9175
rect 21135 -9295 21190 -9175
rect 21310 -9295 21355 -9175
rect 21475 -9295 21520 -9175
rect 21640 -9295 21685 -9175
rect 21805 -9295 21860 -9175
rect 21980 -9295 22025 -9175
rect 22145 -9295 22190 -9175
rect 22310 -9295 22355 -9175
rect 22475 -9295 22530 -9175
rect 22650 -9295 22695 -9175
rect 22815 -9295 22860 -9175
rect 22980 -9295 23025 -9175
rect 23145 -9295 23200 -9175
rect 23320 -9295 23365 -9175
rect 23485 -9295 23530 -9175
rect 23650 -9295 23695 -9175
rect 23815 -9295 23870 -9175
rect 23990 -9295 24015 -9175
rect 18485 -9340 24015 -9295
rect 18485 -9460 18510 -9340
rect 18630 -9460 18675 -9340
rect 18795 -9460 18840 -9340
rect 18960 -9460 19005 -9340
rect 19125 -9460 19180 -9340
rect 19300 -9460 19345 -9340
rect 19465 -9460 19510 -9340
rect 19630 -9460 19675 -9340
rect 19795 -9460 19850 -9340
rect 19970 -9460 20015 -9340
rect 20135 -9460 20180 -9340
rect 20300 -9460 20345 -9340
rect 20465 -9460 20520 -9340
rect 20640 -9460 20685 -9340
rect 20805 -9460 20850 -9340
rect 20970 -9460 21015 -9340
rect 21135 -9460 21190 -9340
rect 21310 -9460 21355 -9340
rect 21475 -9460 21520 -9340
rect 21640 -9460 21685 -9340
rect 21805 -9460 21860 -9340
rect 21980 -9460 22025 -9340
rect 22145 -9460 22190 -9340
rect 22310 -9460 22355 -9340
rect 22475 -9460 22530 -9340
rect 22650 -9460 22695 -9340
rect 22815 -9460 22860 -9340
rect 22980 -9460 23025 -9340
rect 23145 -9460 23200 -9340
rect 23320 -9460 23365 -9340
rect 23485 -9460 23530 -9340
rect 23650 -9460 23695 -9340
rect 23815 -9460 23870 -9340
rect 23990 -9460 24015 -9340
rect 18485 -9505 24015 -9460
rect 18485 -9625 18510 -9505
rect 18630 -9625 18675 -9505
rect 18795 -9625 18840 -9505
rect 18960 -9625 19005 -9505
rect 19125 -9625 19180 -9505
rect 19300 -9625 19345 -9505
rect 19465 -9625 19510 -9505
rect 19630 -9625 19675 -9505
rect 19795 -9625 19850 -9505
rect 19970 -9625 20015 -9505
rect 20135 -9625 20180 -9505
rect 20300 -9625 20345 -9505
rect 20465 -9625 20520 -9505
rect 20640 -9625 20685 -9505
rect 20805 -9625 20850 -9505
rect 20970 -9625 21015 -9505
rect 21135 -9625 21190 -9505
rect 21310 -9625 21355 -9505
rect 21475 -9625 21520 -9505
rect 21640 -9625 21685 -9505
rect 21805 -9625 21860 -9505
rect 21980 -9625 22025 -9505
rect 22145 -9625 22190 -9505
rect 22310 -9625 22355 -9505
rect 22475 -9625 22530 -9505
rect 22650 -9625 22695 -9505
rect 22815 -9625 22860 -9505
rect 22980 -9625 23025 -9505
rect 23145 -9625 23200 -9505
rect 23320 -9625 23365 -9505
rect 23485 -9625 23530 -9505
rect 23650 -9625 23695 -9505
rect 23815 -9625 23870 -9505
rect 23990 -9625 24015 -9505
rect 18485 -9670 24015 -9625
rect 18485 -9790 18510 -9670
rect 18630 -9790 18675 -9670
rect 18795 -9790 18840 -9670
rect 18960 -9790 19005 -9670
rect 19125 -9790 19180 -9670
rect 19300 -9790 19345 -9670
rect 19465 -9790 19510 -9670
rect 19630 -9790 19675 -9670
rect 19795 -9790 19850 -9670
rect 19970 -9790 20015 -9670
rect 20135 -9790 20180 -9670
rect 20300 -9790 20345 -9670
rect 20465 -9790 20520 -9670
rect 20640 -9790 20685 -9670
rect 20805 -9790 20850 -9670
rect 20970 -9790 21015 -9670
rect 21135 -9790 21190 -9670
rect 21310 -9790 21355 -9670
rect 21475 -9790 21520 -9670
rect 21640 -9790 21685 -9670
rect 21805 -9790 21860 -9670
rect 21980 -9790 22025 -9670
rect 22145 -9790 22190 -9670
rect 22310 -9790 22355 -9670
rect 22475 -9790 22530 -9670
rect 22650 -9790 22695 -9670
rect 22815 -9790 22860 -9670
rect 22980 -9790 23025 -9670
rect 23145 -9790 23200 -9670
rect 23320 -9790 23365 -9670
rect 23485 -9790 23530 -9670
rect 23650 -9790 23695 -9670
rect 23815 -9790 23870 -9670
rect 23990 -9790 24015 -9670
rect 18485 -9815 24015 -9790
rect 24175 -4430 24200 -4345
rect 24320 -4430 24365 -4310
rect 24485 -4430 24530 -4310
rect 24650 -4430 24695 -4310
rect 24815 -4430 24870 -4310
rect 24990 -4430 25035 -4310
rect 25155 -4430 25200 -4310
rect 25320 -4430 25365 -4310
rect 25485 -4430 25540 -4310
rect 25660 -4430 25705 -4310
rect 25825 -4430 25870 -4310
rect 25990 -4430 26035 -4310
rect 26155 -4430 26210 -4310
rect 26330 -4430 26375 -4310
rect 26495 -4430 26540 -4310
rect 26660 -4430 26705 -4310
rect 26825 -4430 26880 -4310
rect 27000 -4430 27045 -4310
rect 27165 -4430 27210 -4310
rect 27330 -4430 27375 -4310
rect 27495 -4430 27550 -4310
rect 27670 -4430 27715 -4310
rect 27835 -4430 27880 -4310
rect 28000 -4430 28045 -4310
rect 28165 -4430 28220 -4310
rect 28340 -4430 28385 -4310
rect 28505 -4430 28550 -4310
rect 28670 -4430 28715 -4310
rect 28835 -4430 28890 -4310
rect 29010 -4430 29055 -4310
rect 29175 -4430 29220 -4310
rect 29340 -4430 29385 -4310
rect 29505 -4430 29560 -4310
rect 29680 -4430 29705 -4310
rect 24175 -4485 29705 -4430
rect 24175 -4605 24200 -4485
rect 24320 -4605 24365 -4485
rect 24485 -4605 24530 -4485
rect 24650 -4605 24695 -4485
rect 24815 -4605 24870 -4485
rect 24990 -4605 25035 -4485
rect 25155 -4605 25200 -4485
rect 25320 -4605 25365 -4485
rect 25485 -4605 25540 -4485
rect 25660 -4605 25705 -4485
rect 25825 -4605 25870 -4485
rect 25990 -4605 26035 -4485
rect 26155 -4605 26210 -4485
rect 26330 -4605 26375 -4485
rect 26495 -4605 26540 -4485
rect 26660 -4605 26705 -4485
rect 26825 -4605 26880 -4485
rect 27000 -4605 27045 -4485
rect 27165 -4605 27210 -4485
rect 27330 -4605 27375 -4485
rect 27495 -4605 27550 -4485
rect 27670 -4605 27715 -4485
rect 27835 -4605 27880 -4485
rect 28000 -4605 28045 -4485
rect 28165 -4605 28220 -4485
rect 28340 -4605 28385 -4485
rect 28505 -4605 28550 -4485
rect 28670 -4605 28715 -4485
rect 28835 -4605 28890 -4485
rect 29010 -4605 29055 -4485
rect 29175 -4605 29220 -4485
rect 29340 -4605 29385 -4485
rect 29505 -4605 29560 -4485
rect 29680 -4605 29705 -4485
rect 24175 -4650 29705 -4605
rect 24175 -4770 24200 -4650
rect 24320 -4770 24365 -4650
rect 24485 -4770 24530 -4650
rect 24650 -4770 24695 -4650
rect 24815 -4770 24870 -4650
rect 24990 -4770 25035 -4650
rect 25155 -4770 25200 -4650
rect 25320 -4770 25365 -4650
rect 25485 -4770 25540 -4650
rect 25660 -4770 25705 -4650
rect 25825 -4770 25870 -4650
rect 25990 -4770 26035 -4650
rect 26155 -4770 26210 -4650
rect 26330 -4770 26375 -4650
rect 26495 -4770 26540 -4650
rect 26660 -4770 26705 -4650
rect 26825 -4770 26880 -4650
rect 27000 -4770 27045 -4650
rect 27165 -4770 27210 -4650
rect 27330 -4770 27375 -4650
rect 27495 -4770 27550 -4650
rect 27670 -4770 27715 -4650
rect 27835 -4770 27880 -4650
rect 28000 -4770 28045 -4650
rect 28165 -4770 28220 -4650
rect 28340 -4770 28385 -4650
rect 28505 -4770 28550 -4650
rect 28670 -4770 28715 -4650
rect 28835 -4770 28890 -4650
rect 29010 -4770 29055 -4650
rect 29175 -4770 29220 -4650
rect 29340 -4770 29385 -4650
rect 29505 -4770 29560 -4650
rect 29680 -4770 29705 -4650
rect 24175 -4815 29705 -4770
rect 24175 -4935 24200 -4815
rect 24320 -4935 24365 -4815
rect 24485 -4935 24530 -4815
rect 24650 -4935 24695 -4815
rect 24815 -4935 24870 -4815
rect 24990 -4935 25035 -4815
rect 25155 -4935 25200 -4815
rect 25320 -4935 25365 -4815
rect 25485 -4935 25540 -4815
rect 25660 -4935 25705 -4815
rect 25825 -4935 25870 -4815
rect 25990 -4935 26035 -4815
rect 26155 -4935 26210 -4815
rect 26330 -4935 26375 -4815
rect 26495 -4935 26540 -4815
rect 26660 -4935 26705 -4815
rect 26825 -4935 26880 -4815
rect 27000 -4935 27045 -4815
rect 27165 -4935 27210 -4815
rect 27330 -4935 27375 -4815
rect 27495 -4935 27550 -4815
rect 27670 -4935 27715 -4815
rect 27835 -4935 27880 -4815
rect 28000 -4935 28045 -4815
rect 28165 -4935 28220 -4815
rect 28340 -4935 28385 -4815
rect 28505 -4935 28550 -4815
rect 28670 -4935 28715 -4815
rect 28835 -4935 28890 -4815
rect 29010 -4935 29055 -4815
rect 29175 -4935 29220 -4815
rect 29340 -4935 29385 -4815
rect 29505 -4935 29560 -4815
rect 29680 -4935 29705 -4815
rect 24175 -4980 29705 -4935
rect 24175 -5100 24200 -4980
rect 24320 -5100 24365 -4980
rect 24485 -5100 24530 -4980
rect 24650 -5100 24695 -4980
rect 24815 -5100 24870 -4980
rect 24990 -5100 25035 -4980
rect 25155 -5100 25200 -4980
rect 25320 -5100 25365 -4980
rect 25485 -5100 25540 -4980
rect 25660 -5100 25705 -4980
rect 25825 -5100 25870 -4980
rect 25990 -5100 26035 -4980
rect 26155 -5100 26210 -4980
rect 26330 -5100 26375 -4980
rect 26495 -5100 26540 -4980
rect 26660 -5100 26705 -4980
rect 26825 -5100 26880 -4980
rect 27000 -5100 27045 -4980
rect 27165 -5100 27210 -4980
rect 27330 -5100 27375 -4980
rect 27495 -5100 27550 -4980
rect 27670 -5100 27715 -4980
rect 27835 -5100 27880 -4980
rect 28000 -5100 28045 -4980
rect 28165 -5100 28220 -4980
rect 28340 -5100 28385 -4980
rect 28505 -5100 28550 -4980
rect 28670 -5100 28715 -4980
rect 28835 -5100 28890 -4980
rect 29010 -5100 29055 -4980
rect 29175 -5100 29220 -4980
rect 29340 -5100 29385 -4980
rect 29505 -5100 29560 -4980
rect 29680 -5100 29705 -4980
rect 24175 -5155 29705 -5100
rect 24175 -5275 24200 -5155
rect 24320 -5275 24365 -5155
rect 24485 -5275 24530 -5155
rect 24650 -5275 24695 -5155
rect 24815 -5275 24870 -5155
rect 24990 -5275 25035 -5155
rect 25155 -5275 25200 -5155
rect 25320 -5275 25365 -5155
rect 25485 -5275 25540 -5155
rect 25660 -5275 25705 -5155
rect 25825 -5275 25870 -5155
rect 25990 -5275 26035 -5155
rect 26155 -5275 26210 -5155
rect 26330 -5275 26375 -5155
rect 26495 -5275 26540 -5155
rect 26660 -5275 26705 -5155
rect 26825 -5275 26880 -5155
rect 27000 -5275 27045 -5155
rect 27165 -5275 27210 -5155
rect 27330 -5275 27375 -5155
rect 27495 -5275 27550 -5155
rect 27670 -5275 27715 -5155
rect 27835 -5275 27880 -5155
rect 28000 -5275 28045 -5155
rect 28165 -5275 28220 -5155
rect 28340 -5275 28385 -5155
rect 28505 -5275 28550 -5155
rect 28670 -5275 28715 -5155
rect 28835 -5275 28890 -5155
rect 29010 -5275 29055 -5155
rect 29175 -5275 29220 -5155
rect 29340 -5275 29385 -5155
rect 29505 -5275 29560 -5155
rect 29680 -5275 29705 -5155
rect 24175 -5320 29705 -5275
rect 24175 -5440 24200 -5320
rect 24320 -5440 24365 -5320
rect 24485 -5440 24530 -5320
rect 24650 -5440 24695 -5320
rect 24815 -5440 24870 -5320
rect 24990 -5440 25035 -5320
rect 25155 -5440 25200 -5320
rect 25320 -5440 25365 -5320
rect 25485 -5440 25540 -5320
rect 25660 -5440 25705 -5320
rect 25825 -5440 25870 -5320
rect 25990 -5440 26035 -5320
rect 26155 -5440 26210 -5320
rect 26330 -5440 26375 -5320
rect 26495 -5440 26540 -5320
rect 26660 -5440 26705 -5320
rect 26825 -5440 26880 -5320
rect 27000 -5440 27045 -5320
rect 27165 -5440 27210 -5320
rect 27330 -5440 27375 -5320
rect 27495 -5440 27550 -5320
rect 27670 -5440 27715 -5320
rect 27835 -5440 27880 -5320
rect 28000 -5440 28045 -5320
rect 28165 -5440 28220 -5320
rect 28340 -5440 28385 -5320
rect 28505 -5440 28550 -5320
rect 28670 -5440 28715 -5320
rect 28835 -5440 28890 -5320
rect 29010 -5440 29055 -5320
rect 29175 -5440 29220 -5320
rect 29340 -5440 29385 -5320
rect 29505 -5440 29560 -5320
rect 29680 -5440 29705 -5320
rect 24175 -5485 29705 -5440
rect 24175 -5605 24200 -5485
rect 24320 -5605 24365 -5485
rect 24485 -5605 24530 -5485
rect 24650 -5605 24695 -5485
rect 24815 -5605 24870 -5485
rect 24990 -5605 25035 -5485
rect 25155 -5605 25200 -5485
rect 25320 -5605 25365 -5485
rect 25485 -5605 25540 -5485
rect 25660 -5605 25705 -5485
rect 25825 -5605 25870 -5485
rect 25990 -5605 26035 -5485
rect 26155 -5605 26210 -5485
rect 26330 -5605 26375 -5485
rect 26495 -5605 26540 -5485
rect 26660 -5605 26705 -5485
rect 26825 -5605 26880 -5485
rect 27000 -5605 27045 -5485
rect 27165 -5605 27210 -5485
rect 27330 -5605 27375 -5485
rect 27495 -5605 27550 -5485
rect 27670 -5605 27715 -5485
rect 27835 -5605 27880 -5485
rect 28000 -5605 28045 -5485
rect 28165 -5605 28220 -5485
rect 28340 -5605 28385 -5485
rect 28505 -5605 28550 -5485
rect 28670 -5605 28715 -5485
rect 28835 -5605 28890 -5485
rect 29010 -5605 29055 -5485
rect 29175 -5605 29220 -5485
rect 29340 -5605 29385 -5485
rect 29505 -5605 29560 -5485
rect 29680 -5605 29705 -5485
rect 24175 -5650 29705 -5605
rect 24175 -5770 24200 -5650
rect 24320 -5770 24365 -5650
rect 24485 -5770 24530 -5650
rect 24650 -5770 24695 -5650
rect 24815 -5770 24870 -5650
rect 24990 -5770 25035 -5650
rect 25155 -5770 25200 -5650
rect 25320 -5770 25365 -5650
rect 25485 -5770 25540 -5650
rect 25660 -5770 25705 -5650
rect 25825 -5770 25870 -5650
rect 25990 -5770 26035 -5650
rect 26155 -5770 26210 -5650
rect 26330 -5770 26375 -5650
rect 26495 -5770 26540 -5650
rect 26660 -5770 26705 -5650
rect 26825 -5770 26880 -5650
rect 27000 -5770 27045 -5650
rect 27165 -5770 27210 -5650
rect 27330 -5770 27375 -5650
rect 27495 -5770 27550 -5650
rect 27670 -5770 27715 -5650
rect 27835 -5770 27880 -5650
rect 28000 -5770 28045 -5650
rect 28165 -5770 28220 -5650
rect 28340 -5770 28385 -5650
rect 28505 -5770 28550 -5650
rect 28670 -5770 28715 -5650
rect 28835 -5770 28890 -5650
rect 29010 -5770 29055 -5650
rect 29175 -5770 29220 -5650
rect 29340 -5770 29385 -5650
rect 29505 -5770 29560 -5650
rect 29680 -5770 29705 -5650
rect 24175 -5825 29705 -5770
rect 24175 -5945 24200 -5825
rect 24320 -5945 24365 -5825
rect 24485 -5945 24530 -5825
rect 24650 -5945 24695 -5825
rect 24815 -5945 24870 -5825
rect 24990 -5945 25035 -5825
rect 25155 -5945 25200 -5825
rect 25320 -5945 25365 -5825
rect 25485 -5945 25540 -5825
rect 25660 -5945 25705 -5825
rect 25825 -5945 25870 -5825
rect 25990 -5945 26035 -5825
rect 26155 -5945 26210 -5825
rect 26330 -5945 26375 -5825
rect 26495 -5945 26540 -5825
rect 26660 -5945 26705 -5825
rect 26825 -5945 26880 -5825
rect 27000 -5945 27045 -5825
rect 27165 -5945 27210 -5825
rect 27330 -5945 27375 -5825
rect 27495 -5945 27550 -5825
rect 27670 -5945 27715 -5825
rect 27835 -5945 27880 -5825
rect 28000 -5945 28045 -5825
rect 28165 -5945 28220 -5825
rect 28340 -5945 28385 -5825
rect 28505 -5945 28550 -5825
rect 28670 -5945 28715 -5825
rect 28835 -5945 28890 -5825
rect 29010 -5945 29055 -5825
rect 29175 -5945 29220 -5825
rect 29340 -5945 29385 -5825
rect 29505 -5945 29560 -5825
rect 29680 -5945 29705 -5825
rect 24175 -5990 29705 -5945
rect 24175 -6110 24200 -5990
rect 24320 -6110 24365 -5990
rect 24485 -6110 24530 -5990
rect 24650 -6110 24695 -5990
rect 24815 -6110 24870 -5990
rect 24990 -6110 25035 -5990
rect 25155 -6110 25200 -5990
rect 25320 -6110 25365 -5990
rect 25485 -6110 25540 -5990
rect 25660 -6110 25705 -5990
rect 25825 -6110 25870 -5990
rect 25990 -6110 26035 -5990
rect 26155 -6110 26210 -5990
rect 26330 -6110 26375 -5990
rect 26495 -6110 26540 -5990
rect 26660 -6110 26705 -5990
rect 26825 -6110 26880 -5990
rect 27000 -6110 27045 -5990
rect 27165 -6110 27210 -5990
rect 27330 -6110 27375 -5990
rect 27495 -6110 27550 -5990
rect 27670 -6110 27715 -5990
rect 27835 -6110 27880 -5990
rect 28000 -6110 28045 -5990
rect 28165 -6110 28220 -5990
rect 28340 -6110 28385 -5990
rect 28505 -6110 28550 -5990
rect 28670 -6110 28715 -5990
rect 28835 -6110 28890 -5990
rect 29010 -6110 29055 -5990
rect 29175 -6110 29220 -5990
rect 29340 -6110 29385 -5990
rect 29505 -6110 29560 -5990
rect 29680 -6110 29705 -5990
rect 24175 -6155 29705 -6110
rect 24175 -6275 24200 -6155
rect 24320 -6275 24365 -6155
rect 24485 -6275 24530 -6155
rect 24650 -6275 24695 -6155
rect 24815 -6275 24870 -6155
rect 24990 -6275 25035 -6155
rect 25155 -6275 25200 -6155
rect 25320 -6275 25365 -6155
rect 25485 -6275 25540 -6155
rect 25660 -6275 25705 -6155
rect 25825 -6275 25870 -6155
rect 25990 -6275 26035 -6155
rect 26155 -6275 26210 -6155
rect 26330 -6275 26375 -6155
rect 26495 -6275 26540 -6155
rect 26660 -6275 26705 -6155
rect 26825 -6275 26880 -6155
rect 27000 -6275 27045 -6155
rect 27165 -6275 27210 -6155
rect 27330 -6275 27375 -6155
rect 27495 -6275 27550 -6155
rect 27670 -6275 27715 -6155
rect 27835 -6275 27880 -6155
rect 28000 -6275 28045 -6155
rect 28165 -6275 28220 -6155
rect 28340 -6275 28385 -6155
rect 28505 -6275 28550 -6155
rect 28670 -6275 28715 -6155
rect 28835 -6275 28890 -6155
rect 29010 -6275 29055 -6155
rect 29175 -6275 29220 -6155
rect 29340 -6275 29385 -6155
rect 29505 -6275 29560 -6155
rect 29680 -6275 29705 -6155
rect 24175 -6320 29705 -6275
rect 24175 -6440 24200 -6320
rect 24320 -6440 24365 -6320
rect 24485 -6440 24530 -6320
rect 24650 -6440 24695 -6320
rect 24815 -6440 24870 -6320
rect 24990 -6440 25035 -6320
rect 25155 -6440 25200 -6320
rect 25320 -6440 25365 -6320
rect 25485 -6440 25540 -6320
rect 25660 -6440 25705 -6320
rect 25825 -6440 25870 -6320
rect 25990 -6440 26035 -6320
rect 26155 -6440 26210 -6320
rect 26330 -6440 26375 -6320
rect 26495 -6440 26540 -6320
rect 26660 -6440 26705 -6320
rect 26825 -6440 26880 -6320
rect 27000 -6440 27045 -6320
rect 27165 -6440 27210 -6320
rect 27330 -6440 27375 -6320
rect 27495 -6440 27550 -6320
rect 27670 -6440 27715 -6320
rect 27835 -6440 27880 -6320
rect 28000 -6440 28045 -6320
rect 28165 -6440 28220 -6320
rect 28340 -6440 28385 -6320
rect 28505 -6440 28550 -6320
rect 28670 -6440 28715 -6320
rect 28835 -6440 28890 -6320
rect 29010 -6440 29055 -6320
rect 29175 -6440 29220 -6320
rect 29340 -6440 29385 -6320
rect 29505 -6440 29560 -6320
rect 29680 -6440 29705 -6320
rect 24175 -6495 29705 -6440
rect 24175 -6615 24200 -6495
rect 24320 -6615 24365 -6495
rect 24485 -6615 24530 -6495
rect 24650 -6615 24695 -6495
rect 24815 -6615 24870 -6495
rect 24990 -6615 25035 -6495
rect 25155 -6615 25200 -6495
rect 25320 -6615 25365 -6495
rect 25485 -6615 25540 -6495
rect 25660 -6615 25705 -6495
rect 25825 -6615 25870 -6495
rect 25990 -6615 26035 -6495
rect 26155 -6615 26210 -6495
rect 26330 -6615 26375 -6495
rect 26495 -6615 26540 -6495
rect 26660 -6615 26705 -6495
rect 26825 -6615 26880 -6495
rect 27000 -6615 27045 -6495
rect 27165 -6615 27210 -6495
rect 27330 -6615 27375 -6495
rect 27495 -6615 27550 -6495
rect 27670 -6615 27715 -6495
rect 27835 -6615 27880 -6495
rect 28000 -6615 28045 -6495
rect 28165 -6615 28220 -6495
rect 28340 -6615 28385 -6495
rect 28505 -6615 28550 -6495
rect 28670 -6615 28715 -6495
rect 28835 -6615 28890 -6495
rect 29010 -6615 29055 -6495
rect 29175 -6615 29220 -6495
rect 29340 -6615 29385 -6495
rect 29505 -6615 29560 -6495
rect 29680 -6615 29705 -6495
rect 24175 -6660 29705 -6615
rect 24175 -6780 24200 -6660
rect 24320 -6780 24365 -6660
rect 24485 -6780 24530 -6660
rect 24650 -6780 24695 -6660
rect 24815 -6780 24870 -6660
rect 24990 -6780 25035 -6660
rect 25155 -6780 25200 -6660
rect 25320 -6780 25365 -6660
rect 25485 -6780 25540 -6660
rect 25660 -6780 25705 -6660
rect 25825 -6780 25870 -6660
rect 25990 -6780 26035 -6660
rect 26155 -6780 26210 -6660
rect 26330 -6780 26375 -6660
rect 26495 -6780 26540 -6660
rect 26660 -6780 26705 -6660
rect 26825 -6780 26880 -6660
rect 27000 -6780 27045 -6660
rect 27165 -6780 27210 -6660
rect 27330 -6780 27375 -6660
rect 27495 -6780 27550 -6660
rect 27670 -6780 27715 -6660
rect 27835 -6780 27880 -6660
rect 28000 -6780 28045 -6660
rect 28165 -6780 28220 -6660
rect 28340 -6780 28385 -6660
rect 28505 -6780 28550 -6660
rect 28670 -6780 28715 -6660
rect 28835 -6780 28890 -6660
rect 29010 -6780 29055 -6660
rect 29175 -6780 29220 -6660
rect 29340 -6780 29385 -6660
rect 29505 -6780 29560 -6660
rect 29680 -6780 29705 -6660
rect 24175 -6825 29705 -6780
rect 24175 -6945 24200 -6825
rect 24320 -6945 24365 -6825
rect 24485 -6945 24530 -6825
rect 24650 -6945 24695 -6825
rect 24815 -6945 24870 -6825
rect 24990 -6945 25035 -6825
rect 25155 -6945 25200 -6825
rect 25320 -6945 25365 -6825
rect 25485 -6945 25540 -6825
rect 25660 -6945 25705 -6825
rect 25825 -6945 25870 -6825
rect 25990 -6945 26035 -6825
rect 26155 -6945 26210 -6825
rect 26330 -6945 26375 -6825
rect 26495 -6945 26540 -6825
rect 26660 -6945 26705 -6825
rect 26825 -6945 26880 -6825
rect 27000 -6945 27045 -6825
rect 27165 -6945 27210 -6825
rect 27330 -6945 27375 -6825
rect 27495 -6945 27550 -6825
rect 27670 -6945 27715 -6825
rect 27835 -6945 27880 -6825
rect 28000 -6945 28045 -6825
rect 28165 -6945 28220 -6825
rect 28340 -6945 28385 -6825
rect 28505 -6945 28550 -6825
rect 28670 -6945 28715 -6825
rect 28835 -6945 28890 -6825
rect 29010 -6945 29055 -6825
rect 29175 -6945 29220 -6825
rect 29340 -6945 29385 -6825
rect 29505 -6945 29560 -6825
rect 29680 -6945 29705 -6825
rect 24175 -6990 29705 -6945
rect 24175 -7110 24200 -6990
rect 24320 -7110 24365 -6990
rect 24485 -7110 24530 -6990
rect 24650 -7110 24695 -6990
rect 24815 -7110 24870 -6990
rect 24990 -7110 25035 -6990
rect 25155 -7110 25200 -6990
rect 25320 -7110 25365 -6990
rect 25485 -7110 25540 -6990
rect 25660 -7110 25705 -6990
rect 25825 -7110 25870 -6990
rect 25990 -7110 26035 -6990
rect 26155 -7110 26210 -6990
rect 26330 -7110 26375 -6990
rect 26495 -7110 26540 -6990
rect 26660 -7110 26705 -6990
rect 26825 -7110 26880 -6990
rect 27000 -7110 27045 -6990
rect 27165 -7110 27210 -6990
rect 27330 -7110 27375 -6990
rect 27495 -7110 27550 -6990
rect 27670 -7110 27715 -6990
rect 27835 -7110 27880 -6990
rect 28000 -7110 28045 -6990
rect 28165 -7110 28220 -6990
rect 28340 -7110 28385 -6990
rect 28505 -7110 28550 -6990
rect 28670 -7110 28715 -6990
rect 28835 -7110 28890 -6990
rect 29010 -7110 29055 -6990
rect 29175 -7110 29220 -6990
rect 29340 -7110 29385 -6990
rect 29505 -7110 29560 -6990
rect 29680 -7110 29705 -6990
rect 24175 -7165 29705 -7110
rect 24175 -7285 24200 -7165
rect 24320 -7285 24365 -7165
rect 24485 -7285 24530 -7165
rect 24650 -7285 24695 -7165
rect 24815 -7285 24870 -7165
rect 24990 -7285 25035 -7165
rect 25155 -7285 25200 -7165
rect 25320 -7285 25365 -7165
rect 25485 -7285 25540 -7165
rect 25660 -7285 25705 -7165
rect 25825 -7285 25870 -7165
rect 25990 -7285 26035 -7165
rect 26155 -7285 26210 -7165
rect 26330 -7285 26375 -7165
rect 26495 -7285 26540 -7165
rect 26660 -7285 26705 -7165
rect 26825 -7285 26880 -7165
rect 27000 -7285 27045 -7165
rect 27165 -7285 27210 -7165
rect 27330 -7285 27375 -7165
rect 27495 -7285 27550 -7165
rect 27670 -7285 27715 -7165
rect 27835 -7285 27880 -7165
rect 28000 -7285 28045 -7165
rect 28165 -7285 28220 -7165
rect 28340 -7285 28385 -7165
rect 28505 -7285 28550 -7165
rect 28670 -7285 28715 -7165
rect 28835 -7285 28890 -7165
rect 29010 -7285 29055 -7165
rect 29175 -7285 29220 -7165
rect 29340 -7285 29385 -7165
rect 29505 -7285 29560 -7165
rect 29680 -7285 29705 -7165
rect 24175 -7330 29705 -7285
rect 24175 -7450 24200 -7330
rect 24320 -7450 24365 -7330
rect 24485 -7450 24530 -7330
rect 24650 -7450 24695 -7330
rect 24815 -7450 24870 -7330
rect 24990 -7450 25035 -7330
rect 25155 -7450 25200 -7330
rect 25320 -7450 25365 -7330
rect 25485 -7450 25540 -7330
rect 25660 -7450 25705 -7330
rect 25825 -7450 25870 -7330
rect 25990 -7450 26035 -7330
rect 26155 -7450 26210 -7330
rect 26330 -7450 26375 -7330
rect 26495 -7450 26540 -7330
rect 26660 -7450 26705 -7330
rect 26825 -7450 26880 -7330
rect 27000 -7450 27045 -7330
rect 27165 -7450 27210 -7330
rect 27330 -7450 27375 -7330
rect 27495 -7450 27550 -7330
rect 27670 -7450 27715 -7330
rect 27835 -7450 27880 -7330
rect 28000 -7450 28045 -7330
rect 28165 -7450 28220 -7330
rect 28340 -7450 28385 -7330
rect 28505 -7450 28550 -7330
rect 28670 -7450 28715 -7330
rect 28835 -7450 28890 -7330
rect 29010 -7450 29055 -7330
rect 29175 -7450 29220 -7330
rect 29340 -7450 29385 -7330
rect 29505 -7450 29560 -7330
rect 29680 -7450 29705 -7330
rect 24175 -7495 29705 -7450
rect 24175 -7615 24200 -7495
rect 24320 -7615 24365 -7495
rect 24485 -7615 24530 -7495
rect 24650 -7615 24695 -7495
rect 24815 -7615 24870 -7495
rect 24990 -7615 25035 -7495
rect 25155 -7615 25200 -7495
rect 25320 -7615 25365 -7495
rect 25485 -7615 25540 -7495
rect 25660 -7615 25705 -7495
rect 25825 -7615 25870 -7495
rect 25990 -7615 26035 -7495
rect 26155 -7615 26210 -7495
rect 26330 -7615 26375 -7495
rect 26495 -7615 26540 -7495
rect 26660 -7615 26705 -7495
rect 26825 -7615 26880 -7495
rect 27000 -7615 27045 -7495
rect 27165 -7615 27210 -7495
rect 27330 -7615 27375 -7495
rect 27495 -7615 27550 -7495
rect 27670 -7615 27715 -7495
rect 27835 -7615 27880 -7495
rect 28000 -7615 28045 -7495
rect 28165 -7615 28220 -7495
rect 28340 -7615 28385 -7495
rect 28505 -7615 28550 -7495
rect 28670 -7615 28715 -7495
rect 28835 -7615 28890 -7495
rect 29010 -7615 29055 -7495
rect 29175 -7615 29220 -7495
rect 29340 -7615 29385 -7495
rect 29505 -7615 29560 -7495
rect 29680 -7615 29705 -7495
rect 24175 -7660 29705 -7615
rect 24175 -7780 24200 -7660
rect 24320 -7780 24365 -7660
rect 24485 -7780 24530 -7660
rect 24650 -7780 24695 -7660
rect 24815 -7780 24870 -7660
rect 24990 -7780 25035 -7660
rect 25155 -7780 25200 -7660
rect 25320 -7780 25365 -7660
rect 25485 -7780 25540 -7660
rect 25660 -7780 25705 -7660
rect 25825 -7780 25870 -7660
rect 25990 -7780 26035 -7660
rect 26155 -7780 26210 -7660
rect 26330 -7780 26375 -7660
rect 26495 -7780 26540 -7660
rect 26660 -7780 26705 -7660
rect 26825 -7780 26880 -7660
rect 27000 -7780 27045 -7660
rect 27165 -7780 27210 -7660
rect 27330 -7780 27375 -7660
rect 27495 -7780 27550 -7660
rect 27670 -7780 27715 -7660
rect 27835 -7780 27880 -7660
rect 28000 -7780 28045 -7660
rect 28165 -7780 28220 -7660
rect 28340 -7780 28385 -7660
rect 28505 -7780 28550 -7660
rect 28670 -7780 28715 -7660
rect 28835 -7780 28890 -7660
rect 29010 -7780 29055 -7660
rect 29175 -7780 29220 -7660
rect 29340 -7780 29385 -7660
rect 29505 -7780 29560 -7660
rect 29680 -7780 29705 -7660
rect 24175 -7835 29705 -7780
rect 24175 -7955 24200 -7835
rect 24320 -7955 24365 -7835
rect 24485 -7955 24530 -7835
rect 24650 -7955 24695 -7835
rect 24815 -7955 24870 -7835
rect 24990 -7955 25035 -7835
rect 25155 -7955 25200 -7835
rect 25320 -7955 25365 -7835
rect 25485 -7955 25540 -7835
rect 25660 -7955 25705 -7835
rect 25825 -7955 25870 -7835
rect 25990 -7955 26035 -7835
rect 26155 -7955 26210 -7835
rect 26330 -7955 26375 -7835
rect 26495 -7955 26540 -7835
rect 26660 -7955 26705 -7835
rect 26825 -7955 26880 -7835
rect 27000 -7955 27045 -7835
rect 27165 -7955 27210 -7835
rect 27330 -7955 27375 -7835
rect 27495 -7955 27550 -7835
rect 27670 -7955 27715 -7835
rect 27835 -7955 27880 -7835
rect 28000 -7955 28045 -7835
rect 28165 -7955 28220 -7835
rect 28340 -7955 28385 -7835
rect 28505 -7955 28550 -7835
rect 28670 -7955 28715 -7835
rect 28835 -7955 28890 -7835
rect 29010 -7955 29055 -7835
rect 29175 -7955 29220 -7835
rect 29340 -7955 29385 -7835
rect 29505 -7955 29560 -7835
rect 29680 -7955 29705 -7835
rect 24175 -8000 29705 -7955
rect 24175 -8120 24200 -8000
rect 24320 -8120 24365 -8000
rect 24485 -8120 24530 -8000
rect 24650 -8120 24695 -8000
rect 24815 -8120 24870 -8000
rect 24990 -8120 25035 -8000
rect 25155 -8120 25200 -8000
rect 25320 -8120 25365 -8000
rect 25485 -8120 25540 -8000
rect 25660 -8120 25705 -8000
rect 25825 -8120 25870 -8000
rect 25990 -8120 26035 -8000
rect 26155 -8120 26210 -8000
rect 26330 -8120 26375 -8000
rect 26495 -8120 26540 -8000
rect 26660 -8120 26705 -8000
rect 26825 -8120 26880 -8000
rect 27000 -8120 27045 -8000
rect 27165 -8120 27210 -8000
rect 27330 -8120 27375 -8000
rect 27495 -8120 27550 -8000
rect 27670 -8120 27715 -8000
rect 27835 -8120 27880 -8000
rect 28000 -8120 28045 -8000
rect 28165 -8120 28220 -8000
rect 28340 -8120 28385 -8000
rect 28505 -8120 28550 -8000
rect 28670 -8120 28715 -8000
rect 28835 -8120 28890 -8000
rect 29010 -8120 29055 -8000
rect 29175 -8120 29220 -8000
rect 29340 -8120 29385 -8000
rect 29505 -8120 29560 -8000
rect 29680 -8120 29705 -8000
rect 24175 -8165 29705 -8120
rect 24175 -8285 24200 -8165
rect 24320 -8285 24365 -8165
rect 24485 -8285 24530 -8165
rect 24650 -8285 24695 -8165
rect 24815 -8285 24870 -8165
rect 24990 -8285 25035 -8165
rect 25155 -8285 25200 -8165
rect 25320 -8285 25365 -8165
rect 25485 -8285 25540 -8165
rect 25660 -8285 25705 -8165
rect 25825 -8285 25870 -8165
rect 25990 -8285 26035 -8165
rect 26155 -8285 26210 -8165
rect 26330 -8285 26375 -8165
rect 26495 -8285 26540 -8165
rect 26660 -8285 26705 -8165
rect 26825 -8285 26880 -8165
rect 27000 -8285 27045 -8165
rect 27165 -8285 27210 -8165
rect 27330 -8285 27375 -8165
rect 27495 -8285 27550 -8165
rect 27670 -8285 27715 -8165
rect 27835 -8285 27880 -8165
rect 28000 -8285 28045 -8165
rect 28165 -8285 28220 -8165
rect 28340 -8285 28385 -8165
rect 28505 -8285 28550 -8165
rect 28670 -8285 28715 -8165
rect 28835 -8285 28890 -8165
rect 29010 -8285 29055 -8165
rect 29175 -8285 29220 -8165
rect 29340 -8285 29385 -8165
rect 29505 -8285 29560 -8165
rect 29680 -8285 29705 -8165
rect 24175 -8330 29705 -8285
rect 24175 -8450 24200 -8330
rect 24320 -8450 24365 -8330
rect 24485 -8450 24530 -8330
rect 24650 -8450 24695 -8330
rect 24815 -8450 24870 -8330
rect 24990 -8450 25035 -8330
rect 25155 -8450 25200 -8330
rect 25320 -8450 25365 -8330
rect 25485 -8450 25540 -8330
rect 25660 -8450 25705 -8330
rect 25825 -8450 25870 -8330
rect 25990 -8450 26035 -8330
rect 26155 -8450 26210 -8330
rect 26330 -8450 26375 -8330
rect 26495 -8450 26540 -8330
rect 26660 -8450 26705 -8330
rect 26825 -8450 26880 -8330
rect 27000 -8450 27045 -8330
rect 27165 -8450 27210 -8330
rect 27330 -8450 27375 -8330
rect 27495 -8450 27550 -8330
rect 27670 -8450 27715 -8330
rect 27835 -8450 27880 -8330
rect 28000 -8450 28045 -8330
rect 28165 -8450 28220 -8330
rect 28340 -8450 28385 -8330
rect 28505 -8450 28550 -8330
rect 28670 -8450 28715 -8330
rect 28835 -8450 28890 -8330
rect 29010 -8450 29055 -8330
rect 29175 -8450 29220 -8330
rect 29340 -8450 29385 -8330
rect 29505 -8450 29560 -8330
rect 29680 -8450 29705 -8330
rect 24175 -8505 29705 -8450
rect 24175 -8625 24200 -8505
rect 24320 -8625 24365 -8505
rect 24485 -8625 24530 -8505
rect 24650 -8625 24695 -8505
rect 24815 -8625 24870 -8505
rect 24990 -8625 25035 -8505
rect 25155 -8625 25200 -8505
rect 25320 -8625 25365 -8505
rect 25485 -8625 25540 -8505
rect 25660 -8625 25705 -8505
rect 25825 -8625 25870 -8505
rect 25990 -8625 26035 -8505
rect 26155 -8625 26210 -8505
rect 26330 -8625 26375 -8505
rect 26495 -8625 26540 -8505
rect 26660 -8625 26705 -8505
rect 26825 -8625 26880 -8505
rect 27000 -8625 27045 -8505
rect 27165 -8625 27210 -8505
rect 27330 -8625 27375 -8505
rect 27495 -8625 27550 -8505
rect 27670 -8625 27715 -8505
rect 27835 -8625 27880 -8505
rect 28000 -8625 28045 -8505
rect 28165 -8625 28220 -8505
rect 28340 -8625 28385 -8505
rect 28505 -8625 28550 -8505
rect 28670 -8625 28715 -8505
rect 28835 -8625 28890 -8505
rect 29010 -8625 29055 -8505
rect 29175 -8625 29220 -8505
rect 29340 -8625 29385 -8505
rect 29505 -8625 29560 -8505
rect 29680 -8625 29705 -8505
rect 24175 -8670 29705 -8625
rect 24175 -8790 24200 -8670
rect 24320 -8790 24365 -8670
rect 24485 -8790 24530 -8670
rect 24650 -8790 24695 -8670
rect 24815 -8790 24870 -8670
rect 24990 -8790 25035 -8670
rect 25155 -8790 25200 -8670
rect 25320 -8790 25365 -8670
rect 25485 -8790 25540 -8670
rect 25660 -8790 25705 -8670
rect 25825 -8790 25870 -8670
rect 25990 -8790 26035 -8670
rect 26155 -8790 26210 -8670
rect 26330 -8790 26375 -8670
rect 26495 -8790 26540 -8670
rect 26660 -8790 26705 -8670
rect 26825 -8790 26880 -8670
rect 27000 -8790 27045 -8670
rect 27165 -8790 27210 -8670
rect 27330 -8790 27375 -8670
rect 27495 -8790 27550 -8670
rect 27670 -8790 27715 -8670
rect 27835 -8790 27880 -8670
rect 28000 -8790 28045 -8670
rect 28165 -8790 28220 -8670
rect 28340 -8790 28385 -8670
rect 28505 -8790 28550 -8670
rect 28670 -8790 28715 -8670
rect 28835 -8790 28890 -8670
rect 29010 -8790 29055 -8670
rect 29175 -8790 29220 -8670
rect 29340 -8790 29385 -8670
rect 29505 -8790 29560 -8670
rect 29680 -8790 29705 -8670
rect 24175 -8835 29705 -8790
rect 24175 -8955 24200 -8835
rect 24320 -8955 24365 -8835
rect 24485 -8955 24530 -8835
rect 24650 -8955 24695 -8835
rect 24815 -8955 24870 -8835
rect 24990 -8955 25035 -8835
rect 25155 -8955 25200 -8835
rect 25320 -8955 25365 -8835
rect 25485 -8955 25540 -8835
rect 25660 -8955 25705 -8835
rect 25825 -8955 25870 -8835
rect 25990 -8955 26035 -8835
rect 26155 -8955 26210 -8835
rect 26330 -8955 26375 -8835
rect 26495 -8955 26540 -8835
rect 26660 -8955 26705 -8835
rect 26825 -8955 26880 -8835
rect 27000 -8955 27045 -8835
rect 27165 -8955 27210 -8835
rect 27330 -8955 27375 -8835
rect 27495 -8955 27550 -8835
rect 27670 -8955 27715 -8835
rect 27835 -8955 27880 -8835
rect 28000 -8955 28045 -8835
rect 28165 -8955 28220 -8835
rect 28340 -8955 28385 -8835
rect 28505 -8955 28550 -8835
rect 28670 -8955 28715 -8835
rect 28835 -8955 28890 -8835
rect 29010 -8955 29055 -8835
rect 29175 -8955 29220 -8835
rect 29340 -8955 29385 -8835
rect 29505 -8955 29560 -8835
rect 29680 -8955 29705 -8835
rect 24175 -9000 29705 -8955
rect 24175 -9120 24200 -9000
rect 24320 -9120 24365 -9000
rect 24485 -9120 24530 -9000
rect 24650 -9120 24695 -9000
rect 24815 -9120 24870 -9000
rect 24990 -9120 25035 -9000
rect 25155 -9120 25200 -9000
rect 25320 -9120 25365 -9000
rect 25485 -9120 25540 -9000
rect 25660 -9120 25705 -9000
rect 25825 -9120 25870 -9000
rect 25990 -9120 26035 -9000
rect 26155 -9120 26210 -9000
rect 26330 -9120 26375 -9000
rect 26495 -9120 26540 -9000
rect 26660 -9120 26705 -9000
rect 26825 -9120 26880 -9000
rect 27000 -9120 27045 -9000
rect 27165 -9120 27210 -9000
rect 27330 -9120 27375 -9000
rect 27495 -9120 27550 -9000
rect 27670 -9120 27715 -9000
rect 27835 -9120 27880 -9000
rect 28000 -9120 28045 -9000
rect 28165 -9120 28220 -9000
rect 28340 -9120 28385 -9000
rect 28505 -9120 28550 -9000
rect 28670 -9120 28715 -9000
rect 28835 -9120 28890 -9000
rect 29010 -9120 29055 -9000
rect 29175 -9120 29220 -9000
rect 29340 -9120 29385 -9000
rect 29505 -9120 29560 -9000
rect 29680 -9120 29705 -9000
rect 24175 -9175 29705 -9120
rect 24175 -9295 24200 -9175
rect 24320 -9295 24365 -9175
rect 24485 -9295 24530 -9175
rect 24650 -9295 24695 -9175
rect 24815 -9295 24870 -9175
rect 24990 -9295 25035 -9175
rect 25155 -9295 25200 -9175
rect 25320 -9295 25365 -9175
rect 25485 -9295 25540 -9175
rect 25660 -9295 25705 -9175
rect 25825 -9295 25870 -9175
rect 25990 -9295 26035 -9175
rect 26155 -9295 26210 -9175
rect 26330 -9295 26375 -9175
rect 26495 -9295 26540 -9175
rect 26660 -9295 26705 -9175
rect 26825 -9295 26880 -9175
rect 27000 -9295 27045 -9175
rect 27165 -9295 27210 -9175
rect 27330 -9295 27375 -9175
rect 27495 -9295 27550 -9175
rect 27670 -9295 27715 -9175
rect 27835 -9295 27880 -9175
rect 28000 -9295 28045 -9175
rect 28165 -9295 28220 -9175
rect 28340 -9295 28385 -9175
rect 28505 -9295 28550 -9175
rect 28670 -9295 28715 -9175
rect 28835 -9295 28890 -9175
rect 29010 -9295 29055 -9175
rect 29175 -9295 29220 -9175
rect 29340 -9295 29385 -9175
rect 29505 -9295 29560 -9175
rect 29680 -9295 29705 -9175
rect 24175 -9340 29705 -9295
rect 24175 -9460 24200 -9340
rect 24320 -9460 24365 -9340
rect 24485 -9460 24530 -9340
rect 24650 -9460 24695 -9340
rect 24815 -9460 24870 -9340
rect 24990 -9460 25035 -9340
rect 25155 -9460 25200 -9340
rect 25320 -9460 25365 -9340
rect 25485 -9460 25540 -9340
rect 25660 -9460 25705 -9340
rect 25825 -9460 25870 -9340
rect 25990 -9460 26035 -9340
rect 26155 -9460 26210 -9340
rect 26330 -9460 26375 -9340
rect 26495 -9460 26540 -9340
rect 26660 -9460 26705 -9340
rect 26825 -9460 26880 -9340
rect 27000 -9460 27045 -9340
rect 27165 -9460 27210 -9340
rect 27330 -9460 27375 -9340
rect 27495 -9460 27550 -9340
rect 27670 -9460 27715 -9340
rect 27835 -9460 27880 -9340
rect 28000 -9460 28045 -9340
rect 28165 -9460 28220 -9340
rect 28340 -9460 28385 -9340
rect 28505 -9460 28550 -9340
rect 28670 -9460 28715 -9340
rect 28835 -9460 28890 -9340
rect 29010 -9460 29055 -9340
rect 29175 -9460 29220 -9340
rect 29340 -9460 29385 -9340
rect 29505 -9460 29560 -9340
rect 29680 -9460 29705 -9340
rect 24175 -9505 29705 -9460
rect 24175 -9625 24200 -9505
rect 24320 -9625 24365 -9505
rect 24485 -9625 24530 -9505
rect 24650 -9625 24695 -9505
rect 24815 -9625 24870 -9505
rect 24990 -9625 25035 -9505
rect 25155 -9625 25200 -9505
rect 25320 -9625 25365 -9505
rect 25485 -9625 25540 -9505
rect 25660 -9625 25705 -9505
rect 25825 -9625 25870 -9505
rect 25990 -9625 26035 -9505
rect 26155 -9625 26210 -9505
rect 26330 -9625 26375 -9505
rect 26495 -9625 26540 -9505
rect 26660 -9625 26705 -9505
rect 26825 -9625 26880 -9505
rect 27000 -9625 27045 -9505
rect 27165 -9625 27210 -9505
rect 27330 -9625 27375 -9505
rect 27495 -9625 27550 -9505
rect 27670 -9625 27715 -9505
rect 27835 -9625 27880 -9505
rect 28000 -9625 28045 -9505
rect 28165 -9625 28220 -9505
rect 28340 -9625 28385 -9505
rect 28505 -9625 28550 -9505
rect 28670 -9625 28715 -9505
rect 28835 -9625 28890 -9505
rect 29010 -9625 29055 -9505
rect 29175 -9625 29220 -9505
rect 29340 -9625 29385 -9505
rect 29505 -9625 29560 -9505
rect 29680 -9625 29705 -9505
rect 24175 -9670 29705 -9625
rect 24175 -9790 24200 -9670
rect 24320 -9790 24365 -9670
rect 24485 -9790 24530 -9670
rect 24650 -9790 24695 -9670
rect 24815 -9790 24870 -9670
rect 24990 -9790 25035 -9670
rect 25155 -9790 25200 -9670
rect 25320 -9790 25365 -9670
rect 25485 -9790 25540 -9670
rect 25660 -9790 25705 -9670
rect 25825 -9790 25870 -9670
rect 25990 -9790 26035 -9670
rect 26155 -9790 26210 -9670
rect 26330 -9790 26375 -9670
rect 26495 -9790 26540 -9670
rect 26660 -9790 26705 -9670
rect 26825 -9790 26880 -9670
rect 27000 -9790 27045 -9670
rect 27165 -9790 27210 -9670
rect 27330 -9790 27375 -9670
rect 27495 -9790 27550 -9670
rect 27670 -9790 27715 -9670
rect 27835 -9790 27880 -9670
rect 28000 -9790 28045 -9670
rect 28165 -9790 28220 -9670
rect 28340 -9790 28385 -9670
rect 28505 -9790 28550 -9670
rect 28670 -9790 28715 -9670
rect 28835 -9790 28890 -9670
rect 29010 -9790 29055 -9670
rect 29175 -9790 29220 -9670
rect 29340 -9790 29385 -9670
rect 29505 -9790 29560 -9670
rect 29680 -9790 29705 -9670
rect 24175 -9815 29705 -9790
rect 12635 -9865 12795 -9860
rect 18325 -9865 18485 -9860
rect 24015 -9865 24175 -9860
rect 7105 -9880 29705 -9865
rect 7105 -10000 7170 -9880
rect 7290 -10000 7335 -9880
rect 7455 -10000 7500 -9880
rect 7620 -10000 7665 -9880
rect 7785 -10000 7830 -9880
rect 7950 -10000 7995 -9880
rect 8115 -10000 8160 -9880
rect 8280 -10000 8325 -9880
rect 8445 -10000 8490 -9880
rect 8610 -10000 8655 -9880
rect 8775 -10000 8820 -9880
rect 8940 -10000 8985 -9880
rect 9105 -10000 9150 -9880
rect 9270 -10000 9315 -9880
rect 9435 -10000 9480 -9880
rect 9600 -10000 9645 -9880
rect 9765 -10000 9810 -9880
rect 9930 -10000 9975 -9880
rect 10095 -10000 10140 -9880
rect 10260 -10000 10305 -9880
rect 10425 -10000 10470 -9880
rect 10590 -10000 10635 -9880
rect 10755 -10000 10800 -9880
rect 10920 -10000 10965 -9880
rect 11085 -10000 11130 -9880
rect 11250 -10000 11295 -9880
rect 11415 -10000 11460 -9880
rect 11580 -10000 11625 -9880
rect 11745 -10000 11790 -9880
rect 11910 -10000 11955 -9880
rect 12075 -10000 12120 -9880
rect 12240 -10000 12285 -9880
rect 12405 -10000 12450 -9880
rect 12570 -10000 12860 -9880
rect 12980 -10000 13025 -9880
rect 13145 -10000 13190 -9880
rect 13310 -10000 13355 -9880
rect 13475 -10000 13520 -9880
rect 13640 -10000 13685 -9880
rect 13805 -10000 13850 -9880
rect 13970 -10000 14015 -9880
rect 14135 -10000 14180 -9880
rect 14300 -10000 14345 -9880
rect 14465 -10000 14510 -9880
rect 14630 -10000 14675 -9880
rect 14795 -10000 14840 -9880
rect 14960 -10000 15005 -9880
rect 15125 -10000 15170 -9880
rect 15290 -10000 15335 -9880
rect 15455 -10000 15500 -9880
rect 15620 -10000 15665 -9880
rect 15785 -10000 15830 -9880
rect 15950 -10000 15995 -9880
rect 16115 -10000 16160 -9880
rect 16280 -10000 16325 -9880
rect 16445 -10000 16490 -9880
rect 16610 -10000 16655 -9880
rect 16775 -10000 16820 -9880
rect 16940 -10000 16985 -9880
rect 17105 -10000 17150 -9880
rect 17270 -10000 17315 -9880
rect 17435 -10000 17480 -9880
rect 17600 -10000 17645 -9880
rect 17765 -10000 17810 -9880
rect 17930 -10000 17975 -9880
rect 18095 -10000 18140 -9880
rect 18260 -10000 18550 -9880
rect 18670 -10000 18715 -9880
rect 18835 -10000 18880 -9880
rect 19000 -10000 19045 -9880
rect 19165 -10000 19210 -9880
rect 19330 -10000 19375 -9880
rect 19495 -10000 19540 -9880
rect 19660 -10000 19705 -9880
rect 19825 -10000 19870 -9880
rect 19990 -10000 20035 -9880
rect 20155 -10000 20200 -9880
rect 20320 -10000 20365 -9880
rect 20485 -10000 20530 -9880
rect 20650 -10000 20695 -9880
rect 20815 -10000 20860 -9880
rect 20980 -10000 21025 -9880
rect 21145 -10000 21190 -9880
rect 21310 -10000 21355 -9880
rect 21475 -10000 21520 -9880
rect 21640 -10000 21685 -9880
rect 21805 -10000 21850 -9880
rect 21970 -10000 22015 -9880
rect 22135 -10000 22180 -9880
rect 22300 -10000 22345 -9880
rect 22465 -10000 22510 -9880
rect 22630 -10000 22675 -9880
rect 22795 -10000 22840 -9880
rect 22960 -10000 23005 -9880
rect 23125 -10000 23170 -9880
rect 23290 -10000 23335 -9880
rect 23455 -10000 23500 -9880
rect 23620 -10000 23665 -9880
rect 23785 -10000 23830 -9880
rect 23950 -10000 24240 -9880
rect 24360 -10000 24405 -9880
rect 24525 -10000 24570 -9880
rect 24690 -10000 24735 -9880
rect 24855 -10000 24900 -9880
rect 25020 -10000 25065 -9880
rect 25185 -10000 25230 -9880
rect 25350 -10000 25395 -9880
rect 25515 -10000 25560 -9880
rect 25680 -10000 25725 -9880
rect 25845 -10000 25890 -9880
rect 26010 -10000 26055 -9880
rect 26175 -10000 26220 -9880
rect 26340 -10000 26385 -9880
rect 26505 -10000 26550 -9880
rect 26670 -10000 26715 -9880
rect 26835 -10000 26880 -9880
rect 27000 -10000 27045 -9880
rect 27165 -10000 27210 -9880
rect 27330 -10000 27375 -9880
rect 27495 -10000 27540 -9880
rect 27660 -10000 27705 -9880
rect 27825 -10000 27870 -9880
rect 27990 -10000 28035 -9880
rect 28155 -10000 28200 -9880
rect 28320 -10000 28365 -9880
rect 28485 -10000 28530 -9880
rect 28650 -10000 28695 -9880
rect 28815 -10000 28860 -9880
rect 28980 -10000 29025 -9880
rect 29145 -10000 29190 -9880
rect 29310 -10000 29355 -9880
rect 29475 -10000 29520 -9880
rect 29640 -10000 29705 -9880
rect 7105 -10015 29705 -10000
rect 12635 -10020 12795 -10015
rect 18325 -10020 18485 -10015
rect 24015 -10020 24175 -10015
rect 7105 -10090 12635 -10065
rect 7105 -10210 7130 -10090
rect 7250 -10210 7305 -10090
rect 7425 -10210 7470 -10090
rect 7590 -10210 7635 -10090
rect 7755 -10210 7800 -10090
rect 7920 -10210 7975 -10090
rect 8095 -10210 8140 -10090
rect 8260 -10210 8305 -10090
rect 8425 -10210 8470 -10090
rect 8590 -10210 8645 -10090
rect 8765 -10210 8810 -10090
rect 8930 -10210 8975 -10090
rect 9095 -10210 9140 -10090
rect 9260 -10210 9315 -10090
rect 9435 -10210 9480 -10090
rect 9600 -10210 9645 -10090
rect 9765 -10210 9810 -10090
rect 9930 -10210 9985 -10090
rect 10105 -10210 10150 -10090
rect 10270 -10210 10315 -10090
rect 10435 -10210 10480 -10090
rect 10600 -10210 10655 -10090
rect 10775 -10210 10820 -10090
rect 10940 -10210 10985 -10090
rect 11105 -10210 11150 -10090
rect 11270 -10210 11325 -10090
rect 11445 -10210 11490 -10090
rect 11610 -10210 11655 -10090
rect 11775 -10210 11820 -10090
rect 11940 -10210 11995 -10090
rect 12115 -10210 12160 -10090
rect 12280 -10210 12325 -10090
rect 12445 -10210 12490 -10090
rect 12610 -10210 12635 -10090
rect 7105 -10255 12635 -10210
rect 7105 -10375 7130 -10255
rect 7250 -10375 7305 -10255
rect 7425 -10375 7470 -10255
rect 7590 -10375 7635 -10255
rect 7755 -10375 7800 -10255
rect 7920 -10375 7975 -10255
rect 8095 -10375 8140 -10255
rect 8260 -10375 8305 -10255
rect 8425 -10375 8470 -10255
rect 8590 -10375 8645 -10255
rect 8765 -10375 8810 -10255
rect 8930 -10375 8975 -10255
rect 9095 -10375 9140 -10255
rect 9260 -10375 9315 -10255
rect 9435 -10375 9480 -10255
rect 9600 -10375 9645 -10255
rect 9765 -10375 9810 -10255
rect 9930 -10375 9985 -10255
rect 10105 -10375 10150 -10255
rect 10270 -10375 10315 -10255
rect 10435 -10375 10480 -10255
rect 10600 -10375 10655 -10255
rect 10775 -10375 10820 -10255
rect 10940 -10375 10985 -10255
rect 11105 -10375 11150 -10255
rect 11270 -10375 11325 -10255
rect 11445 -10375 11490 -10255
rect 11610 -10375 11655 -10255
rect 11775 -10375 11820 -10255
rect 11940 -10375 11995 -10255
rect 12115 -10375 12160 -10255
rect 12280 -10375 12325 -10255
rect 12445 -10375 12490 -10255
rect 12610 -10375 12635 -10255
rect 7105 -10420 12635 -10375
rect 7105 -10540 7130 -10420
rect 7250 -10540 7305 -10420
rect 7425 -10540 7470 -10420
rect 7590 -10540 7635 -10420
rect 7755 -10540 7800 -10420
rect 7920 -10540 7975 -10420
rect 8095 -10540 8140 -10420
rect 8260 -10540 8305 -10420
rect 8425 -10540 8470 -10420
rect 8590 -10540 8645 -10420
rect 8765 -10540 8810 -10420
rect 8930 -10540 8975 -10420
rect 9095 -10540 9140 -10420
rect 9260 -10540 9315 -10420
rect 9435 -10540 9480 -10420
rect 9600 -10540 9645 -10420
rect 9765 -10540 9810 -10420
rect 9930 -10540 9985 -10420
rect 10105 -10540 10150 -10420
rect 10270 -10540 10315 -10420
rect 10435 -10540 10480 -10420
rect 10600 -10540 10655 -10420
rect 10775 -10540 10820 -10420
rect 10940 -10540 10985 -10420
rect 11105 -10540 11150 -10420
rect 11270 -10540 11325 -10420
rect 11445 -10540 11490 -10420
rect 11610 -10540 11655 -10420
rect 11775 -10540 11820 -10420
rect 11940 -10540 11995 -10420
rect 12115 -10540 12160 -10420
rect 12280 -10540 12325 -10420
rect 12445 -10540 12490 -10420
rect 12610 -10540 12635 -10420
rect 7105 -10585 12635 -10540
rect 7105 -10705 7130 -10585
rect 7250 -10705 7305 -10585
rect 7425 -10705 7470 -10585
rect 7590 -10705 7635 -10585
rect 7755 -10705 7800 -10585
rect 7920 -10705 7975 -10585
rect 8095 -10705 8140 -10585
rect 8260 -10705 8305 -10585
rect 8425 -10705 8470 -10585
rect 8590 -10705 8645 -10585
rect 8765 -10705 8810 -10585
rect 8930 -10705 8975 -10585
rect 9095 -10705 9140 -10585
rect 9260 -10705 9315 -10585
rect 9435 -10705 9480 -10585
rect 9600 -10705 9645 -10585
rect 9765 -10705 9810 -10585
rect 9930 -10705 9985 -10585
rect 10105 -10705 10150 -10585
rect 10270 -10705 10315 -10585
rect 10435 -10705 10480 -10585
rect 10600 -10705 10655 -10585
rect 10775 -10705 10820 -10585
rect 10940 -10705 10985 -10585
rect 11105 -10705 11150 -10585
rect 11270 -10705 11325 -10585
rect 11445 -10705 11490 -10585
rect 11610 -10705 11655 -10585
rect 11775 -10705 11820 -10585
rect 11940 -10705 11995 -10585
rect 12115 -10705 12160 -10585
rect 12280 -10705 12325 -10585
rect 12445 -10705 12490 -10585
rect 12610 -10705 12635 -10585
rect 7105 -10760 12635 -10705
rect 7105 -10880 7130 -10760
rect 7250 -10880 7305 -10760
rect 7425 -10880 7470 -10760
rect 7590 -10880 7635 -10760
rect 7755 -10880 7800 -10760
rect 7920 -10880 7975 -10760
rect 8095 -10880 8140 -10760
rect 8260 -10880 8305 -10760
rect 8425 -10880 8470 -10760
rect 8590 -10880 8645 -10760
rect 8765 -10880 8810 -10760
rect 8930 -10880 8975 -10760
rect 9095 -10880 9140 -10760
rect 9260 -10880 9315 -10760
rect 9435 -10880 9480 -10760
rect 9600 -10880 9645 -10760
rect 9765 -10880 9810 -10760
rect 9930 -10880 9985 -10760
rect 10105 -10880 10150 -10760
rect 10270 -10880 10315 -10760
rect 10435 -10880 10480 -10760
rect 10600 -10880 10655 -10760
rect 10775 -10880 10820 -10760
rect 10940 -10880 10985 -10760
rect 11105 -10880 11150 -10760
rect 11270 -10880 11325 -10760
rect 11445 -10880 11490 -10760
rect 11610 -10880 11655 -10760
rect 11775 -10880 11820 -10760
rect 11940 -10880 11995 -10760
rect 12115 -10880 12160 -10760
rect 12280 -10880 12325 -10760
rect 12445 -10880 12490 -10760
rect 12610 -10880 12635 -10760
rect 7105 -10925 12635 -10880
rect 7105 -11045 7130 -10925
rect 7250 -11045 7305 -10925
rect 7425 -11045 7470 -10925
rect 7590 -11045 7635 -10925
rect 7755 -11045 7800 -10925
rect 7920 -11045 7975 -10925
rect 8095 -11045 8140 -10925
rect 8260 -11045 8305 -10925
rect 8425 -11045 8470 -10925
rect 8590 -11045 8645 -10925
rect 8765 -11045 8810 -10925
rect 8930 -11045 8975 -10925
rect 9095 -11045 9140 -10925
rect 9260 -11045 9315 -10925
rect 9435 -11045 9480 -10925
rect 9600 -11045 9645 -10925
rect 9765 -11045 9810 -10925
rect 9930 -11045 9985 -10925
rect 10105 -11045 10150 -10925
rect 10270 -11045 10315 -10925
rect 10435 -11045 10480 -10925
rect 10600 -11045 10655 -10925
rect 10775 -11045 10820 -10925
rect 10940 -11045 10985 -10925
rect 11105 -11045 11150 -10925
rect 11270 -11045 11325 -10925
rect 11445 -11045 11490 -10925
rect 11610 -11045 11655 -10925
rect 11775 -11045 11820 -10925
rect 11940 -11045 11995 -10925
rect 12115 -11045 12160 -10925
rect 12280 -11045 12325 -10925
rect 12445 -11045 12490 -10925
rect 12610 -11045 12635 -10925
rect 7105 -11090 12635 -11045
rect 7105 -11210 7130 -11090
rect 7250 -11210 7305 -11090
rect 7425 -11210 7470 -11090
rect 7590 -11210 7635 -11090
rect 7755 -11210 7800 -11090
rect 7920 -11210 7975 -11090
rect 8095 -11210 8140 -11090
rect 8260 -11210 8305 -11090
rect 8425 -11210 8470 -11090
rect 8590 -11210 8645 -11090
rect 8765 -11210 8810 -11090
rect 8930 -11210 8975 -11090
rect 9095 -11210 9140 -11090
rect 9260 -11210 9315 -11090
rect 9435 -11210 9480 -11090
rect 9600 -11210 9645 -11090
rect 9765 -11210 9810 -11090
rect 9930 -11210 9985 -11090
rect 10105 -11210 10150 -11090
rect 10270 -11210 10315 -11090
rect 10435 -11210 10480 -11090
rect 10600 -11210 10655 -11090
rect 10775 -11210 10820 -11090
rect 10940 -11210 10985 -11090
rect 11105 -11210 11150 -11090
rect 11270 -11210 11325 -11090
rect 11445 -11210 11490 -11090
rect 11610 -11210 11655 -11090
rect 11775 -11210 11820 -11090
rect 11940 -11210 11995 -11090
rect 12115 -11210 12160 -11090
rect 12280 -11210 12325 -11090
rect 12445 -11210 12490 -11090
rect 12610 -11210 12635 -11090
rect 7105 -11255 12635 -11210
rect 7105 -11375 7130 -11255
rect 7250 -11375 7305 -11255
rect 7425 -11375 7470 -11255
rect 7590 -11375 7635 -11255
rect 7755 -11375 7800 -11255
rect 7920 -11375 7975 -11255
rect 8095 -11375 8140 -11255
rect 8260 -11375 8305 -11255
rect 8425 -11375 8470 -11255
rect 8590 -11375 8645 -11255
rect 8765 -11375 8810 -11255
rect 8930 -11375 8975 -11255
rect 9095 -11375 9140 -11255
rect 9260 -11375 9315 -11255
rect 9435 -11375 9480 -11255
rect 9600 -11375 9645 -11255
rect 9765 -11375 9810 -11255
rect 9930 -11375 9985 -11255
rect 10105 -11375 10150 -11255
rect 10270 -11375 10315 -11255
rect 10435 -11375 10480 -11255
rect 10600 -11375 10655 -11255
rect 10775 -11375 10820 -11255
rect 10940 -11375 10985 -11255
rect 11105 -11375 11150 -11255
rect 11270 -11375 11325 -11255
rect 11445 -11375 11490 -11255
rect 11610 -11375 11655 -11255
rect 11775 -11375 11820 -11255
rect 11940 -11375 11995 -11255
rect 12115 -11375 12160 -11255
rect 12280 -11375 12325 -11255
rect 12445 -11375 12490 -11255
rect 12610 -11375 12635 -11255
rect 7105 -11430 12635 -11375
rect 7105 -11550 7130 -11430
rect 7250 -11550 7305 -11430
rect 7425 -11550 7470 -11430
rect 7590 -11550 7635 -11430
rect 7755 -11550 7800 -11430
rect 7920 -11550 7975 -11430
rect 8095 -11550 8140 -11430
rect 8260 -11550 8305 -11430
rect 8425 -11550 8470 -11430
rect 8590 -11550 8645 -11430
rect 8765 -11550 8810 -11430
rect 8930 -11550 8975 -11430
rect 9095 -11550 9140 -11430
rect 9260 -11550 9315 -11430
rect 9435 -11550 9480 -11430
rect 9600 -11550 9645 -11430
rect 9765 -11550 9810 -11430
rect 9930 -11550 9985 -11430
rect 10105 -11550 10150 -11430
rect 10270 -11550 10315 -11430
rect 10435 -11550 10480 -11430
rect 10600 -11550 10655 -11430
rect 10775 -11550 10820 -11430
rect 10940 -11550 10985 -11430
rect 11105 -11550 11150 -11430
rect 11270 -11550 11325 -11430
rect 11445 -11550 11490 -11430
rect 11610 -11550 11655 -11430
rect 11775 -11550 11820 -11430
rect 11940 -11550 11995 -11430
rect 12115 -11550 12160 -11430
rect 12280 -11550 12325 -11430
rect 12445 -11550 12490 -11430
rect 12610 -11550 12635 -11430
rect 7105 -11595 12635 -11550
rect 7105 -11715 7130 -11595
rect 7250 -11715 7305 -11595
rect 7425 -11715 7470 -11595
rect 7590 -11715 7635 -11595
rect 7755 -11715 7800 -11595
rect 7920 -11715 7975 -11595
rect 8095 -11715 8140 -11595
rect 8260 -11715 8305 -11595
rect 8425 -11715 8470 -11595
rect 8590 -11715 8645 -11595
rect 8765 -11715 8810 -11595
rect 8930 -11715 8975 -11595
rect 9095 -11715 9140 -11595
rect 9260 -11715 9315 -11595
rect 9435 -11715 9480 -11595
rect 9600 -11715 9645 -11595
rect 9765 -11715 9810 -11595
rect 9930 -11715 9985 -11595
rect 10105 -11715 10150 -11595
rect 10270 -11715 10315 -11595
rect 10435 -11715 10480 -11595
rect 10600 -11715 10655 -11595
rect 10775 -11715 10820 -11595
rect 10940 -11715 10985 -11595
rect 11105 -11715 11150 -11595
rect 11270 -11715 11325 -11595
rect 11445 -11715 11490 -11595
rect 11610 -11715 11655 -11595
rect 11775 -11715 11820 -11595
rect 11940 -11715 11995 -11595
rect 12115 -11715 12160 -11595
rect 12280 -11715 12325 -11595
rect 12445 -11715 12490 -11595
rect 12610 -11715 12635 -11595
rect 7105 -11760 12635 -11715
rect 7105 -11880 7130 -11760
rect 7250 -11880 7305 -11760
rect 7425 -11880 7470 -11760
rect 7590 -11880 7635 -11760
rect 7755 -11880 7800 -11760
rect 7920 -11880 7975 -11760
rect 8095 -11880 8140 -11760
rect 8260 -11880 8305 -11760
rect 8425 -11880 8470 -11760
rect 8590 -11880 8645 -11760
rect 8765 -11880 8810 -11760
rect 8930 -11880 8975 -11760
rect 9095 -11880 9140 -11760
rect 9260 -11880 9315 -11760
rect 9435 -11880 9480 -11760
rect 9600 -11880 9645 -11760
rect 9765 -11880 9810 -11760
rect 9930 -11880 9985 -11760
rect 10105 -11880 10150 -11760
rect 10270 -11880 10315 -11760
rect 10435 -11880 10480 -11760
rect 10600 -11880 10655 -11760
rect 10775 -11880 10820 -11760
rect 10940 -11880 10985 -11760
rect 11105 -11880 11150 -11760
rect 11270 -11880 11325 -11760
rect 11445 -11880 11490 -11760
rect 11610 -11880 11655 -11760
rect 11775 -11880 11820 -11760
rect 11940 -11880 11995 -11760
rect 12115 -11880 12160 -11760
rect 12280 -11880 12325 -11760
rect 12445 -11880 12490 -11760
rect 12610 -11880 12635 -11760
rect 7105 -11925 12635 -11880
rect 7105 -12045 7130 -11925
rect 7250 -12045 7305 -11925
rect 7425 -12045 7470 -11925
rect 7590 -12045 7635 -11925
rect 7755 -12045 7800 -11925
rect 7920 -12045 7975 -11925
rect 8095 -12045 8140 -11925
rect 8260 -12045 8305 -11925
rect 8425 -12045 8470 -11925
rect 8590 -12045 8645 -11925
rect 8765 -12045 8810 -11925
rect 8930 -12045 8975 -11925
rect 9095 -12045 9140 -11925
rect 9260 -12045 9315 -11925
rect 9435 -12045 9480 -11925
rect 9600 -12045 9645 -11925
rect 9765 -12045 9810 -11925
rect 9930 -12045 9985 -11925
rect 10105 -12045 10150 -11925
rect 10270 -12045 10315 -11925
rect 10435 -12045 10480 -11925
rect 10600 -12045 10655 -11925
rect 10775 -12045 10820 -11925
rect 10940 -12045 10985 -11925
rect 11105 -12045 11150 -11925
rect 11270 -12045 11325 -11925
rect 11445 -12045 11490 -11925
rect 11610 -12045 11655 -11925
rect 11775 -12045 11820 -11925
rect 11940 -12045 11995 -11925
rect 12115 -12045 12160 -11925
rect 12280 -12045 12325 -11925
rect 12445 -12045 12490 -11925
rect 12610 -12045 12635 -11925
rect 7105 -12100 12635 -12045
rect 7105 -12220 7130 -12100
rect 7250 -12220 7305 -12100
rect 7425 -12220 7470 -12100
rect 7590 -12220 7635 -12100
rect 7755 -12220 7800 -12100
rect 7920 -12220 7975 -12100
rect 8095 -12220 8140 -12100
rect 8260 -12220 8305 -12100
rect 8425 -12220 8470 -12100
rect 8590 -12220 8645 -12100
rect 8765 -12220 8810 -12100
rect 8930 -12220 8975 -12100
rect 9095 -12220 9140 -12100
rect 9260 -12220 9315 -12100
rect 9435 -12220 9480 -12100
rect 9600 -12220 9645 -12100
rect 9765 -12220 9810 -12100
rect 9930 -12220 9985 -12100
rect 10105 -12220 10150 -12100
rect 10270 -12220 10315 -12100
rect 10435 -12220 10480 -12100
rect 10600 -12220 10655 -12100
rect 10775 -12220 10820 -12100
rect 10940 -12220 10985 -12100
rect 11105 -12220 11150 -12100
rect 11270 -12220 11325 -12100
rect 11445 -12220 11490 -12100
rect 11610 -12220 11655 -12100
rect 11775 -12220 11820 -12100
rect 11940 -12220 11995 -12100
rect 12115 -12220 12160 -12100
rect 12280 -12220 12325 -12100
rect 12445 -12220 12490 -12100
rect 12610 -12220 12635 -12100
rect 7105 -12265 12635 -12220
rect 7105 -12385 7130 -12265
rect 7250 -12385 7305 -12265
rect 7425 -12385 7470 -12265
rect 7590 -12385 7635 -12265
rect 7755 -12385 7800 -12265
rect 7920 -12385 7975 -12265
rect 8095 -12385 8140 -12265
rect 8260 -12385 8305 -12265
rect 8425 -12385 8470 -12265
rect 8590 -12385 8645 -12265
rect 8765 -12385 8810 -12265
rect 8930 -12385 8975 -12265
rect 9095 -12385 9140 -12265
rect 9260 -12385 9315 -12265
rect 9435 -12385 9480 -12265
rect 9600 -12385 9645 -12265
rect 9765 -12385 9810 -12265
rect 9930 -12385 9985 -12265
rect 10105 -12385 10150 -12265
rect 10270 -12385 10315 -12265
rect 10435 -12385 10480 -12265
rect 10600 -12385 10655 -12265
rect 10775 -12385 10820 -12265
rect 10940 -12385 10985 -12265
rect 11105 -12385 11150 -12265
rect 11270 -12385 11325 -12265
rect 11445 -12385 11490 -12265
rect 11610 -12385 11655 -12265
rect 11775 -12385 11820 -12265
rect 11940 -12385 11995 -12265
rect 12115 -12385 12160 -12265
rect 12280 -12385 12325 -12265
rect 12445 -12385 12490 -12265
rect 12610 -12385 12635 -12265
rect 7105 -12430 12635 -12385
rect 7105 -12550 7130 -12430
rect 7250 -12550 7305 -12430
rect 7425 -12550 7470 -12430
rect 7590 -12550 7635 -12430
rect 7755 -12550 7800 -12430
rect 7920 -12550 7975 -12430
rect 8095 -12550 8140 -12430
rect 8260 -12550 8305 -12430
rect 8425 -12550 8470 -12430
rect 8590 -12550 8645 -12430
rect 8765 -12550 8810 -12430
rect 8930 -12550 8975 -12430
rect 9095 -12550 9140 -12430
rect 9260 -12550 9315 -12430
rect 9435 -12550 9480 -12430
rect 9600 -12550 9645 -12430
rect 9765 -12550 9810 -12430
rect 9930 -12550 9985 -12430
rect 10105 -12550 10150 -12430
rect 10270 -12550 10315 -12430
rect 10435 -12550 10480 -12430
rect 10600 -12550 10655 -12430
rect 10775 -12550 10820 -12430
rect 10940 -12550 10985 -12430
rect 11105 -12550 11150 -12430
rect 11270 -12550 11325 -12430
rect 11445 -12550 11490 -12430
rect 11610 -12550 11655 -12430
rect 11775 -12550 11820 -12430
rect 11940 -12550 11995 -12430
rect 12115 -12550 12160 -12430
rect 12280 -12550 12325 -12430
rect 12445 -12550 12490 -12430
rect 12610 -12550 12635 -12430
rect 7105 -12595 12635 -12550
rect 7105 -12715 7130 -12595
rect 7250 -12715 7305 -12595
rect 7425 -12715 7470 -12595
rect 7590 -12715 7635 -12595
rect 7755 -12715 7800 -12595
rect 7920 -12715 7975 -12595
rect 8095 -12715 8140 -12595
rect 8260 -12715 8305 -12595
rect 8425 -12715 8470 -12595
rect 8590 -12715 8645 -12595
rect 8765 -12715 8810 -12595
rect 8930 -12715 8975 -12595
rect 9095 -12715 9140 -12595
rect 9260 -12715 9315 -12595
rect 9435 -12715 9480 -12595
rect 9600 -12715 9645 -12595
rect 9765 -12715 9810 -12595
rect 9930 -12715 9985 -12595
rect 10105 -12715 10150 -12595
rect 10270 -12715 10315 -12595
rect 10435 -12715 10480 -12595
rect 10600 -12715 10655 -12595
rect 10775 -12715 10820 -12595
rect 10940 -12715 10985 -12595
rect 11105 -12715 11150 -12595
rect 11270 -12715 11325 -12595
rect 11445 -12715 11490 -12595
rect 11610 -12715 11655 -12595
rect 11775 -12715 11820 -12595
rect 11940 -12715 11995 -12595
rect 12115 -12715 12160 -12595
rect 12280 -12715 12325 -12595
rect 12445 -12715 12490 -12595
rect 12610 -12715 12635 -12595
rect 7105 -12770 12635 -12715
rect 7105 -12890 7130 -12770
rect 7250 -12890 7305 -12770
rect 7425 -12890 7470 -12770
rect 7590 -12890 7635 -12770
rect 7755 -12890 7800 -12770
rect 7920 -12890 7975 -12770
rect 8095 -12890 8140 -12770
rect 8260 -12890 8305 -12770
rect 8425 -12890 8470 -12770
rect 8590 -12890 8645 -12770
rect 8765 -12890 8810 -12770
rect 8930 -12890 8975 -12770
rect 9095 -12890 9140 -12770
rect 9260 -12890 9315 -12770
rect 9435 -12890 9480 -12770
rect 9600 -12890 9645 -12770
rect 9765 -12890 9810 -12770
rect 9930 -12890 9985 -12770
rect 10105 -12890 10150 -12770
rect 10270 -12890 10315 -12770
rect 10435 -12890 10480 -12770
rect 10600 -12890 10655 -12770
rect 10775 -12890 10820 -12770
rect 10940 -12890 10985 -12770
rect 11105 -12890 11150 -12770
rect 11270 -12890 11325 -12770
rect 11445 -12890 11490 -12770
rect 11610 -12890 11655 -12770
rect 11775 -12890 11820 -12770
rect 11940 -12890 11995 -12770
rect 12115 -12890 12160 -12770
rect 12280 -12890 12325 -12770
rect 12445 -12890 12490 -12770
rect 12610 -12890 12635 -12770
rect 7105 -12935 12635 -12890
rect 7105 -13055 7130 -12935
rect 7250 -13055 7305 -12935
rect 7425 -13055 7470 -12935
rect 7590 -13055 7635 -12935
rect 7755 -13055 7800 -12935
rect 7920 -13055 7975 -12935
rect 8095 -13055 8140 -12935
rect 8260 -13055 8305 -12935
rect 8425 -13055 8470 -12935
rect 8590 -13055 8645 -12935
rect 8765 -13055 8810 -12935
rect 8930 -13055 8975 -12935
rect 9095 -13055 9140 -12935
rect 9260 -13055 9315 -12935
rect 9435 -13055 9480 -12935
rect 9600 -13055 9645 -12935
rect 9765 -13055 9810 -12935
rect 9930 -13055 9985 -12935
rect 10105 -13055 10150 -12935
rect 10270 -13055 10315 -12935
rect 10435 -13055 10480 -12935
rect 10600 -13055 10655 -12935
rect 10775 -13055 10820 -12935
rect 10940 -13055 10985 -12935
rect 11105 -13055 11150 -12935
rect 11270 -13055 11325 -12935
rect 11445 -13055 11490 -12935
rect 11610 -13055 11655 -12935
rect 11775 -13055 11820 -12935
rect 11940 -13055 11995 -12935
rect 12115 -13055 12160 -12935
rect 12280 -13055 12325 -12935
rect 12445 -13055 12490 -12935
rect 12610 -13055 12635 -12935
rect 7105 -13100 12635 -13055
rect 7105 -13220 7130 -13100
rect 7250 -13220 7305 -13100
rect 7425 -13220 7470 -13100
rect 7590 -13220 7635 -13100
rect 7755 -13220 7800 -13100
rect 7920 -13220 7975 -13100
rect 8095 -13220 8140 -13100
rect 8260 -13220 8305 -13100
rect 8425 -13220 8470 -13100
rect 8590 -13220 8645 -13100
rect 8765 -13220 8810 -13100
rect 8930 -13220 8975 -13100
rect 9095 -13220 9140 -13100
rect 9260 -13220 9315 -13100
rect 9435 -13220 9480 -13100
rect 9600 -13220 9645 -13100
rect 9765 -13220 9810 -13100
rect 9930 -13220 9985 -13100
rect 10105 -13220 10150 -13100
rect 10270 -13220 10315 -13100
rect 10435 -13220 10480 -13100
rect 10600 -13220 10655 -13100
rect 10775 -13220 10820 -13100
rect 10940 -13220 10985 -13100
rect 11105 -13220 11150 -13100
rect 11270 -13220 11325 -13100
rect 11445 -13220 11490 -13100
rect 11610 -13220 11655 -13100
rect 11775 -13220 11820 -13100
rect 11940 -13220 11995 -13100
rect 12115 -13220 12160 -13100
rect 12280 -13220 12325 -13100
rect 12445 -13220 12490 -13100
rect 12610 -13220 12635 -13100
rect 7105 -13265 12635 -13220
rect 7105 -13385 7130 -13265
rect 7250 -13385 7305 -13265
rect 7425 -13385 7470 -13265
rect 7590 -13385 7635 -13265
rect 7755 -13385 7800 -13265
rect 7920 -13385 7975 -13265
rect 8095 -13385 8140 -13265
rect 8260 -13385 8305 -13265
rect 8425 -13385 8470 -13265
rect 8590 -13385 8645 -13265
rect 8765 -13385 8810 -13265
rect 8930 -13385 8975 -13265
rect 9095 -13385 9140 -13265
rect 9260 -13385 9315 -13265
rect 9435 -13385 9480 -13265
rect 9600 -13385 9645 -13265
rect 9765 -13385 9810 -13265
rect 9930 -13385 9985 -13265
rect 10105 -13385 10150 -13265
rect 10270 -13385 10315 -13265
rect 10435 -13385 10480 -13265
rect 10600 -13385 10655 -13265
rect 10775 -13385 10820 -13265
rect 10940 -13385 10985 -13265
rect 11105 -13385 11150 -13265
rect 11270 -13385 11325 -13265
rect 11445 -13385 11490 -13265
rect 11610 -13385 11655 -13265
rect 11775 -13385 11820 -13265
rect 11940 -13385 11995 -13265
rect 12115 -13385 12160 -13265
rect 12280 -13385 12325 -13265
rect 12445 -13385 12490 -13265
rect 12610 -13385 12635 -13265
rect 7105 -13440 12635 -13385
rect 7105 -13560 7130 -13440
rect 7250 -13560 7305 -13440
rect 7425 -13560 7470 -13440
rect 7590 -13560 7635 -13440
rect 7755 -13560 7800 -13440
rect 7920 -13560 7975 -13440
rect 8095 -13560 8140 -13440
rect 8260 -13560 8305 -13440
rect 8425 -13560 8470 -13440
rect 8590 -13560 8645 -13440
rect 8765 -13560 8810 -13440
rect 8930 -13560 8975 -13440
rect 9095 -13560 9140 -13440
rect 9260 -13560 9315 -13440
rect 9435 -13560 9480 -13440
rect 9600 -13560 9645 -13440
rect 9765 -13560 9810 -13440
rect 9930 -13560 9985 -13440
rect 10105 -13560 10150 -13440
rect 10270 -13560 10315 -13440
rect 10435 -13560 10480 -13440
rect 10600 -13560 10655 -13440
rect 10775 -13560 10820 -13440
rect 10940 -13560 10985 -13440
rect 11105 -13560 11150 -13440
rect 11270 -13560 11325 -13440
rect 11445 -13560 11490 -13440
rect 11610 -13560 11655 -13440
rect 11775 -13560 11820 -13440
rect 11940 -13560 11995 -13440
rect 12115 -13560 12160 -13440
rect 12280 -13560 12325 -13440
rect 12445 -13560 12490 -13440
rect 12610 -13560 12635 -13440
rect 7105 -13605 12635 -13560
rect 7105 -13725 7130 -13605
rect 7250 -13725 7305 -13605
rect 7425 -13725 7470 -13605
rect 7590 -13725 7635 -13605
rect 7755 -13725 7800 -13605
rect 7920 -13725 7975 -13605
rect 8095 -13725 8140 -13605
rect 8260 -13725 8305 -13605
rect 8425 -13725 8470 -13605
rect 8590 -13725 8645 -13605
rect 8765 -13725 8810 -13605
rect 8930 -13725 8975 -13605
rect 9095 -13725 9140 -13605
rect 9260 -13725 9315 -13605
rect 9435 -13725 9480 -13605
rect 9600 -13725 9645 -13605
rect 9765 -13725 9810 -13605
rect 9930 -13725 9985 -13605
rect 10105 -13725 10150 -13605
rect 10270 -13725 10315 -13605
rect 10435 -13725 10480 -13605
rect 10600 -13725 10655 -13605
rect 10775 -13725 10820 -13605
rect 10940 -13725 10985 -13605
rect 11105 -13725 11150 -13605
rect 11270 -13725 11325 -13605
rect 11445 -13725 11490 -13605
rect 11610 -13725 11655 -13605
rect 11775 -13725 11820 -13605
rect 11940 -13725 11995 -13605
rect 12115 -13725 12160 -13605
rect 12280 -13725 12325 -13605
rect 12445 -13725 12490 -13605
rect 12610 -13725 12635 -13605
rect 7105 -13770 12635 -13725
rect 7105 -13890 7130 -13770
rect 7250 -13890 7305 -13770
rect 7425 -13890 7470 -13770
rect 7590 -13890 7635 -13770
rect 7755 -13890 7800 -13770
rect 7920 -13890 7975 -13770
rect 8095 -13890 8140 -13770
rect 8260 -13890 8305 -13770
rect 8425 -13890 8470 -13770
rect 8590 -13890 8645 -13770
rect 8765 -13890 8810 -13770
rect 8930 -13890 8975 -13770
rect 9095 -13890 9140 -13770
rect 9260 -13890 9315 -13770
rect 9435 -13890 9480 -13770
rect 9600 -13890 9645 -13770
rect 9765 -13890 9810 -13770
rect 9930 -13890 9985 -13770
rect 10105 -13890 10150 -13770
rect 10270 -13890 10315 -13770
rect 10435 -13890 10480 -13770
rect 10600 -13890 10655 -13770
rect 10775 -13890 10820 -13770
rect 10940 -13890 10985 -13770
rect 11105 -13890 11150 -13770
rect 11270 -13890 11325 -13770
rect 11445 -13890 11490 -13770
rect 11610 -13890 11655 -13770
rect 11775 -13890 11820 -13770
rect 11940 -13890 11995 -13770
rect 12115 -13890 12160 -13770
rect 12280 -13890 12325 -13770
rect 12445 -13890 12490 -13770
rect 12610 -13890 12635 -13770
rect 7105 -13935 12635 -13890
rect 7105 -14055 7130 -13935
rect 7250 -14055 7305 -13935
rect 7425 -14055 7470 -13935
rect 7590 -14055 7635 -13935
rect 7755 -14055 7800 -13935
rect 7920 -14055 7975 -13935
rect 8095 -14055 8140 -13935
rect 8260 -14055 8305 -13935
rect 8425 -14055 8470 -13935
rect 8590 -14055 8645 -13935
rect 8765 -14055 8810 -13935
rect 8930 -14055 8975 -13935
rect 9095 -14055 9140 -13935
rect 9260 -14055 9315 -13935
rect 9435 -14055 9480 -13935
rect 9600 -14055 9645 -13935
rect 9765 -14055 9810 -13935
rect 9930 -14055 9985 -13935
rect 10105 -14055 10150 -13935
rect 10270 -14055 10315 -13935
rect 10435 -14055 10480 -13935
rect 10600 -14055 10655 -13935
rect 10775 -14055 10820 -13935
rect 10940 -14055 10985 -13935
rect 11105 -14055 11150 -13935
rect 11270 -14055 11325 -13935
rect 11445 -14055 11490 -13935
rect 11610 -14055 11655 -13935
rect 11775 -14055 11820 -13935
rect 11940 -14055 11995 -13935
rect 12115 -14055 12160 -13935
rect 12280 -14055 12325 -13935
rect 12445 -14055 12490 -13935
rect 12610 -14055 12635 -13935
rect 7105 -14110 12635 -14055
rect 7105 -14230 7130 -14110
rect 7250 -14230 7305 -14110
rect 7425 -14230 7470 -14110
rect 7590 -14230 7635 -14110
rect 7755 -14230 7800 -14110
rect 7920 -14230 7975 -14110
rect 8095 -14230 8140 -14110
rect 8260 -14230 8305 -14110
rect 8425 -14230 8470 -14110
rect 8590 -14230 8645 -14110
rect 8765 -14230 8810 -14110
rect 8930 -14230 8975 -14110
rect 9095 -14230 9140 -14110
rect 9260 -14230 9315 -14110
rect 9435 -14230 9480 -14110
rect 9600 -14230 9645 -14110
rect 9765 -14230 9810 -14110
rect 9930 -14230 9985 -14110
rect 10105 -14230 10150 -14110
rect 10270 -14230 10315 -14110
rect 10435 -14230 10480 -14110
rect 10600 -14230 10655 -14110
rect 10775 -14230 10820 -14110
rect 10940 -14230 10985 -14110
rect 11105 -14230 11150 -14110
rect 11270 -14230 11325 -14110
rect 11445 -14230 11490 -14110
rect 11610 -14230 11655 -14110
rect 11775 -14230 11820 -14110
rect 11940 -14230 11995 -14110
rect 12115 -14230 12160 -14110
rect 12280 -14230 12325 -14110
rect 12445 -14230 12490 -14110
rect 12610 -14230 12635 -14110
rect 7105 -14275 12635 -14230
rect 7105 -14395 7130 -14275
rect 7250 -14395 7305 -14275
rect 7425 -14395 7470 -14275
rect 7590 -14395 7635 -14275
rect 7755 -14395 7800 -14275
rect 7920 -14395 7975 -14275
rect 8095 -14395 8140 -14275
rect 8260 -14395 8305 -14275
rect 8425 -14395 8470 -14275
rect 8590 -14395 8645 -14275
rect 8765 -14395 8810 -14275
rect 8930 -14395 8975 -14275
rect 9095 -14395 9140 -14275
rect 9260 -14395 9315 -14275
rect 9435 -14395 9480 -14275
rect 9600 -14395 9645 -14275
rect 9765 -14395 9810 -14275
rect 9930 -14395 9985 -14275
rect 10105 -14395 10150 -14275
rect 10270 -14395 10315 -14275
rect 10435 -14395 10480 -14275
rect 10600 -14395 10655 -14275
rect 10775 -14395 10820 -14275
rect 10940 -14395 10985 -14275
rect 11105 -14395 11150 -14275
rect 11270 -14395 11325 -14275
rect 11445 -14395 11490 -14275
rect 11610 -14395 11655 -14275
rect 11775 -14395 11820 -14275
rect 11940 -14395 11995 -14275
rect 12115 -14395 12160 -14275
rect 12280 -14395 12325 -14275
rect 12445 -14395 12490 -14275
rect 12610 -14395 12635 -14275
rect 7105 -14440 12635 -14395
rect 7105 -14560 7130 -14440
rect 7250 -14560 7305 -14440
rect 7425 -14560 7470 -14440
rect 7590 -14560 7635 -14440
rect 7755 -14560 7800 -14440
rect 7920 -14560 7975 -14440
rect 8095 -14560 8140 -14440
rect 8260 -14560 8305 -14440
rect 8425 -14560 8470 -14440
rect 8590 -14560 8645 -14440
rect 8765 -14560 8810 -14440
rect 8930 -14560 8975 -14440
rect 9095 -14560 9140 -14440
rect 9260 -14560 9315 -14440
rect 9435 -14560 9480 -14440
rect 9600 -14560 9645 -14440
rect 9765 -14560 9810 -14440
rect 9930 -14560 9985 -14440
rect 10105 -14560 10150 -14440
rect 10270 -14560 10315 -14440
rect 10435 -14560 10480 -14440
rect 10600 -14560 10655 -14440
rect 10775 -14560 10820 -14440
rect 10940 -14560 10985 -14440
rect 11105 -14560 11150 -14440
rect 11270 -14560 11325 -14440
rect 11445 -14560 11490 -14440
rect 11610 -14560 11655 -14440
rect 11775 -14560 11820 -14440
rect 11940 -14560 11995 -14440
rect 12115 -14560 12160 -14440
rect 12280 -14560 12325 -14440
rect 12445 -14560 12490 -14440
rect 12610 -14560 12635 -14440
rect 7105 -14605 12635 -14560
rect 7105 -14725 7130 -14605
rect 7250 -14725 7305 -14605
rect 7425 -14725 7470 -14605
rect 7590 -14725 7635 -14605
rect 7755 -14725 7800 -14605
rect 7920 -14725 7975 -14605
rect 8095 -14725 8140 -14605
rect 8260 -14725 8305 -14605
rect 8425 -14725 8470 -14605
rect 8590 -14725 8645 -14605
rect 8765 -14725 8810 -14605
rect 8930 -14725 8975 -14605
rect 9095 -14725 9140 -14605
rect 9260 -14725 9315 -14605
rect 9435 -14725 9480 -14605
rect 9600 -14725 9645 -14605
rect 9765 -14725 9810 -14605
rect 9930 -14725 9985 -14605
rect 10105 -14725 10150 -14605
rect 10270 -14725 10315 -14605
rect 10435 -14725 10480 -14605
rect 10600 -14725 10655 -14605
rect 10775 -14725 10820 -14605
rect 10940 -14725 10985 -14605
rect 11105 -14725 11150 -14605
rect 11270 -14725 11325 -14605
rect 11445 -14725 11490 -14605
rect 11610 -14725 11655 -14605
rect 11775 -14725 11820 -14605
rect 11940 -14725 11995 -14605
rect 12115 -14725 12160 -14605
rect 12280 -14725 12325 -14605
rect 12445 -14725 12490 -14605
rect 12610 -14725 12635 -14605
rect 7105 -14780 12635 -14725
rect 7105 -14900 7130 -14780
rect 7250 -14900 7305 -14780
rect 7425 -14900 7470 -14780
rect 7590 -14900 7635 -14780
rect 7755 -14900 7800 -14780
rect 7920 -14900 7975 -14780
rect 8095 -14900 8140 -14780
rect 8260 -14900 8305 -14780
rect 8425 -14900 8470 -14780
rect 8590 -14900 8645 -14780
rect 8765 -14900 8810 -14780
rect 8930 -14900 8975 -14780
rect 9095 -14900 9140 -14780
rect 9260 -14900 9315 -14780
rect 9435 -14900 9480 -14780
rect 9600 -14900 9645 -14780
rect 9765 -14900 9810 -14780
rect 9930 -14900 9985 -14780
rect 10105 -14900 10150 -14780
rect 10270 -14900 10315 -14780
rect 10435 -14900 10480 -14780
rect 10600 -14900 10655 -14780
rect 10775 -14900 10820 -14780
rect 10940 -14900 10985 -14780
rect 11105 -14900 11150 -14780
rect 11270 -14900 11325 -14780
rect 11445 -14900 11490 -14780
rect 11610 -14900 11655 -14780
rect 11775 -14900 11820 -14780
rect 11940 -14900 11995 -14780
rect 12115 -14900 12160 -14780
rect 12280 -14900 12325 -14780
rect 12445 -14900 12490 -14780
rect 12610 -14900 12635 -14780
rect 7105 -14945 12635 -14900
rect 7105 -15065 7130 -14945
rect 7250 -15065 7305 -14945
rect 7425 -15065 7470 -14945
rect 7590 -15065 7635 -14945
rect 7755 -15065 7800 -14945
rect 7920 -15065 7975 -14945
rect 8095 -15065 8140 -14945
rect 8260 -15065 8305 -14945
rect 8425 -15065 8470 -14945
rect 8590 -15065 8645 -14945
rect 8765 -15065 8810 -14945
rect 8930 -15065 8975 -14945
rect 9095 -15065 9140 -14945
rect 9260 -15065 9315 -14945
rect 9435 -15065 9480 -14945
rect 9600 -15065 9645 -14945
rect 9765 -15065 9810 -14945
rect 9930 -15065 9985 -14945
rect 10105 -15065 10150 -14945
rect 10270 -15065 10315 -14945
rect 10435 -15065 10480 -14945
rect 10600 -15065 10655 -14945
rect 10775 -15065 10820 -14945
rect 10940 -15065 10985 -14945
rect 11105 -15065 11150 -14945
rect 11270 -15065 11325 -14945
rect 11445 -15065 11490 -14945
rect 11610 -15065 11655 -14945
rect 11775 -15065 11820 -14945
rect 11940 -15065 11995 -14945
rect 12115 -15065 12160 -14945
rect 12280 -15065 12325 -14945
rect 12445 -15065 12490 -14945
rect 12610 -15065 12635 -14945
rect 7105 -15110 12635 -15065
rect 7105 -15230 7130 -15110
rect 7250 -15230 7305 -15110
rect 7425 -15230 7470 -15110
rect 7590 -15230 7635 -15110
rect 7755 -15230 7800 -15110
rect 7920 -15230 7975 -15110
rect 8095 -15230 8140 -15110
rect 8260 -15230 8305 -15110
rect 8425 -15230 8470 -15110
rect 8590 -15230 8645 -15110
rect 8765 -15230 8810 -15110
rect 8930 -15230 8975 -15110
rect 9095 -15230 9140 -15110
rect 9260 -15230 9315 -15110
rect 9435 -15230 9480 -15110
rect 9600 -15230 9645 -15110
rect 9765 -15230 9810 -15110
rect 9930 -15230 9985 -15110
rect 10105 -15230 10150 -15110
rect 10270 -15230 10315 -15110
rect 10435 -15230 10480 -15110
rect 10600 -15230 10655 -15110
rect 10775 -15230 10820 -15110
rect 10940 -15230 10985 -15110
rect 11105 -15230 11150 -15110
rect 11270 -15230 11325 -15110
rect 11445 -15230 11490 -15110
rect 11610 -15230 11655 -15110
rect 11775 -15230 11820 -15110
rect 11940 -15230 11995 -15110
rect 12115 -15230 12160 -15110
rect 12280 -15230 12325 -15110
rect 12445 -15230 12490 -15110
rect 12610 -15230 12635 -15110
rect 7105 -15275 12635 -15230
rect 7105 -15395 7130 -15275
rect 7250 -15395 7305 -15275
rect 7425 -15395 7470 -15275
rect 7590 -15395 7635 -15275
rect 7755 -15395 7800 -15275
rect 7920 -15395 7975 -15275
rect 8095 -15395 8140 -15275
rect 8260 -15395 8305 -15275
rect 8425 -15395 8470 -15275
rect 8590 -15395 8645 -15275
rect 8765 -15395 8810 -15275
rect 8930 -15395 8975 -15275
rect 9095 -15395 9140 -15275
rect 9260 -15395 9315 -15275
rect 9435 -15395 9480 -15275
rect 9600 -15395 9645 -15275
rect 9765 -15395 9810 -15275
rect 9930 -15395 9985 -15275
rect 10105 -15395 10150 -15275
rect 10270 -15395 10315 -15275
rect 10435 -15395 10480 -15275
rect 10600 -15395 10655 -15275
rect 10775 -15395 10820 -15275
rect 10940 -15395 10985 -15275
rect 11105 -15395 11150 -15275
rect 11270 -15395 11325 -15275
rect 11445 -15395 11490 -15275
rect 11610 -15395 11655 -15275
rect 11775 -15395 11820 -15275
rect 11940 -15395 11995 -15275
rect 12115 -15395 12160 -15275
rect 12280 -15395 12325 -15275
rect 12445 -15395 12490 -15275
rect 12610 -15395 12635 -15275
rect 7105 -15450 12635 -15395
rect 7105 -15570 7130 -15450
rect 7250 -15570 7305 -15450
rect 7425 -15570 7470 -15450
rect 7590 -15570 7635 -15450
rect 7755 -15570 7800 -15450
rect 7920 -15570 7975 -15450
rect 8095 -15570 8140 -15450
rect 8260 -15570 8305 -15450
rect 8425 -15570 8470 -15450
rect 8590 -15570 8645 -15450
rect 8765 -15570 8810 -15450
rect 8930 -15570 8975 -15450
rect 9095 -15570 9140 -15450
rect 9260 -15570 9315 -15450
rect 9435 -15570 9480 -15450
rect 9600 -15570 9645 -15450
rect 9765 -15570 9810 -15450
rect 9930 -15570 9985 -15450
rect 10105 -15570 10150 -15450
rect 10270 -15570 10315 -15450
rect 10435 -15570 10480 -15450
rect 10600 -15570 10655 -15450
rect 10775 -15570 10820 -15450
rect 10940 -15570 10985 -15450
rect 11105 -15570 11150 -15450
rect 11270 -15570 11325 -15450
rect 11445 -15570 11490 -15450
rect 11610 -15570 11655 -15450
rect 11775 -15570 11820 -15450
rect 11940 -15570 11995 -15450
rect 12115 -15570 12160 -15450
rect 12280 -15570 12325 -15450
rect 12445 -15570 12490 -15450
rect 12610 -15535 12635 -15450
rect 12795 -10090 18325 -10065
rect 12795 -10210 12820 -10090
rect 12940 -10210 12995 -10090
rect 13115 -10210 13160 -10090
rect 13280 -10210 13325 -10090
rect 13445 -10210 13490 -10090
rect 13610 -10210 13665 -10090
rect 13785 -10210 13830 -10090
rect 13950 -10210 13995 -10090
rect 14115 -10210 14160 -10090
rect 14280 -10210 14335 -10090
rect 14455 -10210 14500 -10090
rect 14620 -10210 14665 -10090
rect 14785 -10210 14830 -10090
rect 14950 -10210 15005 -10090
rect 15125 -10210 15170 -10090
rect 15290 -10210 15335 -10090
rect 15455 -10210 15500 -10090
rect 15620 -10210 15675 -10090
rect 15795 -10210 15840 -10090
rect 15960 -10210 16005 -10090
rect 16125 -10210 16170 -10090
rect 16290 -10210 16345 -10090
rect 16465 -10210 16510 -10090
rect 16630 -10210 16675 -10090
rect 16795 -10210 16840 -10090
rect 16960 -10210 17015 -10090
rect 17135 -10210 17180 -10090
rect 17300 -10210 17345 -10090
rect 17465 -10210 17510 -10090
rect 17630 -10210 17685 -10090
rect 17805 -10210 17850 -10090
rect 17970 -10210 18015 -10090
rect 18135 -10210 18180 -10090
rect 18300 -10210 18325 -10090
rect 12795 -10255 18325 -10210
rect 12795 -10375 12820 -10255
rect 12940 -10375 12995 -10255
rect 13115 -10375 13160 -10255
rect 13280 -10375 13325 -10255
rect 13445 -10375 13490 -10255
rect 13610 -10375 13665 -10255
rect 13785 -10375 13830 -10255
rect 13950 -10375 13995 -10255
rect 14115 -10375 14160 -10255
rect 14280 -10375 14335 -10255
rect 14455 -10375 14500 -10255
rect 14620 -10375 14665 -10255
rect 14785 -10375 14830 -10255
rect 14950 -10375 15005 -10255
rect 15125 -10375 15170 -10255
rect 15290 -10375 15335 -10255
rect 15455 -10375 15500 -10255
rect 15620 -10375 15675 -10255
rect 15795 -10375 15840 -10255
rect 15960 -10375 16005 -10255
rect 16125 -10375 16170 -10255
rect 16290 -10375 16345 -10255
rect 16465 -10375 16510 -10255
rect 16630 -10375 16675 -10255
rect 16795 -10375 16840 -10255
rect 16960 -10375 17015 -10255
rect 17135 -10375 17180 -10255
rect 17300 -10375 17345 -10255
rect 17465 -10375 17510 -10255
rect 17630 -10375 17685 -10255
rect 17805 -10375 17850 -10255
rect 17970 -10375 18015 -10255
rect 18135 -10375 18180 -10255
rect 18300 -10375 18325 -10255
rect 12795 -10420 18325 -10375
rect 12795 -10540 12820 -10420
rect 12940 -10540 12995 -10420
rect 13115 -10540 13160 -10420
rect 13280 -10540 13325 -10420
rect 13445 -10540 13490 -10420
rect 13610 -10540 13665 -10420
rect 13785 -10540 13830 -10420
rect 13950 -10540 13995 -10420
rect 14115 -10540 14160 -10420
rect 14280 -10540 14335 -10420
rect 14455 -10540 14500 -10420
rect 14620 -10540 14665 -10420
rect 14785 -10540 14830 -10420
rect 14950 -10540 15005 -10420
rect 15125 -10540 15170 -10420
rect 15290 -10540 15335 -10420
rect 15455 -10540 15500 -10420
rect 15620 -10540 15675 -10420
rect 15795 -10540 15840 -10420
rect 15960 -10540 16005 -10420
rect 16125 -10540 16170 -10420
rect 16290 -10540 16345 -10420
rect 16465 -10540 16510 -10420
rect 16630 -10540 16675 -10420
rect 16795 -10540 16840 -10420
rect 16960 -10540 17015 -10420
rect 17135 -10540 17180 -10420
rect 17300 -10540 17345 -10420
rect 17465 -10540 17510 -10420
rect 17630 -10540 17685 -10420
rect 17805 -10540 17850 -10420
rect 17970 -10540 18015 -10420
rect 18135 -10540 18180 -10420
rect 18300 -10540 18325 -10420
rect 12795 -10585 18325 -10540
rect 12795 -10705 12820 -10585
rect 12940 -10705 12995 -10585
rect 13115 -10705 13160 -10585
rect 13280 -10705 13325 -10585
rect 13445 -10705 13490 -10585
rect 13610 -10705 13665 -10585
rect 13785 -10705 13830 -10585
rect 13950 -10705 13995 -10585
rect 14115 -10705 14160 -10585
rect 14280 -10705 14335 -10585
rect 14455 -10705 14500 -10585
rect 14620 -10705 14665 -10585
rect 14785 -10705 14830 -10585
rect 14950 -10705 15005 -10585
rect 15125 -10705 15170 -10585
rect 15290 -10705 15335 -10585
rect 15455 -10705 15500 -10585
rect 15620 -10705 15675 -10585
rect 15795 -10705 15840 -10585
rect 15960 -10705 16005 -10585
rect 16125 -10705 16170 -10585
rect 16290 -10705 16345 -10585
rect 16465 -10705 16510 -10585
rect 16630 -10705 16675 -10585
rect 16795 -10705 16840 -10585
rect 16960 -10705 17015 -10585
rect 17135 -10705 17180 -10585
rect 17300 -10705 17345 -10585
rect 17465 -10705 17510 -10585
rect 17630 -10705 17685 -10585
rect 17805 -10705 17850 -10585
rect 17970 -10705 18015 -10585
rect 18135 -10705 18180 -10585
rect 18300 -10705 18325 -10585
rect 12795 -10760 18325 -10705
rect 12795 -10880 12820 -10760
rect 12940 -10880 12995 -10760
rect 13115 -10880 13160 -10760
rect 13280 -10880 13325 -10760
rect 13445 -10880 13490 -10760
rect 13610 -10880 13665 -10760
rect 13785 -10880 13830 -10760
rect 13950 -10880 13995 -10760
rect 14115 -10880 14160 -10760
rect 14280 -10880 14335 -10760
rect 14455 -10880 14500 -10760
rect 14620 -10880 14665 -10760
rect 14785 -10880 14830 -10760
rect 14950 -10880 15005 -10760
rect 15125 -10880 15170 -10760
rect 15290 -10880 15335 -10760
rect 15455 -10880 15500 -10760
rect 15620 -10880 15675 -10760
rect 15795 -10880 15840 -10760
rect 15960 -10880 16005 -10760
rect 16125 -10880 16170 -10760
rect 16290 -10880 16345 -10760
rect 16465 -10880 16510 -10760
rect 16630 -10880 16675 -10760
rect 16795 -10880 16840 -10760
rect 16960 -10880 17015 -10760
rect 17135 -10880 17180 -10760
rect 17300 -10880 17345 -10760
rect 17465 -10880 17510 -10760
rect 17630 -10880 17685 -10760
rect 17805 -10880 17850 -10760
rect 17970 -10880 18015 -10760
rect 18135 -10880 18180 -10760
rect 18300 -10880 18325 -10760
rect 12795 -10925 18325 -10880
rect 12795 -11045 12820 -10925
rect 12940 -11045 12995 -10925
rect 13115 -11045 13160 -10925
rect 13280 -11045 13325 -10925
rect 13445 -11045 13490 -10925
rect 13610 -11045 13665 -10925
rect 13785 -11045 13830 -10925
rect 13950 -11045 13995 -10925
rect 14115 -11045 14160 -10925
rect 14280 -11045 14335 -10925
rect 14455 -11045 14500 -10925
rect 14620 -11045 14665 -10925
rect 14785 -11045 14830 -10925
rect 14950 -11045 15005 -10925
rect 15125 -11045 15170 -10925
rect 15290 -11045 15335 -10925
rect 15455 -11045 15500 -10925
rect 15620 -11045 15675 -10925
rect 15795 -11045 15840 -10925
rect 15960 -11045 16005 -10925
rect 16125 -11045 16170 -10925
rect 16290 -11045 16345 -10925
rect 16465 -11045 16510 -10925
rect 16630 -11045 16675 -10925
rect 16795 -11045 16840 -10925
rect 16960 -11045 17015 -10925
rect 17135 -11045 17180 -10925
rect 17300 -11045 17345 -10925
rect 17465 -11045 17510 -10925
rect 17630 -11045 17685 -10925
rect 17805 -11045 17850 -10925
rect 17970 -11045 18015 -10925
rect 18135 -11045 18180 -10925
rect 18300 -11045 18325 -10925
rect 12795 -11090 18325 -11045
rect 12795 -11210 12820 -11090
rect 12940 -11210 12995 -11090
rect 13115 -11210 13160 -11090
rect 13280 -11210 13325 -11090
rect 13445 -11210 13490 -11090
rect 13610 -11210 13665 -11090
rect 13785 -11210 13830 -11090
rect 13950 -11210 13995 -11090
rect 14115 -11210 14160 -11090
rect 14280 -11210 14335 -11090
rect 14455 -11210 14500 -11090
rect 14620 -11210 14665 -11090
rect 14785 -11210 14830 -11090
rect 14950 -11210 15005 -11090
rect 15125 -11210 15170 -11090
rect 15290 -11210 15335 -11090
rect 15455 -11210 15500 -11090
rect 15620 -11210 15675 -11090
rect 15795 -11210 15840 -11090
rect 15960 -11210 16005 -11090
rect 16125 -11210 16170 -11090
rect 16290 -11210 16345 -11090
rect 16465 -11210 16510 -11090
rect 16630 -11210 16675 -11090
rect 16795 -11210 16840 -11090
rect 16960 -11210 17015 -11090
rect 17135 -11210 17180 -11090
rect 17300 -11210 17345 -11090
rect 17465 -11210 17510 -11090
rect 17630 -11210 17685 -11090
rect 17805 -11210 17850 -11090
rect 17970 -11210 18015 -11090
rect 18135 -11210 18180 -11090
rect 18300 -11210 18325 -11090
rect 12795 -11255 18325 -11210
rect 12795 -11375 12820 -11255
rect 12940 -11375 12995 -11255
rect 13115 -11375 13160 -11255
rect 13280 -11375 13325 -11255
rect 13445 -11375 13490 -11255
rect 13610 -11375 13665 -11255
rect 13785 -11375 13830 -11255
rect 13950 -11375 13995 -11255
rect 14115 -11375 14160 -11255
rect 14280 -11375 14335 -11255
rect 14455 -11375 14500 -11255
rect 14620 -11375 14665 -11255
rect 14785 -11375 14830 -11255
rect 14950 -11375 15005 -11255
rect 15125 -11375 15170 -11255
rect 15290 -11375 15335 -11255
rect 15455 -11375 15500 -11255
rect 15620 -11375 15675 -11255
rect 15795 -11375 15840 -11255
rect 15960 -11375 16005 -11255
rect 16125 -11375 16170 -11255
rect 16290 -11375 16345 -11255
rect 16465 -11375 16510 -11255
rect 16630 -11375 16675 -11255
rect 16795 -11375 16840 -11255
rect 16960 -11375 17015 -11255
rect 17135 -11375 17180 -11255
rect 17300 -11375 17345 -11255
rect 17465 -11375 17510 -11255
rect 17630 -11375 17685 -11255
rect 17805 -11375 17850 -11255
rect 17970 -11375 18015 -11255
rect 18135 -11375 18180 -11255
rect 18300 -11375 18325 -11255
rect 12795 -11430 18325 -11375
rect 12795 -11550 12820 -11430
rect 12940 -11550 12995 -11430
rect 13115 -11550 13160 -11430
rect 13280 -11550 13325 -11430
rect 13445 -11550 13490 -11430
rect 13610 -11550 13665 -11430
rect 13785 -11550 13830 -11430
rect 13950 -11550 13995 -11430
rect 14115 -11550 14160 -11430
rect 14280 -11550 14335 -11430
rect 14455 -11550 14500 -11430
rect 14620 -11550 14665 -11430
rect 14785 -11550 14830 -11430
rect 14950 -11550 15005 -11430
rect 15125 -11550 15170 -11430
rect 15290 -11550 15335 -11430
rect 15455 -11550 15500 -11430
rect 15620 -11550 15675 -11430
rect 15795 -11550 15840 -11430
rect 15960 -11550 16005 -11430
rect 16125 -11550 16170 -11430
rect 16290 -11550 16345 -11430
rect 16465 -11550 16510 -11430
rect 16630 -11550 16675 -11430
rect 16795 -11550 16840 -11430
rect 16960 -11550 17015 -11430
rect 17135 -11550 17180 -11430
rect 17300 -11550 17345 -11430
rect 17465 -11550 17510 -11430
rect 17630 -11550 17685 -11430
rect 17805 -11550 17850 -11430
rect 17970 -11550 18015 -11430
rect 18135 -11550 18180 -11430
rect 18300 -11550 18325 -11430
rect 12795 -11595 18325 -11550
rect 12795 -11715 12820 -11595
rect 12940 -11715 12995 -11595
rect 13115 -11715 13160 -11595
rect 13280 -11715 13325 -11595
rect 13445 -11715 13490 -11595
rect 13610 -11715 13665 -11595
rect 13785 -11715 13830 -11595
rect 13950 -11715 13995 -11595
rect 14115 -11715 14160 -11595
rect 14280 -11715 14335 -11595
rect 14455 -11715 14500 -11595
rect 14620 -11715 14665 -11595
rect 14785 -11715 14830 -11595
rect 14950 -11715 15005 -11595
rect 15125 -11715 15170 -11595
rect 15290 -11715 15335 -11595
rect 15455 -11715 15500 -11595
rect 15620 -11715 15675 -11595
rect 15795 -11715 15840 -11595
rect 15960 -11715 16005 -11595
rect 16125 -11715 16170 -11595
rect 16290 -11715 16345 -11595
rect 16465 -11715 16510 -11595
rect 16630 -11715 16675 -11595
rect 16795 -11715 16840 -11595
rect 16960 -11715 17015 -11595
rect 17135 -11715 17180 -11595
rect 17300 -11715 17345 -11595
rect 17465 -11715 17510 -11595
rect 17630 -11715 17685 -11595
rect 17805 -11715 17850 -11595
rect 17970 -11715 18015 -11595
rect 18135 -11715 18180 -11595
rect 18300 -11715 18325 -11595
rect 12795 -11760 18325 -11715
rect 12795 -11880 12820 -11760
rect 12940 -11880 12995 -11760
rect 13115 -11880 13160 -11760
rect 13280 -11880 13325 -11760
rect 13445 -11880 13490 -11760
rect 13610 -11880 13665 -11760
rect 13785 -11880 13830 -11760
rect 13950 -11880 13995 -11760
rect 14115 -11880 14160 -11760
rect 14280 -11880 14335 -11760
rect 14455 -11880 14500 -11760
rect 14620 -11880 14665 -11760
rect 14785 -11880 14830 -11760
rect 14950 -11880 15005 -11760
rect 15125 -11880 15170 -11760
rect 15290 -11880 15335 -11760
rect 15455 -11880 15500 -11760
rect 15620 -11880 15675 -11760
rect 15795 -11880 15840 -11760
rect 15960 -11880 16005 -11760
rect 16125 -11880 16170 -11760
rect 16290 -11880 16345 -11760
rect 16465 -11880 16510 -11760
rect 16630 -11880 16675 -11760
rect 16795 -11880 16840 -11760
rect 16960 -11880 17015 -11760
rect 17135 -11880 17180 -11760
rect 17300 -11880 17345 -11760
rect 17465 -11880 17510 -11760
rect 17630 -11880 17685 -11760
rect 17805 -11880 17850 -11760
rect 17970 -11880 18015 -11760
rect 18135 -11880 18180 -11760
rect 18300 -11880 18325 -11760
rect 12795 -11925 18325 -11880
rect 12795 -12045 12820 -11925
rect 12940 -12045 12995 -11925
rect 13115 -12045 13160 -11925
rect 13280 -12045 13325 -11925
rect 13445 -12045 13490 -11925
rect 13610 -12045 13665 -11925
rect 13785 -12045 13830 -11925
rect 13950 -12045 13995 -11925
rect 14115 -12045 14160 -11925
rect 14280 -12045 14335 -11925
rect 14455 -12045 14500 -11925
rect 14620 -12045 14665 -11925
rect 14785 -12045 14830 -11925
rect 14950 -12045 15005 -11925
rect 15125 -12045 15170 -11925
rect 15290 -12045 15335 -11925
rect 15455 -12045 15500 -11925
rect 15620 -12045 15675 -11925
rect 15795 -12045 15840 -11925
rect 15960 -12045 16005 -11925
rect 16125 -12045 16170 -11925
rect 16290 -12045 16345 -11925
rect 16465 -12045 16510 -11925
rect 16630 -12045 16675 -11925
rect 16795 -12045 16840 -11925
rect 16960 -12045 17015 -11925
rect 17135 -12045 17180 -11925
rect 17300 -12045 17345 -11925
rect 17465 -12045 17510 -11925
rect 17630 -12045 17685 -11925
rect 17805 -12045 17850 -11925
rect 17970 -12045 18015 -11925
rect 18135 -12045 18180 -11925
rect 18300 -12045 18325 -11925
rect 12795 -12100 18325 -12045
rect 12795 -12220 12820 -12100
rect 12940 -12220 12995 -12100
rect 13115 -12220 13160 -12100
rect 13280 -12220 13325 -12100
rect 13445 -12220 13490 -12100
rect 13610 -12220 13665 -12100
rect 13785 -12220 13830 -12100
rect 13950 -12220 13995 -12100
rect 14115 -12220 14160 -12100
rect 14280 -12220 14335 -12100
rect 14455 -12220 14500 -12100
rect 14620 -12220 14665 -12100
rect 14785 -12220 14830 -12100
rect 14950 -12220 15005 -12100
rect 15125 -12220 15170 -12100
rect 15290 -12220 15335 -12100
rect 15455 -12220 15500 -12100
rect 15620 -12220 15675 -12100
rect 15795 -12220 15840 -12100
rect 15960 -12220 16005 -12100
rect 16125 -12220 16170 -12100
rect 16290 -12220 16345 -12100
rect 16465 -12220 16510 -12100
rect 16630 -12220 16675 -12100
rect 16795 -12220 16840 -12100
rect 16960 -12220 17015 -12100
rect 17135 -12220 17180 -12100
rect 17300 -12220 17345 -12100
rect 17465 -12220 17510 -12100
rect 17630 -12220 17685 -12100
rect 17805 -12220 17850 -12100
rect 17970 -12220 18015 -12100
rect 18135 -12220 18180 -12100
rect 18300 -12220 18325 -12100
rect 12795 -12265 18325 -12220
rect 12795 -12385 12820 -12265
rect 12940 -12385 12995 -12265
rect 13115 -12385 13160 -12265
rect 13280 -12385 13325 -12265
rect 13445 -12385 13490 -12265
rect 13610 -12385 13665 -12265
rect 13785 -12385 13830 -12265
rect 13950 -12385 13995 -12265
rect 14115 -12385 14160 -12265
rect 14280 -12385 14335 -12265
rect 14455 -12385 14500 -12265
rect 14620 -12385 14665 -12265
rect 14785 -12385 14830 -12265
rect 14950 -12385 15005 -12265
rect 15125 -12385 15170 -12265
rect 15290 -12385 15335 -12265
rect 15455 -12385 15500 -12265
rect 15620 -12385 15675 -12265
rect 15795 -12385 15840 -12265
rect 15960 -12385 16005 -12265
rect 16125 -12385 16170 -12265
rect 16290 -12385 16345 -12265
rect 16465 -12385 16510 -12265
rect 16630 -12385 16675 -12265
rect 16795 -12385 16840 -12265
rect 16960 -12385 17015 -12265
rect 17135 -12385 17180 -12265
rect 17300 -12385 17345 -12265
rect 17465 -12385 17510 -12265
rect 17630 -12385 17685 -12265
rect 17805 -12385 17850 -12265
rect 17970 -12385 18015 -12265
rect 18135 -12385 18180 -12265
rect 18300 -12385 18325 -12265
rect 12795 -12430 18325 -12385
rect 12795 -12550 12820 -12430
rect 12940 -12550 12995 -12430
rect 13115 -12550 13160 -12430
rect 13280 -12550 13325 -12430
rect 13445 -12550 13490 -12430
rect 13610 -12550 13665 -12430
rect 13785 -12550 13830 -12430
rect 13950 -12550 13995 -12430
rect 14115 -12550 14160 -12430
rect 14280 -12550 14335 -12430
rect 14455 -12550 14500 -12430
rect 14620 -12550 14665 -12430
rect 14785 -12550 14830 -12430
rect 14950 -12550 15005 -12430
rect 15125 -12550 15170 -12430
rect 15290 -12550 15335 -12430
rect 15455 -12550 15500 -12430
rect 15620 -12550 15675 -12430
rect 15795 -12550 15840 -12430
rect 15960 -12550 16005 -12430
rect 16125 -12550 16170 -12430
rect 16290 -12550 16345 -12430
rect 16465 -12550 16510 -12430
rect 16630 -12550 16675 -12430
rect 16795 -12550 16840 -12430
rect 16960 -12550 17015 -12430
rect 17135 -12550 17180 -12430
rect 17300 -12550 17345 -12430
rect 17465 -12550 17510 -12430
rect 17630 -12550 17685 -12430
rect 17805 -12550 17850 -12430
rect 17970 -12550 18015 -12430
rect 18135 -12550 18180 -12430
rect 18300 -12550 18325 -12430
rect 12795 -12595 18325 -12550
rect 12795 -12715 12820 -12595
rect 12940 -12715 12995 -12595
rect 13115 -12715 13160 -12595
rect 13280 -12715 13325 -12595
rect 13445 -12715 13490 -12595
rect 13610 -12715 13665 -12595
rect 13785 -12715 13830 -12595
rect 13950 -12715 13995 -12595
rect 14115 -12715 14160 -12595
rect 14280 -12715 14335 -12595
rect 14455 -12715 14500 -12595
rect 14620 -12715 14665 -12595
rect 14785 -12715 14830 -12595
rect 14950 -12715 15005 -12595
rect 15125 -12715 15170 -12595
rect 15290 -12715 15335 -12595
rect 15455 -12715 15500 -12595
rect 15620 -12715 15675 -12595
rect 15795 -12715 15840 -12595
rect 15960 -12715 16005 -12595
rect 16125 -12715 16170 -12595
rect 16290 -12715 16345 -12595
rect 16465 -12715 16510 -12595
rect 16630 -12715 16675 -12595
rect 16795 -12715 16840 -12595
rect 16960 -12715 17015 -12595
rect 17135 -12715 17180 -12595
rect 17300 -12715 17345 -12595
rect 17465 -12715 17510 -12595
rect 17630 -12715 17685 -12595
rect 17805 -12715 17850 -12595
rect 17970 -12715 18015 -12595
rect 18135 -12715 18180 -12595
rect 18300 -12715 18325 -12595
rect 12795 -12770 18325 -12715
rect 12795 -12890 12820 -12770
rect 12940 -12890 12995 -12770
rect 13115 -12890 13160 -12770
rect 13280 -12890 13325 -12770
rect 13445 -12890 13490 -12770
rect 13610 -12890 13665 -12770
rect 13785 -12890 13830 -12770
rect 13950 -12890 13995 -12770
rect 14115 -12890 14160 -12770
rect 14280 -12890 14335 -12770
rect 14455 -12890 14500 -12770
rect 14620 -12890 14665 -12770
rect 14785 -12890 14830 -12770
rect 14950 -12890 15005 -12770
rect 15125 -12890 15170 -12770
rect 15290 -12890 15335 -12770
rect 15455 -12890 15500 -12770
rect 15620 -12890 15675 -12770
rect 15795 -12890 15840 -12770
rect 15960 -12890 16005 -12770
rect 16125 -12890 16170 -12770
rect 16290 -12890 16345 -12770
rect 16465 -12890 16510 -12770
rect 16630 -12890 16675 -12770
rect 16795 -12890 16840 -12770
rect 16960 -12890 17015 -12770
rect 17135 -12890 17180 -12770
rect 17300 -12890 17345 -12770
rect 17465 -12890 17510 -12770
rect 17630 -12890 17685 -12770
rect 17805 -12890 17850 -12770
rect 17970 -12890 18015 -12770
rect 18135 -12890 18180 -12770
rect 18300 -12890 18325 -12770
rect 12795 -12935 18325 -12890
rect 12795 -13055 12820 -12935
rect 12940 -13055 12995 -12935
rect 13115 -13055 13160 -12935
rect 13280 -13055 13325 -12935
rect 13445 -13055 13490 -12935
rect 13610 -13055 13665 -12935
rect 13785 -13055 13830 -12935
rect 13950 -13055 13995 -12935
rect 14115 -13055 14160 -12935
rect 14280 -13055 14335 -12935
rect 14455 -13055 14500 -12935
rect 14620 -13055 14665 -12935
rect 14785 -13055 14830 -12935
rect 14950 -13055 15005 -12935
rect 15125 -13055 15170 -12935
rect 15290 -13055 15335 -12935
rect 15455 -13055 15500 -12935
rect 15620 -13055 15675 -12935
rect 15795 -13055 15840 -12935
rect 15960 -13055 16005 -12935
rect 16125 -13055 16170 -12935
rect 16290 -13055 16345 -12935
rect 16465 -13055 16510 -12935
rect 16630 -13055 16675 -12935
rect 16795 -13055 16840 -12935
rect 16960 -13055 17015 -12935
rect 17135 -13055 17180 -12935
rect 17300 -13055 17345 -12935
rect 17465 -13055 17510 -12935
rect 17630 -13055 17685 -12935
rect 17805 -13055 17850 -12935
rect 17970 -13055 18015 -12935
rect 18135 -13055 18180 -12935
rect 18300 -13055 18325 -12935
rect 12795 -13100 18325 -13055
rect 12795 -13220 12820 -13100
rect 12940 -13220 12995 -13100
rect 13115 -13220 13160 -13100
rect 13280 -13220 13325 -13100
rect 13445 -13220 13490 -13100
rect 13610 -13220 13665 -13100
rect 13785 -13220 13830 -13100
rect 13950 -13220 13995 -13100
rect 14115 -13220 14160 -13100
rect 14280 -13220 14335 -13100
rect 14455 -13220 14500 -13100
rect 14620 -13220 14665 -13100
rect 14785 -13220 14830 -13100
rect 14950 -13220 15005 -13100
rect 15125 -13220 15170 -13100
rect 15290 -13220 15335 -13100
rect 15455 -13220 15500 -13100
rect 15620 -13220 15675 -13100
rect 15795 -13220 15840 -13100
rect 15960 -13220 16005 -13100
rect 16125 -13220 16170 -13100
rect 16290 -13220 16345 -13100
rect 16465 -13220 16510 -13100
rect 16630 -13220 16675 -13100
rect 16795 -13220 16840 -13100
rect 16960 -13220 17015 -13100
rect 17135 -13220 17180 -13100
rect 17300 -13220 17345 -13100
rect 17465 -13220 17510 -13100
rect 17630 -13220 17685 -13100
rect 17805 -13220 17850 -13100
rect 17970 -13220 18015 -13100
rect 18135 -13220 18180 -13100
rect 18300 -13220 18325 -13100
rect 12795 -13265 18325 -13220
rect 12795 -13385 12820 -13265
rect 12940 -13385 12995 -13265
rect 13115 -13385 13160 -13265
rect 13280 -13385 13325 -13265
rect 13445 -13385 13490 -13265
rect 13610 -13385 13665 -13265
rect 13785 -13385 13830 -13265
rect 13950 -13385 13995 -13265
rect 14115 -13385 14160 -13265
rect 14280 -13385 14335 -13265
rect 14455 -13385 14500 -13265
rect 14620 -13385 14665 -13265
rect 14785 -13385 14830 -13265
rect 14950 -13385 15005 -13265
rect 15125 -13385 15170 -13265
rect 15290 -13385 15335 -13265
rect 15455 -13385 15500 -13265
rect 15620 -13385 15675 -13265
rect 15795 -13385 15840 -13265
rect 15960 -13385 16005 -13265
rect 16125 -13385 16170 -13265
rect 16290 -13385 16345 -13265
rect 16465 -13385 16510 -13265
rect 16630 -13385 16675 -13265
rect 16795 -13385 16840 -13265
rect 16960 -13385 17015 -13265
rect 17135 -13385 17180 -13265
rect 17300 -13385 17345 -13265
rect 17465 -13385 17510 -13265
rect 17630 -13385 17685 -13265
rect 17805 -13385 17850 -13265
rect 17970 -13385 18015 -13265
rect 18135 -13385 18180 -13265
rect 18300 -13385 18325 -13265
rect 12795 -13440 18325 -13385
rect 12795 -13560 12820 -13440
rect 12940 -13560 12995 -13440
rect 13115 -13560 13160 -13440
rect 13280 -13560 13325 -13440
rect 13445 -13560 13490 -13440
rect 13610 -13560 13665 -13440
rect 13785 -13560 13830 -13440
rect 13950 -13560 13995 -13440
rect 14115 -13560 14160 -13440
rect 14280 -13560 14335 -13440
rect 14455 -13560 14500 -13440
rect 14620 -13560 14665 -13440
rect 14785 -13560 14830 -13440
rect 14950 -13560 15005 -13440
rect 15125 -13560 15170 -13440
rect 15290 -13560 15335 -13440
rect 15455 -13560 15500 -13440
rect 15620 -13560 15675 -13440
rect 15795 -13560 15840 -13440
rect 15960 -13560 16005 -13440
rect 16125 -13560 16170 -13440
rect 16290 -13560 16345 -13440
rect 16465 -13560 16510 -13440
rect 16630 -13560 16675 -13440
rect 16795 -13560 16840 -13440
rect 16960 -13560 17015 -13440
rect 17135 -13560 17180 -13440
rect 17300 -13560 17345 -13440
rect 17465 -13560 17510 -13440
rect 17630 -13560 17685 -13440
rect 17805 -13560 17850 -13440
rect 17970 -13560 18015 -13440
rect 18135 -13560 18180 -13440
rect 18300 -13560 18325 -13440
rect 12795 -13605 18325 -13560
rect 12795 -13725 12820 -13605
rect 12940 -13725 12995 -13605
rect 13115 -13725 13160 -13605
rect 13280 -13725 13325 -13605
rect 13445 -13725 13490 -13605
rect 13610 -13725 13665 -13605
rect 13785 -13725 13830 -13605
rect 13950 -13725 13995 -13605
rect 14115 -13725 14160 -13605
rect 14280 -13725 14335 -13605
rect 14455 -13725 14500 -13605
rect 14620 -13725 14665 -13605
rect 14785 -13725 14830 -13605
rect 14950 -13725 15005 -13605
rect 15125 -13725 15170 -13605
rect 15290 -13725 15335 -13605
rect 15455 -13725 15500 -13605
rect 15620 -13725 15675 -13605
rect 15795 -13725 15840 -13605
rect 15960 -13725 16005 -13605
rect 16125 -13725 16170 -13605
rect 16290 -13725 16345 -13605
rect 16465 -13725 16510 -13605
rect 16630 -13725 16675 -13605
rect 16795 -13725 16840 -13605
rect 16960 -13725 17015 -13605
rect 17135 -13725 17180 -13605
rect 17300 -13725 17345 -13605
rect 17465 -13725 17510 -13605
rect 17630 -13725 17685 -13605
rect 17805 -13725 17850 -13605
rect 17970 -13725 18015 -13605
rect 18135 -13725 18180 -13605
rect 18300 -13725 18325 -13605
rect 12795 -13770 18325 -13725
rect 12795 -13890 12820 -13770
rect 12940 -13890 12995 -13770
rect 13115 -13890 13160 -13770
rect 13280 -13890 13325 -13770
rect 13445 -13890 13490 -13770
rect 13610 -13890 13665 -13770
rect 13785 -13890 13830 -13770
rect 13950 -13890 13995 -13770
rect 14115 -13890 14160 -13770
rect 14280 -13890 14335 -13770
rect 14455 -13890 14500 -13770
rect 14620 -13890 14665 -13770
rect 14785 -13890 14830 -13770
rect 14950 -13890 15005 -13770
rect 15125 -13890 15170 -13770
rect 15290 -13890 15335 -13770
rect 15455 -13890 15500 -13770
rect 15620 -13890 15675 -13770
rect 15795 -13890 15840 -13770
rect 15960 -13890 16005 -13770
rect 16125 -13890 16170 -13770
rect 16290 -13890 16345 -13770
rect 16465 -13890 16510 -13770
rect 16630 -13890 16675 -13770
rect 16795 -13890 16840 -13770
rect 16960 -13890 17015 -13770
rect 17135 -13890 17180 -13770
rect 17300 -13890 17345 -13770
rect 17465 -13890 17510 -13770
rect 17630 -13890 17685 -13770
rect 17805 -13890 17850 -13770
rect 17970 -13890 18015 -13770
rect 18135 -13890 18180 -13770
rect 18300 -13890 18325 -13770
rect 12795 -13935 18325 -13890
rect 12795 -14055 12820 -13935
rect 12940 -14055 12995 -13935
rect 13115 -14055 13160 -13935
rect 13280 -14055 13325 -13935
rect 13445 -14055 13490 -13935
rect 13610 -14055 13665 -13935
rect 13785 -14055 13830 -13935
rect 13950 -14055 13995 -13935
rect 14115 -14055 14160 -13935
rect 14280 -14055 14335 -13935
rect 14455 -14055 14500 -13935
rect 14620 -14055 14665 -13935
rect 14785 -14055 14830 -13935
rect 14950 -14055 15005 -13935
rect 15125 -14055 15170 -13935
rect 15290 -14055 15335 -13935
rect 15455 -14055 15500 -13935
rect 15620 -14055 15675 -13935
rect 15795 -14055 15840 -13935
rect 15960 -14055 16005 -13935
rect 16125 -14055 16170 -13935
rect 16290 -14055 16345 -13935
rect 16465 -14055 16510 -13935
rect 16630 -14055 16675 -13935
rect 16795 -14055 16840 -13935
rect 16960 -14055 17015 -13935
rect 17135 -14055 17180 -13935
rect 17300 -14055 17345 -13935
rect 17465 -14055 17510 -13935
rect 17630 -14055 17685 -13935
rect 17805 -14055 17850 -13935
rect 17970 -14055 18015 -13935
rect 18135 -14055 18180 -13935
rect 18300 -14055 18325 -13935
rect 12795 -14110 18325 -14055
rect 12795 -14230 12820 -14110
rect 12940 -14230 12995 -14110
rect 13115 -14230 13160 -14110
rect 13280 -14230 13325 -14110
rect 13445 -14230 13490 -14110
rect 13610 -14230 13665 -14110
rect 13785 -14230 13830 -14110
rect 13950 -14230 13995 -14110
rect 14115 -14230 14160 -14110
rect 14280 -14230 14335 -14110
rect 14455 -14230 14500 -14110
rect 14620 -14230 14665 -14110
rect 14785 -14230 14830 -14110
rect 14950 -14230 15005 -14110
rect 15125 -14230 15170 -14110
rect 15290 -14230 15335 -14110
rect 15455 -14230 15500 -14110
rect 15620 -14230 15675 -14110
rect 15795 -14230 15840 -14110
rect 15960 -14230 16005 -14110
rect 16125 -14230 16170 -14110
rect 16290 -14230 16345 -14110
rect 16465 -14230 16510 -14110
rect 16630 -14230 16675 -14110
rect 16795 -14230 16840 -14110
rect 16960 -14230 17015 -14110
rect 17135 -14230 17180 -14110
rect 17300 -14230 17345 -14110
rect 17465 -14230 17510 -14110
rect 17630 -14230 17685 -14110
rect 17805 -14230 17850 -14110
rect 17970 -14230 18015 -14110
rect 18135 -14230 18180 -14110
rect 18300 -14230 18325 -14110
rect 12795 -14275 18325 -14230
rect 12795 -14395 12820 -14275
rect 12940 -14395 12995 -14275
rect 13115 -14395 13160 -14275
rect 13280 -14395 13325 -14275
rect 13445 -14395 13490 -14275
rect 13610 -14395 13665 -14275
rect 13785 -14395 13830 -14275
rect 13950 -14395 13995 -14275
rect 14115 -14395 14160 -14275
rect 14280 -14395 14335 -14275
rect 14455 -14395 14500 -14275
rect 14620 -14395 14665 -14275
rect 14785 -14395 14830 -14275
rect 14950 -14395 15005 -14275
rect 15125 -14395 15170 -14275
rect 15290 -14395 15335 -14275
rect 15455 -14395 15500 -14275
rect 15620 -14395 15675 -14275
rect 15795 -14395 15840 -14275
rect 15960 -14395 16005 -14275
rect 16125 -14395 16170 -14275
rect 16290 -14395 16345 -14275
rect 16465 -14395 16510 -14275
rect 16630 -14395 16675 -14275
rect 16795 -14395 16840 -14275
rect 16960 -14395 17015 -14275
rect 17135 -14395 17180 -14275
rect 17300 -14395 17345 -14275
rect 17465 -14395 17510 -14275
rect 17630 -14395 17685 -14275
rect 17805 -14395 17850 -14275
rect 17970 -14395 18015 -14275
rect 18135 -14395 18180 -14275
rect 18300 -14395 18325 -14275
rect 12795 -14440 18325 -14395
rect 12795 -14560 12820 -14440
rect 12940 -14560 12995 -14440
rect 13115 -14560 13160 -14440
rect 13280 -14560 13325 -14440
rect 13445 -14560 13490 -14440
rect 13610 -14560 13665 -14440
rect 13785 -14560 13830 -14440
rect 13950 -14560 13995 -14440
rect 14115 -14560 14160 -14440
rect 14280 -14560 14335 -14440
rect 14455 -14560 14500 -14440
rect 14620 -14560 14665 -14440
rect 14785 -14560 14830 -14440
rect 14950 -14560 15005 -14440
rect 15125 -14560 15170 -14440
rect 15290 -14560 15335 -14440
rect 15455 -14560 15500 -14440
rect 15620 -14560 15675 -14440
rect 15795 -14560 15840 -14440
rect 15960 -14560 16005 -14440
rect 16125 -14560 16170 -14440
rect 16290 -14560 16345 -14440
rect 16465 -14560 16510 -14440
rect 16630 -14560 16675 -14440
rect 16795 -14560 16840 -14440
rect 16960 -14560 17015 -14440
rect 17135 -14560 17180 -14440
rect 17300 -14560 17345 -14440
rect 17465 -14560 17510 -14440
rect 17630 -14560 17685 -14440
rect 17805 -14560 17850 -14440
rect 17970 -14560 18015 -14440
rect 18135 -14560 18180 -14440
rect 18300 -14560 18325 -14440
rect 12795 -14605 18325 -14560
rect 12795 -14725 12820 -14605
rect 12940 -14725 12995 -14605
rect 13115 -14725 13160 -14605
rect 13280 -14725 13325 -14605
rect 13445 -14725 13490 -14605
rect 13610 -14725 13665 -14605
rect 13785 -14725 13830 -14605
rect 13950 -14725 13995 -14605
rect 14115 -14725 14160 -14605
rect 14280 -14725 14335 -14605
rect 14455 -14725 14500 -14605
rect 14620 -14725 14665 -14605
rect 14785 -14725 14830 -14605
rect 14950 -14725 15005 -14605
rect 15125 -14725 15170 -14605
rect 15290 -14725 15335 -14605
rect 15455 -14725 15500 -14605
rect 15620 -14725 15675 -14605
rect 15795 -14725 15840 -14605
rect 15960 -14725 16005 -14605
rect 16125 -14725 16170 -14605
rect 16290 -14725 16345 -14605
rect 16465 -14725 16510 -14605
rect 16630 -14725 16675 -14605
rect 16795 -14725 16840 -14605
rect 16960 -14725 17015 -14605
rect 17135 -14725 17180 -14605
rect 17300 -14725 17345 -14605
rect 17465 -14725 17510 -14605
rect 17630 -14725 17685 -14605
rect 17805 -14725 17850 -14605
rect 17970 -14725 18015 -14605
rect 18135 -14725 18180 -14605
rect 18300 -14725 18325 -14605
rect 12795 -14780 18325 -14725
rect 12795 -14900 12820 -14780
rect 12940 -14900 12995 -14780
rect 13115 -14900 13160 -14780
rect 13280 -14900 13325 -14780
rect 13445 -14900 13490 -14780
rect 13610 -14900 13665 -14780
rect 13785 -14900 13830 -14780
rect 13950 -14900 13995 -14780
rect 14115 -14900 14160 -14780
rect 14280 -14900 14335 -14780
rect 14455 -14900 14500 -14780
rect 14620 -14900 14665 -14780
rect 14785 -14900 14830 -14780
rect 14950 -14900 15005 -14780
rect 15125 -14900 15170 -14780
rect 15290 -14900 15335 -14780
rect 15455 -14900 15500 -14780
rect 15620 -14900 15675 -14780
rect 15795 -14900 15840 -14780
rect 15960 -14900 16005 -14780
rect 16125 -14900 16170 -14780
rect 16290 -14900 16345 -14780
rect 16465 -14900 16510 -14780
rect 16630 -14900 16675 -14780
rect 16795 -14900 16840 -14780
rect 16960 -14900 17015 -14780
rect 17135 -14900 17180 -14780
rect 17300 -14900 17345 -14780
rect 17465 -14900 17510 -14780
rect 17630 -14900 17685 -14780
rect 17805 -14900 17850 -14780
rect 17970 -14900 18015 -14780
rect 18135 -14900 18180 -14780
rect 18300 -14900 18325 -14780
rect 12795 -14945 18325 -14900
rect 12795 -15065 12820 -14945
rect 12940 -15065 12995 -14945
rect 13115 -15065 13160 -14945
rect 13280 -15065 13325 -14945
rect 13445 -15065 13490 -14945
rect 13610 -15065 13665 -14945
rect 13785 -15065 13830 -14945
rect 13950 -15065 13995 -14945
rect 14115 -15065 14160 -14945
rect 14280 -15065 14335 -14945
rect 14455 -15065 14500 -14945
rect 14620 -15065 14665 -14945
rect 14785 -15065 14830 -14945
rect 14950 -15065 15005 -14945
rect 15125 -15065 15170 -14945
rect 15290 -15065 15335 -14945
rect 15455 -15065 15500 -14945
rect 15620 -15065 15675 -14945
rect 15795 -15065 15840 -14945
rect 15960 -15065 16005 -14945
rect 16125 -15065 16170 -14945
rect 16290 -15065 16345 -14945
rect 16465 -15065 16510 -14945
rect 16630 -15065 16675 -14945
rect 16795 -15065 16840 -14945
rect 16960 -15065 17015 -14945
rect 17135 -15065 17180 -14945
rect 17300 -15065 17345 -14945
rect 17465 -15065 17510 -14945
rect 17630 -15065 17685 -14945
rect 17805 -15065 17850 -14945
rect 17970 -15065 18015 -14945
rect 18135 -15065 18180 -14945
rect 18300 -15065 18325 -14945
rect 12795 -15110 18325 -15065
rect 12795 -15230 12820 -15110
rect 12940 -15230 12995 -15110
rect 13115 -15230 13160 -15110
rect 13280 -15230 13325 -15110
rect 13445 -15230 13490 -15110
rect 13610 -15230 13665 -15110
rect 13785 -15230 13830 -15110
rect 13950 -15230 13995 -15110
rect 14115 -15230 14160 -15110
rect 14280 -15230 14335 -15110
rect 14455 -15230 14500 -15110
rect 14620 -15230 14665 -15110
rect 14785 -15230 14830 -15110
rect 14950 -15230 15005 -15110
rect 15125 -15230 15170 -15110
rect 15290 -15230 15335 -15110
rect 15455 -15230 15500 -15110
rect 15620 -15230 15675 -15110
rect 15795 -15230 15840 -15110
rect 15960 -15230 16005 -15110
rect 16125 -15230 16170 -15110
rect 16290 -15230 16345 -15110
rect 16465 -15230 16510 -15110
rect 16630 -15230 16675 -15110
rect 16795 -15230 16840 -15110
rect 16960 -15230 17015 -15110
rect 17135 -15230 17180 -15110
rect 17300 -15230 17345 -15110
rect 17465 -15230 17510 -15110
rect 17630 -15230 17685 -15110
rect 17805 -15230 17850 -15110
rect 17970 -15230 18015 -15110
rect 18135 -15230 18180 -15110
rect 18300 -15230 18325 -15110
rect 12795 -15275 18325 -15230
rect 12795 -15395 12820 -15275
rect 12940 -15395 12995 -15275
rect 13115 -15395 13160 -15275
rect 13280 -15395 13325 -15275
rect 13445 -15395 13490 -15275
rect 13610 -15395 13665 -15275
rect 13785 -15395 13830 -15275
rect 13950 -15395 13995 -15275
rect 14115 -15395 14160 -15275
rect 14280 -15395 14335 -15275
rect 14455 -15395 14500 -15275
rect 14620 -15395 14665 -15275
rect 14785 -15395 14830 -15275
rect 14950 -15395 15005 -15275
rect 15125 -15395 15170 -15275
rect 15290 -15395 15335 -15275
rect 15455 -15395 15500 -15275
rect 15620 -15395 15675 -15275
rect 15795 -15395 15840 -15275
rect 15960 -15395 16005 -15275
rect 16125 -15395 16170 -15275
rect 16290 -15395 16345 -15275
rect 16465 -15395 16510 -15275
rect 16630 -15395 16675 -15275
rect 16795 -15395 16840 -15275
rect 16960 -15395 17015 -15275
rect 17135 -15395 17180 -15275
rect 17300 -15395 17345 -15275
rect 17465 -15395 17510 -15275
rect 17630 -15395 17685 -15275
rect 17805 -15395 17850 -15275
rect 17970 -15395 18015 -15275
rect 18135 -15395 18180 -15275
rect 18300 -15395 18325 -15275
rect 12795 -15450 18325 -15395
rect 12795 -15535 12820 -15450
rect 12610 -15570 12820 -15535
rect 12940 -15570 12995 -15450
rect 13115 -15570 13160 -15450
rect 13280 -15570 13325 -15450
rect 13445 -15570 13490 -15450
rect 13610 -15570 13665 -15450
rect 13785 -15570 13830 -15450
rect 13950 -15570 13995 -15450
rect 14115 -15570 14160 -15450
rect 14280 -15570 14335 -15450
rect 14455 -15570 14500 -15450
rect 14620 -15570 14665 -15450
rect 14785 -15570 14830 -15450
rect 14950 -15570 15005 -15450
rect 15125 -15570 15170 -15450
rect 15290 -15570 15335 -15450
rect 15455 -15570 15500 -15450
rect 15620 -15570 15675 -15450
rect 15795 -15570 15840 -15450
rect 15960 -15570 16005 -15450
rect 16125 -15570 16170 -15450
rect 16290 -15570 16345 -15450
rect 16465 -15570 16510 -15450
rect 16630 -15570 16675 -15450
rect 16795 -15570 16840 -15450
rect 16960 -15570 17015 -15450
rect 17135 -15570 17180 -15450
rect 17300 -15570 17345 -15450
rect 17465 -15570 17510 -15450
rect 17630 -15570 17685 -15450
rect 17805 -15570 17850 -15450
rect 17970 -15570 18015 -15450
rect 18135 -15570 18180 -15450
rect 18300 -15535 18325 -15450
rect 18485 -10090 24015 -10065
rect 18485 -10210 18510 -10090
rect 18630 -10210 18685 -10090
rect 18805 -10210 18850 -10090
rect 18970 -10210 19015 -10090
rect 19135 -10210 19180 -10090
rect 19300 -10210 19355 -10090
rect 19475 -10210 19520 -10090
rect 19640 -10210 19685 -10090
rect 19805 -10210 19850 -10090
rect 19970 -10210 20025 -10090
rect 20145 -10210 20190 -10090
rect 20310 -10210 20355 -10090
rect 20475 -10210 20520 -10090
rect 20640 -10210 20695 -10090
rect 20815 -10210 20860 -10090
rect 20980 -10210 21025 -10090
rect 21145 -10210 21190 -10090
rect 21310 -10210 21365 -10090
rect 21485 -10210 21530 -10090
rect 21650 -10210 21695 -10090
rect 21815 -10210 21860 -10090
rect 21980 -10210 22035 -10090
rect 22155 -10210 22200 -10090
rect 22320 -10210 22365 -10090
rect 22485 -10210 22530 -10090
rect 22650 -10210 22705 -10090
rect 22825 -10210 22870 -10090
rect 22990 -10210 23035 -10090
rect 23155 -10210 23200 -10090
rect 23320 -10210 23375 -10090
rect 23495 -10210 23540 -10090
rect 23660 -10210 23705 -10090
rect 23825 -10210 23870 -10090
rect 23990 -10210 24015 -10090
rect 18485 -10255 24015 -10210
rect 18485 -10375 18510 -10255
rect 18630 -10375 18685 -10255
rect 18805 -10375 18850 -10255
rect 18970 -10375 19015 -10255
rect 19135 -10375 19180 -10255
rect 19300 -10375 19355 -10255
rect 19475 -10375 19520 -10255
rect 19640 -10375 19685 -10255
rect 19805 -10375 19850 -10255
rect 19970 -10375 20025 -10255
rect 20145 -10375 20190 -10255
rect 20310 -10375 20355 -10255
rect 20475 -10375 20520 -10255
rect 20640 -10375 20695 -10255
rect 20815 -10375 20860 -10255
rect 20980 -10375 21025 -10255
rect 21145 -10375 21190 -10255
rect 21310 -10375 21365 -10255
rect 21485 -10375 21530 -10255
rect 21650 -10375 21695 -10255
rect 21815 -10375 21860 -10255
rect 21980 -10375 22035 -10255
rect 22155 -10375 22200 -10255
rect 22320 -10375 22365 -10255
rect 22485 -10375 22530 -10255
rect 22650 -10375 22705 -10255
rect 22825 -10375 22870 -10255
rect 22990 -10375 23035 -10255
rect 23155 -10375 23200 -10255
rect 23320 -10375 23375 -10255
rect 23495 -10375 23540 -10255
rect 23660 -10375 23705 -10255
rect 23825 -10375 23870 -10255
rect 23990 -10375 24015 -10255
rect 18485 -10420 24015 -10375
rect 18485 -10540 18510 -10420
rect 18630 -10540 18685 -10420
rect 18805 -10540 18850 -10420
rect 18970 -10540 19015 -10420
rect 19135 -10540 19180 -10420
rect 19300 -10540 19355 -10420
rect 19475 -10540 19520 -10420
rect 19640 -10540 19685 -10420
rect 19805 -10540 19850 -10420
rect 19970 -10540 20025 -10420
rect 20145 -10540 20190 -10420
rect 20310 -10540 20355 -10420
rect 20475 -10540 20520 -10420
rect 20640 -10540 20695 -10420
rect 20815 -10540 20860 -10420
rect 20980 -10540 21025 -10420
rect 21145 -10540 21190 -10420
rect 21310 -10540 21365 -10420
rect 21485 -10540 21530 -10420
rect 21650 -10540 21695 -10420
rect 21815 -10540 21860 -10420
rect 21980 -10540 22035 -10420
rect 22155 -10540 22200 -10420
rect 22320 -10540 22365 -10420
rect 22485 -10540 22530 -10420
rect 22650 -10540 22705 -10420
rect 22825 -10540 22870 -10420
rect 22990 -10540 23035 -10420
rect 23155 -10540 23200 -10420
rect 23320 -10540 23375 -10420
rect 23495 -10540 23540 -10420
rect 23660 -10540 23705 -10420
rect 23825 -10540 23870 -10420
rect 23990 -10540 24015 -10420
rect 18485 -10585 24015 -10540
rect 18485 -10705 18510 -10585
rect 18630 -10705 18685 -10585
rect 18805 -10705 18850 -10585
rect 18970 -10705 19015 -10585
rect 19135 -10705 19180 -10585
rect 19300 -10705 19355 -10585
rect 19475 -10705 19520 -10585
rect 19640 -10705 19685 -10585
rect 19805 -10705 19850 -10585
rect 19970 -10705 20025 -10585
rect 20145 -10705 20190 -10585
rect 20310 -10705 20355 -10585
rect 20475 -10705 20520 -10585
rect 20640 -10705 20695 -10585
rect 20815 -10705 20860 -10585
rect 20980 -10705 21025 -10585
rect 21145 -10705 21190 -10585
rect 21310 -10705 21365 -10585
rect 21485 -10705 21530 -10585
rect 21650 -10705 21695 -10585
rect 21815 -10705 21860 -10585
rect 21980 -10705 22035 -10585
rect 22155 -10705 22200 -10585
rect 22320 -10705 22365 -10585
rect 22485 -10705 22530 -10585
rect 22650 -10705 22705 -10585
rect 22825 -10705 22870 -10585
rect 22990 -10705 23035 -10585
rect 23155 -10705 23200 -10585
rect 23320 -10705 23375 -10585
rect 23495 -10705 23540 -10585
rect 23660 -10705 23705 -10585
rect 23825 -10705 23870 -10585
rect 23990 -10705 24015 -10585
rect 18485 -10760 24015 -10705
rect 18485 -10880 18510 -10760
rect 18630 -10880 18685 -10760
rect 18805 -10880 18850 -10760
rect 18970 -10880 19015 -10760
rect 19135 -10880 19180 -10760
rect 19300 -10880 19355 -10760
rect 19475 -10880 19520 -10760
rect 19640 -10880 19685 -10760
rect 19805 -10880 19850 -10760
rect 19970 -10880 20025 -10760
rect 20145 -10880 20190 -10760
rect 20310 -10880 20355 -10760
rect 20475 -10880 20520 -10760
rect 20640 -10880 20695 -10760
rect 20815 -10880 20860 -10760
rect 20980 -10880 21025 -10760
rect 21145 -10880 21190 -10760
rect 21310 -10880 21365 -10760
rect 21485 -10880 21530 -10760
rect 21650 -10880 21695 -10760
rect 21815 -10880 21860 -10760
rect 21980 -10880 22035 -10760
rect 22155 -10880 22200 -10760
rect 22320 -10880 22365 -10760
rect 22485 -10880 22530 -10760
rect 22650 -10880 22705 -10760
rect 22825 -10880 22870 -10760
rect 22990 -10880 23035 -10760
rect 23155 -10880 23200 -10760
rect 23320 -10880 23375 -10760
rect 23495 -10880 23540 -10760
rect 23660 -10880 23705 -10760
rect 23825 -10880 23870 -10760
rect 23990 -10880 24015 -10760
rect 18485 -10925 24015 -10880
rect 18485 -11045 18510 -10925
rect 18630 -11045 18685 -10925
rect 18805 -11045 18850 -10925
rect 18970 -11045 19015 -10925
rect 19135 -11045 19180 -10925
rect 19300 -11045 19355 -10925
rect 19475 -11045 19520 -10925
rect 19640 -11045 19685 -10925
rect 19805 -11045 19850 -10925
rect 19970 -11045 20025 -10925
rect 20145 -11045 20190 -10925
rect 20310 -11045 20355 -10925
rect 20475 -11045 20520 -10925
rect 20640 -11045 20695 -10925
rect 20815 -11045 20860 -10925
rect 20980 -11045 21025 -10925
rect 21145 -11045 21190 -10925
rect 21310 -11045 21365 -10925
rect 21485 -11045 21530 -10925
rect 21650 -11045 21695 -10925
rect 21815 -11045 21860 -10925
rect 21980 -11045 22035 -10925
rect 22155 -11045 22200 -10925
rect 22320 -11045 22365 -10925
rect 22485 -11045 22530 -10925
rect 22650 -11045 22705 -10925
rect 22825 -11045 22870 -10925
rect 22990 -11045 23035 -10925
rect 23155 -11045 23200 -10925
rect 23320 -11045 23375 -10925
rect 23495 -11045 23540 -10925
rect 23660 -11045 23705 -10925
rect 23825 -11045 23870 -10925
rect 23990 -11045 24015 -10925
rect 18485 -11090 24015 -11045
rect 18485 -11210 18510 -11090
rect 18630 -11210 18685 -11090
rect 18805 -11210 18850 -11090
rect 18970 -11210 19015 -11090
rect 19135 -11210 19180 -11090
rect 19300 -11210 19355 -11090
rect 19475 -11210 19520 -11090
rect 19640 -11210 19685 -11090
rect 19805 -11210 19850 -11090
rect 19970 -11210 20025 -11090
rect 20145 -11210 20190 -11090
rect 20310 -11210 20355 -11090
rect 20475 -11210 20520 -11090
rect 20640 -11210 20695 -11090
rect 20815 -11210 20860 -11090
rect 20980 -11210 21025 -11090
rect 21145 -11210 21190 -11090
rect 21310 -11210 21365 -11090
rect 21485 -11210 21530 -11090
rect 21650 -11210 21695 -11090
rect 21815 -11210 21860 -11090
rect 21980 -11210 22035 -11090
rect 22155 -11210 22200 -11090
rect 22320 -11210 22365 -11090
rect 22485 -11210 22530 -11090
rect 22650 -11210 22705 -11090
rect 22825 -11210 22870 -11090
rect 22990 -11210 23035 -11090
rect 23155 -11210 23200 -11090
rect 23320 -11210 23375 -11090
rect 23495 -11210 23540 -11090
rect 23660 -11210 23705 -11090
rect 23825 -11210 23870 -11090
rect 23990 -11210 24015 -11090
rect 18485 -11255 24015 -11210
rect 18485 -11375 18510 -11255
rect 18630 -11375 18685 -11255
rect 18805 -11375 18850 -11255
rect 18970 -11375 19015 -11255
rect 19135 -11375 19180 -11255
rect 19300 -11375 19355 -11255
rect 19475 -11375 19520 -11255
rect 19640 -11375 19685 -11255
rect 19805 -11375 19850 -11255
rect 19970 -11375 20025 -11255
rect 20145 -11375 20190 -11255
rect 20310 -11375 20355 -11255
rect 20475 -11375 20520 -11255
rect 20640 -11375 20695 -11255
rect 20815 -11375 20860 -11255
rect 20980 -11375 21025 -11255
rect 21145 -11375 21190 -11255
rect 21310 -11375 21365 -11255
rect 21485 -11375 21530 -11255
rect 21650 -11375 21695 -11255
rect 21815 -11375 21860 -11255
rect 21980 -11375 22035 -11255
rect 22155 -11375 22200 -11255
rect 22320 -11375 22365 -11255
rect 22485 -11375 22530 -11255
rect 22650 -11375 22705 -11255
rect 22825 -11375 22870 -11255
rect 22990 -11375 23035 -11255
rect 23155 -11375 23200 -11255
rect 23320 -11375 23375 -11255
rect 23495 -11375 23540 -11255
rect 23660 -11375 23705 -11255
rect 23825 -11375 23870 -11255
rect 23990 -11375 24015 -11255
rect 18485 -11430 24015 -11375
rect 18485 -11550 18510 -11430
rect 18630 -11550 18685 -11430
rect 18805 -11550 18850 -11430
rect 18970 -11550 19015 -11430
rect 19135 -11550 19180 -11430
rect 19300 -11550 19355 -11430
rect 19475 -11550 19520 -11430
rect 19640 -11550 19685 -11430
rect 19805 -11550 19850 -11430
rect 19970 -11550 20025 -11430
rect 20145 -11550 20190 -11430
rect 20310 -11550 20355 -11430
rect 20475 -11550 20520 -11430
rect 20640 -11550 20695 -11430
rect 20815 -11550 20860 -11430
rect 20980 -11550 21025 -11430
rect 21145 -11550 21190 -11430
rect 21310 -11550 21365 -11430
rect 21485 -11550 21530 -11430
rect 21650 -11550 21695 -11430
rect 21815 -11550 21860 -11430
rect 21980 -11550 22035 -11430
rect 22155 -11550 22200 -11430
rect 22320 -11550 22365 -11430
rect 22485 -11550 22530 -11430
rect 22650 -11550 22705 -11430
rect 22825 -11550 22870 -11430
rect 22990 -11550 23035 -11430
rect 23155 -11550 23200 -11430
rect 23320 -11550 23375 -11430
rect 23495 -11550 23540 -11430
rect 23660 -11550 23705 -11430
rect 23825 -11550 23870 -11430
rect 23990 -11550 24015 -11430
rect 18485 -11595 24015 -11550
rect 18485 -11715 18510 -11595
rect 18630 -11715 18685 -11595
rect 18805 -11715 18850 -11595
rect 18970 -11715 19015 -11595
rect 19135 -11715 19180 -11595
rect 19300 -11715 19355 -11595
rect 19475 -11715 19520 -11595
rect 19640 -11715 19685 -11595
rect 19805 -11715 19850 -11595
rect 19970 -11715 20025 -11595
rect 20145 -11715 20190 -11595
rect 20310 -11715 20355 -11595
rect 20475 -11715 20520 -11595
rect 20640 -11715 20695 -11595
rect 20815 -11715 20860 -11595
rect 20980 -11715 21025 -11595
rect 21145 -11715 21190 -11595
rect 21310 -11715 21365 -11595
rect 21485 -11715 21530 -11595
rect 21650 -11715 21695 -11595
rect 21815 -11715 21860 -11595
rect 21980 -11715 22035 -11595
rect 22155 -11715 22200 -11595
rect 22320 -11715 22365 -11595
rect 22485 -11715 22530 -11595
rect 22650 -11715 22705 -11595
rect 22825 -11715 22870 -11595
rect 22990 -11715 23035 -11595
rect 23155 -11715 23200 -11595
rect 23320 -11715 23375 -11595
rect 23495 -11715 23540 -11595
rect 23660 -11715 23705 -11595
rect 23825 -11715 23870 -11595
rect 23990 -11715 24015 -11595
rect 18485 -11760 24015 -11715
rect 18485 -11880 18510 -11760
rect 18630 -11880 18685 -11760
rect 18805 -11880 18850 -11760
rect 18970 -11880 19015 -11760
rect 19135 -11880 19180 -11760
rect 19300 -11880 19355 -11760
rect 19475 -11880 19520 -11760
rect 19640 -11880 19685 -11760
rect 19805 -11880 19850 -11760
rect 19970 -11880 20025 -11760
rect 20145 -11880 20190 -11760
rect 20310 -11880 20355 -11760
rect 20475 -11880 20520 -11760
rect 20640 -11880 20695 -11760
rect 20815 -11880 20860 -11760
rect 20980 -11880 21025 -11760
rect 21145 -11880 21190 -11760
rect 21310 -11880 21365 -11760
rect 21485 -11880 21530 -11760
rect 21650 -11880 21695 -11760
rect 21815 -11880 21860 -11760
rect 21980 -11880 22035 -11760
rect 22155 -11880 22200 -11760
rect 22320 -11880 22365 -11760
rect 22485 -11880 22530 -11760
rect 22650 -11880 22705 -11760
rect 22825 -11880 22870 -11760
rect 22990 -11880 23035 -11760
rect 23155 -11880 23200 -11760
rect 23320 -11880 23375 -11760
rect 23495 -11880 23540 -11760
rect 23660 -11880 23705 -11760
rect 23825 -11880 23870 -11760
rect 23990 -11880 24015 -11760
rect 18485 -11925 24015 -11880
rect 18485 -12045 18510 -11925
rect 18630 -12045 18685 -11925
rect 18805 -12045 18850 -11925
rect 18970 -12045 19015 -11925
rect 19135 -12045 19180 -11925
rect 19300 -12045 19355 -11925
rect 19475 -12045 19520 -11925
rect 19640 -12045 19685 -11925
rect 19805 -12045 19850 -11925
rect 19970 -12045 20025 -11925
rect 20145 -12045 20190 -11925
rect 20310 -12045 20355 -11925
rect 20475 -12045 20520 -11925
rect 20640 -12045 20695 -11925
rect 20815 -12045 20860 -11925
rect 20980 -12045 21025 -11925
rect 21145 -12045 21190 -11925
rect 21310 -12045 21365 -11925
rect 21485 -12045 21530 -11925
rect 21650 -12045 21695 -11925
rect 21815 -12045 21860 -11925
rect 21980 -12045 22035 -11925
rect 22155 -12045 22200 -11925
rect 22320 -12045 22365 -11925
rect 22485 -12045 22530 -11925
rect 22650 -12045 22705 -11925
rect 22825 -12045 22870 -11925
rect 22990 -12045 23035 -11925
rect 23155 -12045 23200 -11925
rect 23320 -12045 23375 -11925
rect 23495 -12045 23540 -11925
rect 23660 -12045 23705 -11925
rect 23825 -12045 23870 -11925
rect 23990 -12045 24015 -11925
rect 18485 -12100 24015 -12045
rect 18485 -12220 18510 -12100
rect 18630 -12220 18685 -12100
rect 18805 -12220 18850 -12100
rect 18970 -12220 19015 -12100
rect 19135 -12220 19180 -12100
rect 19300 -12220 19355 -12100
rect 19475 -12220 19520 -12100
rect 19640 -12220 19685 -12100
rect 19805 -12220 19850 -12100
rect 19970 -12220 20025 -12100
rect 20145 -12220 20190 -12100
rect 20310 -12220 20355 -12100
rect 20475 -12220 20520 -12100
rect 20640 -12220 20695 -12100
rect 20815 -12220 20860 -12100
rect 20980 -12220 21025 -12100
rect 21145 -12220 21190 -12100
rect 21310 -12220 21365 -12100
rect 21485 -12220 21530 -12100
rect 21650 -12220 21695 -12100
rect 21815 -12220 21860 -12100
rect 21980 -12220 22035 -12100
rect 22155 -12220 22200 -12100
rect 22320 -12220 22365 -12100
rect 22485 -12220 22530 -12100
rect 22650 -12220 22705 -12100
rect 22825 -12220 22870 -12100
rect 22990 -12220 23035 -12100
rect 23155 -12220 23200 -12100
rect 23320 -12220 23375 -12100
rect 23495 -12220 23540 -12100
rect 23660 -12220 23705 -12100
rect 23825 -12220 23870 -12100
rect 23990 -12220 24015 -12100
rect 18485 -12265 24015 -12220
rect 18485 -12385 18510 -12265
rect 18630 -12385 18685 -12265
rect 18805 -12385 18850 -12265
rect 18970 -12385 19015 -12265
rect 19135 -12385 19180 -12265
rect 19300 -12385 19355 -12265
rect 19475 -12385 19520 -12265
rect 19640 -12385 19685 -12265
rect 19805 -12385 19850 -12265
rect 19970 -12385 20025 -12265
rect 20145 -12385 20190 -12265
rect 20310 -12385 20355 -12265
rect 20475 -12385 20520 -12265
rect 20640 -12385 20695 -12265
rect 20815 -12385 20860 -12265
rect 20980 -12385 21025 -12265
rect 21145 -12385 21190 -12265
rect 21310 -12385 21365 -12265
rect 21485 -12385 21530 -12265
rect 21650 -12385 21695 -12265
rect 21815 -12385 21860 -12265
rect 21980 -12385 22035 -12265
rect 22155 -12385 22200 -12265
rect 22320 -12385 22365 -12265
rect 22485 -12385 22530 -12265
rect 22650 -12385 22705 -12265
rect 22825 -12385 22870 -12265
rect 22990 -12385 23035 -12265
rect 23155 -12385 23200 -12265
rect 23320 -12385 23375 -12265
rect 23495 -12385 23540 -12265
rect 23660 -12385 23705 -12265
rect 23825 -12385 23870 -12265
rect 23990 -12385 24015 -12265
rect 18485 -12430 24015 -12385
rect 18485 -12550 18510 -12430
rect 18630 -12550 18685 -12430
rect 18805 -12550 18850 -12430
rect 18970 -12550 19015 -12430
rect 19135 -12550 19180 -12430
rect 19300 -12550 19355 -12430
rect 19475 -12550 19520 -12430
rect 19640 -12550 19685 -12430
rect 19805 -12550 19850 -12430
rect 19970 -12550 20025 -12430
rect 20145 -12550 20190 -12430
rect 20310 -12550 20355 -12430
rect 20475 -12550 20520 -12430
rect 20640 -12550 20695 -12430
rect 20815 -12550 20860 -12430
rect 20980 -12550 21025 -12430
rect 21145 -12550 21190 -12430
rect 21310 -12550 21365 -12430
rect 21485 -12550 21530 -12430
rect 21650 -12550 21695 -12430
rect 21815 -12550 21860 -12430
rect 21980 -12550 22035 -12430
rect 22155 -12550 22200 -12430
rect 22320 -12550 22365 -12430
rect 22485 -12550 22530 -12430
rect 22650 -12550 22705 -12430
rect 22825 -12550 22870 -12430
rect 22990 -12550 23035 -12430
rect 23155 -12550 23200 -12430
rect 23320 -12550 23375 -12430
rect 23495 -12550 23540 -12430
rect 23660 -12550 23705 -12430
rect 23825 -12550 23870 -12430
rect 23990 -12550 24015 -12430
rect 18485 -12595 24015 -12550
rect 18485 -12715 18510 -12595
rect 18630 -12715 18685 -12595
rect 18805 -12715 18850 -12595
rect 18970 -12715 19015 -12595
rect 19135 -12715 19180 -12595
rect 19300 -12715 19355 -12595
rect 19475 -12715 19520 -12595
rect 19640 -12715 19685 -12595
rect 19805 -12715 19850 -12595
rect 19970 -12715 20025 -12595
rect 20145 -12715 20190 -12595
rect 20310 -12715 20355 -12595
rect 20475 -12715 20520 -12595
rect 20640 -12715 20695 -12595
rect 20815 -12715 20860 -12595
rect 20980 -12715 21025 -12595
rect 21145 -12715 21190 -12595
rect 21310 -12715 21365 -12595
rect 21485 -12715 21530 -12595
rect 21650 -12715 21695 -12595
rect 21815 -12715 21860 -12595
rect 21980 -12715 22035 -12595
rect 22155 -12715 22200 -12595
rect 22320 -12715 22365 -12595
rect 22485 -12715 22530 -12595
rect 22650 -12715 22705 -12595
rect 22825 -12715 22870 -12595
rect 22990 -12715 23035 -12595
rect 23155 -12715 23200 -12595
rect 23320 -12715 23375 -12595
rect 23495 -12715 23540 -12595
rect 23660 -12715 23705 -12595
rect 23825 -12715 23870 -12595
rect 23990 -12715 24015 -12595
rect 18485 -12770 24015 -12715
rect 18485 -12890 18510 -12770
rect 18630 -12890 18685 -12770
rect 18805 -12890 18850 -12770
rect 18970 -12890 19015 -12770
rect 19135 -12890 19180 -12770
rect 19300 -12890 19355 -12770
rect 19475 -12890 19520 -12770
rect 19640 -12890 19685 -12770
rect 19805 -12890 19850 -12770
rect 19970 -12890 20025 -12770
rect 20145 -12890 20190 -12770
rect 20310 -12890 20355 -12770
rect 20475 -12890 20520 -12770
rect 20640 -12890 20695 -12770
rect 20815 -12890 20860 -12770
rect 20980 -12890 21025 -12770
rect 21145 -12890 21190 -12770
rect 21310 -12890 21365 -12770
rect 21485 -12890 21530 -12770
rect 21650 -12890 21695 -12770
rect 21815 -12890 21860 -12770
rect 21980 -12890 22035 -12770
rect 22155 -12890 22200 -12770
rect 22320 -12890 22365 -12770
rect 22485 -12890 22530 -12770
rect 22650 -12890 22705 -12770
rect 22825 -12890 22870 -12770
rect 22990 -12890 23035 -12770
rect 23155 -12890 23200 -12770
rect 23320 -12890 23375 -12770
rect 23495 -12890 23540 -12770
rect 23660 -12890 23705 -12770
rect 23825 -12890 23870 -12770
rect 23990 -12890 24015 -12770
rect 18485 -12935 24015 -12890
rect 18485 -13055 18510 -12935
rect 18630 -13055 18685 -12935
rect 18805 -13055 18850 -12935
rect 18970 -13055 19015 -12935
rect 19135 -13055 19180 -12935
rect 19300 -13055 19355 -12935
rect 19475 -13055 19520 -12935
rect 19640 -13055 19685 -12935
rect 19805 -13055 19850 -12935
rect 19970 -13055 20025 -12935
rect 20145 -13055 20190 -12935
rect 20310 -13055 20355 -12935
rect 20475 -13055 20520 -12935
rect 20640 -13055 20695 -12935
rect 20815 -13055 20860 -12935
rect 20980 -13055 21025 -12935
rect 21145 -13055 21190 -12935
rect 21310 -13055 21365 -12935
rect 21485 -13055 21530 -12935
rect 21650 -13055 21695 -12935
rect 21815 -13055 21860 -12935
rect 21980 -13055 22035 -12935
rect 22155 -13055 22200 -12935
rect 22320 -13055 22365 -12935
rect 22485 -13055 22530 -12935
rect 22650 -13055 22705 -12935
rect 22825 -13055 22870 -12935
rect 22990 -13055 23035 -12935
rect 23155 -13055 23200 -12935
rect 23320 -13055 23375 -12935
rect 23495 -13055 23540 -12935
rect 23660 -13055 23705 -12935
rect 23825 -13055 23870 -12935
rect 23990 -13055 24015 -12935
rect 18485 -13100 24015 -13055
rect 18485 -13220 18510 -13100
rect 18630 -13220 18685 -13100
rect 18805 -13220 18850 -13100
rect 18970 -13220 19015 -13100
rect 19135 -13220 19180 -13100
rect 19300 -13220 19355 -13100
rect 19475 -13220 19520 -13100
rect 19640 -13220 19685 -13100
rect 19805 -13220 19850 -13100
rect 19970 -13220 20025 -13100
rect 20145 -13220 20190 -13100
rect 20310 -13220 20355 -13100
rect 20475 -13220 20520 -13100
rect 20640 -13220 20695 -13100
rect 20815 -13220 20860 -13100
rect 20980 -13220 21025 -13100
rect 21145 -13220 21190 -13100
rect 21310 -13220 21365 -13100
rect 21485 -13220 21530 -13100
rect 21650 -13220 21695 -13100
rect 21815 -13220 21860 -13100
rect 21980 -13220 22035 -13100
rect 22155 -13220 22200 -13100
rect 22320 -13220 22365 -13100
rect 22485 -13220 22530 -13100
rect 22650 -13220 22705 -13100
rect 22825 -13220 22870 -13100
rect 22990 -13220 23035 -13100
rect 23155 -13220 23200 -13100
rect 23320 -13220 23375 -13100
rect 23495 -13220 23540 -13100
rect 23660 -13220 23705 -13100
rect 23825 -13220 23870 -13100
rect 23990 -13220 24015 -13100
rect 18485 -13265 24015 -13220
rect 18485 -13385 18510 -13265
rect 18630 -13385 18685 -13265
rect 18805 -13385 18850 -13265
rect 18970 -13385 19015 -13265
rect 19135 -13385 19180 -13265
rect 19300 -13385 19355 -13265
rect 19475 -13385 19520 -13265
rect 19640 -13385 19685 -13265
rect 19805 -13385 19850 -13265
rect 19970 -13385 20025 -13265
rect 20145 -13385 20190 -13265
rect 20310 -13385 20355 -13265
rect 20475 -13385 20520 -13265
rect 20640 -13385 20695 -13265
rect 20815 -13385 20860 -13265
rect 20980 -13385 21025 -13265
rect 21145 -13385 21190 -13265
rect 21310 -13385 21365 -13265
rect 21485 -13385 21530 -13265
rect 21650 -13385 21695 -13265
rect 21815 -13385 21860 -13265
rect 21980 -13385 22035 -13265
rect 22155 -13385 22200 -13265
rect 22320 -13385 22365 -13265
rect 22485 -13385 22530 -13265
rect 22650 -13385 22705 -13265
rect 22825 -13385 22870 -13265
rect 22990 -13385 23035 -13265
rect 23155 -13385 23200 -13265
rect 23320 -13385 23375 -13265
rect 23495 -13385 23540 -13265
rect 23660 -13385 23705 -13265
rect 23825 -13385 23870 -13265
rect 23990 -13385 24015 -13265
rect 18485 -13440 24015 -13385
rect 18485 -13560 18510 -13440
rect 18630 -13560 18685 -13440
rect 18805 -13560 18850 -13440
rect 18970 -13560 19015 -13440
rect 19135 -13560 19180 -13440
rect 19300 -13560 19355 -13440
rect 19475 -13560 19520 -13440
rect 19640 -13560 19685 -13440
rect 19805 -13560 19850 -13440
rect 19970 -13560 20025 -13440
rect 20145 -13560 20190 -13440
rect 20310 -13560 20355 -13440
rect 20475 -13560 20520 -13440
rect 20640 -13560 20695 -13440
rect 20815 -13560 20860 -13440
rect 20980 -13560 21025 -13440
rect 21145 -13560 21190 -13440
rect 21310 -13560 21365 -13440
rect 21485 -13560 21530 -13440
rect 21650 -13560 21695 -13440
rect 21815 -13560 21860 -13440
rect 21980 -13560 22035 -13440
rect 22155 -13560 22200 -13440
rect 22320 -13560 22365 -13440
rect 22485 -13560 22530 -13440
rect 22650 -13560 22705 -13440
rect 22825 -13560 22870 -13440
rect 22990 -13560 23035 -13440
rect 23155 -13560 23200 -13440
rect 23320 -13560 23375 -13440
rect 23495 -13560 23540 -13440
rect 23660 -13560 23705 -13440
rect 23825 -13560 23870 -13440
rect 23990 -13560 24015 -13440
rect 18485 -13605 24015 -13560
rect 18485 -13725 18510 -13605
rect 18630 -13725 18685 -13605
rect 18805 -13725 18850 -13605
rect 18970 -13725 19015 -13605
rect 19135 -13725 19180 -13605
rect 19300 -13725 19355 -13605
rect 19475 -13725 19520 -13605
rect 19640 -13725 19685 -13605
rect 19805 -13725 19850 -13605
rect 19970 -13725 20025 -13605
rect 20145 -13725 20190 -13605
rect 20310 -13725 20355 -13605
rect 20475 -13725 20520 -13605
rect 20640 -13725 20695 -13605
rect 20815 -13725 20860 -13605
rect 20980 -13725 21025 -13605
rect 21145 -13725 21190 -13605
rect 21310 -13725 21365 -13605
rect 21485 -13725 21530 -13605
rect 21650 -13725 21695 -13605
rect 21815 -13725 21860 -13605
rect 21980 -13725 22035 -13605
rect 22155 -13725 22200 -13605
rect 22320 -13725 22365 -13605
rect 22485 -13725 22530 -13605
rect 22650 -13725 22705 -13605
rect 22825 -13725 22870 -13605
rect 22990 -13725 23035 -13605
rect 23155 -13725 23200 -13605
rect 23320 -13725 23375 -13605
rect 23495 -13725 23540 -13605
rect 23660 -13725 23705 -13605
rect 23825 -13725 23870 -13605
rect 23990 -13725 24015 -13605
rect 18485 -13770 24015 -13725
rect 18485 -13890 18510 -13770
rect 18630 -13890 18685 -13770
rect 18805 -13890 18850 -13770
rect 18970 -13890 19015 -13770
rect 19135 -13890 19180 -13770
rect 19300 -13890 19355 -13770
rect 19475 -13890 19520 -13770
rect 19640 -13890 19685 -13770
rect 19805 -13890 19850 -13770
rect 19970 -13890 20025 -13770
rect 20145 -13890 20190 -13770
rect 20310 -13890 20355 -13770
rect 20475 -13890 20520 -13770
rect 20640 -13890 20695 -13770
rect 20815 -13890 20860 -13770
rect 20980 -13890 21025 -13770
rect 21145 -13890 21190 -13770
rect 21310 -13890 21365 -13770
rect 21485 -13890 21530 -13770
rect 21650 -13890 21695 -13770
rect 21815 -13890 21860 -13770
rect 21980 -13890 22035 -13770
rect 22155 -13890 22200 -13770
rect 22320 -13890 22365 -13770
rect 22485 -13890 22530 -13770
rect 22650 -13890 22705 -13770
rect 22825 -13890 22870 -13770
rect 22990 -13890 23035 -13770
rect 23155 -13890 23200 -13770
rect 23320 -13890 23375 -13770
rect 23495 -13890 23540 -13770
rect 23660 -13890 23705 -13770
rect 23825 -13890 23870 -13770
rect 23990 -13890 24015 -13770
rect 18485 -13935 24015 -13890
rect 18485 -14055 18510 -13935
rect 18630 -14055 18685 -13935
rect 18805 -14055 18850 -13935
rect 18970 -14055 19015 -13935
rect 19135 -14055 19180 -13935
rect 19300 -14055 19355 -13935
rect 19475 -14055 19520 -13935
rect 19640 -14055 19685 -13935
rect 19805 -14055 19850 -13935
rect 19970 -14055 20025 -13935
rect 20145 -14055 20190 -13935
rect 20310 -14055 20355 -13935
rect 20475 -14055 20520 -13935
rect 20640 -14055 20695 -13935
rect 20815 -14055 20860 -13935
rect 20980 -14055 21025 -13935
rect 21145 -14055 21190 -13935
rect 21310 -14055 21365 -13935
rect 21485 -14055 21530 -13935
rect 21650 -14055 21695 -13935
rect 21815 -14055 21860 -13935
rect 21980 -14055 22035 -13935
rect 22155 -14055 22200 -13935
rect 22320 -14055 22365 -13935
rect 22485 -14055 22530 -13935
rect 22650 -14055 22705 -13935
rect 22825 -14055 22870 -13935
rect 22990 -14055 23035 -13935
rect 23155 -14055 23200 -13935
rect 23320 -14055 23375 -13935
rect 23495 -14055 23540 -13935
rect 23660 -14055 23705 -13935
rect 23825 -14055 23870 -13935
rect 23990 -14055 24015 -13935
rect 18485 -14110 24015 -14055
rect 18485 -14230 18510 -14110
rect 18630 -14230 18685 -14110
rect 18805 -14230 18850 -14110
rect 18970 -14230 19015 -14110
rect 19135 -14230 19180 -14110
rect 19300 -14230 19355 -14110
rect 19475 -14230 19520 -14110
rect 19640 -14230 19685 -14110
rect 19805 -14230 19850 -14110
rect 19970 -14230 20025 -14110
rect 20145 -14230 20190 -14110
rect 20310 -14230 20355 -14110
rect 20475 -14230 20520 -14110
rect 20640 -14230 20695 -14110
rect 20815 -14230 20860 -14110
rect 20980 -14230 21025 -14110
rect 21145 -14230 21190 -14110
rect 21310 -14230 21365 -14110
rect 21485 -14230 21530 -14110
rect 21650 -14230 21695 -14110
rect 21815 -14230 21860 -14110
rect 21980 -14230 22035 -14110
rect 22155 -14230 22200 -14110
rect 22320 -14230 22365 -14110
rect 22485 -14230 22530 -14110
rect 22650 -14230 22705 -14110
rect 22825 -14230 22870 -14110
rect 22990 -14230 23035 -14110
rect 23155 -14230 23200 -14110
rect 23320 -14230 23375 -14110
rect 23495 -14230 23540 -14110
rect 23660 -14230 23705 -14110
rect 23825 -14230 23870 -14110
rect 23990 -14230 24015 -14110
rect 18485 -14275 24015 -14230
rect 18485 -14395 18510 -14275
rect 18630 -14395 18685 -14275
rect 18805 -14395 18850 -14275
rect 18970 -14395 19015 -14275
rect 19135 -14395 19180 -14275
rect 19300 -14395 19355 -14275
rect 19475 -14395 19520 -14275
rect 19640 -14395 19685 -14275
rect 19805 -14395 19850 -14275
rect 19970 -14395 20025 -14275
rect 20145 -14395 20190 -14275
rect 20310 -14395 20355 -14275
rect 20475 -14395 20520 -14275
rect 20640 -14395 20695 -14275
rect 20815 -14395 20860 -14275
rect 20980 -14395 21025 -14275
rect 21145 -14395 21190 -14275
rect 21310 -14395 21365 -14275
rect 21485 -14395 21530 -14275
rect 21650 -14395 21695 -14275
rect 21815 -14395 21860 -14275
rect 21980 -14395 22035 -14275
rect 22155 -14395 22200 -14275
rect 22320 -14395 22365 -14275
rect 22485 -14395 22530 -14275
rect 22650 -14395 22705 -14275
rect 22825 -14395 22870 -14275
rect 22990 -14395 23035 -14275
rect 23155 -14395 23200 -14275
rect 23320 -14395 23375 -14275
rect 23495 -14395 23540 -14275
rect 23660 -14395 23705 -14275
rect 23825 -14395 23870 -14275
rect 23990 -14395 24015 -14275
rect 18485 -14440 24015 -14395
rect 18485 -14560 18510 -14440
rect 18630 -14560 18685 -14440
rect 18805 -14560 18850 -14440
rect 18970 -14560 19015 -14440
rect 19135 -14560 19180 -14440
rect 19300 -14560 19355 -14440
rect 19475 -14560 19520 -14440
rect 19640 -14560 19685 -14440
rect 19805 -14560 19850 -14440
rect 19970 -14560 20025 -14440
rect 20145 -14560 20190 -14440
rect 20310 -14560 20355 -14440
rect 20475 -14560 20520 -14440
rect 20640 -14560 20695 -14440
rect 20815 -14560 20860 -14440
rect 20980 -14560 21025 -14440
rect 21145 -14560 21190 -14440
rect 21310 -14560 21365 -14440
rect 21485 -14560 21530 -14440
rect 21650 -14560 21695 -14440
rect 21815 -14560 21860 -14440
rect 21980 -14560 22035 -14440
rect 22155 -14560 22200 -14440
rect 22320 -14560 22365 -14440
rect 22485 -14560 22530 -14440
rect 22650 -14560 22705 -14440
rect 22825 -14560 22870 -14440
rect 22990 -14560 23035 -14440
rect 23155 -14560 23200 -14440
rect 23320 -14560 23375 -14440
rect 23495 -14560 23540 -14440
rect 23660 -14560 23705 -14440
rect 23825 -14560 23870 -14440
rect 23990 -14560 24015 -14440
rect 18485 -14605 24015 -14560
rect 18485 -14725 18510 -14605
rect 18630 -14725 18685 -14605
rect 18805 -14725 18850 -14605
rect 18970 -14725 19015 -14605
rect 19135 -14725 19180 -14605
rect 19300 -14725 19355 -14605
rect 19475 -14725 19520 -14605
rect 19640 -14725 19685 -14605
rect 19805 -14725 19850 -14605
rect 19970 -14725 20025 -14605
rect 20145 -14725 20190 -14605
rect 20310 -14725 20355 -14605
rect 20475 -14725 20520 -14605
rect 20640 -14725 20695 -14605
rect 20815 -14725 20860 -14605
rect 20980 -14725 21025 -14605
rect 21145 -14725 21190 -14605
rect 21310 -14725 21365 -14605
rect 21485 -14725 21530 -14605
rect 21650 -14725 21695 -14605
rect 21815 -14725 21860 -14605
rect 21980 -14725 22035 -14605
rect 22155 -14725 22200 -14605
rect 22320 -14725 22365 -14605
rect 22485 -14725 22530 -14605
rect 22650 -14725 22705 -14605
rect 22825 -14725 22870 -14605
rect 22990 -14725 23035 -14605
rect 23155 -14725 23200 -14605
rect 23320 -14725 23375 -14605
rect 23495 -14725 23540 -14605
rect 23660 -14725 23705 -14605
rect 23825 -14725 23870 -14605
rect 23990 -14725 24015 -14605
rect 18485 -14780 24015 -14725
rect 18485 -14900 18510 -14780
rect 18630 -14900 18685 -14780
rect 18805 -14900 18850 -14780
rect 18970 -14900 19015 -14780
rect 19135 -14900 19180 -14780
rect 19300 -14900 19355 -14780
rect 19475 -14900 19520 -14780
rect 19640 -14900 19685 -14780
rect 19805 -14900 19850 -14780
rect 19970 -14900 20025 -14780
rect 20145 -14900 20190 -14780
rect 20310 -14900 20355 -14780
rect 20475 -14900 20520 -14780
rect 20640 -14900 20695 -14780
rect 20815 -14900 20860 -14780
rect 20980 -14900 21025 -14780
rect 21145 -14900 21190 -14780
rect 21310 -14900 21365 -14780
rect 21485 -14900 21530 -14780
rect 21650 -14900 21695 -14780
rect 21815 -14900 21860 -14780
rect 21980 -14900 22035 -14780
rect 22155 -14900 22200 -14780
rect 22320 -14900 22365 -14780
rect 22485 -14900 22530 -14780
rect 22650 -14900 22705 -14780
rect 22825 -14900 22870 -14780
rect 22990 -14900 23035 -14780
rect 23155 -14900 23200 -14780
rect 23320 -14900 23375 -14780
rect 23495 -14900 23540 -14780
rect 23660 -14900 23705 -14780
rect 23825 -14900 23870 -14780
rect 23990 -14900 24015 -14780
rect 18485 -14945 24015 -14900
rect 18485 -15065 18510 -14945
rect 18630 -15065 18685 -14945
rect 18805 -15065 18850 -14945
rect 18970 -15065 19015 -14945
rect 19135 -15065 19180 -14945
rect 19300 -15065 19355 -14945
rect 19475 -15065 19520 -14945
rect 19640 -15065 19685 -14945
rect 19805 -15065 19850 -14945
rect 19970 -15065 20025 -14945
rect 20145 -15065 20190 -14945
rect 20310 -15065 20355 -14945
rect 20475 -15065 20520 -14945
rect 20640 -15065 20695 -14945
rect 20815 -15065 20860 -14945
rect 20980 -15065 21025 -14945
rect 21145 -15065 21190 -14945
rect 21310 -15065 21365 -14945
rect 21485 -15065 21530 -14945
rect 21650 -15065 21695 -14945
rect 21815 -15065 21860 -14945
rect 21980 -15065 22035 -14945
rect 22155 -15065 22200 -14945
rect 22320 -15065 22365 -14945
rect 22485 -15065 22530 -14945
rect 22650 -15065 22705 -14945
rect 22825 -15065 22870 -14945
rect 22990 -15065 23035 -14945
rect 23155 -15065 23200 -14945
rect 23320 -15065 23375 -14945
rect 23495 -15065 23540 -14945
rect 23660 -15065 23705 -14945
rect 23825 -15065 23870 -14945
rect 23990 -15065 24015 -14945
rect 18485 -15110 24015 -15065
rect 18485 -15230 18510 -15110
rect 18630 -15230 18685 -15110
rect 18805 -15230 18850 -15110
rect 18970 -15230 19015 -15110
rect 19135 -15230 19180 -15110
rect 19300 -15230 19355 -15110
rect 19475 -15230 19520 -15110
rect 19640 -15230 19685 -15110
rect 19805 -15230 19850 -15110
rect 19970 -15230 20025 -15110
rect 20145 -15230 20190 -15110
rect 20310 -15230 20355 -15110
rect 20475 -15230 20520 -15110
rect 20640 -15230 20695 -15110
rect 20815 -15230 20860 -15110
rect 20980 -15230 21025 -15110
rect 21145 -15230 21190 -15110
rect 21310 -15230 21365 -15110
rect 21485 -15230 21530 -15110
rect 21650 -15230 21695 -15110
rect 21815 -15230 21860 -15110
rect 21980 -15230 22035 -15110
rect 22155 -15230 22200 -15110
rect 22320 -15230 22365 -15110
rect 22485 -15230 22530 -15110
rect 22650 -15230 22705 -15110
rect 22825 -15230 22870 -15110
rect 22990 -15230 23035 -15110
rect 23155 -15230 23200 -15110
rect 23320 -15230 23375 -15110
rect 23495 -15230 23540 -15110
rect 23660 -15230 23705 -15110
rect 23825 -15230 23870 -15110
rect 23990 -15230 24015 -15110
rect 18485 -15275 24015 -15230
rect 18485 -15395 18510 -15275
rect 18630 -15395 18685 -15275
rect 18805 -15395 18850 -15275
rect 18970 -15395 19015 -15275
rect 19135 -15395 19180 -15275
rect 19300 -15395 19355 -15275
rect 19475 -15395 19520 -15275
rect 19640 -15395 19685 -15275
rect 19805 -15395 19850 -15275
rect 19970 -15395 20025 -15275
rect 20145 -15395 20190 -15275
rect 20310 -15395 20355 -15275
rect 20475 -15395 20520 -15275
rect 20640 -15395 20695 -15275
rect 20815 -15395 20860 -15275
rect 20980 -15395 21025 -15275
rect 21145 -15395 21190 -15275
rect 21310 -15395 21365 -15275
rect 21485 -15395 21530 -15275
rect 21650 -15395 21695 -15275
rect 21815 -15395 21860 -15275
rect 21980 -15395 22035 -15275
rect 22155 -15395 22200 -15275
rect 22320 -15395 22365 -15275
rect 22485 -15395 22530 -15275
rect 22650 -15395 22705 -15275
rect 22825 -15395 22870 -15275
rect 22990 -15395 23035 -15275
rect 23155 -15395 23200 -15275
rect 23320 -15395 23375 -15275
rect 23495 -15395 23540 -15275
rect 23660 -15395 23705 -15275
rect 23825 -15395 23870 -15275
rect 23990 -15395 24015 -15275
rect 18485 -15450 24015 -15395
rect 18485 -15535 18510 -15450
rect 18300 -15570 18510 -15535
rect 18630 -15570 18685 -15450
rect 18805 -15570 18850 -15450
rect 18970 -15570 19015 -15450
rect 19135 -15570 19180 -15450
rect 19300 -15570 19355 -15450
rect 19475 -15570 19520 -15450
rect 19640 -15570 19685 -15450
rect 19805 -15570 19850 -15450
rect 19970 -15570 20025 -15450
rect 20145 -15570 20190 -15450
rect 20310 -15570 20355 -15450
rect 20475 -15570 20520 -15450
rect 20640 -15570 20695 -15450
rect 20815 -15570 20860 -15450
rect 20980 -15570 21025 -15450
rect 21145 -15570 21190 -15450
rect 21310 -15570 21365 -15450
rect 21485 -15570 21530 -15450
rect 21650 -15570 21695 -15450
rect 21815 -15570 21860 -15450
rect 21980 -15570 22035 -15450
rect 22155 -15570 22200 -15450
rect 22320 -15570 22365 -15450
rect 22485 -15570 22530 -15450
rect 22650 -15570 22705 -15450
rect 22825 -15570 22870 -15450
rect 22990 -15570 23035 -15450
rect 23155 -15570 23200 -15450
rect 23320 -15570 23375 -15450
rect 23495 -15570 23540 -15450
rect 23660 -15570 23705 -15450
rect 23825 -15570 23870 -15450
rect 23990 -15535 24015 -15450
rect 24175 -10090 29705 -10065
rect 24175 -10210 24200 -10090
rect 24320 -10210 24375 -10090
rect 24495 -10210 24540 -10090
rect 24660 -10210 24705 -10090
rect 24825 -10210 24870 -10090
rect 24990 -10210 25045 -10090
rect 25165 -10210 25210 -10090
rect 25330 -10210 25375 -10090
rect 25495 -10210 25540 -10090
rect 25660 -10210 25715 -10090
rect 25835 -10210 25880 -10090
rect 26000 -10210 26045 -10090
rect 26165 -10210 26210 -10090
rect 26330 -10210 26385 -10090
rect 26505 -10210 26550 -10090
rect 26670 -10210 26715 -10090
rect 26835 -10210 26880 -10090
rect 27000 -10210 27055 -10090
rect 27175 -10210 27220 -10090
rect 27340 -10210 27385 -10090
rect 27505 -10210 27550 -10090
rect 27670 -10210 27725 -10090
rect 27845 -10210 27890 -10090
rect 28010 -10210 28055 -10090
rect 28175 -10210 28220 -10090
rect 28340 -10210 28395 -10090
rect 28515 -10210 28560 -10090
rect 28680 -10210 28725 -10090
rect 28845 -10210 28890 -10090
rect 29010 -10210 29065 -10090
rect 29185 -10210 29230 -10090
rect 29350 -10210 29395 -10090
rect 29515 -10210 29560 -10090
rect 29680 -10210 29705 -10090
rect 24175 -10255 29705 -10210
rect 24175 -10375 24200 -10255
rect 24320 -10375 24375 -10255
rect 24495 -10375 24540 -10255
rect 24660 -10375 24705 -10255
rect 24825 -10375 24870 -10255
rect 24990 -10375 25045 -10255
rect 25165 -10375 25210 -10255
rect 25330 -10375 25375 -10255
rect 25495 -10375 25540 -10255
rect 25660 -10375 25715 -10255
rect 25835 -10375 25880 -10255
rect 26000 -10375 26045 -10255
rect 26165 -10375 26210 -10255
rect 26330 -10375 26385 -10255
rect 26505 -10375 26550 -10255
rect 26670 -10375 26715 -10255
rect 26835 -10375 26880 -10255
rect 27000 -10375 27055 -10255
rect 27175 -10375 27220 -10255
rect 27340 -10375 27385 -10255
rect 27505 -10375 27550 -10255
rect 27670 -10375 27725 -10255
rect 27845 -10375 27890 -10255
rect 28010 -10375 28055 -10255
rect 28175 -10375 28220 -10255
rect 28340 -10375 28395 -10255
rect 28515 -10375 28560 -10255
rect 28680 -10375 28725 -10255
rect 28845 -10375 28890 -10255
rect 29010 -10375 29065 -10255
rect 29185 -10375 29230 -10255
rect 29350 -10375 29395 -10255
rect 29515 -10375 29560 -10255
rect 29680 -10375 29705 -10255
rect 24175 -10420 29705 -10375
rect 24175 -10540 24200 -10420
rect 24320 -10540 24375 -10420
rect 24495 -10540 24540 -10420
rect 24660 -10540 24705 -10420
rect 24825 -10540 24870 -10420
rect 24990 -10540 25045 -10420
rect 25165 -10540 25210 -10420
rect 25330 -10540 25375 -10420
rect 25495 -10540 25540 -10420
rect 25660 -10540 25715 -10420
rect 25835 -10540 25880 -10420
rect 26000 -10540 26045 -10420
rect 26165 -10540 26210 -10420
rect 26330 -10540 26385 -10420
rect 26505 -10540 26550 -10420
rect 26670 -10540 26715 -10420
rect 26835 -10540 26880 -10420
rect 27000 -10540 27055 -10420
rect 27175 -10540 27220 -10420
rect 27340 -10540 27385 -10420
rect 27505 -10540 27550 -10420
rect 27670 -10540 27725 -10420
rect 27845 -10540 27890 -10420
rect 28010 -10540 28055 -10420
rect 28175 -10540 28220 -10420
rect 28340 -10540 28395 -10420
rect 28515 -10540 28560 -10420
rect 28680 -10540 28725 -10420
rect 28845 -10540 28890 -10420
rect 29010 -10540 29065 -10420
rect 29185 -10540 29230 -10420
rect 29350 -10540 29395 -10420
rect 29515 -10540 29560 -10420
rect 29680 -10540 29705 -10420
rect 24175 -10585 29705 -10540
rect 24175 -10705 24200 -10585
rect 24320 -10705 24375 -10585
rect 24495 -10705 24540 -10585
rect 24660 -10705 24705 -10585
rect 24825 -10705 24870 -10585
rect 24990 -10705 25045 -10585
rect 25165 -10705 25210 -10585
rect 25330 -10705 25375 -10585
rect 25495 -10705 25540 -10585
rect 25660 -10705 25715 -10585
rect 25835 -10705 25880 -10585
rect 26000 -10705 26045 -10585
rect 26165 -10705 26210 -10585
rect 26330 -10705 26385 -10585
rect 26505 -10705 26550 -10585
rect 26670 -10705 26715 -10585
rect 26835 -10705 26880 -10585
rect 27000 -10705 27055 -10585
rect 27175 -10705 27220 -10585
rect 27340 -10705 27385 -10585
rect 27505 -10705 27550 -10585
rect 27670 -10705 27725 -10585
rect 27845 -10705 27890 -10585
rect 28010 -10705 28055 -10585
rect 28175 -10705 28220 -10585
rect 28340 -10705 28395 -10585
rect 28515 -10705 28560 -10585
rect 28680 -10705 28725 -10585
rect 28845 -10705 28890 -10585
rect 29010 -10705 29065 -10585
rect 29185 -10705 29230 -10585
rect 29350 -10705 29395 -10585
rect 29515 -10705 29560 -10585
rect 29680 -10705 29705 -10585
rect 24175 -10760 29705 -10705
rect 24175 -10880 24200 -10760
rect 24320 -10880 24375 -10760
rect 24495 -10880 24540 -10760
rect 24660 -10880 24705 -10760
rect 24825 -10880 24870 -10760
rect 24990 -10880 25045 -10760
rect 25165 -10880 25210 -10760
rect 25330 -10880 25375 -10760
rect 25495 -10880 25540 -10760
rect 25660 -10880 25715 -10760
rect 25835 -10880 25880 -10760
rect 26000 -10880 26045 -10760
rect 26165 -10880 26210 -10760
rect 26330 -10880 26385 -10760
rect 26505 -10880 26550 -10760
rect 26670 -10880 26715 -10760
rect 26835 -10880 26880 -10760
rect 27000 -10880 27055 -10760
rect 27175 -10880 27220 -10760
rect 27340 -10880 27385 -10760
rect 27505 -10880 27550 -10760
rect 27670 -10880 27725 -10760
rect 27845 -10880 27890 -10760
rect 28010 -10880 28055 -10760
rect 28175 -10880 28220 -10760
rect 28340 -10880 28395 -10760
rect 28515 -10880 28560 -10760
rect 28680 -10880 28725 -10760
rect 28845 -10880 28890 -10760
rect 29010 -10880 29065 -10760
rect 29185 -10880 29230 -10760
rect 29350 -10880 29395 -10760
rect 29515 -10880 29560 -10760
rect 29680 -10880 29705 -10760
rect 24175 -10925 29705 -10880
rect 24175 -11045 24200 -10925
rect 24320 -11045 24375 -10925
rect 24495 -11045 24540 -10925
rect 24660 -11045 24705 -10925
rect 24825 -11045 24870 -10925
rect 24990 -11045 25045 -10925
rect 25165 -11045 25210 -10925
rect 25330 -11045 25375 -10925
rect 25495 -11045 25540 -10925
rect 25660 -11045 25715 -10925
rect 25835 -11045 25880 -10925
rect 26000 -11045 26045 -10925
rect 26165 -11045 26210 -10925
rect 26330 -11045 26385 -10925
rect 26505 -11045 26550 -10925
rect 26670 -11045 26715 -10925
rect 26835 -11045 26880 -10925
rect 27000 -11045 27055 -10925
rect 27175 -11045 27220 -10925
rect 27340 -11045 27385 -10925
rect 27505 -11045 27550 -10925
rect 27670 -11045 27725 -10925
rect 27845 -11045 27890 -10925
rect 28010 -11045 28055 -10925
rect 28175 -11045 28220 -10925
rect 28340 -11045 28395 -10925
rect 28515 -11045 28560 -10925
rect 28680 -11045 28725 -10925
rect 28845 -11045 28890 -10925
rect 29010 -11045 29065 -10925
rect 29185 -11045 29230 -10925
rect 29350 -11045 29395 -10925
rect 29515 -11045 29560 -10925
rect 29680 -11045 29705 -10925
rect 24175 -11090 29705 -11045
rect 24175 -11210 24200 -11090
rect 24320 -11210 24375 -11090
rect 24495 -11210 24540 -11090
rect 24660 -11210 24705 -11090
rect 24825 -11210 24870 -11090
rect 24990 -11210 25045 -11090
rect 25165 -11210 25210 -11090
rect 25330 -11210 25375 -11090
rect 25495 -11210 25540 -11090
rect 25660 -11210 25715 -11090
rect 25835 -11210 25880 -11090
rect 26000 -11210 26045 -11090
rect 26165 -11210 26210 -11090
rect 26330 -11210 26385 -11090
rect 26505 -11210 26550 -11090
rect 26670 -11210 26715 -11090
rect 26835 -11210 26880 -11090
rect 27000 -11210 27055 -11090
rect 27175 -11210 27220 -11090
rect 27340 -11210 27385 -11090
rect 27505 -11210 27550 -11090
rect 27670 -11210 27725 -11090
rect 27845 -11210 27890 -11090
rect 28010 -11210 28055 -11090
rect 28175 -11210 28220 -11090
rect 28340 -11210 28395 -11090
rect 28515 -11210 28560 -11090
rect 28680 -11210 28725 -11090
rect 28845 -11210 28890 -11090
rect 29010 -11210 29065 -11090
rect 29185 -11210 29230 -11090
rect 29350 -11210 29395 -11090
rect 29515 -11210 29560 -11090
rect 29680 -11210 29705 -11090
rect 24175 -11255 29705 -11210
rect 24175 -11375 24200 -11255
rect 24320 -11375 24375 -11255
rect 24495 -11375 24540 -11255
rect 24660 -11375 24705 -11255
rect 24825 -11375 24870 -11255
rect 24990 -11375 25045 -11255
rect 25165 -11375 25210 -11255
rect 25330 -11375 25375 -11255
rect 25495 -11375 25540 -11255
rect 25660 -11375 25715 -11255
rect 25835 -11375 25880 -11255
rect 26000 -11375 26045 -11255
rect 26165 -11375 26210 -11255
rect 26330 -11375 26385 -11255
rect 26505 -11375 26550 -11255
rect 26670 -11375 26715 -11255
rect 26835 -11375 26880 -11255
rect 27000 -11375 27055 -11255
rect 27175 -11375 27220 -11255
rect 27340 -11375 27385 -11255
rect 27505 -11375 27550 -11255
rect 27670 -11375 27725 -11255
rect 27845 -11375 27890 -11255
rect 28010 -11375 28055 -11255
rect 28175 -11375 28220 -11255
rect 28340 -11375 28395 -11255
rect 28515 -11375 28560 -11255
rect 28680 -11375 28725 -11255
rect 28845 -11375 28890 -11255
rect 29010 -11375 29065 -11255
rect 29185 -11375 29230 -11255
rect 29350 -11375 29395 -11255
rect 29515 -11375 29560 -11255
rect 29680 -11375 29705 -11255
rect 24175 -11430 29705 -11375
rect 24175 -11550 24200 -11430
rect 24320 -11550 24375 -11430
rect 24495 -11550 24540 -11430
rect 24660 -11550 24705 -11430
rect 24825 -11550 24870 -11430
rect 24990 -11550 25045 -11430
rect 25165 -11550 25210 -11430
rect 25330 -11550 25375 -11430
rect 25495 -11550 25540 -11430
rect 25660 -11550 25715 -11430
rect 25835 -11550 25880 -11430
rect 26000 -11550 26045 -11430
rect 26165 -11550 26210 -11430
rect 26330 -11550 26385 -11430
rect 26505 -11550 26550 -11430
rect 26670 -11550 26715 -11430
rect 26835 -11550 26880 -11430
rect 27000 -11550 27055 -11430
rect 27175 -11550 27220 -11430
rect 27340 -11550 27385 -11430
rect 27505 -11550 27550 -11430
rect 27670 -11550 27725 -11430
rect 27845 -11550 27890 -11430
rect 28010 -11550 28055 -11430
rect 28175 -11550 28220 -11430
rect 28340 -11550 28395 -11430
rect 28515 -11550 28560 -11430
rect 28680 -11550 28725 -11430
rect 28845 -11550 28890 -11430
rect 29010 -11550 29065 -11430
rect 29185 -11550 29230 -11430
rect 29350 -11550 29395 -11430
rect 29515 -11550 29560 -11430
rect 29680 -11550 29705 -11430
rect 24175 -11595 29705 -11550
rect 24175 -11715 24200 -11595
rect 24320 -11715 24375 -11595
rect 24495 -11715 24540 -11595
rect 24660 -11715 24705 -11595
rect 24825 -11715 24870 -11595
rect 24990 -11715 25045 -11595
rect 25165 -11715 25210 -11595
rect 25330 -11715 25375 -11595
rect 25495 -11715 25540 -11595
rect 25660 -11715 25715 -11595
rect 25835 -11715 25880 -11595
rect 26000 -11715 26045 -11595
rect 26165 -11715 26210 -11595
rect 26330 -11715 26385 -11595
rect 26505 -11715 26550 -11595
rect 26670 -11715 26715 -11595
rect 26835 -11715 26880 -11595
rect 27000 -11715 27055 -11595
rect 27175 -11715 27220 -11595
rect 27340 -11715 27385 -11595
rect 27505 -11715 27550 -11595
rect 27670 -11715 27725 -11595
rect 27845 -11715 27890 -11595
rect 28010 -11715 28055 -11595
rect 28175 -11715 28220 -11595
rect 28340 -11715 28395 -11595
rect 28515 -11715 28560 -11595
rect 28680 -11715 28725 -11595
rect 28845 -11715 28890 -11595
rect 29010 -11715 29065 -11595
rect 29185 -11715 29230 -11595
rect 29350 -11715 29395 -11595
rect 29515 -11715 29560 -11595
rect 29680 -11715 29705 -11595
rect 24175 -11760 29705 -11715
rect 24175 -11880 24200 -11760
rect 24320 -11880 24375 -11760
rect 24495 -11880 24540 -11760
rect 24660 -11880 24705 -11760
rect 24825 -11880 24870 -11760
rect 24990 -11880 25045 -11760
rect 25165 -11880 25210 -11760
rect 25330 -11880 25375 -11760
rect 25495 -11880 25540 -11760
rect 25660 -11880 25715 -11760
rect 25835 -11880 25880 -11760
rect 26000 -11880 26045 -11760
rect 26165 -11880 26210 -11760
rect 26330 -11880 26385 -11760
rect 26505 -11880 26550 -11760
rect 26670 -11880 26715 -11760
rect 26835 -11880 26880 -11760
rect 27000 -11880 27055 -11760
rect 27175 -11880 27220 -11760
rect 27340 -11880 27385 -11760
rect 27505 -11880 27550 -11760
rect 27670 -11880 27725 -11760
rect 27845 -11880 27890 -11760
rect 28010 -11880 28055 -11760
rect 28175 -11880 28220 -11760
rect 28340 -11880 28395 -11760
rect 28515 -11880 28560 -11760
rect 28680 -11880 28725 -11760
rect 28845 -11880 28890 -11760
rect 29010 -11880 29065 -11760
rect 29185 -11880 29230 -11760
rect 29350 -11880 29395 -11760
rect 29515 -11880 29560 -11760
rect 29680 -11880 29705 -11760
rect 24175 -11925 29705 -11880
rect 24175 -12045 24200 -11925
rect 24320 -12045 24375 -11925
rect 24495 -12045 24540 -11925
rect 24660 -12045 24705 -11925
rect 24825 -12045 24870 -11925
rect 24990 -12045 25045 -11925
rect 25165 -12045 25210 -11925
rect 25330 -12045 25375 -11925
rect 25495 -12045 25540 -11925
rect 25660 -12045 25715 -11925
rect 25835 -12045 25880 -11925
rect 26000 -12045 26045 -11925
rect 26165 -12045 26210 -11925
rect 26330 -12045 26385 -11925
rect 26505 -12045 26550 -11925
rect 26670 -12045 26715 -11925
rect 26835 -12045 26880 -11925
rect 27000 -12045 27055 -11925
rect 27175 -12045 27220 -11925
rect 27340 -12045 27385 -11925
rect 27505 -12045 27550 -11925
rect 27670 -12045 27725 -11925
rect 27845 -12045 27890 -11925
rect 28010 -12045 28055 -11925
rect 28175 -12045 28220 -11925
rect 28340 -12045 28395 -11925
rect 28515 -12045 28560 -11925
rect 28680 -12045 28725 -11925
rect 28845 -12045 28890 -11925
rect 29010 -12045 29065 -11925
rect 29185 -12045 29230 -11925
rect 29350 -12045 29395 -11925
rect 29515 -12045 29560 -11925
rect 29680 -12045 29705 -11925
rect 24175 -12100 29705 -12045
rect 24175 -12220 24200 -12100
rect 24320 -12220 24375 -12100
rect 24495 -12220 24540 -12100
rect 24660 -12220 24705 -12100
rect 24825 -12220 24870 -12100
rect 24990 -12220 25045 -12100
rect 25165 -12220 25210 -12100
rect 25330 -12220 25375 -12100
rect 25495 -12220 25540 -12100
rect 25660 -12220 25715 -12100
rect 25835 -12220 25880 -12100
rect 26000 -12220 26045 -12100
rect 26165 -12220 26210 -12100
rect 26330 -12220 26385 -12100
rect 26505 -12220 26550 -12100
rect 26670 -12220 26715 -12100
rect 26835 -12220 26880 -12100
rect 27000 -12220 27055 -12100
rect 27175 -12220 27220 -12100
rect 27340 -12220 27385 -12100
rect 27505 -12220 27550 -12100
rect 27670 -12220 27725 -12100
rect 27845 -12220 27890 -12100
rect 28010 -12220 28055 -12100
rect 28175 -12220 28220 -12100
rect 28340 -12220 28395 -12100
rect 28515 -12220 28560 -12100
rect 28680 -12220 28725 -12100
rect 28845 -12220 28890 -12100
rect 29010 -12220 29065 -12100
rect 29185 -12220 29230 -12100
rect 29350 -12220 29395 -12100
rect 29515 -12220 29560 -12100
rect 29680 -12220 29705 -12100
rect 24175 -12265 29705 -12220
rect 24175 -12385 24200 -12265
rect 24320 -12385 24375 -12265
rect 24495 -12385 24540 -12265
rect 24660 -12385 24705 -12265
rect 24825 -12385 24870 -12265
rect 24990 -12385 25045 -12265
rect 25165 -12385 25210 -12265
rect 25330 -12385 25375 -12265
rect 25495 -12385 25540 -12265
rect 25660 -12385 25715 -12265
rect 25835 -12385 25880 -12265
rect 26000 -12385 26045 -12265
rect 26165 -12385 26210 -12265
rect 26330 -12385 26385 -12265
rect 26505 -12385 26550 -12265
rect 26670 -12385 26715 -12265
rect 26835 -12385 26880 -12265
rect 27000 -12385 27055 -12265
rect 27175 -12385 27220 -12265
rect 27340 -12385 27385 -12265
rect 27505 -12385 27550 -12265
rect 27670 -12385 27725 -12265
rect 27845 -12385 27890 -12265
rect 28010 -12385 28055 -12265
rect 28175 -12385 28220 -12265
rect 28340 -12385 28395 -12265
rect 28515 -12385 28560 -12265
rect 28680 -12385 28725 -12265
rect 28845 -12385 28890 -12265
rect 29010 -12385 29065 -12265
rect 29185 -12385 29230 -12265
rect 29350 -12385 29395 -12265
rect 29515 -12385 29560 -12265
rect 29680 -12385 29705 -12265
rect 24175 -12430 29705 -12385
rect 24175 -12550 24200 -12430
rect 24320 -12550 24375 -12430
rect 24495 -12550 24540 -12430
rect 24660 -12550 24705 -12430
rect 24825 -12550 24870 -12430
rect 24990 -12550 25045 -12430
rect 25165 -12550 25210 -12430
rect 25330 -12550 25375 -12430
rect 25495 -12550 25540 -12430
rect 25660 -12550 25715 -12430
rect 25835 -12550 25880 -12430
rect 26000 -12550 26045 -12430
rect 26165 -12550 26210 -12430
rect 26330 -12550 26385 -12430
rect 26505 -12550 26550 -12430
rect 26670 -12550 26715 -12430
rect 26835 -12550 26880 -12430
rect 27000 -12550 27055 -12430
rect 27175 -12550 27220 -12430
rect 27340 -12550 27385 -12430
rect 27505 -12550 27550 -12430
rect 27670 -12550 27725 -12430
rect 27845 -12550 27890 -12430
rect 28010 -12550 28055 -12430
rect 28175 -12550 28220 -12430
rect 28340 -12550 28395 -12430
rect 28515 -12550 28560 -12430
rect 28680 -12550 28725 -12430
rect 28845 -12550 28890 -12430
rect 29010 -12550 29065 -12430
rect 29185 -12550 29230 -12430
rect 29350 -12550 29395 -12430
rect 29515 -12550 29560 -12430
rect 29680 -12550 29705 -12430
rect 24175 -12595 29705 -12550
rect 24175 -12715 24200 -12595
rect 24320 -12715 24375 -12595
rect 24495 -12715 24540 -12595
rect 24660 -12715 24705 -12595
rect 24825 -12715 24870 -12595
rect 24990 -12715 25045 -12595
rect 25165 -12715 25210 -12595
rect 25330 -12715 25375 -12595
rect 25495 -12715 25540 -12595
rect 25660 -12715 25715 -12595
rect 25835 -12715 25880 -12595
rect 26000 -12715 26045 -12595
rect 26165 -12715 26210 -12595
rect 26330 -12715 26385 -12595
rect 26505 -12715 26550 -12595
rect 26670 -12715 26715 -12595
rect 26835 -12715 26880 -12595
rect 27000 -12715 27055 -12595
rect 27175 -12715 27220 -12595
rect 27340 -12715 27385 -12595
rect 27505 -12715 27550 -12595
rect 27670 -12715 27725 -12595
rect 27845 -12715 27890 -12595
rect 28010 -12715 28055 -12595
rect 28175 -12715 28220 -12595
rect 28340 -12715 28395 -12595
rect 28515 -12715 28560 -12595
rect 28680 -12715 28725 -12595
rect 28845 -12715 28890 -12595
rect 29010 -12715 29065 -12595
rect 29185 -12715 29230 -12595
rect 29350 -12715 29395 -12595
rect 29515 -12715 29560 -12595
rect 29680 -12715 29705 -12595
rect 24175 -12770 29705 -12715
rect 24175 -12890 24200 -12770
rect 24320 -12890 24375 -12770
rect 24495 -12890 24540 -12770
rect 24660 -12890 24705 -12770
rect 24825 -12890 24870 -12770
rect 24990 -12890 25045 -12770
rect 25165 -12890 25210 -12770
rect 25330 -12890 25375 -12770
rect 25495 -12890 25540 -12770
rect 25660 -12890 25715 -12770
rect 25835 -12890 25880 -12770
rect 26000 -12890 26045 -12770
rect 26165 -12890 26210 -12770
rect 26330 -12890 26385 -12770
rect 26505 -12890 26550 -12770
rect 26670 -12890 26715 -12770
rect 26835 -12890 26880 -12770
rect 27000 -12890 27055 -12770
rect 27175 -12890 27220 -12770
rect 27340 -12890 27385 -12770
rect 27505 -12890 27550 -12770
rect 27670 -12890 27725 -12770
rect 27845 -12890 27890 -12770
rect 28010 -12890 28055 -12770
rect 28175 -12890 28220 -12770
rect 28340 -12890 28395 -12770
rect 28515 -12890 28560 -12770
rect 28680 -12890 28725 -12770
rect 28845 -12890 28890 -12770
rect 29010 -12890 29065 -12770
rect 29185 -12890 29230 -12770
rect 29350 -12890 29395 -12770
rect 29515 -12890 29560 -12770
rect 29680 -12890 29705 -12770
rect 24175 -12935 29705 -12890
rect 24175 -13055 24200 -12935
rect 24320 -13055 24375 -12935
rect 24495 -13055 24540 -12935
rect 24660 -13055 24705 -12935
rect 24825 -13055 24870 -12935
rect 24990 -13055 25045 -12935
rect 25165 -13055 25210 -12935
rect 25330 -13055 25375 -12935
rect 25495 -13055 25540 -12935
rect 25660 -13055 25715 -12935
rect 25835 -13055 25880 -12935
rect 26000 -13055 26045 -12935
rect 26165 -13055 26210 -12935
rect 26330 -13055 26385 -12935
rect 26505 -13055 26550 -12935
rect 26670 -13055 26715 -12935
rect 26835 -13055 26880 -12935
rect 27000 -13055 27055 -12935
rect 27175 -13055 27220 -12935
rect 27340 -13055 27385 -12935
rect 27505 -13055 27550 -12935
rect 27670 -13055 27725 -12935
rect 27845 -13055 27890 -12935
rect 28010 -13055 28055 -12935
rect 28175 -13055 28220 -12935
rect 28340 -13055 28395 -12935
rect 28515 -13055 28560 -12935
rect 28680 -13055 28725 -12935
rect 28845 -13055 28890 -12935
rect 29010 -13055 29065 -12935
rect 29185 -13055 29230 -12935
rect 29350 -13055 29395 -12935
rect 29515 -13055 29560 -12935
rect 29680 -13055 29705 -12935
rect 24175 -13100 29705 -13055
rect 24175 -13220 24200 -13100
rect 24320 -13220 24375 -13100
rect 24495 -13220 24540 -13100
rect 24660 -13220 24705 -13100
rect 24825 -13220 24870 -13100
rect 24990 -13220 25045 -13100
rect 25165 -13220 25210 -13100
rect 25330 -13220 25375 -13100
rect 25495 -13220 25540 -13100
rect 25660 -13220 25715 -13100
rect 25835 -13220 25880 -13100
rect 26000 -13220 26045 -13100
rect 26165 -13220 26210 -13100
rect 26330 -13220 26385 -13100
rect 26505 -13220 26550 -13100
rect 26670 -13220 26715 -13100
rect 26835 -13220 26880 -13100
rect 27000 -13220 27055 -13100
rect 27175 -13220 27220 -13100
rect 27340 -13220 27385 -13100
rect 27505 -13220 27550 -13100
rect 27670 -13220 27725 -13100
rect 27845 -13220 27890 -13100
rect 28010 -13220 28055 -13100
rect 28175 -13220 28220 -13100
rect 28340 -13220 28395 -13100
rect 28515 -13220 28560 -13100
rect 28680 -13220 28725 -13100
rect 28845 -13220 28890 -13100
rect 29010 -13220 29065 -13100
rect 29185 -13220 29230 -13100
rect 29350 -13220 29395 -13100
rect 29515 -13220 29560 -13100
rect 29680 -13220 29705 -13100
rect 24175 -13265 29705 -13220
rect 24175 -13385 24200 -13265
rect 24320 -13385 24375 -13265
rect 24495 -13385 24540 -13265
rect 24660 -13385 24705 -13265
rect 24825 -13385 24870 -13265
rect 24990 -13385 25045 -13265
rect 25165 -13385 25210 -13265
rect 25330 -13385 25375 -13265
rect 25495 -13385 25540 -13265
rect 25660 -13385 25715 -13265
rect 25835 -13385 25880 -13265
rect 26000 -13385 26045 -13265
rect 26165 -13385 26210 -13265
rect 26330 -13385 26385 -13265
rect 26505 -13385 26550 -13265
rect 26670 -13385 26715 -13265
rect 26835 -13385 26880 -13265
rect 27000 -13385 27055 -13265
rect 27175 -13385 27220 -13265
rect 27340 -13385 27385 -13265
rect 27505 -13385 27550 -13265
rect 27670 -13385 27725 -13265
rect 27845 -13385 27890 -13265
rect 28010 -13385 28055 -13265
rect 28175 -13385 28220 -13265
rect 28340 -13385 28395 -13265
rect 28515 -13385 28560 -13265
rect 28680 -13385 28725 -13265
rect 28845 -13385 28890 -13265
rect 29010 -13385 29065 -13265
rect 29185 -13385 29230 -13265
rect 29350 -13385 29395 -13265
rect 29515 -13385 29560 -13265
rect 29680 -13385 29705 -13265
rect 24175 -13440 29705 -13385
rect 24175 -13560 24200 -13440
rect 24320 -13560 24375 -13440
rect 24495 -13560 24540 -13440
rect 24660 -13560 24705 -13440
rect 24825 -13560 24870 -13440
rect 24990 -13560 25045 -13440
rect 25165 -13560 25210 -13440
rect 25330 -13560 25375 -13440
rect 25495 -13560 25540 -13440
rect 25660 -13560 25715 -13440
rect 25835 -13560 25880 -13440
rect 26000 -13560 26045 -13440
rect 26165 -13560 26210 -13440
rect 26330 -13560 26385 -13440
rect 26505 -13560 26550 -13440
rect 26670 -13560 26715 -13440
rect 26835 -13560 26880 -13440
rect 27000 -13560 27055 -13440
rect 27175 -13560 27220 -13440
rect 27340 -13560 27385 -13440
rect 27505 -13560 27550 -13440
rect 27670 -13560 27725 -13440
rect 27845 -13560 27890 -13440
rect 28010 -13560 28055 -13440
rect 28175 -13560 28220 -13440
rect 28340 -13560 28395 -13440
rect 28515 -13560 28560 -13440
rect 28680 -13560 28725 -13440
rect 28845 -13560 28890 -13440
rect 29010 -13560 29065 -13440
rect 29185 -13560 29230 -13440
rect 29350 -13560 29395 -13440
rect 29515 -13560 29560 -13440
rect 29680 -13560 29705 -13440
rect 24175 -13605 29705 -13560
rect 24175 -13725 24200 -13605
rect 24320 -13725 24375 -13605
rect 24495 -13725 24540 -13605
rect 24660 -13725 24705 -13605
rect 24825 -13725 24870 -13605
rect 24990 -13725 25045 -13605
rect 25165 -13725 25210 -13605
rect 25330 -13725 25375 -13605
rect 25495 -13725 25540 -13605
rect 25660 -13725 25715 -13605
rect 25835 -13725 25880 -13605
rect 26000 -13725 26045 -13605
rect 26165 -13725 26210 -13605
rect 26330 -13725 26385 -13605
rect 26505 -13725 26550 -13605
rect 26670 -13725 26715 -13605
rect 26835 -13725 26880 -13605
rect 27000 -13725 27055 -13605
rect 27175 -13725 27220 -13605
rect 27340 -13725 27385 -13605
rect 27505 -13725 27550 -13605
rect 27670 -13725 27725 -13605
rect 27845 -13725 27890 -13605
rect 28010 -13725 28055 -13605
rect 28175 -13725 28220 -13605
rect 28340 -13725 28395 -13605
rect 28515 -13725 28560 -13605
rect 28680 -13725 28725 -13605
rect 28845 -13725 28890 -13605
rect 29010 -13725 29065 -13605
rect 29185 -13725 29230 -13605
rect 29350 -13725 29395 -13605
rect 29515 -13725 29560 -13605
rect 29680 -13725 29705 -13605
rect 24175 -13770 29705 -13725
rect 24175 -13890 24200 -13770
rect 24320 -13890 24375 -13770
rect 24495 -13890 24540 -13770
rect 24660 -13890 24705 -13770
rect 24825 -13890 24870 -13770
rect 24990 -13890 25045 -13770
rect 25165 -13890 25210 -13770
rect 25330 -13890 25375 -13770
rect 25495 -13890 25540 -13770
rect 25660 -13890 25715 -13770
rect 25835 -13890 25880 -13770
rect 26000 -13890 26045 -13770
rect 26165 -13890 26210 -13770
rect 26330 -13890 26385 -13770
rect 26505 -13890 26550 -13770
rect 26670 -13890 26715 -13770
rect 26835 -13890 26880 -13770
rect 27000 -13890 27055 -13770
rect 27175 -13890 27220 -13770
rect 27340 -13890 27385 -13770
rect 27505 -13890 27550 -13770
rect 27670 -13890 27725 -13770
rect 27845 -13890 27890 -13770
rect 28010 -13890 28055 -13770
rect 28175 -13890 28220 -13770
rect 28340 -13890 28395 -13770
rect 28515 -13890 28560 -13770
rect 28680 -13890 28725 -13770
rect 28845 -13890 28890 -13770
rect 29010 -13890 29065 -13770
rect 29185 -13890 29230 -13770
rect 29350 -13890 29395 -13770
rect 29515 -13890 29560 -13770
rect 29680 -13890 29705 -13770
rect 24175 -13935 29705 -13890
rect 24175 -14055 24200 -13935
rect 24320 -14055 24375 -13935
rect 24495 -14055 24540 -13935
rect 24660 -14055 24705 -13935
rect 24825 -14055 24870 -13935
rect 24990 -14055 25045 -13935
rect 25165 -14055 25210 -13935
rect 25330 -14055 25375 -13935
rect 25495 -14055 25540 -13935
rect 25660 -14055 25715 -13935
rect 25835 -14055 25880 -13935
rect 26000 -14055 26045 -13935
rect 26165 -14055 26210 -13935
rect 26330 -14055 26385 -13935
rect 26505 -14055 26550 -13935
rect 26670 -14055 26715 -13935
rect 26835 -14055 26880 -13935
rect 27000 -14055 27055 -13935
rect 27175 -14055 27220 -13935
rect 27340 -14055 27385 -13935
rect 27505 -14055 27550 -13935
rect 27670 -14055 27725 -13935
rect 27845 -14055 27890 -13935
rect 28010 -14055 28055 -13935
rect 28175 -14055 28220 -13935
rect 28340 -14055 28395 -13935
rect 28515 -14055 28560 -13935
rect 28680 -14055 28725 -13935
rect 28845 -14055 28890 -13935
rect 29010 -14055 29065 -13935
rect 29185 -14055 29230 -13935
rect 29350 -14055 29395 -13935
rect 29515 -14055 29560 -13935
rect 29680 -14055 29705 -13935
rect 24175 -14110 29705 -14055
rect 24175 -14230 24200 -14110
rect 24320 -14230 24375 -14110
rect 24495 -14230 24540 -14110
rect 24660 -14230 24705 -14110
rect 24825 -14230 24870 -14110
rect 24990 -14230 25045 -14110
rect 25165 -14230 25210 -14110
rect 25330 -14230 25375 -14110
rect 25495 -14230 25540 -14110
rect 25660 -14230 25715 -14110
rect 25835 -14230 25880 -14110
rect 26000 -14230 26045 -14110
rect 26165 -14230 26210 -14110
rect 26330 -14230 26385 -14110
rect 26505 -14230 26550 -14110
rect 26670 -14230 26715 -14110
rect 26835 -14230 26880 -14110
rect 27000 -14230 27055 -14110
rect 27175 -14230 27220 -14110
rect 27340 -14230 27385 -14110
rect 27505 -14230 27550 -14110
rect 27670 -14230 27725 -14110
rect 27845 -14230 27890 -14110
rect 28010 -14230 28055 -14110
rect 28175 -14230 28220 -14110
rect 28340 -14230 28395 -14110
rect 28515 -14230 28560 -14110
rect 28680 -14230 28725 -14110
rect 28845 -14230 28890 -14110
rect 29010 -14230 29065 -14110
rect 29185 -14230 29230 -14110
rect 29350 -14230 29395 -14110
rect 29515 -14230 29560 -14110
rect 29680 -14230 29705 -14110
rect 24175 -14275 29705 -14230
rect 24175 -14395 24200 -14275
rect 24320 -14395 24375 -14275
rect 24495 -14395 24540 -14275
rect 24660 -14395 24705 -14275
rect 24825 -14395 24870 -14275
rect 24990 -14395 25045 -14275
rect 25165 -14395 25210 -14275
rect 25330 -14395 25375 -14275
rect 25495 -14395 25540 -14275
rect 25660 -14395 25715 -14275
rect 25835 -14395 25880 -14275
rect 26000 -14395 26045 -14275
rect 26165 -14395 26210 -14275
rect 26330 -14395 26385 -14275
rect 26505 -14395 26550 -14275
rect 26670 -14395 26715 -14275
rect 26835 -14395 26880 -14275
rect 27000 -14395 27055 -14275
rect 27175 -14395 27220 -14275
rect 27340 -14395 27385 -14275
rect 27505 -14395 27550 -14275
rect 27670 -14395 27725 -14275
rect 27845 -14395 27890 -14275
rect 28010 -14395 28055 -14275
rect 28175 -14395 28220 -14275
rect 28340 -14395 28395 -14275
rect 28515 -14395 28560 -14275
rect 28680 -14395 28725 -14275
rect 28845 -14395 28890 -14275
rect 29010 -14395 29065 -14275
rect 29185 -14395 29230 -14275
rect 29350 -14395 29395 -14275
rect 29515 -14395 29560 -14275
rect 29680 -14395 29705 -14275
rect 24175 -14440 29705 -14395
rect 24175 -14560 24200 -14440
rect 24320 -14560 24375 -14440
rect 24495 -14560 24540 -14440
rect 24660 -14560 24705 -14440
rect 24825 -14560 24870 -14440
rect 24990 -14560 25045 -14440
rect 25165 -14560 25210 -14440
rect 25330 -14560 25375 -14440
rect 25495 -14560 25540 -14440
rect 25660 -14560 25715 -14440
rect 25835 -14560 25880 -14440
rect 26000 -14560 26045 -14440
rect 26165 -14560 26210 -14440
rect 26330 -14560 26385 -14440
rect 26505 -14560 26550 -14440
rect 26670 -14560 26715 -14440
rect 26835 -14560 26880 -14440
rect 27000 -14560 27055 -14440
rect 27175 -14560 27220 -14440
rect 27340 -14560 27385 -14440
rect 27505 -14560 27550 -14440
rect 27670 -14560 27725 -14440
rect 27845 -14560 27890 -14440
rect 28010 -14560 28055 -14440
rect 28175 -14560 28220 -14440
rect 28340 -14560 28395 -14440
rect 28515 -14560 28560 -14440
rect 28680 -14560 28725 -14440
rect 28845 -14560 28890 -14440
rect 29010 -14560 29065 -14440
rect 29185 -14560 29230 -14440
rect 29350 -14560 29395 -14440
rect 29515 -14560 29560 -14440
rect 29680 -14560 29705 -14440
rect 24175 -14605 29705 -14560
rect 24175 -14725 24200 -14605
rect 24320 -14725 24375 -14605
rect 24495 -14725 24540 -14605
rect 24660 -14725 24705 -14605
rect 24825 -14725 24870 -14605
rect 24990 -14725 25045 -14605
rect 25165 -14725 25210 -14605
rect 25330 -14725 25375 -14605
rect 25495 -14725 25540 -14605
rect 25660 -14725 25715 -14605
rect 25835 -14725 25880 -14605
rect 26000 -14725 26045 -14605
rect 26165 -14725 26210 -14605
rect 26330 -14725 26385 -14605
rect 26505 -14725 26550 -14605
rect 26670 -14725 26715 -14605
rect 26835 -14725 26880 -14605
rect 27000 -14725 27055 -14605
rect 27175 -14725 27220 -14605
rect 27340 -14725 27385 -14605
rect 27505 -14725 27550 -14605
rect 27670 -14725 27725 -14605
rect 27845 -14725 27890 -14605
rect 28010 -14725 28055 -14605
rect 28175 -14725 28220 -14605
rect 28340 -14725 28395 -14605
rect 28515 -14725 28560 -14605
rect 28680 -14725 28725 -14605
rect 28845 -14725 28890 -14605
rect 29010 -14725 29065 -14605
rect 29185 -14725 29230 -14605
rect 29350 -14725 29395 -14605
rect 29515 -14725 29560 -14605
rect 29680 -14725 29705 -14605
rect 24175 -14780 29705 -14725
rect 24175 -14900 24200 -14780
rect 24320 -14900 24375 -14780
rect 24495 -14900 24540 -14780
rect 24660 -14900 24705 -14780
rect 24825 -14900 24870 -14780
rect 24990 -14900 25045 -14780
rect 25165 -14900 25210 -14780
rect 25330 -14900 25375 -14780
rect 25495 -14900 25540 -14780
rect 25660 -14900 25715 -14780
rect 25835 -14900 25880 -14780
rect 26000 -14900 26045 -14780
rect 26165 -14900 26210 -14780
rect 26330 -14900 26385 -14780
rect 26505 -14900 26550 -14780
rect 26670 -14900 26715 -14780
rect 26835 -14900 26880 -14780
rect 27000 -14900 27055 -14780
rect 27175 -14900 27220 -14780
rect 27340 -14900 27385 -14780
rect 27505 -14900 27550 -14780
rect 27670 -14900 27725 -14780
rect 27845 -14900 27890 -14780
rect 28010 -14900 28055 -14780
rect 28175 -14900 28220 -14780
rect 28340 -14900 28395 -14780
rect 28515 -14900 28560 -14780
rect 28680 -14900 28725 -14780
rect 28845 -14900 28890 -14780
rect 29010 -14900 29065 -14780
rect 29185 -14900 29230 -14780
rect 29350 -14900 29395 -14780
rect 29515 -14900 29560 -14780
rect 29680 -14900 29705 -14780
rect 24175 -14945 29705 -14900
rect 24175 -15065 24200 -14945
rect 24320 -15065 24375 -14945
rect 24495 -15065 24540 -14945
rect 24660 -15065 24705 -14945
rect 24825 -15065 24870 -14945
rect 24990 -15065 25045 -14945
rect 25165 -15065 25210 -14945
rect 25330 -15065 25375 -14945
rect 25495 -15065 25540 -14945
rect 25660 -15065 25715 -14945
rect 25835 -15065 25880 -14945
rect 26000 -15065 26045 -14945
rect 26165 -15065 26210 -14945
rect 26330 -15065 26385 -14945
rect 26505 -15065 26550 -14945
rect 26670 -15065 26715 -14945
rect 26835 -15065 26880 -14945
rect 27000 -15065 27055 -14945
rect 27175 -15065 27220 -14945
rect 27340 -15065 27385 -14945
rect 27505 -15065 27550 -14945
rect 27670 -15065 27725 -14945
rect 27845 -15065 27890 -14945
rect 28010 -15065 28055 -14945
rect 28175 -15065 28220 -14945
rect 28340 -15065 28395 -14945
rect 28515 -15065 28560 -14945
rect 28680 -15065 28725 -14945
rect 28845 -15065 28890 -14945
rect 29010 -15065 29065 -14945
rect 29185 -15065 29230 -14945
rect 29350 -15065 29395 -14945
rect 29515 -15065 29560 -14945
rect 29680 -15065 29705 -14945
rect 24175 -15110 29705 -15065
rect 24175 -15230 24200 -15110
rect 24320 -15230 24375 -15110
rect 24495 -15230 24540 -15110
rect 24660 -15230 24705 -15110
rect 24825 -15230 24870 -15110
rect 24990 -15230 25045 -15110
rect 25165 -15230 25210 -15110
rect 25330 -15230 25375 -15110
rect 25495 -15230 25540 -15110
rect 25660 -15230 25715 -15110
rect 25835 -15230 25880 -15110
rect 26000 -15230 26045 -15110
rect 26165 -15230 26210 -15110
rect 26330 -15230 26385 -15110
rect 26505 -15230 26550 -15110
rect 26670 -15230 26715 -15110
rect 26835 -15230 26880 -15110
rect 27000 -15230 27055 -15110
rect 27175 -15230 27220 -15110
rect 27340 -15230 27385 -15110
rect 27505 -15230 27550 -15110
rect 27670 -15230 27725 -15110
rect 27845 -15230 27890 -15110
rect 28010 -15230 28055 -15110
rect 28175 -15230 28220 -15110
rect 28340 -15230 28395 -15110
rect 28515 -15230 28560 -15110
rect 28680 -15230 28725 -15110
rect 28845 -15230 28890 -15110
rect 29010 -15230 29065 -15110
rect 29185 -15230 29230 -15110
rect 29350 -15230 29395 -15110
rect 29515 -15230 29560 -15110
rect 29680 -15230 29705 -15110
rect 24175 -15275 29705 -15230
rect 24175 -15395 24200 -15275
rect 24320 -15395 24375 -15275
rect 24495 -15395 24540 -15275
rect 24660 -15395 24705 -15275
rect 24825 -15395 24870 -15275
rect 24990 -15395 25045 -15275
rect 25165 -15395 25210 -15275
rect 25330 -15395 25375 -15275
rect 25495 -15395 25540 -15275
rect 25660 -15395 25715 -15275
rect 25835 -15395 25880 -15275
rect 26000 -15395 26045 -15275
rect 26165 -15395 26210 -15275
rect 26330 -15395 26385 -15275
rect 26505 -15395 26550 -15275
rect 26670 -15395 26715 -15275
rect 26835 -15395 26880 -15275
rect 27000 -15395 27055 -15275
rect 27175 -15395 27220 -15275
rect 27340 -15395 27385 -15275
rect 27505 -15395 27550 -15275
rect 27670 -15395 27725 -15275
rect 27845 -15395 27890 -15275
rect 28010 -15395 28055 -15275
rect 28175 -15395 28220 -15275
rect 28340 -15395 28395 -15275
rect 28515 -15395 28560 -15275
rect 28680 -15395 28725 -15275
rect 28845 -15395 28890 -15275
rect 29010 -15395 29065 -15275
rect 29185 -15395 29230 -15275
rect 29350 -15395 29395 -15275
rect 29515 -15395 29560 -15275
rect 29680 -15395 29705 -15275
rect 24175 -15450 29705 -15395
rect 24175 -15535 24200 -15450
rect 23990 -15570 24200 -15535
rect 24320 -15570 24375 -15450
rect 24495 -15570 24540 -15450
rect 24660 -15570 24705 -15450
rect 24825 -15570 24870 -15450
rect 24990 -15570 25045 -15450
rect 25165 -15570 25210 -15450
rect 25330 -15570 25375 -15450
rect 25495 -15570 25540 -15450
rect 25660 -15570 25715 -15450
rect 25835 -15570 25880 -15450
rect 26000 -15570 26045 -15450
rect 26165 -15570 26210 -15450
rect 26330 -15570 26385 -15450
rect 26505 -15570 26550 -15450
rect 26670 -15570 26715 -15450
rect 26835 -15570 26880 -15450
rect 27000 -15570 27055 -15450
rect 27175 -15570 27220 -15450
rect 27340 -15570 27385 -15450
rect 27505 -15570 27550 -15450
rect 27670 -15570 27725 -15450
rect 27845 -15570 27890 -15450
rect 28010 -15570 28055 -15450
rect 28175 -15570 28220 -15450
rect 28340 -15570 28395 -15450
rect 28515 -15570 28560 -15450
rect 28680 -15570 28725 -15450
rect 28845 -15570 28890 -15450
rect 29010 -15570 29065 -15450
rect 29185 -15570 29230 -15450
rect 29350 -15570 29395 -15450
rect 29515 -15570 29560 -15450
rect 29680 -15570 29705 -15450
rect 7105 -15595 29705 -15570
<< via4 >>
rect 7170 1470 7290 1590
rect 7335 1470 7455 1590
rect 7500 1470 7620 1590
rect 7665 1470 7785 1590
rect 7830 1470 7950 1590
rect 7995 1470 8115 1590
rect 8160 1470 8280 1590
rect 8325 1470 8445 1590
rect 8490 1470 8610 1590
rect 8655 1470 8775 1590
rect 8820 1470 8940 1590
rect 8985 1470 9105 1590
rect 9150 1470 9270 1590
rect 9315 1470 9435 1590
rect 9480 1470 9600 1590
rect 9645 1470 9765 1590
rect 9810 1470 9930 1590
rect 9975 1470 10095 1590
rect 10140 1470 10260 1590
rect 10305 1470 10425 1590
rect 10470 1470 10590 1590
rect 10635 1470 10755 1590
rect 10800 1470 10920 1590
rect 10965 1470 11085 1590
rect 11130 1470 11250 1590
rect 11295 1470 11415 1590
rect 11460 1470 11580 1590
rect 11625 1470 11745 1590
rect 11790 1470 11910 1590
rect 11955 1470 12075 1590
rect 12120 1470 12240 1590
rect 12285 1470 12405 1590
rect 12450 1470 12570 1590
rect 12860 1470 12980 1590
rect 13025 1470 13145 1590
rect 13190 1470 13310 1590
rect 13355 1470 13475 1590
rect 13520 1470 13640 1590
rect 13685 1470 13805 1590
rect 13850 1470 13970 1590
rect 14015 1470 14135 1590
rect 14180 1470 14300 1590
rect 14345 1470 14465 1590
rect 14510 1470 14630 1590
rect 14675 1470 14795 1590
rect 14840 1470 14960 1590
rect 15005 1470 15125 1590
rect 15170 1470 15290 1590
rect 15335 1470 15455 1590
rect 15500 1470 15620 1590
rect 15665 1470 15785 1590
rect 15830 1470 15950 1590
rect 15995 1470 16115 1590
rect 16160 1470 16280 1590
rect 16325 1470 16445 1590
rect 16490 1470 16610 1590
rect 16655 1470 16775 1590
rect 16820 1470 16940 1590
rect 16985 1470 17105 1590
rect 17150 1470 17270 1590
rect 17315 1470 17435 1590
rect 17480 1470 17600 1590
rect 17645 1470 17765 1590
rect 17810 1470 17930 1590
rect 17975 1470 18095 1590
rect 18140 1470 18260 1590
rect 18550 1470 18670 1590
rect 18715 1470 18835 1590
rect 18880 1470 19000 1590
rect 19045 1470 19165 1590
rect 19210 1470 19330 1590
rect 19375 1470 19495 1590
rect 19540 1470 19660 1590
rect 19705 1470 19825 1590
rect 19870 1470 19990 1590
rect 20035 1470 20155 1590
rect 20200 1470 20320 1590
rect 20365 1470 20485 1590
rect 20530 1470 20650 1590
rect 20695 1470 20815 1590
rect 20860 1470 20980 1590
rect 21025 1470 21145 1590
rect 21190 1470 21310 1590
rect 21355 1470 21475 1590
rect 21520 1470 21640 1590
rect 21685 1470 21805 1590
rect 21850 1470 21970 1590
rect 22015 1470 22135 1590
rect 22180 1470 22300 1590
rect 22345 1470 22465 1590
rect 22510 1470 22630 1590
rect 22675 1470 22795 1590
rect 22840 1470 22960 1590
rect 23005 1470 23125 1590
rect 23170 1470 23290 1590
rect 23335 1470 23455 1590
rect 23500 1470 23620 1590
rect 23665 1470 23785 1590
rect 23830 1470 23950 1590
rect 24240 1470 24360 1590
rect 24405 1470 24525 1590
rect 24570 1470 24690 1590
rect 24735 1470 24855 1590
rect 24900 1470 25020 1590
rect 25065 1470 25185 1590
rect 25230 1470 25350 1590
rect 25395 1470 25515 1590
rect 25560 1470 25680 1590
rect 25725 1470 25845 1590
rect 25890 1470 26010 1590
rect 26055 1470 26175 1590
rect 26220 1470 26340 1590
rect 26385 1470 26505 1590
rect 26550 1470 26670 1590
rect 26715 1470 26835 1590
rect 26880 1470 27000 1590
rect 27045 1470 27165 1590
rect 27210 1470 27330 1590
rect 27375 1470 27495 1590
rect 27540 1470 27660 1590
rect 27705 1470 27825 1590
rect 27870 1470 27990 1590
rect 28035 1470 28155 1590
rect 28200 1470 28320 1590
rect 28365 1470 28485 1590
rect 28530 1470 28650 1590
rect 28695 1470 28815 1590
rect 28860 1470 28980 1590
rect 29025 1470 29145 1590
rect 29190 1470 29310 1590
rect 29355 1470 29475 1590
rect 29520 1470 29640 1590
rect 7170 -10000 7290 -9880
rect 7335 -10000 7455 -9880
rect 7500 -10000 7620 -9880
rect 7665 -10000 7785 -9880
rect 7830 -10000 7950 -9880
rect 7995 -10000 8115 -9880
rect 8160 -10000 8280 -9880
rect 8325 -10000 8445 -9880
rect 8490 -10000 8610 -9880
rect 8655 -10000 8775 -9880
rect 8820 -10000 8940 -9880
rect 8985 -10000 9105 -9880
rect 9150 -10000 9270 -9880
rect 9315 -10000 9435 -9880
rect 9480 -10000 9600 -9880
rect 9645 -10000 9765 -9880
rect 9810 -10000 9930 -9880
rect 9975 -10000 10095 -9880
rect 10140 -10000 10260 -9880
rect 10305 -10000 10425 -9880
rect 10470 -10000 10590 -9880
rect 10635 -10000 10755 -9880
rect 10800 -10000 10920 -9880
rect 10965 -10000 11085 -9880
rect 11130 -10000 11250 -9880
rect 11295 -10000 11415 -9880
rect 11460 -10000 11580 -9880
rect 11625 -10000 11745 -9880
rect 11790 -10000 11910 -9880
rect 11955 -10000 12075 -9880
rect 12120 -10000 12240 -9880
rect 12285 -10000 12405 -9880
rect 12450 -10000 12570 -9880
rect 12860 -10000 12980 -9880
rect 13025 -10000 13145 -9880
rect 13190 -10000 13310 -9880
rect 13355 -10000 13475 -9880
rect 13520 -10000 13640 -9880
rect 13685 -10000 13805 -9880
rect 13850 -10000 13970 -9880
rect 14015 -10000 14135 -9880
rect 14180 -10000 14300 -9880
rect 14345 -10000 14465 -9880
rect 14510 -10000 14630 -9880
rect 14675 -10000 14795 -9880
rect 14840 -10000 14960 -9880
rect 15005 -10000 15125 -9880
rect 15170 -10000 15290 -9880
rect 15335 -10000 15455 -9880
rect 15500 -10000 15620 -9880
rect 15665 -10000 15785 -9880
rect 15830 -10000 15950 -9880
rect 15995 -10000 16115 -9880
rect 16160 -10000 16280 -9880
rect 16325 -10000 16445 -9880
rect 16490 -10000 16610 -9880
rect 16655 -10000 16775 -9880
rect 16820 -10000 16940 -9880
rect 16985 -10000 17105 -9880
rect 17150 -10000 17270 -9880
rect 17315 -10000 17435 -9880
rect 17480 -10000 17600 -9880
rect 17645 -10000 17765 -9880
rect 17810 -10000 17930 -9880
rect 17975 -10000 18095 -9880
rect 18140 -10000 18260 -9880
rect 18550 -10000 18670 -9880
rect 18715 -10000 18835 -9880
rect 18880 -10000 19000 -9880
rect 19045 -10000 19165 -9880
rect 19210 -10000 19330 -9880
rect 19375 -10000 19495 -9880
rect 19540 -10000 19660 -9880
rect 19705 -10000 19825 -9880
rect 19870 -10000 19990 -9880
rect 20035 -10000 20155 -9880
rect 20200 -10000 20320 -9880
rect 20365 -10000 20485 -9880
rect 20530 -10000 20650 -9880
rect 20695 -10000 20815 -9880
rect 20860 -10000 20980 -9880
rect 21025 -10000 21145 -9880
rect 21190 -10000 21310 -9880
rect 21355 -10000 21475 -9880
rect 21520 -10000 21640 -9880
rect 21685 -10000 21805 -9880
rect 21850 -10000 21970 -9880
rect 22015 -10000 22135 -9880
rect 22180 -10000 22300 -9880
rect 22345 -10000 22465 -9880
rect 22510 -10000 22630 -9880
rect 22675 -10000 22795 -9880
rect 22840 -10000 22960 -9880
rect 23005 -10000 23125 -9880
rect 23170 -10000 23290 -9880
rect 23335 -10000 23455 -9880
rect 23500 -10000 23620 -9880
rect 23665 -10000 23785 -9880
rect 23830 -10000 23950 -9880
rect 24240 -10000 24360 -9880
rect 24405 -10000 24525 -9880
rect 24570 -10000 24690 -9880
rect 24735 -10000 24855 -9880
rect 24900 -10000 25020 -9880
rect 25065 -10000 25185 -9880
rect 25230 -10000 25350 -9880
rect 25395 -10000 25515 -9880
rect 25560 -10000 25680 -9880
rect 25725 -10000 25845 -9880
rect 25890 -10000 26010 -9880
rect 26055 -10000 26175 -9880
rect 26220 -10000 26340 -9880
rect 26385 -10000 26505 -9880
rect 26550 -10000 26670 -9880
rect 26715 -10000 26835 -9880
rect 26880 -10000 27000 -9880
rect 27045 -10000 27165 -9880
rect 27210 -10000 27330 -9880
rect 27375 -10000 27495 -9880
rect 27540 -10000 27660 -9880
rect 27705 -10000 27825 -9880
rect 27870 -10000 27990 -9880
rect 28035 -10000 28155 -9880
rect 28200 -10000 28320 -9880
rect 28365 -10000 28485 -9880
rect 28530 -10000 28650 -9880
rect 28695 -10000 28815 -9880
rect 28860 -10000 28980 -9880
rect 29025 -10000 29145 -9880
rect 29190 -10000 29310 -9880
rect 29355 -10000 29475 -9880
rect 29520 -10000 29640 -9880
<< mimcap2 >>
rect 7120 7160 12620 7170
rect 7120 7040 7130 7160
rect 7250 7040 7295 7160
rect 7415 7040 7460 7160
rect 7580 7040 7625 7160
rect 7745 7040 7800 7160
rect 7920 7040 7965 7160
rect 8085 7040 8130 7160
rect 8250 7040 8295 7160
rect 8415 7040 8470 7160
rect 8590 7040 8635 7160
rect 8755 7040 8800 7160
rect 8920 7040 8965 7160
rect 9085 7040 9140 7160
rect 9260 7040 9305 7160
rect 9425 7040 9470 7160
rect 9590 7040 9635 7160
rect 9755 7040 9810 7160
rect 9930 7040 9975 7160
rect 10095 7040 10140 7160
rect 10260 7040 10305 7160
rect 10425 7040 10480 7160
rect 10600 7040 10645 7160
rect 10765 7040 10810 7160
rect 10930 7040 10975 7160
rect 11095 7040 11150 7160
rect 11270 7040 11315 7160
rect 11435 7040 11480 7160
rect 11600 7040 11645 7160
rect 11765 7040 11820 7160
rect 11940 7040 11985 7160
rect 12105 7040 12150 7160
rect 12270 7040 12315 7160
rect 12435 7040 12490 7160
rect 12610 7040 12620 7160
rect 7120 6985 12620 7040
rect 7120 6865 7130 6985
rect 7250 6865 7295 6985
rect 7415 6865 7460 6985
rect 7580 6865 7625 6985
rect 7745 6865 7800 6985
rect 7920 6865 7965 6985
rect 8085 6865 8130 6985
rect 8250 6865 8295 6985
rect 8415 6865 8470 6985
rect 8590 6865 8635 6985
rect 8755 6865 8800 6985
rect 8920 6865 8965 6985
rect 9085 6865 9140 6985
rect 9260 6865 9305 6985
rect 9425 6865 9470 6985
rect 9590 6865 9635 6985
rect 9755 6865 9810 6985
rect 9930 6865 9975 6985
rect 10095 6865 10140 6985
rect 10260 6865 10305 6985
rect 10425 6865 10480 6985
rect 10600 6865 10645 6985
rect 10765 6865 10810 6985
rect 10930 6865 10975 6985
rect 11095 6865 11150 6985
rect 11270 6865 11315 6985
rect 11435 6865 11480 6985
rect 11600 6865 11645 6985
rect 11765 6865 11820 6985
rect 11940 6865 11985 6985
rect 12105 6865 12150 6985
rect 12270 6865 12315 6985
rect 12435 6865 12490 6985
rect 12610 6865 12620 6985
rect 7120 6820 12620 6865
rect 7120 6700 7130 6820
rect 7250 6700 7295 6820
rect 7415 6700 7460 6820
rect 7580 6700 7625 6820
rect 7745 6700 7800 6820
rect 7920 6700 7965 6820
rect 8085 6700 8130 6820
rect 8250 6700 8295 6820
rect 8415 6700 8470 6820
rect 8590 6700 8635 6820
rect 8755 6700 8800 6820
rect 8920 6700 8965 6820
rect 9085 6700 9140 6820
rect 9260 6700 9305 6820
rect 9425 6700 9470 6820
rect 9590 6700 9635 6820
rect 9755 6700 9810 6820
rect 9930 6700 9975 6820
rect 10095 6700 10140 6820
rect 10260 6700 10305 6820
rect 10425 6700 10480 6820
rect 10600 6700 10645 6820
rect 10765 6700 10810 6820
rect 10930 6700 10975 6820
rect 11095 6700 11150 6820
rect 11270 6700 11315 6820
rect 11435 6700 11480 6820
rect 11600 6700 11645 6820
rect 11765 6700 11820 6820
rect 11940 6700 11985 6820
rect 12105 6700 12150 6820
rect 12270 6700 12315 6820
rect 12435 6700 12490 6820
rect 12610 6700 12620 6820
rect 7120 6655 12620 6700
rect 7120 6535 7130 6655
rect 7250 6535 7295 6655
rect 7415 6535 7460 6655
rect 7580 6535 7625 6655
rect 7745 6535 7800 6655
rect 7920 6535 7965 6655
rect 8085 6535 8130 6655
rect 8250 6535 8295 6655
rect 8415 6535 8470 6655
rect 8590 6535 8635 6655
rect 8755 6535 8800 6655
rect 8920 6535 8965 6655
rect 9085 6535 9140 6655
rect 9260 6535 9305 6655
rect 9425 6535 9470 6655
rect 9590 6535 9635 6655
rect 9755 6535 9810 6655
rect 9930 6535 9975 6655
rect 10095 6535 10140 6655
rect 10260 6535 10305 6655
rect 10425 6535 10480 6655
rect 10600 6535 10645 6655
rect 10765 6535 10810 6655
rect 10930 6535 10975 6655
rect 11095 6535 11150 6655
rect 11270 6535 11315 6655
rect 11435 6535 11480 6655
rect 11600 6535 11645 6655
rect 11765 6535 11820 6655
rect 11940 6535 11985 6655
rect 12105 6535 12150 6655
rect 12270 6535 12315 6655
rect 12435 6535 12490 6655
rect 12610 6535 12620 6655
rect 7120 6490 12620 6535
rect 7120 6370 7130 6490
rect 7250 6370 7295 6490
rect 7415 6370 7460 6490
rect 7580 6370 7625 6490
rect 7745 6370 7800 6490
rect 7920 6370 7965 6490
rect 8085 6370 8130 6490
rect 8250 6370 8295 6490
rect 8415 6370 8470 6490
rect 8590 6370 8635 6490
rect 8755 6370 8800 6490
rect 8920 6370 8965 6490
rect 9085 6370 9140 6490
rect 9260 6370 9305 6490
rect 9425 6370 9470 6490
rect 9590 6370 9635 6490
rect 9755 6370 9810 6490
rect 9930 6370 9975 6490
rect 10095 6370 10140 6490
rect 10260 6370 10305 6490
rect 10425 6370 10480 6490
rect 10600 6370 10645 6490
rect 10765 6370 10810 6490
rect 10930 6370 10975 6490
rect 11095 6370 11150 6490
rect 11270 6370 11315 6490
rect 11435 6370 11480 6490
rect 11600 6370 11645 6490
rect 11765 6370 11820 6490
rect 11940 6370 11985 6490
rect 12105 6370 12150 6490
rect 12270 6370 12315 6490
rect 12435 6370 12490 6490
rect 12610 6370 12620 6490
rect 7120 6315 12620 6370
rect 7120 6195 7130 6315
rect 7250 6195 7295 6315
rect 7415 6195 7460 6315
rect 7580 6195 7625 6315
rect 7745 6195 7800 6315
rect 7920 6195 7965 6315
rect 8085 6195 8130 6315
rect 8250 6195 8295 6315
rect 8415 6195 8470 6315
rect 8590 6195 8635 6315
rect 8755 6195 8800 6315
rect 8920 6195 8965 6315
rect 9085 6195 9140 6315
rect 9260 6195 9305 6315
rect 9425 6195 9470 6315
rect 9590 6195 9635 6315
rect 9755 6195 9810 6315
rect 9930 6195 9975 6315
rect 10095 6195 10140 6315
rect 10260 6195 10305 6315
rect 10425 6195 10480 6315
rect 10600 6195 10645 6315
rect 10765 6195 10810 6315
rect 10930 6195 10975 6315
rect 11095 6195 11150 6315
rect 11270 6195 11315 6315
rect 11435 6195 11480 6315
rect 11600 6195 11645 6315
rect 11765 6195 11820 6315
rect 11940 6195 11985 6315
rect 12105 6195 12150 6315
rect 12270 6195 12315 6315
rect 12435 6195 12490 6315
rect 12610 6195 12620 6315
rect 7120 6150 12620 6195
rect 7120 6030 7130 6150
rect 7250 6030 7295 6150
rect 7415 6030 7460 6150
rect 7580 6030 7625 6150
rect 7745 6030 7800 6150
rect 7920 6030 7965 6150
rect 8085 6030 8130 6150
rect 8250 6030 8295 6150
rect 8415 6030 8470 6150
rect 8590 6030 8635 6150
rect 8755 6030 8800 6150
rect 8920 6030 8965 6150
rect 9085 6030 9140 6150
rect 9260 6030 9305 6150
rect 9425 6030 9470 6150
rect 9590 6030 9635 6150
rect 9755 6030 9810 6150
rect 9930 6030 9975 6150
rect 10095 6030 10140 6150
rect 10260 6030 10305 6150
rect 10425 6030 10480 6150
rect 10600 6030 10645 6150
rect 10765 6030 10810 6150
rect 10930 6030 10975 6150
rect 11095 6030 11150 6150
rect 11270 6030 11315 6150
rect 11435 6030 11480 6150
rect 11600 6030 11645 6150
rect 11765 6030 11820 6150
rect 11940 6030 11985 6150
rect 12105 6030 12150 6150
rect 12270 6030 12315 6150
rect 12435 6030 12490 6150
rect 12610 6030 12620 6150
rect 7120 5985 12620 6030
rect 7120 5865 7130 5985
rect 7250 5865 7295 5985
rect 7415 5865 7460 5985
rect 7580 5865 7625 5985
rect 7745 5865 7800 5985
rect 7920 5865 7965 5985
rect 8085 5865 8130 5985
rect 8250 5865 8295 5985
rect 8415 5865 8470 5985
rect 8590 5865 8635 5985
rect 8755 5865 8800 5985
rect 8920 5865 8965 5985
rect 9085 5865 9140 5985
rect 9260 5865 9305 5985
rect 9425 5865 9470 5985
rect 9590 5865 9635 5985
rect 9755 5865 9810 5985
rect 9930 5865 9975 5985
rect 10095 5865 10140 5985
rect 10260 5865 10305 5985
rect 10425 5865 10480 5985
rect 10600 5865 10645 5985
rect 10765 5865 10810 5985
rect 10930 5865 10975 5985
rect 11095 5865 11150 5985
rect 11270 5865 11315 5985
rect 11435 5865 11480 5985
rect 11600 5865 11645 5985
rect 11765 5865 11820 5985
rect 11940 5865 11985 5985
rect 12105 5865 12150 5985
rect 12270 5865 12315 5985
rect 12435 5865 12490 5985
rect 12610 5865 12620 5985
rect 7120 5820 12620 5865
rect 7120 5700 7130 5820
rect 7250 5700 7295 5820
rect 7415 5700 7460 5820
rect 7580 5700 7625 5820
rect 7745 5700 7800 5820
rect 7920 5700 7965 5820
rect 8085 5700 8130 5820
rect 8250 5700 8295 5820
rect 8415 5700 8470 5820
rect 8590 5700 8635 5820
rect 8755 5700 8800 5820
rect 8920 5700 8965 5820
rect 9085 5700 9140 5820
rect 9260 5700 9305 5820
rect 9425 5700 9470 5820
rect 9590 5700 9635 5820
rect 9755 5700 9810 5820
rect 9930 5700 9975 5820
rect 10095 5700 10140 5820
rect 10260 5700 10305 5820
rect 10425 5700 10480 5820
rect 10600 5700 10645 5820
rect 10765 5700 10810 5820
rect 10930 5700 10975 5820
rect 11095 5700 11150 5820
rect 11270 5700 11315 5820
rect 11435 5700 11480 5820
rect 11600 5700 11645 5820
rect 11765 5700 11820 5820
rect 11940 5700 11985 5820
rect 12105 5700 12150 5820
rect 12270 5700 12315 5820
rect 12435 5700 12490 5820
rect 12610 5700 12620 5820
rect 7120 5645 12620 5700
rect 7120 5525 7130 5645
rect 7250 5525 7295 5645
rect 7415 5525 7460 5645
rect 7580 5525 7625 5645
rect 7745 5525 7800 5645
rect 7920 5525 7965 5645
rect 8085 5525 8130 5645
rect 8250 5525 8295 5645
rect 8415 5525 8470 5645
rect 8590 5525 8635 5645
rect 8755 5525 8800 5645
rect 8920 5525 8965 5645
rect 9085 5525 9140 5645
rect 9260 5525 9305 5645
rect 9425 5525 9470 5645
rect 9590 5525 9635 5645
rect 9755 5525 9810 5645
rect 9930 5525 9975 5645
rect 10095 5525 10140 5645
rect 10260 5525 10305 5645
rect 10425 5525 10480 5645
rect 10600 5525 10645 5645
rect 10765 5525 10810 5645
rect 10930 5525 10975 5645
rect 11095 5525 11150 5645
rect 11270 5525 11315 5645
rect 11435 5525 11480 5645
rect 11600 5525 11645 5645
rect 11765 5525 11820 5645
rect 11940 5525 11985 5645
rect 12105 5525 12150 5645
rect 12270 5525 12315 5645
rect 12435 5525 12490 5645
rect 12610 5525 12620 5645
rect 7120 5480 12620 5525
rect 7120 5360 7130 5480
rect 7250 5360 7295 5480
rect 7415 5360 7460 5480
rect 7580 5360 7625 5480
rect 7745 5360 7800 5480
rect 7920 5360 7965 5480
rect 8085 5360 8130 5480
rect 8250 5360 8295 5480
rect 8415 5360 8470 5480
rect 8590 5360 8635 5480
rect 8755 5360 8800 5480
rect 8920 5360 8965 5480
rect 9085 5360 9140 5480
rect 9260 5360 9305 5480
rect 9425 5360 9470 5480
rect 9590 5360 9635 5480
rect 9755 5360 9810 5480
rect 9930 5360 9975 5480
rect 10095 5360 10140 5480
rect 10260 5360 10305 5480
rect 10425 5360 10480 5480
rect 10600 5360 10645 5480
rect 10765 5360 10810 5480
rect 10930 5360 10975 5480
rect 11095 5360 11150 5480
rect 11270 5360 11315 5480
rect 11435 5360 11480 5480
rect 11600 5360 11645 5480
rect 11765 5360 11820 5480
rect 11940 5360 11985 5480
rect 12105 5360 12150 5480
rect 12270 5360 12315 5480
rect 12435 5360 12490 5480
rect 12610 5360 12620 5480
rect 7120 5315 12620 5360
rect 7120 5195 7130 5315
rect 7250 5195 7295 5315
rect 7415 5195 7460 5315
rect 7580 5195 7625 5315
rect 7745 5195 7800 5315
rect 7920 5195 7965 5315
rect 8085 5195 8130 5315
rect 8250 5195 8295 5315
rect 8415 5195 8470 5315
rect 8590 5195 8635 5315
rect 8755 5195 8800 5315
rect 8920 5195 8965 5315
rect 9085 5195 9140 5315
rect 9260 5195 9305 5315
rect 9425 5195 9470 5315
rect 9590 5195 9635 5315
rect 9755 5195 9810 5315
rect 9930 5195 9975 5315
rect 10095 5195 10140 5315
rect 10260 5195 10305 5315
rect 10425 5195 10480 5315
rect 10600 5195 10645 5315
rect 10765 5195 10810 5315
rect 10930 5195 10975 5315
rect 11095 5195 11150 5315
rect 11270 5195 11315 5315
rect 11435 5195 11480 5315
rect 11600 5195 11645 5315
rect 11765 5195 11820 5315
rect 11940 5195 11985 5315
rect 12105 5195 12150 5315
rect 12270 5195 12315 5315
rect 12435 5195 12490 5315
rect 12610 5195 12620 5315
rect 7120 5150 12620 5195
rect 7120 5030 7130 5150
rect 7250 5030 7295 5150
rect 7415 5030 7460 5150
rect 7580 5030 7625 5150
rect 7745 5030 7800 5150
rect 7920 5030 7965 5150
rect 8085 5030 8130 5150
rect 8250 5030 8295 5150
rect 8415 5030 8470 5150
rect 8590 5030 8635 5150
rect 8755 5030 8800 5150
rect 8920 5030 8965 5150
rect 9085 5030 9140 5150
rect 9260 5030 9305 5150
rect 9425 5030 9470 5150
rect 9590 5030 9635 5150
rect 9755 5030 9810 5150
rect 9930 5030 9975 5150
rect 10095 5030 10140 5150
rect 10260 5030 10305 5150
rect 10425 5030 10480 5150
rect 10600 5030 10645 5150
rect 10765 5030 10810 5150
rect 10930 5030 10975 5150
rect 11095 5030 11150 5150
rect 11270 5030 11315 5150
rect 11435 5030 11480 5150
rect 11600 5030 11645 5150
rect 11765 5030 11820 5150
rect 11940 5030 11985 5150
rect 12105 5030 12150 5150
rect 12270 5030 12315 5150
rect 12435 5030 12490 5150
rect 12610 5030 12620 5150
rect 7120 4975 12620 5030
rect 7120 4855 7130 4975
rect 7250 4855 7295 4975
rect 7415 4855 7460 4975
rect 7580 4855 7625 4975
rect 7745 4855 7800 4975
rect 7920 4855 7965 4975
rect 8085 4855 8130 4975
rect 8250 4855 8295 4975
rect 8415 4855 8470 4975
rect 8590 4855 8635 4975
rect 8755 4855 8800 4975
rect 8920 4855 8965 4975
rect 9085 4855 9140 4975
rect 9260 4855 9305 4975
rect 9425 4855 9470 4975
rect 9590 4855 9635 4975
rect 9755 4855 9810 4975
rect 9930 4855 9975 4975
rect 10095 4855 10140 4975
rect 10260 4855 10305 4975
rect 10425 4855 10480 4975
rect 10600 4855 10645 4975
rect 10765 4855 10810 4975
rect 10930 4855 10975 4975
rect 11095 4855 11150 4975
rect 11270 4855 11315 4975
rect 11435 4855 11480 4975
rect 11600 4855 11645 4975
rect 11765 4855 11820 4975
rect 11940 4855 11985 4975
rect 12105 4855 12150 4975
rect 12270 4855 12315 4975
rect 12435 4855 12490 4975
rect 12610 4855 12620 4975
rect 7120 4810 12620 4855
rect 7120 4690 7130 4810
rect 7250 4690 7295 4810
rect 7415 4690 7460 4810
rect 7580 4690 7625 4810
rect 7745 4690 7800 4810
rect 7920 4690 7965 4810
rect 8085 4690 8130 4810
rect 8250 4690 8295 4810
rect 8415 4690 8470 4810
rect 8590 4690 8635 4810
rect 8755 4690 8800 4810
rect 8920 4690 8965 4810
rect 9085 4690 9140 4810
rect 9260 4690 9305 4810
rect 9425 4690 9470 4810
rect 9590 4690 9635 4810
rect 9755 4690 9810 4810
rect 9930 4690 9975 4810
rect 10095 4690 10140 4810
rect 10260 4690 10305 4810
rect 10425 4690 10480 4810
rect 10600 4690 10645 4810
rect 10765 4690 10810 4810
rect 10930 4690 10975 4810
rect 11095 4690 11150 4810
rect 11270 4690 11315 4810
rect 11435 4690 11480 4810
rect 11600 4690 11645 4810
rect 11765 4690 11820 4810
rect 11940 4690 11985 4810
rect 12105 4690 12150 4810
rect 12270 4690 12315 4810
rect 12435 4690 12490 4810
rect 12610 4690 12620 4810
rect 7120 4645 12620 4690
rect 7120 4525 7130 4645
rect 7250 4525 7295 4645
rect 7415 4525 7460 4645
rect 7580 4525 7625 4645
rect 7745 4525 7800 4645
rect 7920 4525 7965 4645
rect 8085 4525 8130 4645
rect 8250 4525 8295 4645
rect 8415 4525 8470 4645
rect 8590 4525 8635 4645
rect 8755 4525 8800 4645
rect 8920 4525 8965 4645
rect 9085 4525 9140 4645
rect 9260 4525 9305 4645
rect 9425 4525 9470 4645
rect 9590 4525 9635 4645
rect 9755 4525 9810 4645
rect 9930 4525 9975 4645
rect 10095 4525 10140 4645
rect 10260 4525 10305 4645
rect 10425 4525 10480 4645
rect 10600 4525 10645 4645
rect 10765 4525 10810 4645
rect 10930 4525 10975 4645
rect 11095 4525 11150 4645
rect 11270 4525 11315 4645
rect 11435 4525 11480 4645
rect 11600 4525 11645 4645
rect 11765 4525 11820 4645
rect 11940 4525 11985 4645
rect 12105 4525 12150 4645
rect 12270 4525 12315 4645
rect 12435 4525 12490 4645
rect 12610 4525 12620 4645
rect 7120 4480 12620 4525
rect 7120 4360 7130 4480
rect 7250 4360 7295 4480
rect 7415 4360 7460 4480
rect 7580 4360 7625 4480
rect 7745 4360 7800 4480
rect 7920 4360 7965 4480
rect 8085 4360 8130 4480
rect 8250 4360 8295 4480
rect 8415 4360 8470 4480
rect 8590 4360 8635 4480
rect 8755 4360 8800 4480
rect 8920 4360 8965 4480
rect 9085 4360 9140 4480
rect 9260 4360 9305 4480
rect 9425 4360 9470 4480
rect 9590 4360 9635 4480
rect 9755 4360 9810 4480
rect 9930 4360 9975 4480
rect 10095 4360 10140 4480
rect 10260 4360 10305 4480
rect 10425 4360 10480 4480
rect 10600 4360 10645 4480
rect 10765 4360 10810 4480
rect 10930 4360 10975 4480
rect 11095 4360 11150 4480
rect 11270 4360 11315 4480
rect 11435 4360 11480 4480
rect 11600 4360 11645 4480
rect 11765 4360 11820 4480
rect 11940 4360 11985 4480
rect 12105 4360 12150 4480
rect 12270 4360 12315 4480
rect 12435 4360 12490 4480
rect 12610 4360 12620 4480
rect 7120 4305 12620 4360
rect 7120 4185 7130 4305
rect 7250 4185 7295 4305
rect 7415 4185 7460 4305
rect 7580 4185 7625 4305
rect 7745 4185 7800 4305
rect 7920 4185 7965 4305
rect 8085 4185 8130 4305
rect 8250 4185 8295 4305
rect 8415 4185 8470 4305
rect 8590 4185 8635 4305
rect 8755 4185 8800 4305
rect 8920 4185 8965 4305
rect 9085 4185 9140 4305
rect 9260 4185 9305 4305
rect 9425 4185 9470 4305
rect 9590 4185 9635 4305
rect 9755 4185 9810 4305
rect 9930 4185 9975 4305
rect 10095 4185 10140 4305
rect 10260 4185 10305 4305
rect 10425 4185 10480 4305
rect 10600 4185 10645 4305
rect 10765 4185 10810 4305
rect 10930 4185 10975 4305
rect 11095 4185 11150 4305
rect 11270 4185 11315 4305
rect 11435 4185 11480 4305
rect 11600 4185 11645 4305
rect 11765 4185 11820 4305
rect 11940 4185 11985 4305
rect 12105 4185 12150 4305
rect 12270 4185 12315 4305
rect 12435 4185 12490 4305
rect 12610 4185 12620 4305
rect 7120 4140 12620 4185
rect 7120 4020 7130 4140
rect 7250 4020 7295 4140
rect 7415 4020 7460 4140
rect 7580 4020 7625 4140
rect 7745 4020 7800 4140
rect 7920 4020 7965 4140
rect 8085 4020 8130 4140
rect 8250 4020 8295 4140
rect 8415 4020 8470 4140
rect 8590 4020 8635 4140
rect 8755 4020 8800 4140
rect 8920 4020 8965 4140
rect 9085 4020 9140 4140
rect 9260 4020 9305 4140
rect 9425 4020 9470 4140
rect 9590 4020 9635 4140
rect 9755 4020 9810 4140
rect 9930 4020 9975 4140
rect 10095 4020 10140 4140
rect 10260 4020 10305 4140
rect 10425 4020 10480 4140
rect 10600 4020 10645 4140
rect 10765 4020 10810 4140
rect 10930 4020 10975 4140
rect 11095 4020 11150 4140
rect 11270 4020 11315 4140
rect 11435 4020 11480 4140
rect 11600 4020 11645 4140
rect 11765 4020 11820 4140
rect 11940 4020 11985 4140
rect 12105 4020 12150 4140
rect 12270 4020 12315 4140
rect 12435 4020 12490 4140
rect 12610 4020 12620 4140
rect 7120 3975 12620 4020
rect 7120 3855 7130 3975
rect 7250 3855 7295 3975
rect 7415 3855 7460 3975
rect 7580 3855 7625 3975
rect 7745 3855 7800 3975
rect 7920 3855 7965 3975
rect 8085 3855 8130 3975
rect 8250 3855 8295 3975
rect 8415 3855 8470 3975
rect 8590 3855 8635 3975
rect 8755 3855 8800 3975
rect 8920 3855 8965 3975
rect 9085 3855 9140 3975
rect 9260 3855 9305 3975
rect 9425 3855 9470 3975
rect 9590 3855 9635 3975
rect 9755 3855 9810 3975
rect 9930 3855 9975 3975
rect 10095 3855 10140 3975
rect 10260 3855 10305 3975
rect 10425 3855 10480 3975
rect 10600 3855 10645 3975
rect 10765 3855 10810 3975
rect 10930 3855 10975 3975
rect 11095 3855 11150 3975
rect 11270 3855 11315 3975
rect 11435 3855 11480 3975
rect 11600 3855 11645 3975
rect 11765 3855 11820 3975
rect 11940 3855 11985 3975
rect 12105 3855 12150 3975
rect 12270 3855 12315 3975
rect 12435 3855 12490 3975
rect 12610 3855 12620 3975
rect 7120 3810 12620 3855
rect 7120 3690 7130 3810
rect 7250 3690 7295 3810
rect 7415 3690 7460 3810
rect 7580 3690 7625 3810
rect 7745 3690 7800 3810
rect 7920 3690 7965 3810
rect 8085 3690 8130 3810
rect 8250 3690 8295 3810
rect 8415 3690 8470 3810
rect 8590 3690 8635 3810
rect 8755 3690 8800 3810
rect 8920 3690 8965 3810
rect 9085 3690 9140 3810
rect 9260 3690 9305 3810
rect 9425 3690 9470 3810
rect 9590 3690 9635 3810
rect 9755 3690 9810 3810
rect 9930 3690 9975 3810
rect 10095 3690 10140 3810
rect 10260 3690 10305 3810
rect 10425 3690 10480 3810
rect 10600 3690 10645 3810
rect 10765 3690 10810 3810
rect 10930 3690 10975 3810
rect 11095 3690 11150 3810
rect 11270 3690 11315 3810
rect 11435 3690 11480 3810
rect 11600 3690 11645 3810
rect 11765 3690 11820 3810
rect 11940 3690 11985 3810
rect 12105 3690 12150 3810
rect 12270 3690 12315 3810
rect 12435 3690 12490 3810
rect 12610 3690 12620 3810
rect 7120 3635 12620 3690
rect 7120 3515 7130 3635
rect 7250 3515 7295 3635
rect 7415 3515 7460 3635
rect 7580 3515 7625 3635
rect 7745 3515 7800 3635
rect 7920 3515 7965 3635
rect 8085 3515 8130 3635
rect 8250 3515 8295 3635
rect 8415 3515 8470 3635
rect 8590 3515 8635 3635
rect 8755 3515 8800 3635
rect 8920 3515 8965 3635
rect 9085 3515 9140 3635
rect 9260 3515 9305 3635
rect 9425 3515 9470 3635
rect 9590 3515 9635 3635
rect 9755 3515 9810 3635
rect 9930 3515 9975 3635
rect 10095 3515 10140 3635
rect 10260 3515 10305 3635
rect 10425 3515 10480 3635
rect 10600 3515 10645 3635
rect 10765 3515 10810 3635
rect 10930 3515 10975 3635
rect 11095 3515 11150 3635
rect 11270 3515 11315 3635
rect 11435 3515 11480 3635
rect 11600 3515 11645 3635
rect 11765 3515 11820 3635
rect 11940 3515 11985 3635
rect 12105 3515 12150 3635
rect 12270 3515 12315 3635
rect 12435 3515 12490 3635
rect 12610 3515 12620 3635
rect 7120 3470 12620 3515
rect 7120 3350 7130 3470
rect 7250 3350 7295 3470
rect 7415 3350 7460 3470
rect 7580 3350 7625 3470
rect 7745 3350 7800 3470
rect 7920 3350 7965 3470
rect 8085 3350 8130 3470
rect 8250 3350 8295 3470
rect 8415 3350 8470 3470
rect 8590 3350 8635 3470
rect 8755 3350 8800 3470
rect 8920 3350 8965 3470
rect 9085 3350 9140 3470
rect 9260 3350 9305 3470
rect 9425 3350 9470 3470
rect 9590 3350 9635 3470
rect 9755 3350 9810 3470
rect 9930 3350 9975 3470
rect 10095 3350 10140 3470
rect 10260 3350 10305 3470
rect 10425 3350 10480 3470
rect 10600 3350 10645 3470
rect 10765 3350 10810 3470
rect 10930 3350 10975 3470
rect 11095 3350 11150 3470
rect 11270 3350 11315 3470
rect 11435 3350 11480 3470
rect 11600 3350 11645 3470
rect 11765 3350 11820 3470
rect 11940 3350 11985 3470
rect 12105 3350 12150 3470
rect 12270 3350 12315 3470
rect 12435 3350 12490 3470
rect 12610 3350 12620 3470
rect 7120 3305 12620 3350
rect 7120 3185 7130 3305
rect 7250 3185 7295 3305
rect 7415 3185 7460 3305
rect 7580 3185 7625 3305
rect 7745 3185 7800 3305
rect 7920 3185 7965 3305
rect 8085 3185 8130 3305
rect 8250 3185 8295 3305
rect 8415 3185 8470 3305
rect 8590 3185 8635 3305
rect 8755 3185 8800 3305
rect 8920 3185 8965 3305
rect 9085 3185 9140 3305
rect 9260 3185 9305 3305
rect 9425 3185 9470 3305
rect 9590 3185 9635 3305
rect 9755 3185 9810 3305
rect 9930 3185 9975 3305
rect 10095 3185 10140 3305
rect 10260 3185 10305 3305
rect 10425 3185 10480 3305
rect 10600 3185 10645 3305
rect 10765 3185 10810 3305
rect 10930 3185 10975 3305
rect 11095 3185 11150 3305
rect 11270 3185 11315 3305
rect 11435 3185 11480 3305
rect 11600 3185 11645 3305
rect 11765 3185 11820 3305
rect 11940 3185 11985 3305
rect 12105 3185 12150 3305
rect 12270 3185 12315 3305
rect 12435 3185 12490 3305
rect 12610 3185 12620 3305
rect 7120 3140 12620 3185
rect 7120 3020 7130 3140
rect 7250 3020 7295 3140
rect 7415 3020 7460 3140
rect 7580 3020 7625 3140
rect 7745 3020 7800 3140
rect 7920 3020 7965 3140
rect 8085 3020 8130 3140
rect 8250 3020 8295 3140
rect 8415 3020 8470 3140
rect 8590 3020 8635 3140
rect 8755 3020 8800 3140
rect 8920 3020 8965 3140
rect 9085 3020 9140 3140
rect 9260 3020 9305 3140
rect 9425 3020 9470 3140
rect 9590 3020 9635 3140
rect 9755 3020 9810 3140
rect 9930 3020 9975 3140
rect 10095 3020 10140 3140
rect 10260 3020 10305 3140
rect 10425 3020 10480 3140
rect 10600 3020 10645 3140
rect 10765 3020 10810 3140
rect 10930 3020 10975 3140
rect 11095 3020 11150 3140
rect 11270 3020 11315 3140
rect 11435 3020 11480 3140
rect 11600 3020 11645 3140
rect 11765 3020 11820 3140
rect 11940 3020 11985 3140
rect 12105 3020 12150 3140
rect 12270 3020 12315 3140
rect 12435 3020 12490 3140
rect 12610 3020 12620 3140
rect 7120 2965 12620 3020
rect 7120 2845 7130 2965
rect 7250 2845 7295 2965
rect 7415 2845 7460 2965
rect 7580 2845 7625 2965
rect 7745 2845 7800 2965
rect 7920 2845 7965 2965
rect 8085 2845 8130 2965
rect 8250 2845 8295 2965
rect 8415 2845 8470 2965
rect 8590 2845 8635 2965
rect 8755 2845 8800 2965
rect 8920 2845 8965 2965
rect 9085 2845 9140 2965
rect 9260 2845 9305 2965
rect 9425 2845 9470 2965
rect 9590 2845 9635 2965
rect 9755 2845 9810 2965
rect 9930 2845 9975 2965
rect 10095 2845 10140 2965
rect 10260 2845 10305 2965
rect 10425 2845 10480 2965
rect 10600 2845 10645 2965
rect 10765 2845 10810 2965
rect 10930 2845 10975 2965
rect 11095 2845 11150 2965
rect 11270 2845 11315 2965
rect 11435 2845 11480 2965
rect 11600 2845 11645 2965
rect 11765 2845 11820 2965
rect 11940 2845 11985 2965
rect 12105 2845 12150 2965
rect 12270 2845 12315 2965
rect 12435 2845 12490 2965
rect 12610 2845 12620 2965
rect 7120 2800 12620 2845
rect 7120 2680 7130 2800
rect 7250 2680 7295 2800
rect 7415 2680 7460 2800
rect 7580 2680 7625 2800
rect 7745 2680 7800 2800
rect 7920 2680 7965 2800
rect 8085 2680 8130 2800
rect 8250 2680 8295 2800
rect 8415 2680 8470 2800
rect 8590 2680 8635 2800
rect 8755 2680 8800 2800
rect 8920 2680 8965 2800
rect 9085 2680 9140 2800
rect 9260 2680 9305 2800
rect 9425 2680 9470 2800
rect 9590 2680 9635 2800
rect 9755 2680 9810 2800
rect 9930 2680 9975 2800
rect 10095 2680 10140 2800
rect 10260 2680 10305 2800
rect 10425 2680 10480 2800
rect 10600 2680 10645 2800
rect 10765 2680 10810 2800
rect 10930 2680 10975 2800
rect 11095 2680 11150 2800
rect 11270 2680 11315 2800
rect 11435 2680 11480 2800
rect 11600 2680 11645 2800
rect 11765 2680 11820 2800
rect 11940 2680 11985 2800
rect 12105 2680 12150 2800
rect 12270 2680 12315 2800
rect 12435 2680 12490 2800
rect 12610 2680 12620 2800
rect 7120 2635 12620 2680
rect 7120 2515 7130 2635
rect 7250 2515 7295 2635
rect 7415 2515 7460 2635
rect 7580 2515 7625 2635
rect 7745 2515 7800 2635
rect 7920 2515 7965 2635
rect 8085 2515 8130 2635
rect 8250 2515 8295 2635
rect 8415 2515 8470 2635
rect 8590 2515 8635 2635
rect 8755 2515 8800 2635
rect 8920 2515 8965 2635
rect 9085 2515 9140 2635
rect 9260 2515 9305 2635
rect 9425 2515 9470 2635
rect 9590 2515 9635 2635
rect 9755 2515 9810 2635
rect 9930 2515 9975 2635
rect 10095 2515 10140 2635
rect 10260 2515 10305 2635
rect 10425 2515 10480 2635
rect 10600 2515 10645 2635
rect 10765 2515 10810 2635
rect 10930 2515 10975 2635
rect 11095 2515 11150 2635
rect 11270 2515 11315 2635
rect 11435 2515 11480 2635
rect 11600 2515 11645 2635
rect 11765 2515 11820 2635
rect 11940 2515 11985 2635
rect 12105 2515 12150 2635
rect 12270 2515 12315 2635
rect 12435 2515 12490 2635
rect 12610 2515 12620 2635
rect 7120 2470 12620 2515
rect 7120 2350 7130 2470
rect 7250 2350 7295 2470
rect 7415 2350 7460 2470
rect 7580 2350 7625 2470
rect 7745 2350 7800 2470
rect 7920 2350 7965 2470
rect 8085 2350 8130 2470
rect 8250 2350 8295 2470
rect 8415 2350 8470 2470
rect 8590 2350 8635 2470
rect 8755 2350 8800 2470
rect 8920 2350 8965 2470
rect 9085 2350 9140 2470
rect 9260 2350 9305 2470
rect 9425 2350 9470 2470
rect 9590 2350 9635 2470
rect 9755 2350 9810 2470
rect 9930 2350 9975 2470
rect 10095 2350 10140 2470
rect 10260 2350 10305 2470
rect 10425 2350 10480 2470
rect 10600 2350 10645 2470
rect 10765 2350 10810 2470
rect 10930 2350 10975 2470
rect 11095 2350 11150 2470
rect 11270 2350 11315 2470
rect 11435 2350 11480 2470
rect 11600 2350 11645 2470
rect 11765 2350 11820 2470
rect 11940 2350 11985 2470
rect 12105 2350 12150 2470
rect 12270 2350 12315 2470
rect 12435 2350 12490 2470
rect 12610 2350 12620 2470
rect 7120 2295 12620 2350
rect 7120 2175 7130 2295
rect 7250 2175 7295 2295
rect 7415 2175 7460 2295
rect 7580 2175 7625 2295
rect 7745 2175 7800 2295
rect 7920 2175 7965 2295
rect 8085 2175 8130 2295
rect 8250 2175 8295 2295
rect 8415 2175 8470 2295
rect 8590 2175 8635 2295
rect 8755 2175 8800 2295
rect 8920 2175 8965 2295
rect 9085 2175 9140 2295
rect 9260 2175 9305 2295
rect 9425 2175 9470 2295
rect 9590 2175 9635 2295
rect 9755 2175 9810 2295
rect 9930 2175 9975 2295
rect 10095 2175 10140 2295
rect 10260 2175 10305 2295
rect 10425 2175 10480 2295
rect 10600 2175 10645 2295
rect 10765 2175 10810 2295
rect 10930 2175 10975 2295
rect 11095 2175 11150 2295
rect 11270 2175 11315 2295
rect 11435 2175 11480 2295
rect 11600 2175 11645 2295
rect 11765 2175 11820 2295
rect 11940 2175 11985 2295
rect 12105 2175 12150 2295
rect 12270 2175 12315 2295
rect 12435 2175 12490 2295
rect 12610 2175 12620 2295
rect 7120 2130 12620 2175
rect 7120 2010 7130 2130
rect 7250 2010 7295 2130
rect 7415 2010 7460 2130
rect 7580 2010 7625 2130
rect 7745 2010 7800 2130
rect 7920 2010 7965 2130
rect 8085 2010 8130 2130
rect 8250 2010 8295 2130
rect 8415 2010 8470 2130
rect 8590 2010 8635 2130
rect 8755 2010 8800 2130
rect 8920 2010 8965 2130
rect 9085 2010 9140 2130
rect 9260 2010 9305 2130
rect 9425 2010 9470 2130
rect 9590 2010 9635 2130
rect 9755 2010 9810 2130
rect 9930 2010 9975 2130
rect 10095 2010 10140 2130
rect 10260 2010 10305 2130
rect 10425 2010 10480 2130
rect 10600 2010 10645 2130
rect 10765 2010 10810 2130
rect 10930 2010 10975 2130
rect 11095 2010 11150 2130
rect 11270 2010 11315 2130
rect 11435 2010 11480 2130
rect 11600 2010 11645 2130
rect 11765 2010 11820 2130
rect 11940 2010 11985 2130
rect 12105 2010 12150 2130
rect 12270 2010 12315 2130
rect 12435 2010 12490 2130
rect 12610 2010 12620 2130
rect 7120 1965 12620 2010
rect 7120 1845 7130 1965
rect 7250 1845 7295 1965
rect 7415 1845 7460 1965
rect 7580 1845 7625 1965
rect 7745 1845 7800 1965
rect 7920 1845 7965 1965
rect 8085 1845 8130 1965
rect 8250 1845 8295 1965
rect 8415 1845 8470 1965
rect 8590 1845 8635 1965
rect 8755 1845 8800 1965
rect 8920 1845 8965 1965
rect 9085 1845 9140 1965
rect 9260 1845 9305 1965
rect 9425 1845 9470 1965
rect 9590 1845 9635 1965
rect 9755 1845 9810 1965
rect 9930 1845 9975 1965
rect 10095 1845 10140 1965
rect 10260 1845 10305 1965
rect 10425 1845 10480 1965
rect 10600 1845 10645 1965
rect 10765 1845 10810 1965
rect 10930 1845 10975 1965
rect 11095 1845 11150 1965
rect 11270 1845 11315 1965
rect 11435 1845 11480 1965
rect 11600 1845 11645 1965
rect 11765 1845 11820 1965
rect 11940 1845 11985 1965
rect 12105 1845 12150 1965
rect 12270 1845 12315 1965
rect 12435 1845 12490 1965
rect 12610 1845 12620 1965
rect 7120 1800 12620 1845
rect 7120 1680 7130 1800
rect 7250 1680 7295 1800
rect 7415 1680 7460 1800
rect 7580 1680 7625 1800
rect 7745 1680 7800 1800
rect 7920 1680 7965 1800
rect 8085 1680 8130 1800
rect 8250 1680 8295 1800
rect 8415 1680 8470 1800
rect 8590 1680 8635 1800
rect 8755 1680 8800 1800
rect 8920 1680 8965 1800
rect 9085 1680 9140 1800
rect 9260 1680 9305 1800
rect 9425 1680 9470 1800
rect 9590 1680 9635 1800
rect 9755 1680 9810 1800
rect 9930 1680 9975 1800
rect 10095 1680 10140 1800
rect 10260 1680 10305 1800
rect 10425 1680 10480 1800
rect 10600 1680 10645 1800
rect 10765 1680 10810 1800
rect 10930 1680 10975 1800
rect 11095 1680 11150 1800
rect 11270 1680 11315 1800
rect 11435 1680 11480 1800
rect 11600 1680 11645 1800
rect 11765 1680 11820 1800
rect 11940 1680 11985 1800
rect 12105 1680 12150 1800
rect 12270 1680 12315 1800
rect 12435 1680 12490 1800
rect 12610 1680 12620 1800
rect 7120 1670 12620 1680
rect 12810 7160 18310 7170
rect 12810 7040 12820 7160
rect 12940 7040 12985 7160
rect 13105 7040 13150 7160
rect 13270 7040 13315 7160
rect 13435 7040 13490 7160
rect 13610 7040 13655 7160
rect 13775 7040 13820 7160
rect 13940 7040 13985 7160
rect 14105 7040 14160 7160
rect 14280 7040 14325 7160
rect 14445 7040 14490 7160
rect 14610 7040 14655 7160
rect 14775 7040 14830 7160
rect 14950 7040 14995 7160
rect 15115 7040 15160 7160
rect 15280 7040 15325 7160
rect 15445 7040 15500 7160
rect 15620 7040 15665 7160
rect 15785 7040 15830 7160
rect 15950 7040 15995 7160
rect 16115 7040 16170 7160
rect 16290 7040 16335 7160
rect 16455 7040 16500 7160
rect 16620 7040 16665 7160
rect 16785 7040 16840 7160
rect 16960 7040 17005 7160
rect 17125 7040 17170 7160
rect 17290 7040 17335 7160
rect 17455 7040 17510 7160
rect 17630 7040 17675 7160
rect 17795 7040 17840 7160
rect 17960 7040 18005 7160
rect 18125 7040 18180 7160
rect 18300 7040 18310 7160
rect 12810 6985 18310 7040
rect 12810 6865 12820 6985
rect 12940 6865 12985 6985
rect 13105 6865 13150 6985
rect 13270 6865 13315 6985
rect 13435 6865 13490 6985
rect 13610 6865 13655 6985
rect 13775 6865 13820 6985
rect 13940 6865 13985 6985
rect 14105 6865 14160 6985
rect 14280 6865 14325 6985
rect 14445 6865 14490 6985
rect 14610 6865 14655 6985
rect 14775 6865 14830 6985
rect 14950 6865 14995 6985
rect 15115 6865 15160 6985
rect 15280 6865 15325 6985
rect 15445 6865 15500 6985
rect 15620 6865 15665 6985
rect 15785 6865 15830 6985
rect 15950 6865 15995 6985
rect 16115 6865 16170 6985
rect 16290 6865 16335 6985
rect 16455 6865 16500 6985
rect 16620 6865 16665 6985
rect 16785 6865 16840 6985
rect 16960 6865 17005 6985
rect 17125 6865 17170 6985
rect 17290 6865 17335 6985
rect 17455 6865 17510 6985
rect 17630 6865 17675 6985
rect 17795 6865 17840 6985
rect 17960 6865 18005 6985
rect 18125 6865 18180 6985
rect 18300 6865 18310 6985
rect 12810 6820 18310 6865
rect 12810 6700 12820 6820
rect 12940 6700 12985 6820
rect 13105 6700 13150 6820
rect 13270 6700 13315 6820
rect 13435 6700 13490 6820
rect 13610 6700 13655 6820
rect 13775 6700 13820 6820
rect 13940 6700 13985 6820
rect 14105 6700 14160 6820
rect 14280 6700 14325 6820
rect 14445 6700 14490 6820
rect 14610 6700 14655 6820
rect 14775 6700 14830 6820
rect 14950 6700 14995 6820
rect 15115 6700 15160 6820
rect 15280 6700 15325 6820
rect 15445 6700 15500 6820
rect 15620 6700 15665 6820
rect 15785 6700 15830 6820
rect 15950 6700 15995 6820
rect 16115 6700 16170 6820
rect 16290 6700 16335 6820
rect 16455 6700 16500 6820
rect 16620 6700 16665 6820
rect 16785 6700 16840 6820
rect 16960 6700 17005 6820
rect 17125 6700 17170 6820
rect 17290 6700 17335 6820
rect 17455 6700 17510 6820
rect 17630 6700 17675 6820
rect 17795 6700 17840 6820
rect 17960 6700 18005 6820
rect 18125 6700 18180 6820
rect 18300 6700 18310 6820
rect 12810 6655 18310 6700
rect 12810 6535 12820 6655
rect 12940 6535 12985 6655
rect 13105 6535 13150 6655
rect 13270 6535 13315 6655
rect 13435 6535 13490 6655
rect 13610 6535 13655 6655
rect 13775 6535 13820 6655
rect 13940 6535 13985 6655
rect 14105 6535 14160 6655
rect 14280 6535 14325 6655
rect 14445 6535 14490 6655
rect 14610 6535 14655 6655
rect 14775 6535 14830 6655
rect 14950 6535 14995 6655
rect 15115 6535 15160 6655
rect 15280 6535 15325 6655
rect 15445 6535 15500 6655
rect 15620 6535 15665 6655
rect 15785 6535 15830 6655
rect 15950 6535 15995 6655
rect 16115 6535 16170 6655
rect 16290 6535 16335 6655
rect 16455 6535 16500 6655
rect 16620 6535 16665 6655
rect 16785 6535 16840 6655
rect 16960 6535 17005 6655
rect 17125 6535 17170 6655
rect 17290 6535 17335 6655
rect 17455 6535 17510 6655
rect 17630 6535 17675 6655
rect 17795 6535 17840 6655
rect 17960 6535 18005 6655
rect 18125 6535 18180 6655
rect 18300 6535 18310 6655
rect 12810 6490 18310 6535
rect 12810 6370 12820 6490
rect 12940 6370 12985 6490
rect 13105 6370 13150 6490
rect 13270 6370 13315 6490
rect 13435 6370 13490 6490
rect 13610 6370 13655 6490
rect 13775 6370 13820 6490
rect 13940 6370 13985 6490
rect 14105 6370 14160 6490
rect 14280 6370 14325 6490
rect 14445 6370 14490 6490
rect 14610 6370 14655 6490
rect 14775 6370 14830 6490
rect 14950 6370 14995 6490
rect 15115 6370 15160 6490
rect 15280 6370 15325 6490
rect 15445 6370 15500 6490
rect 15620 6370 15665 6490
rect 15785 6370 15830 6490
rect 15950 6370 15995 6490
rect 16115 6370 16170 6490
rect 16290 6370 16335 6490
rect 16455 6370 16500 6490
rect 16620 6370 16665 6490
rect 16785 6370 16840 6490
rect 16960 6370 17005 6490
rect 17125 6370 17170 6490
rect 17290 6370 17335 6490
rect 17455 6370 17510 6490
rect 17630 6370 17675 6490
rect 17795 6370 17840 6490
rect 17960 6370 18005 6490
rect 18125 6370 18180 6490
rect 18300 6370 18310 6490
rect 12810 6315 18310 6370
rect 12810 6195 12820 6315
rect 12940 6195 12985 6315
rect 13105 6195 13150 6315
rect 13270 6195 13315 6315
rect 13435 6195 13490 6315
rect 13610 6195 13655 6315
rect 13775 6195 13820 6315
rect 13940 6195 13985 6315
rect 14105 6195 14160 6315
rect 14280 6195 14325 6315
rect 14445 6195 14490 6315
rect 14610 6195 14655 6315
rect 14775 6195 14830 6315
rect 14950 6195 14995 6315
rect 15115 6195 15160 6315
rect 15280 6195 15325 6315
rect 15445 6195 15500 6315
rect 15620 6195 15665 6315
rect 15785 6195 15830 6315
rect 15950 6195 15995 6315
rect 16115 6195 16170 6315
rect 16290 6195 16335 6315
rect 16455 6195 16500 6315
rect 16620 6195 16665 6315
rect 16785 6195 16840 6315
rect 16960 6195 17005 6315
rect 17125 6195 17170 6315
rect 17290 6195 17335 6315
rect 17455 6195 17510 6315
rect 17630 6195 17675 6315
rect 17795 6195 17840 6315
rect 17960 6195 18005 6315
rect 18125 6195 18180 6315
rect 18300 6195 18310 6315
rect 12810 6150 18310 6195
rect 12810 6030 12820 6150
rect 12940 6030 12985 6150
rect 13105 6030 13150 6150
rect 13270 6030 13315 6150
rect 13435 6030 13490 6150
rect 13610 6030 13655 6150
rect 13775 6030 13820 6150
rect 13940 6030 13985 6150
rect 14105 6030 14160 6150
rect 14280 6030 14325 6150
rect 14445 6030 14490 6150
rect 14610 6030 14655 6150
rect 14775 6030 14830 6150
rect 14950 6030 14995 6150
rect 15115 6030 15160 6150
rect 15280 6030 15325 6150
rect 15445 6030 15500 6150
rect 15620 6030 15665 6150
rect 15785 6030 15830 6150
rect 15950 6030 15995 6150
rect 16115 6030 16170 6150
rect 16290 6030 16335 6150
rect 16455 6030 16500 6150
rect 16620 6030 16665 6150
rect 16785 6030 16840 6150
rect 16960 6030 17005 6150
rect 17125 6030 17170 6150
rect 17290 6030 17335 6150
rect 17455 6030 17510 6150
rect 17630 6030 17675 6150
rect 17795 6030 17840 6150
rect 17960 6030 18005 6150
rect 18125 6030 18180 6150
rect 18300 6030 18310 6150
rect 12810 5985 18310 6030
rect 12810 5865 12820 5985
rect 12940 5865 12985 5985
rect 13105 5865 13150 5985
rect 13270 5865 13315 5985
rect 13435 5865 13490 5985
rect 13610 5865 13655 5985
rect 13775 5865 13820 5985
rect 13940 5865 13985 5985
rect 14105 5865 14160 5985
rect 14280 5865 14325 5985
rect 14445 5865 14490 5985
rect 14610 5865 14655 5985
rect 14775 5865 14830 5985
rect 14950 5865 14995 5985
rect 15115 5865 15160 5985
rect 15280 5865 15325 5985
rect 15445 5865 15500 5985
rect 15620 5865 15665 5985
rect 15785 5865 15830 5985
rect 15950 5865 15995 5985
rect 16115 5865 16170 5985
rect 16290 5865 16335 5985
rect 16455 5865 16500 5985
rect 16620 5865 16665 5985
rect 16785 5865 16840 5985
rect 16960 5865 17005 5985
rect 17125 5865 17170 5985
rect 17290 5865 17335 5985
rect 17455 5865 17510 5985
rect 17630 5865 17675 5985
rect 17795 5865 17840 5985
rect 17960 5865 18005 5985
rect 18125 5865 18180 5985
rect 18300 5865 18310 5985
rect 12810 5820 18310 5865
rect 12810 5700 12820 5820
rect 12940 5700 12985 5820
rect 13105 5700 13150 5820
rect 13270 5700 13315 5820
rect 13435 5700 13490 5820
rect 13610 5700 13655 5820
rect 13775 5700 13820 5820
rect 13940 5700 13985 5820
rect 14105 5700 14160 5820
rect 14280 5700 14325 5820
rect 14445 5700 14490 5820
rect 14610 5700 14655 5820
rect 14775 5700 14830 5820
rect 14950 5700 14995 5820
rect 15115 5700 15160 5820
rect 15280 5700 15325 5820
rect 15445 5700 15500 5820
rect 15620 5700 15665 5820
rect 15785 5700 15830 5820
rect 15950 5700 15995 5820
rect 16115 5700 16170 5820
rect 16290 5700 16335 5820
rect 16455 5700 16500 5820
rect 16620 5700 16665 5820
rect 16785 5700 16840 5820
rect 16960 5700 17005 5820
rect 17125 5700 17170 5820
rect 17290 5700 17335 5820
rect 17455 5700 17510 5820
rect 17630 5700 17675 5820
rect 17795 5700 17840 5820
rect 17960 5700 18005 5820
rect 18125 5700 18180 5820
rect 18300 5700 18310 5820
rect 12810 5645 18310 5700
rect 12810 5525 12820 5645
rect 12940 5525 12985 5645
rect 13105 5525 13150 5645
rect 13270 5525 13315 5645
rect 13435 5525 13490 5645
rect 13610 5525 13655 5645
rect 13775 5525 13820 5645
rect 13940 5525 13985 5645
rect 14105 5525 14160 5645
rect 14280 5525 14325 5645
rect 14445 5525 14490 5645
rect 14610 5525 14655 5645
rect 14775 5525 14830 5645
rect 14950 5525 14995 5645
rect 15115 5525 15160 5645
rect 15280 5525 15325 5645
rect 15445 5525 15500 5645
rect 15620 5525 15665 5645
rect 15785 5525 15830 5645
rect 15950 5525 15995 5645
rect 16115 5525 16170 5645
rect 16290 5525 16335 5645
rect 16455 5525 16500 5645
rect 16620 5525 16665 5645
rect 16785 5525 16840 5645
rect 16960 5525 17005 5645
rect 17125 5525 17170 5645
rect 17290 5525 17335 5645
rect 17455 5525 17510 5645
rect 17630 5525 17675 5645
rect 17795 5525 17840 5645
rect 17960 5525 18005 5645
rect 18125 5525 18180 5645
rect 18300 5525 18310 5645
rect 12810 5480 18310 5525
rect 12810 5360 12820 5480
rect 12940 5360 12985 5480
rect 13105 5360 13150 5480
rect 13270 5360 13315 5480
rect 13435 5360 13490 5480
rect 13610 5360 13655 5480
rect 13775 5360 13820 5480
rect 13940 5360 13985 5480
rect 14105 5360 14160 5480
rect 14280 5360 14325 5480
rect 14445 5360 14490 5480
rect 14610 5360 14655 5480
rect 14775 5360 14830 5480
rect 14950 5360 14995 5480
rect 15115 5360 15160 5480
rect 15280 5360 15325 5480
rect 15445 5360 15500 5480
rect 15620 5360 15665 5480
rect 15785 5360 15830 5480
rect 15950 5360 15995 5480
rect 16115 5360 16170 5480
rect 16290 5360 16335 5480
rect 16455 5360 16500 5480
rect 16620 5360 16665 5480
rect 16785 5360 16840 5480
rect 16960 5360 17005 5480
rect 17125 5360 17170 5480
rect 17290 5360 17335 5480
rect 17455 5360 17510 5480
rect 17630 5360 17675 5480
rect 17795 5360 17840 5480
rect 17960 5360 18005 5480
rect 18125 5360 18180 5480
rect 18300 5360 18310 5480
rect 12810 5315 18310 5360
rect 12810 5195 12820 5315
rect 12940 5195 12985 5315
rect 13105 5195 13150 5315
rect 13270 5195 13315 5315
rect 13435 5195 13490 5315
rect 13610 5195 13655 5315
rect 13775 5195 13820 5315
rect 13940 5195 13985 5315
rect 14105 5195 14160 5315
rect 14280 5195 14325 5315
rect 14445 5195 14490 5315
rect 14610 5195 14655 5315
rect 14775 5195 14830 5315
rect 14950 5195 14995 5315
rect 15115 5195 15160 5315
rect 15280 5195 15325 5315
rect 15445 5195 15500 5315
rect 15620 5195 15665 5315
rect 15785 5195 15830 5315
rect 15950 5195 15995 5315
rect 16115 5195 16170 5315
rect 16290 5195 16335 5315
rect 16455 5195 16500 5315
rect 16620 5195 16665 5315
rect 16785 5195 16840 5315
rect 16960 5195 17005 5315
rect 17125 5195 17170 5315
rect 17290 5195 17335 5315
rect 17455 5195 17510 5315
rect 17630 5195 17675 5315
rect 17795 5195 17840 5315
rect 17960 5195 18005 5315
rect 18125 5195 18180 5315
rect 18300 5195 18310 5315
rect 12810 5150 18310 5195
rect 12810 5030 12820 5150
rect 12940 5030 12985 5150
rect 13105 5030 13150 5150
rect 13270 5030 13315 5150
rect 13435 5030 13490 5150
rect 13610 5030 13655 5150
rect 13775 5030 13820 5150
rect 13940 5030 13985 5150
rect 14105 5030 14160 5150
rect 14280 5030 14325 5150
rect 14445 5030 14490 5150
rect 14610 5030 14655 5150
rect 14775 5030 14830 5150
rect 14950 5030 14995 5150
rect 15115 5030 15160 5150
rect 15280 5030 15325 5150
rect 15445 5030 15500 5150
rect 15620 5030 15665 5150
rect 15785 5030 15830 5150
rect 15950 5030 15995 5150
rect 16115 5030 16170 5150
rect 16290 5030 16335 5150
rect 16455 5030 16500 5150
rect 16620 5030 16665 5150
rect 16785 5030 16840 5150
rect 16960 5030 17005 5150
rect 17125 5030 17170 5150
rect 17290 5030 17335 5150
rect 17455 5030 17510 5150
rect 17630 5030 17675 5150
rect 17795 5030 17840 5150
rect 17960 5030 18005 5150
rect 18125 5030 18180 5150
rect 18300 5030 18310 5150
rect 12810 4975 18310 5030
rect 12810 4855 12820 4975
rect 12940 4855 12985 4975
rect 13105 4855 13150 4975
rect 13270 4855 13315 4975
rect 13435 4855 13490 4975
rect 13610 4855 13655 4975
rect 13775 4855 13820 4975
rect 13940 4855 13985 4975
rect 14105 4855 14160 4975
rect 14280 4855 14325 4975
rect 14445 4855 14490 4975
rect 14610 4855 14655 4975
rect 14775 4855 14830 4975
rect 14950 4855 14995 4975
rect 15115 4855 15160 4975
rect 15280 4855 15325 4975
rect 15445 4855 15500 4975
rect 15620 4855 15665 4975
rect 15785 4855 15830 4975
rect 15950 4855 15995 4975
rect 16115 4855 16170 4975
rect 16290 4855 16335 4975
rect 16455 4855 16500 4975
rect 16620 4855 16665 4975
rect 16785 4855 16840 4975
rect 16960 4855 17005 4975
rect 17125 4855 17170 4975
rect 17290 4855 17335 4975
rect 17455 4855 17510 4975
rect 17630 4855 17675 4975
rect 17795 4855 17840 4975
rect 17960 4855 18005 4975
rect 18125 4855 18180 4975
rect 18300 4855 18310 4975
rect 12810 4810 18310 4855
rect 12810 4690 12820 4810
rect 12940 4690 12985 4810
rect 13105 4690 13150 4810
rect 13270 4690 13315 4810
rect 13435 4690 13490 4810
rect 13610 4690 13655 4810
rect 13775 4690 13820 4810
rect 13940 4690 13985 4810
rect 14105 4690 14160 4810
rect 14280 4690 14325 4810
rect 14445 4690 14490 4810
rect 14610 4690 14655 4810
rect 14775 4690 14830 4810
rect 14950 4690 14995 4810
rect 15115 4690 15160 4810
rect 15280 4690 15325 4810
rect 15445 4690 15500 4810
rect 15620 4690 15665 4810
rect 15785 4690 15830 4810
rect 15950 4690 15995 4810
rect 16115 4690 16170 4810
rect 16290 4690 16335 4810
rect 16455 4690 16500 4810
rect 16620 4690 16665 4810
rect 16785 4690 16840 4810
rect 16960 4690 17005 4810
rect 17125 4690 17170 4810
rect 17290 4690 17335 4810
rect 17455 4690 17510 4810
rect 17630 4690 17675 4810
rect 17795 4690 17840 4810
rect 17960 4690 18005 4810
rect 18125 4690 18180 4810
rect 18300 4690 18310 4810
rect 12810 4645 18310 4690
rect 12810 4525 12820 4645
rect 12940 4525 12985 4645
rect 13105 4525 13150 4645
rect 13270 4525 13315 4645
rect 13435 4525 13490 4645
rect 13610 4525 13655 4645
rect 13775 4525 13820 4645
rect 13940 4525 13985 4645
rect 14105 4525 14160 4645
rect 14280 4525 14325 4645
rect 14445 4525 14490 4645
rect 14610 4525 14655 4645
rect 14775 4525 14830 4645
rect 14950 4525 14995 4645
rect 15115 4525 15160 4645
rect 15280 4525 15325 4645
rect 15445 4525 15500 4645
rect 15620 4525 15665 4645
rect 15785 4525 15830 4645
rect 15950 4525 15995 4645
rect 16115 4525 16170 4645
rect 16290 4525 16335 4645
rect 16455 4525 16500 4645
rect 16620 4525 16665 4645
rect 16785 4525 16840 4645
rect 16960 4525 17005 4645
rect 17125 4525 17170 4645
rect 17290 4525 17335 4645
rect 17455 4525 17510 4645
rect 17630 4525 17675 4645
rect 17795 4525 17840 4645
rect 17960 4525 18005 4645
rect 18125 4525 18180 4645
rect 18300 4525 18310 4645
rect 12810 4480 18310 4525
rect 12810 4360 12820 4480
rect 12940 4360 12985 4480
rect 13105 4360 13150 4480
rect 13270 4360 13315 4480
rect 13435 4360 13490 4480
rect 13610 4360 13655 4480
rect 13775 4360 13820 4480
rect 13940 4360 13985 4480
rect 14105 4360 14160 4480
rect 14280 4360 14325 4480
rect 14445 4360 14490 4480
rect 14610 4360 14655 4480
rect 14775 4360 14830 4480
rect 14950 4360 14995 4480
rect 15115 4360 15160 4480
rect 15280 4360 15325 4480
rect 15445 4360 15500 4480
rect 15620 4360 15665 4480
rect 15785 4360 15830 4480
rect 15950 4360 15995 4480
rect 16115 4360 16170 4480
rect 16290 4360 16335 4480
rect 16455 4360 16500 4480
rect 16620 4360 16665 4480
rect 16785 4360 16840 4480
rect 16960 4360 17005 4480
rect 17125 4360 17170 4480
rect 17290 4360 17335 4480
rect 17455 4360 17510 4480
rect 17630 4360 17675 4480
rect 17795 4360 17840 4480
rect 17960 4360 18005 4480
rect 18125 4360 18180 4480
rect 18300 4360 18310 4480
rect 12810 4305 18310 4360
rect 12810 4185 12820 4305
rect 12940 4185 12985 4305
rect 13105 4185 13150 4305
rect 13270 4185 13315 4305
rect 13435 4185 13490 4305
rect 13610 4185 13655 4305
rect 13775 4185 13820 4305
rect 13940 4185 13985 4305
rect 14105 4185 14160 4305
rect 14280 4185 14325 4305
rect 14445 4185 14490 4305
rect 14610 4185 14655 4305
rect 14775 4185 14830 4305
rect 14950 4185 14995 4305
rect 15115 4185 15160 4305
rect 15280 4185 15325 4305
rect 15445 4185 15500 4305
rect 15620 4185 15665 4305
rect 15785 4185 15830 4305
rect 15950 4185 15995 4305
rect 16115 4185 16170 4305
rect 16290 4185 16335 4305
rect 16455 4185 16500 4305
rect 16620 4185 16665 4305
rect 16785 4185 16840 4305
rect 16960 4185 17005 4305
rect 17125 4185 17170 4305
rect 17290 4185 17335 4305
rect 17455 4185 17510 4305
rect 17630 4185 17675 4305
rect 17795 4185 17840 4305
rect 17960 4185 18005 4305
rect 18125 4185 18180 4305
rect 18300 4185 18310 4305
rect 12810 4140 18310 4185
rect 12810 4020 12820 4140
rect 12940 4020 12985 4140
rect 13105 4020 13150 4140
rect 13270 4020 13315 4140
rect 13435 4020 13490 4140
rect 13610 4020 13655 4140
rect 13775 4020 13820 4140
rect 13940 4020 13985 4140
rect 14105 4020 14160 4140
rect 14280 4020 14325 4140
rect 14445 4020 14490 4140
rect 14610 4020 14655 4140
rect 14775 4020 14830 4140
rect 14950 4020 14995 4140
rect 15115 4020 15160 4140
rect 15280 4020 15325 4140
rect 15445 4020 15500 4140
rect 15620 4020 15665 4140
rect 15785 4020 15830 4140
rect 15950 4020 15995 4140
rect 16115 4020 16170 4140
rect 16290 4020 16335 4140
rect 16455 4020 16500 4140
rect 16620 4020 16665 4140
rect 16785 4020 16840 4140
rect 16960 4020 17005 4140
rect 17125 4020 17170 4140
rect 17290 4020 17335 4140
rect 17455 4020 17510 4140
rect 17630 4020 17675 4140
rect 17795 4020 17840 4140
rect 17960 4020 18005 4140
rect 18125 4020 18180 4140
rect 18300 4020 18310 4140
rect 12810 3975 18310 4020
rect 12810 3855 12820 3975
rect 12940 3855 12985 3975
rect 13105 3855 13150 3975
rect 13270 3855 13315 3975
rect 13435 3855 13490 3975
rect 13610 3855 13655 3975
rect 13775 3855 13820 3975
rect 13940 3855 13985 3975
rect 14105 3855 14160 3975
rect 14280 3855 14325 3975
rect 14445 3855 14490 3975
rect 14610 3855 14655 3975
rect 14775 3855 14830 3975
rect 14950 3855 14995 3975
rect 15115 3855 15160 3975
rect 15280 3855 15325 3975
rect 15445 3855 15500 3975
rect 15620 3855 15665 3975
rect 15785 3855 15830 3975
rect 15950 3855 15995 3975
rect 16115 3855 16170 3975
rect 16290 3855 16335 3975
rect 16455 3855 16500 3975
rect 16620 3855 16665 3975
rect 16785 3855 16840 3975
rect 16960 3855 17005 3975
rect 17125 3855 17170 3975
rect 17290 3855 17335 3975
rect 17455 3855 17510 3975
rect 17630 3855 17675 3975
rect 17795 3855 17840 3975
rect 17960 3855 18005 3975
rect 18125 3855 18180 3975
rect 18300 3855 18310 3975
rect 12810 3810 18310 3855
rect 12810 3690 12820 3810
rect 12940 3690 12985 3810
rect 13105 3690 13150 3810
rect 13270 3690 13315 3810
rect 13435 3690 13490 3810
rect 13610 3690 13655 3810
rect 13775 3690 13820 3810
rect 13940 3690 13985 3810
rect 14105 3690 14160 3810
rect 14280 3690 14325 3810
rect 14445 3690 14490 3810
rect 14610 3690 14655 3810
rect 14775 3690 14830 3810
rect 14950 3690 14995 3810
rect 15115 3690 15160 3810
rect 15280 3690 15325 3810
rect 15445 3690 15500 3810
rect 15620 3690 15665 3810
rect 15785 3690 15830 3810
rect 15950 3690 15995 3810
rect 16115 3690 16170 3810
rect 16290 3690 16335 3810
rect 16455 3690 16500 3810
rect 16620 3690 16665 3810
rect 16785 3690 16840 3810
rect 16960 3690 17005 3810
rect 17125 3690 17170 3810
rect 17290 3690 17335 3810
rect 17455 3690 17510 3810
rect 17630 3690 17675 3810
rect 17795 3690 17840 3810
rect 17960 3690 18005 3810
rect 18125 3690 18180 3810
rect 18300 3690 18310 3810
rect 12810 3635 18310 3690
rect 12810 3515 12820 3635
rect 12940 3515 12985 3635
rect 13105 3515 13150 3635
rect 13270 3515 13315 3635
rect 13435 3515 13490 3635
rect 13610 3515 13655 3635
rect 13775 3515 13820 3635
rect 13940 3515 13985 3635
rect 14105 3515 14160 3635
rect 14280 3515 14325 3635
rect 14445 3515 14490 3635
rect 14610 3515 14655 3635
rect 14775 3515 14830 3635
rect 14950 3515 14995 3635
rect 15115 3515 15160 3635
rect 15280 3515 15325 3635
rect 15445 3515 15500 3635
rect 15620 3515 15665 3635
rect 15785 3515 15830 3635
rect 15950 3515 15995 3635
rect 16115 3515 16170 3635
rect 16290 3515 16335 3635
rect 16455 3515 16500 3635
rect 16620 3515 16665 3635
rect 16785 3515 16840 3635
rect 16960 3515 17005 3635
rect 17125 3515 17170 3635
rect 17290 3515 17335 3635
rect 17455 3515 17510 3635
rect 17630 3515 17675 3635
rect 17795 3515 17840 3635
rect 17960 3515 18005 3635
rect 18125 3515 18180 3635
rect 18300 3515 18310 3635
rect 12810 3470 18310 3515
rect 12810 3350 12820 3470
rect 12940 3350 12985 3470
rect 13105 3350 13150 3470
rect 13270 3350 13315 3470
rect 13435 3350 13490 3470
rect 13610 3350 13655 3470
rect 13775 3350 13820 3470
rect 13940 3350 13985 3470
rect 14105 3350 14160 3470
rect 14280 3350 14325 3470
rect 14445 3350 14490 3470
rect 14610 3350 14655 3470
rect 14775 3350 14830 3470
rect 14950 3350 14995 3470
rect 15115 3350 15160 3470
rect 15280 3350 15325 3470
rect 15445 3350 15500 3470
rect 15620 3350 15665 3470
rect 15785 3350 15830 3470
rect 15950 3350 15995 3470
rect 16115 3350 16170 3470
rect 16290 3350 16335 3470
rect 16455 3350 16500 3470
rect 16620 3350 16665 3470
rect 16785 3350 16840 3470
rect 16960 3350 17005 3470
rect 17125 3350 17170 3470
rect 17290 3350 17335 3470
rect 17455 3350 17510 3470
rect 17630 3350 17675 3470
rect 17795 3350 17840 3470
rect 17960 3350 18005 3470
rect 18125 3350 18180 3470
rect 18300 3350 18310 3470
rect 12810 3305 18310 3350
rect 12810 3185 12820 3305
rect 12940 3185 12985 3305
rect 13105 3185 13150 3305
rect 13270 3185 13315 3305
rect 13435 3185 13490 3305
rect 13610 3185 13655 3305
rect 13775 3185 13820 3305
rect 13940 3185 13985 3305
rect 14105 3185 14160 3305
rect 14280 3185 14325 3305
rect 14445 3185 14490 3305
rect 14610 3185 14655 3305
rect 14775 3185 14830 3305
rect 14950 3185 14995 3305
rect 15115 3185 15160 3305
rect 15280 3185 15325 3305
rect 15445 3185 15500 3305
rect 15620 3185 15665 3305
rect 15785 3185 15830 3305
rect 15950 3185 15995 3305
rect 16115 3185 16170 3305
rect 16290 3185 16335 3305
rect 16455 3185 16500 3305
rect 16620 3185 16665 3305
rect 16785 3185 16840 3305
rect 16960 3185 17005 3305
rect 17125 3185 17170 3305
rect 17290 3185 17335 3305
rect 17455 3185 17510 3305
rect 17630 3185 17675 3305
rect 17795 3185 17840 3305
rect 17960 3185 18005 3305
rect 18125 3185 18180 3305
rect 18300 3185 18310 3305
rect 12810 3140 18310 3185
rect 12810 3020 12820 3140
rect 12940 3020 12985 3140
rect 13105 3020 13150 3140
rect 13270 3020 13315 3140
rect 13435 3020 13490 3140
rect 13610 3020 13655 3140
rect 13775 3020 13820 3140
rect 13940 3020 13985 3140
rect 14105 3020 14160 3140
rect 14280 3020 14325 3140
rect 14445 3020 14490 3140
rect 14610 3020 14655 3140
rect 14775 3020 14830 3140
rect 14950 3020 14995 3140
rect 15115 3020 15160 3140
rect 15280 3020 15325 3140
rect 15445 3020 15500 3140
rect 15620 3020 15665 3140
rect 15785 3020 15830 3140
rect 15950 3020 15995 3140
rect 16115 3020 16170 3140
rect 16290 3020 16335 3140
rect 16455 3020 16500 3140
rect 16620 3020 16665 3140
rect 16785 3020 16840 3140
rect 16960 3020 17005 3140
rect 17125 3020 17170 3140
rect 17290 3020 17335 3140
rect 17455 3020 17510 3140
rect 17630 3020 17675 3140
rect 17795 3020 17840 3140
rect 17960 3020 18005 3140
rect 18125 3020 18180 3140
rect 18300 3020 18310 3140
rect 12810 2965 18310 3020
rect 12810 2845 12820 2965
rect 12940 2845 12985 2965
rect 13105 2845 13150 2965
rect 13270 2845 13315 2965
rect 13435 2845 13490 2965
rect 13610 2845 13655 2965
rect 13775 2845 13820 2965
rect 13940 2845 13985 2965
rect 14105 2845 14160 2965
rect 14280 2845 14325 2965
rect 14445 2845 14490 2965
rect 14610 2845 14655 2965
rect 14775 2845 14830 2965
rect 14950 2845 14995 2965
rect 15115 2845 15160 2965
rect 15280 2845 15325 2965
rect 15445 2845 15500 2965
rect 15620 2845 15665 2965
rect 15785 2845 15830 2965
rect 15950 2845 15995 2965
rect 16115 2845 16170 2965
rect 16290 2845 16335 2965
rect 16455 2845 16500 2965
rect 16620 2845 16665 2965
rect 16785 2845 16840 2965
rect 16960 2845 17005 2965
rect 17125 2845 17170 2965
rect 17290 2845 17335 2965
rect 17455 2845 17510 2965
rect 17630 2845 17675 2965
rect 17795 2845 17840 2965
rect 17960 2845 18005 2965
rect 18125 2845 18180 2965
rect 18300 2845 18310 2965
rect 12810 2800 18310 2845
rect 12810 2680 12820 2800
rect 12940 2680 12985 2800
rect 13105 2680 13150 2800
rect 13270 2680 13315 2800
rect 13435 2680 13490 2800
rect 13610 2680 13655 2800
rect 13775 2680 13820 2800
rect 13940 2680 13985 2800
rect 14105 2680 14160 2800
rect 14280 2680 14325 2800
rect 14445 2680 14490 2800
rect 14610 2680 14655 2800
rect 14775 2680 14830 2800
rect 14950 2680 14995 2800
rect 15115 2680 15160 2800
rect 15280 2680 15325 2800
rect 15445 2680 15500 2800
rect 15620 2680 15665 2800
rect 15785 2680 15830 2800
rect 15950 2680 15995 2800
rect 16115 2680 16170 2800
rect 16290 2680 16335 2800
rect 16455 2680 16500 2800
rect 16620 2680 16665 2800
rect 16785 2680 16840 2800
rect 16960 2680 17005 2800
rect 17125 2680 17170 2800
rect 17290 2680 17335 2800
rect 17455 2680 17510 2800
rect 17630 2680 17675 2800
rect 17795 2680 17840 2800
rect 17960 2680 18005 2800
rect 18125 2680 18180 2800
rect 18300 2680 18310 2800
rect 12810 2635 18310 2680
rect 12810 2515 12820 2635
rect 12940 2515 12985 2635
rect 13105 2515 13150 2635
rect 13270 2515 13315 2635
rect 13435 2515 13490 2635
rect 13610 2515 13655 2635
rect 13775 2515 13820 2635
rect 13940 2515 13985 2635
rect 14105 2515 14160 2635
rect 14280 2515 14325 2635
rect 14445 2515 14490 2635
rect 14610 2515 14655 2635
rect 14775 2515 14830 2635
rect 14950 2515 14995 2635
rect 15115 2515 15160 2635
rect 15280 2515 15325 2635
rect 15445 2515 15500 2635
rect 15620 2515 15665 2635
rect 15785 2515 15830 2635
rect 15950 2515 15995 2635
rect 16115 2515 16170 2635
rect 16290 2515 16335 2635
rect 16455 2515 16500 2635
rect 16620 2515 16665 2635
rect 16785 2515 16840 2635
rect 16960 2515 17005 2635
rect 17125 2515 17170 2635
rect 17290 2515 17335 2635
rect 17455 2515 17510 2635
rect 17630 2515 17675 2635
rect 17795 2515 17840 2635
rect 17960 2515 18005 2635
rect 18125 2515 18180 2635
rect 18300 2515 18310 2635
rect 12810 2470 18310 2515
rect 12810 2350 12820 2470
rect 12940 2350 12985 2470
rect 13105 2350 13150 2470
rect 13270 2350 13315 2470
rect 13435 2350 13490 2470
rect 13610 2350 13655 2470
rect 13775 2350 13820 2470
rect 13940 2350 13985 2470
rect 14105 2350 14160 2470
rect 14280 2350 14325 2470
rect 14445 2350 14490 2470
rect 14610 2350 14655 2470
rect 14775 2350 14830 2470
rect 14950 2350 14995 2470
rect 15115 2350 15160 2470
rect 15280 2350 15325 2470
rect 15445 2350 15500 2470
rect 15620 2350 15665 2470
rect 15785 2350 15830 2470
rect 15950 2350 15995 2470
rect 16115 2350 16170 2470
rect 16290 2350 16335 2470
rect 16455 2350 16500 2470
rect 16620 2350 16665 2470
rect 16785 2350 16840 2470
rect 16960 2350 17005 2470
rect 17125 2350 17170 2470
rect 17290 2350 17335 2470
rect 17455 2350 17510 2470
rect 17630 2350 17675 2470
rect 17795 2350 17840 2470
rect 17960 2350 18005 2470
rect 18125 2350 18180 2470
rect 18300 2350 18310 2470
rect 12810 2295 18310 2350
rect 12810 2175 12820 2295
rect 12940 2175 12985 2295
rect 13105 2175 13150 2295
rect 13270 2175 13315 2295
rect 13435 2175 13490 2295
rect 13610 2175 13655 2295
rect 13775 2175 13820 2295
rect 13940 2175 13985 2295
rect 14105 2175 14160 2295
rect 14280 2175 14325 2295
rect 14445 2175 14490 2295
rect 14610 2175 14655 2295
rect 14775 2175 14830 2295
rect 14950 2175 14995 2295
rect 15115 2175 15160 2295
rect 15280 2175 15325 2295
rect 15445 2175 15500 2295
rect 15620 2175 15665 2295
rect 15785 2175 15830 2295
rect 15950 2175 15995 2295
rect 16115 2175 16170 2295
rect 16290 2175 16335 2295
rect 16455 2175 16500 2295
rect 16620 2175 16665 2295
rect 16785 2175 16840 2295
rect 16960 2175 17005 2295
rect 17125 2175 17170 2295
rect 17290 2175 17335 2295
rect 17455 2175 17510 2295
rect 17630 2175 17675 2295
rect 17795 2175 17840 2295
rect 17960 2175 18005 2295
rect 18125 2175 18180 2295
rect 18300 2175 18310 2295
rect 12810 2130 18310 2175
rect 12810 2010 12820 2130
rect 12940 2010 12985 2130
rect 13105 2010 13150 2130
rect 13270 2010 13315 2130
rect 13435 2010 13490 2130
rect 13610 2010 13655 2130
rect 13775 2010 13820 2130
rect 13940 2010 13985 2130
rect 14105 2010 14160 2130
rect 14280 2010 14325 2130
rect 14445 2010 14490 2130
rect 14610 2010 14655 2130
rect 14775 2010 14830 2130
rect 14950 2010 14995 2130
rect 15115 2010 15160 2130
rect 15280 2010 15325 2130
rect 15445 2010 15500 2130
rect 15620 2010 15665 2130
rect 15785 2010 15830 2130
rect 15950 2010 15995 2130
rect 16115 2010 16170 2130
rect 16290 2010 16335 2130
rect 16455 2010 16500 2130
rect 16620 2010 16665 2130
rect 16785 2010 16840 2130
rect 16960 2010 17005 2130
rect 17125 2010 17170 2130
rect 17290 2010 17335 2130
rect 17455 2010 17510 2130
rect 17630 2010 17675 2130
rect 17795 2010 17840 2130
rect 17960 2010 18005 2130
rect 18125 2010 18180 2130
rect 18300 2010 18310 2130
rect 12810 1965 18310 2010
rect 12810 1845 12820 1965
rect 12940 1845 12985 1965
rect 13105 1845 13150 1965
rect 13270 1845 13315 1965
rect 13435 1845 13490 1965
rect 13610 1845 13655 1965
rect 13775 1845 13820 1965
rect 13940 1845 13985 1965
rect 14105 1845 14160 1965
rect 14280 1845 14325 1965
rect 14445 1845 14490 1965
rect 14610 1845 14655 1965
rect 14775 1845 14830 1965
rect 14950 1845 14995 1965
rect 15115 1845 15160 1965
rect 15280 1845 15325 1965
rect 15445 1845 15500 1965
rect 15620 1845 15665 1965
rect 15785 1845 15830 1965
rect 15950 1845 15995 1965
rect 16115 1845 16170 1965
rect 16290 1845 16335 1965
rect 16455 1845 16500 1965
rect 16620 1845 16665 1965
rect 16785 1845 16840 1965
rect 16960 1845 17005 1965
rect 17125 1845 17170 1965
rect 17290 1845 17335 1965
rect 17455 1845 17510 1965
rect 17630 1845 17675 1965
rect 17795 1845 17840 1965
rect 17960 1845 18005 1965
rect 18125 1845 18180 1965
rect 18300 1845 18310 1965
rect 12810 1800 18310 1845
rect 12810 1680 12820 1800
rect 12940 1680 12985 1800
rect 13105 1680 13150 1800
rect 13270 1680 13315 1800
rect 13435 1680 13490 1800
rect 13610 1680 13655 1800
rect 13775 1680 13820 1800
rect 13940 1680 13985 1800
rect 14105 1680 14160 1800
rect 14280 1680 14325 1800
rect 14445 1680 14490 1800
rect 14610 1680 14655 1800
rect 14775 1680 14830 1800
rect 14950 1680 14995 1800
rect 15115 1680 15160 1800
rect 15280 1680 15325 1800
rect 15445 1680 15500 1800
rect 15620 1680 15665 1800
rect 15785 1680 15830 1800
rect 15950 1680 15995 1800
rect 16115 1680 16170 1800
rect 16290 1680 16335 1800
rect 16455 1680 16500 1800
rect 16620 1680 16665 1800
rect 16785 1680 16840 1800
rect 16960 1680 17005 1800
rect 17125 1680 17170 1800
rect 17290 1680 17335 1800
rect 17455 1680 17510 1800
rect 17630 1680 17675 1800
rect 17795 1680 17840 1800
rect 17960 1680 18005 1800
rect 18125 1680 18180 1800
rect 18300 1680 18310 1800
rect 12810 1670 18310 1680
rect 18500 7160 24000 7170
rect 18500 7040 18510 7160
rect 18630 7040 18675 7160
rect 18795 7040 18840 7160
rect 18960 7040 19005 7160
rect 19125 7040 19180 7160
rect 19300 7040 19345 7160
rect 19465 7040 19510 7160
rect 19630 7040 19675 7160
rect 19795 7040 19850 7160
rect 19970 7040 20015 7160
rect 20135 7040 20180 7160
rect 20300 7040 20345 7160
rect 20465 7040 20520 7160
rect 20640 7040 20685 7160
rect 20805 7040 20850 7160
rect 20970 7040 21015 7160
rect 21135 7040 21190 7160
rect 21310 7040 21355 7160
rect 21475 7040 21520 7160
rect 21640 7040 21685 7160
rect 21805 7040 21860 7160
rect 21980 7040 22025 7160
rect 22145 7040 22190 7160
rect 22310 7040 22355 7160
rect 22475 7040 22530 7160
rect 22650 7040 22695 7160
rect 22815 7040 22860 7160
rect 22980 7040 23025 7160
rect 23145 7040 23200 7160
rect 23320 7040 23365 7160
rect 23485 7040 23530 7160
rect 23650 7040 23695 7160
rect 23815 7040 23870 7160
rect 23990 7040 24000 7160
rect 18500 6985 24000 7040
rect 18500 6865 18510 6985
rect 18630 6865 18675 6985
rect 18795 6865 18840 6985
rect 18960 6865 19005 6985
rect 19125 6865 19180 6985
rect 19300 6865 19345 6985
rect 19465 6865 19510 6985
rect 19630 6865 19675 6985
rect 19795 6865 19850 6985
rect 19970 6865 20015 6985
rect 20135 6865 20180 6985
rect 20300 6865 20345 6985
rect 20465 6865 20520 6985
rect 20640 6865 20685 6985
rect 20805 6865 20850 6985
rect 20970 6865 21015 6985
rect 21135 6865 21190 6985
rect 21310 6865 21355 6985
rect 21475 6865 21520 6985
rect 21640 6865 21685 6985
rect 21805 6865 21860 6985
rect 21980 6865 22025 6985
rect 22145 6865 22190 6985
rect 22310 6865 22355 6985
rect 22475 6865 22530 6985
rect 22650 6865 22695 6985
rect 22815 6865 22860 6985
rect 22980 6865 23025 6985
rect 23145 6865 23200 6985
rect 23320 6865 23365 6985
rect 23485 6865 23530 6985
rect 23650 6865 23695 6985
rect 23815 6865 23870 6985
rect 23990 6865 24000 6985
rect 18500 6820 24000 6865
rect 18500 6700 18510 6820
rect 18630 6700 18675 6820
rect 18795 6700 18840 6820
rect 18960 6700 19005 6820
rect 19125 6700 19180 6820
rect 19300 6700 19345 6820
rect 19465 6700 19510 6820
rect 19630 6700 19675 6820
rect 19795 6700 19850 6820
rect 19970 6700 20015 6820
rect 20135 6700 20180 6820
rect 20300 6700 20345 6820
rect 20465 6700 20520 6820
rect 20640 6700 20685 6820
rect 20805 6700 20850 6820
rect 20970 6700 21015 6820
rect 21135 6700 21190 6820
rect 21310 6700 21355 6820
rect 21475 6700 21520 6820
rect 21640 6700 21685 6820
rect 21805 6700 21860 6820
rect 21980 6700 22025 6820
rect 22145 6700 22190 6820
rect 22310 6700 22355 6820
rect 22475 6700 22530 6820
rect 22650 6700 22695 6820
rect 22815 6700 22860 6820
rect 22980 6700 23025 6820
rect 23145 6700 23200 6820
rect 23320 6700 23365 6820
rect 23485 6700 23530 6820
rect 23650 6700 23695 6820
rect 23815 6700 23870 6820
rect 23990 6700 24000 6820
rect 18500 6655 24000 6700
rect 18500 6535 18510 6655
rect 18630 6535 18675 6655
rect 18795 6535 18840 6655
rect 18960 6535 19005 6655
rect 19125 6535 19180 6655
rect 19300 6535 19345 6655
rect 19465 6535 19510 6655
rect 19630 6535 19675 6655
rect 19795 6535 19850 6655
rect 19970 6535 20015 6655
rect 20135 6535 20180 6655
rect 20300 6535 20345 6655
rect 20465 6535 20520 6655
rect 20640 6535 20685 6655
rect 20805 6535 20850 6655
rect 20970 6535 21015 6655
rect 21135 6535 21190 6655
rect 21310 6535 21355 6655
rect 21475 6535 21520 6655
rect 21640 6535 21685 6655
rect 21805 6535 21860 6655
rect 21980 6535 22025 6655
rect 22145 6535 22190 6655
rect 22310 6535 22355 6655
rect 22475 6535 22530 6655
rect 22650 6535 22695 6655
rect 22815 6535 22860 6655
rect 22980 6535 23025 6655
rect 23145 6535 23200 6655
rect 23320 6535 23365 6655
rect 23485 6535 23530 6655
rect 23650 6535 23695 6655
rect 23815 6535 23870 6655
rect 23990 6535 24000 6655
rect 18500 6490 24000 6535
rect 18500 6370 18510 6490
rect 18630 6370 18675 6490
rect 18795 6370 18840 6490
rect 18960 6370 19005 6490
rect 19125 6370 19180 6490
rect 19300 6370 19345 6490
rect 19465 6370 19510 6490
rect 19630 6370 19675 6490
rect 19795 6370 19850 6490
rect 19970 6370 20015 6490
rect 20135 6370 20180 6490
rect 20300 6370 20345 6490
rect 20465 6370 20520 6490
rect 20640 6370 20685 6490
rect 20805 6370 20850 6490
rect 20970 6370 21015 6490
rect 21135 6370 21190 6490
rect 21310 6370 21355 6490
rect 21475 6370 21520 6490
rect 21640 6370 21685 6490
rect 21805 6370 21860 6490
rect 21980 6370 22025 6490
rect 22145 6370 22190 6490
rect 22310 6370 22355 6490
rect 22475 6370 22530 6490
rect 22650 6370 22695 6490
rect 22815 6370 22860 6490
rect 22980 6370 23025 6490
rect 23145 6370 23200 6490
rect 23320 6370 23365 6490
rect 23485 6370 23530 6490
rect 23650 6370 23695 6490
rect 23815 6370 23870 6490
rect 23990 6370 24000 6490
rect 18500 6315 24000 6370
rect 18500 6195 18510 6315
rect 18630 6195 18675 6315
rect 18795 6195 18840 6315
rect 18960 6195 19005 6315
rect 19125 6195 19180 6315
rect 19300 6195 19345 6315
rect 19465 6195 19510 6315
rect 19630 6195 19675 6315
rect 19795 6195 19850 6315
rect 19970 6195 20015 6315
rect 20135 6195 20180 6315
rect 20300 6195 20345 6315
rect 20465 6195 20520 6315
rect 20640 6195 20685 6315
rect 20805 6195 20850 6315
rect 20970 6195 21015 6315
rect 21135 6195 21190 6315
rect 21310 6195 21355 6315
rect 21475 6195 21520 6315
rect 21640 6195 21685 6315
rect 21805 6195 21860 6315
rect 21980 6195 22025 6315
rect 22145 6195 22190 6315
rect 22310 6195 22355 6315
rect 22475 6195 22530 6315
rect 22650 6195 22695 6315
rect 22815 6195 22860 6315
rect 22980 6195 23025 6315
rect 23145 6195 23200 6315
rect 23320 6195 23365 6315
rect 23485 6195 23530 6315
rect 23650 6195 23695 6315
rect 23815 6195 23870 6315
rect 23990 6195 24000 6315
rect 18500 6150 24000 6195
rect 18500 6030 18510 6150
rect 18630 6030 18675 6150
rect 18795 6030 18840 6150
rect 18960 6030 19005 6150
rect 19125 6030 19180 6150
rect 19300 6030 19345 6150
rect 19465 6030 19510 6150
rect 19630 6030 19675 6150
rect 19795 6030 19850 6150
rect 19970 6030 20015 6150
rect 20135 6030 20180 6150
rect 20300 6030 20345 6150
rect 20465 6030 20520 6150
rect 20640 6030 20685 6150
rect 20805 6030 20850 6150
rect 20970 6030 21015 6150
rect 21135 6030 21190 6150
rect 21310 6030 21355 6150
rect 21475 6030 21520 6150
rect 21640 6030 21685 6150
rect 21805 6030 21860 6150
rect 21980 6030 22025 6150
rect 22145 6030 22190 6150
rect 22310 6030 22355 6150
rect 22475 6030 22530 6150
rect 22650 6030 22695 6150
rect 22815 6030 22860 6150
rect 22980 6030 23025 6150
rect 23145 6030 23200 6150
rect 23320 6030 23365 6150
rect 23485 6030 23530 6150
rect 23650 6030 23695 6150
rect 23815 6030 23870 6150
rect 23990 6030 24000 6150
rect 18500 5985 24000 6030
rect 18500 5865 18510 5985
rect 18630 5865 18675 5985
rect 18795 5865 18840 5985
rect 18960 5865 19005 5985
rect 19125 5865 19180 5985
rect 19300 5865 19345 5985
rect 19465 5865 19510 5985
rect 19630 5865 19675 5985
rect 19795 5865 19850 5985
rect 19970 5865 20015 5985
rect 20135 5865 20180 5985
rect 20300 5865 20345 5985
rect 20465 5865 20520 5985
rect 20640 5865 20685 5985
rect 20805 5865 20850 5985
rect 20970 5865 21015 5985
rect 21135 5865 21190 5985
rect 21310 5865 21355 5985
rect 21475 5865 21520 5985
rect 21640 5865 21685 5985
rect 21805 5865 21860 5985
rect 21980 5865 22025 5985
rect 22145 5865 22190 5985
rect 22310 5865 22355 5985
rect 22475 5865 22530 5985
rect 22650 5865 22695 5985
rect 22815 5865 22860 5985
rect 22980 5865 23025 5985
rect 23145 5865 23200 5985
rect 23320 5865 23365 5985
rect 23485 5865 23530 5985
rect 23650 5865 23695 5985
rect 23815 5865 23870 5985
rect 23990 5865 24000 5985
rect 18500 5820 24000 5865
rect 18500 5700 18510 5820
rect 18630 5700 18675 5820
rect 18795 5700 18840 5820
rect 18960 5700 19005 5820
rect 19125 5700 19180 5820
rect 19300 5700 19345 5820
rect 19465 5700 19510 5820
rect 19630 5700 19675 5820
rect 19795 5700 19850 5820
rect 19970 5700 20015 5820
rect 20135 5700 20180 5820
rect 20300 5700 20345 5820
rect 20465 5700 20520 5820
rect 20640 5700 20685 5820
rect 20805 5700 20850 5820
rect 20970 5700 21015 5820
rect 21135 5700 21190 5820
rect 21310 5700 21355 5820
rect 21475 5700 21520 5820
rect 21640 5700 21685 5820
rect 21805 5700 21860 5820
rect 21980 5700 22025 5820
rect 22145 5700 22190 5820
rect 22310 5700 22355 5820
rect 22475 5700 22530 5820
rect 22650 5700 22695 5820
rect 22815 5700 22860 5820
rect 22980 5700 23025 5820
rect 23145 5700 23200 5820
rect 23320 5700 23365 5820
rect 23485 5700 23530 5820
rect 23650 5700 23695 5820
rect 23815 5700 23870 5820
rect 23990 5700 24000 5820
rect 18500 5645 24000 5700
rect 18500 5525 18510 5645
rect 18630 5525 18675 5645
rect 18795 5525 18840 5645
rect 18960 5525 19005 5645
rect 19125 5525 19180 5645
rect 19300 5525 19345 5645
rect 19465 5525 19510 5645
rect 19630 5525 19675 5645
rect 19795 5525 19850 5645
rect 19970 5525 20015 5645
rect 20135 5525 20180 5645
rect 20300 5525 20345 5645
rect 20465 5525 20520 5645
rect 20640 5525 20685 5645
rect 20805 5525 20850 5645
rect 20970 5525 21015 5645
rect 21135 5525 21190 5645
rect 21310 5525 21355 5645
rect 21475 5525 21520 5645
rect 21640 5525 21685 5645
rect 21805 5525 21860 5645
rect 21980 5525 22025 5645
rect 22145 5525 22190 5645
rect 22310 5525 22355 5645
rect 22475 5525 22530 5645
rect 22650 5525 22695 5645
rect 22815 5525 22860 5645
rect 22980 5525 23025 5645
rect 23145 5525 23200 5645
rect 23320 5525 23365 5645
rect 23485 5525 23530 5645
rect 23650 5525 23695 5645
rect 23815 5525 23870 5645
rect 23990 5525 24000 5645
rect 18500 5480 24000 5525
rect 18500 5360 18510 5480
rect 18630 5360 18675 5480
rect 18795 5360 18840 5480
rect 18960 5360 19005 5480
rect 19125 5360 19180 5480
rect 19300 5360 19345 5480
rect 19465 5360 19510 5480
rect 19630 5360 19675 5480
rect 19795 5360 19850 5480
rect 19970 5360 20015 5480
rect 20135 5360 20180 5480
rect 20300 5360 20345 5480
rect 20465 5360 20520 5480
rect 20640 5360 20685 5480
rect 20805 5360 20850 5480
rect 20970 5360 21015 5480
rect 21135 5360 21190 5480
rect 21310 5360 21355 5480
rect 21475 5360 21520 5480
rect 21640 5360 21685 5480
rect 21805 5360 21860 5480
rect 21980 5360 22025 5480
rect 22145 5360 22190 5480
rect 22310 5360 22355 5480
rect 22475 5360 22530 5480
rect 22650 5360 22695 5480
rect 22815 5360 22860 5480
rect 22980 5360 23025 5480
rect 23145 5360 23200 5480
rect 23320 5360 23365 5480
rect 23485 5360 23530 5480
rect 23650 5360 23695 5480
rect 23815 5360 23870 5480
rect 23990 5360 24000 5480
rect 18500 5315 24000 5360
rect 18500 5195 18510 5315
rect 18630 5195 18675 5315
rect 18795 5195 18840 5315
rect 18960 5195 19005 5315
rect 19125 5195 19180 5315
rect 19300 5195 19345 5315
rect 19465 5195 19510 5315
rect 19630 5195 19675 5315
rect 19795 5195 19850 5315
rect 19970 5195 20015 5315
rect 20135 5195 20180 5315
rect 20300 5195 20345 5315
rect 20465 5195 20520 5315
rect 20640 5195 20685 5315
rect 20805 5195 20850 5315
rect 20970 5195 21015 5315
rect 21135 5195 21190 5315
rect 21310 5195 21355 5315
rect 21475 5195 21520 5315
rect 21640 5195 21685 5315
rect 21805 5195 21860 5315
rect 21980 5195 22025 5315
rect 22145 5195 22190 5315
rect 22310 5195 22355 5315
rect 22475 5195 22530 5315
rect 22650 5195 22695 5315
rect 22815 5195 22860 5315
rect 22980 5195 23025 5315
rect 23145 5195 23200 5315
rect 23320 5195 23365 5315
rect 23485 5195 23530 5315
rect 23650 5195 23695 5315
rect 23815 5195 23870 5315
rect 23990 5195 24000 5315
rect 18500 5150 24000 5195
rect 18500 5030 18510 5150
rect 18630 5030 18675 5150
rect 18795 5030 18840 5150
rect 18960 5030 19005 5150
rect 19125 5030 19180 5150
rect 19300 5030 19345 5150
rect 19465 5030 19510 5150
rect 19630 5030 19675 5150
rect 19795 5030 19850 5150
rect 19970 5030 20015 5150
rect 20135 5030 20180 5150
rect 20300 5030 20345 5150
rect 20465 5030 20520 5150
rect 20640 5030 20685 5150
rect 20805 5030 20850 5150
rect 20970 5030 21015 5150
rect 21135 5030 21190 5150
rect 21310 5030 21355 5150
rect 21475 5030 21520 5150
rect 21640 5030 21685 5150
rect 21805 5030 21860 5150
rect 21980 5030 22025 5150
rect 22145 5030 22190 5150
rect 22310 5030 22355 5150
rect 22475 5030 22530 5150
rect 22650 5030 22695 5150
rect 22815 5030 22860 5150
rect 22980 5030 23025 5150
rect 23145 5030 23200 5150
rect 23320 5030 23365 5150
rect 23485 5030 23530 5150
rect 23650 5030 23695 5150
rect 23815 5030 23870 5150
rect 23990 5030 24000 5150
rect 18500 4975 24000 5030
rect 18500 4855 18510 4975
rect 18630 4855 18675 4975
rect 18795 4855 18840 4975
rect 18960 4855 19005 4975
rect 19125 4855 19180 4975
rect 19300 4855 19345 4975
rect 19465 4855 19510 4975
rect 19630 4855 19675 4975
rect 19795 4855 19850 4975
rect 19970 4855 20015 4975
rect 20135 4855 20180 4975
rect 20300 4855 20345 4975
rect 20465 4855 20520 4975
rect 20640 4855 20685 4975
rect 20805 4855 20850 4975
rect 20970 4855 21015 4975
rect 21135 4855 21190 4975
rect 21310 4855 21355 4975
rect 21475 4855 21520 4975
rect 21640 4855 21685 4975
rect 21805 4855 21860 4975
rect 21980 4855 22025 4975
rect 22145 4855 22190 4975
rect 22310 4855 22355 4975
rect 22475 4855 22530 4975
rect 22650 4855 22695 4975
rect 22815 4855 22860 4975
rect 22980 4855 23025 4975
rect 23145 4855 23200 4975
rect 23320 4855 23365 4975
rect 23485 4855 23530 4975
rect 23650 4855 23695 4975
rect 23815 4855 23870 4975
rect 23990 4855 24000 4975
rect 18500 4810 24000 4855
rect 18500 4690 18510 4810
rect 18630 4690 18675 4810
rect 18795 4690 18840 4810
rect 18960 4690 19005 4810
rect 19125 4690 19180 4810
rect 19300 4690 19345 4810
rect 19465 4690 19510 4810
rect 19630 4690 19675 4810
rect 19795 4690 19850 4810
rect 19970 4690 20015 4810
rect 20135 4690 20180 4810
rect 20300 4690 20345 4810
rect 20465 4690 20520 4810
rect 20640 4690 20685 4810
rect 20805 4690 20850 4810
rect 20970 4690 21015 4810
rect 21135 4690 21190 4810
rect 21310 4690 21355 4810
rect 21475 4690 21520 4810
rect 21640 4690 21685 4810
rect 21805 4690 21860 4810
rect 21980 4690 22025 4810
rect 22145 4690 22190 4810
rect 22310 4690 22355 4810
rect 22475 4690 22530 4810
rect 22650 4690 22695 4810
rect 22815 4690 22860 4810
rect 22980 4690 23025 4810
rect 23145 4690 23200 4810
rect 23320 4690 23365 4810
rect 23485 4690 23530 4810
rect 23650 4690 23695 4810
rect 23815 4690 23870 4810
rect 23990 4690 24000 4810
rect 18500 4645 24000 4690
rect 18500 4525 18510 4645
rect 18630 4525 18675 4645
rect 18795 4525 18840 4645
rect 18960 4525 19005 4645
rect 19125 4525 19180 4645
rect 19300 4525 19345 4645
rect 19465 4525 19510 4645
rect 19630 4525 19675 4645
rect 19795 4525 19850 4645
rect 19970 4525 20015 4645
rect 20135 4525 20180 4645
rect 20300 4525 20345 4645
rect 20465 4525 20520 4645
rect 20640 4525 20685 4645
rect 20805 4525 20850 4645
rect 20970 4525 21015 4645
rect 21135 4525 21190 4645
rect 21310 4525 21355 4645
rect 21475 4525 21520 4645
rect 21640 4525 21685 4645
rect 21805 4525 21860 4645
rect 21980 4525 22025 4645
rect 22145 4525 22190 4645
rect 22310 4525 22355 4645
rect 22475 4525 22530 4645
rect 22650 4525 22695 4645
rect 22815 4525 22860 4645
rect 22980 4525 23025 4645
rect 23145 4525 23200 4645
rect 23320 4525 23365 4645
rect 23485 4525 23530 4645
rect 23650 4525 23695 4645
rect 23815 4525 23870 4645
rect 23990 4525 24000 4645
rect 18500 4480 24000 4525
rect 18500 4360 18510 4480
rect 18630 4360 18675 4480
rect 18795 4360 18840 4480
rect 18960 4360 19005 4480
rect 19125 4360 19180 4480
rect 19300 4360 19345 4480
rect 19465 4360 19510 4480
rect 19630 4360 19675 4480
rect 19795 4360 19850 4480
rect 19970 4360 20015 4480
rect 20135 4360 20180 4480
rect 20300 4360 20345 4480
rect 20465 4360 20520 4480
rect 20640 4360 20685 4480
rect 20805 4360 20850 4480
rect 20970 4360 21015 4480
rect 21135 4360 21190 4480
rect 21310 4360 21355 4480
rect 21475 4360 21520 4480
rect 21640 4360 21685 4480
rect 21805 4360 21860 4480
rect 21980 4360 22025 4480
rect 22145 4360 22190 4480
rect 22310 4360 22355 4480
rect 22475 4360 22530 4480
rect 22650 4360 22695 4480
rect 22815 4360 22860 4480
rect 22980 4360 23025 4480
rect 23145 4360 23200 4480
rect 23320 4360 23365 4480
rect 23485 4360 23530 4480
rect 23650 4360 23695 4480
rect 23815 4360 23870 4480
rect 23990 4360 24000 4480
rect 18500 4305 24000 4360
rect 18500 4185 18510 4305
rect 18630 4185 18675 4305
rect 18795 4185 18840 4305
rect 18960 4185 19005 4305
rect 19125 4185 19180 4305
rect 19300 4185 19345 4305
rect 19465 4185 19510 4305
rect 19630 4185 19675 4305
rect 19795 4185 19850 4305
rect 19970 4185 20015 4305
rect 20135 4185 20180 4305
rect 20300 4185 20345 4305
rect 20465 4185 20520 4305
rect 20640 4185 20685 4305
rect 20805 4185 20850 4305
rect 20970 4185 21015 4305
rect 21135 4185 21190 4305
rect 21310 4185 21355 4305
rect 21475 4185 21520 4305
rect 21640 4185 21685 4305
rect 21805 4185 21860 4305
rect 21980 4185 22025 4305
rect 22145 4185 22190 4305
rect 22310 4185 22355 4305
rect 22475 4185 22530 4305
rect 22650 4185 22695 4305
rect 22815 4185 22860 4305
rect 22980 4185 23025 4305
rect 23145 4185 23200 4305
rect 23320 4185 23365 4305
rect 23485 4185 23530 4305
rect 23650 4185 23695 4305
rect 23815 4185 23870 4305
rect 23990 4185 24000 4305
rect 18500 4140 24000 4185
rect 18500 4020 18510 4140
rect 18630 4020 18675 4140
rect 18795 4020 18840 4140
rect 18960 4020 19005 4140
rect 19125 4020 19180 4140
rect 19300 4020 19345 4140
rect 19465 4020 19510 4140
rect 19630 4020 19675 4140
rect 19795 4020 19850 4140
rect 19970 4020 20015 4140
rect 20135 4020 20180 4140
rect 20300 4020 20345 4140
rect 20465 4020 20520 4140
rect 20640 4020 20685 4140
rect 20805 4020 20850 4140
rect 20970 4020 21015 4140
rect 21135 4020 21190 4140
rect 21310 4020 21355 4140
rect 21475 4020 21520 4140
rect 21640 4020 21685 4140
rect 21805 4020 21860 4140
rect 21980 4020 22025 4140
rect 22145 4020 22190 4140
rect 22310 4020 22355 4140
rect 22475 4020 22530 4140
rect 22650 4020 22695 4140
rect 22815 4020 22860 4140
rect 22980 4020 23025 4140
rect 23145 4020 23200 4140
rect 23320 4020 23365 4140
rect 23485 4020 23530 4140
rect 23650 4020 23695 4140
rect 23815 4020 23870 4140
rect 23990 4020 24000 4140
rect 18500 3975 24000 4020
rect 18500 3855 18510 3975
rect 18630 3855 18675 3975
rect 18795 3855 18840 3975
rect 18960 3855 19005 3975
rect 19125 3855 19180 3975
rect 19300 3855 19345 3975
rect 19465 3855 19510 3975
rect 19630 3855 19675 3975
rect 19795 3855 19850 3975
rect 19970 3855 20015 3975
rect 20135 3855 20180 3975
rect 20300 3855 20345 3975
rect 20465 3855 20520 3975
rect 20640 3855 20685 3975
rect 20805 3855 20850 3975
rect 20970 3855 21015 3975
rect 21135 3855 21190 3975
rect 21310 3855 21355 3975
rect 21475 3855 21520 3975
rect 21640 3855 21685 3975
rect 21805 3855 21860 3975
rect 21980 3855 22025 3975
rect 22145 3855 22190 3975
rect 22310 3855 22355 3975
rect 22475 3855 22530 3975
rect 22650 3855 22695 3975
rect 22815 3855 22860 3975
rect 22980 3855 23025 3975
rect 23145 3855 23200 3975
rect 23320 3855 23365 3975
rect 23485 3855 23530 3975
rect 23650 3855 23695 3975
rect 23815 3855 23870 3975
rect 23990 3855 24000 3975
rect 18500 3810 24000 3855
rect 18500 3690 18510 3810
rect 18630 3690 18675 3810
rect 18795 3690 18840 3810
rect 18960 3690 19005 3810
rect 19125 3690 19180 3810
rect 19300 3690 19345 3810
rect 19465 3690 19510 3810
rect 19630 3690 19675 3810
rect 19795 3690 19850 3810
rect 19970 3690 20015 3810
rect 20135 3690 20180 3810
rect 20300 3690 20345 3810
rect 20465 3690 20520 3810
rect 20640 3690 20685 3810
rect 20805 3690 20850 3810
rect 20970 3690 21015 3810
rect 21135 3690 21190 3810
rect 21310 3690 21355 3810
rect 21475 3690 21520 3810
rect 21640 3690 21685 3810
rect 21805 3690 21860 3810
rect 21980 3690 22025 3810
rect 22145 3690 22190 3810
rect 22310 3690 22355 3810
rect 22475 3690 22530 3810
rect 22650 3690 22695 3810
rect 22815 3690 22860 3810
rect 22980 3690 23025 3810
rect 23145 3690 23200 3810
rect 23320 3690 23365 3810
rect 23485 3690 23530 3810
rect 23650 3690 23695 3810
rect 23815 3690 23870 3810
rect 23990 3690 24000 3810
rect 18500 3635 24000 3690
rect 18500 3515 18510 3635
rect 18630 3515 18675 3635
rect 18795 3515 18840 3635
rect 18960 3515 19005 3635
rect 19125 3515 19180 3635
rect 19300 3515 19345 3635
rect 19465 3515 19510 3635
rect 19630 3515 19675 3635
rect 19795 3515 19850 3635
rect 19970 3515 20015 3635
rect 20135 3515 20180 3635
rect 20300 3515 20345 3635
rect 20465 3515 20520 3635
rect 20640 3515 20685 3635
rect 20805 3515 20850 3635
rect 20970 3515 21015 3635
rect 21135 3515 21190 3635
rect 21310 3515 21355 3635
rect 21475 3515 21520 3635
rect 21640 3515 21685 3635
rect 21805 3515 21860 3635
rect 21980 3515 22025 3635
rect 22145 3515 22190 3635
rect 22310 3515 22355 3635
rect 22475 3515 22530 3635
rect 22650 3515 22695 3635
rect 22815 3515 22860 3635
rect 22980 3515 23025 3635
rect 23145 3515 23200 3635
rect 23320 3515 23365 3635
rect 23485 3515 23530 3635
rect 23650 3515 23695 3635
rect 23815 3515 23870 3635
rect 23990 3515 24000 3635
rect 18500 3470 24000 3515
rect 18500 3350 18510 3470
rect 18630 3350 18675 3470
rect 18795 3350 18840 3470
rect 18960 3350 19005 3470
rect 19125 3350 19180 3470
rect 19300 3350 19345 3470
rect 19465 3350 19510 3470
rect 19630 3350 19675 3470
rect 19795 3350 19850 3470
rect 19970 3350 20015 3470
rect 20135 3350 20180 3470
rect 20300 3350 20345 3470
rect 20465 3350 20520 3470
rect 20640 3350 20685 3470
rect 20805 3350 20850 3470
rect 20970 3350 21015 3470
rect 21135 3350 21190 3470
rect 21310 3350 21355 3470
rect 21475 3350 21520 3470
rect 21640 3350 21685 3470
rect 21805 3350 21860 3470
rect 21980 3350 22025 3470
rect 22145 3350 22190 3470
rect 22310 3350 22355 3470
rect 22475 3350 22530 3470
rect 22650 3350 22695 3470
rect 22815 3350 22860 3470
rect 22980 3350 23025 3470
rect 23145 3350 23200 3470
rect 23320 3350 23365 3470
rect 23485 3350 23530 3470
rect 23650 3350 23695 3470
rect 23815 3350 23870 3470
rect 23990 3350 24000 3470
rect 18500 3305 24000 3350
rect 18500 3185 18510 3305
rect 18630 3185 18675 3305
rect 18795 3185 18840 3305
rect 18960 3185 19005 3305
rect 19125 3185 19180 3305
rect 19300 3185 19345 3305
rect 19465 3185 19510 3305
rect 19630 3185 19675 3305
rect 19795 3185 19850 3305
rect 19970 3185 20015 3305
rect 20135 3185 20180 3305
rect 20300 3185 20345 3305
rect 20465 3185 20520 3305
rect 20640 3185 20685 3305
rect 20805 3185 20850 3305
rect 20970 3185 21015 3305
rect 21135 3185 21190 3305
rect 21310 3185 21355 3305
rect 21475 3185 21520 3305
rect 21640 3185 21685 3305
rect 21805 3185 21860 3305
rect 21980 3185 22025 3305
rect 22145 3185 22190 3305
rect 22310 3185 22355 3305
rect 22475 3185 22530 3305
rect 22650 3185 22695 3305
rect 22815 3185 22860 3305
rect 22980 3185 23025 3305
rect 23145 3185 23200 3305
rect 23320 3185 23365 3305
rect 23485 3185 23530 3305
rect 23650 3185 23695 3305
rect 23815 3185 23870 3305
rect 23990 3185 24000 3305
rect 18500 3140 24000 3185
rect 18500 3020 18510 3140
rect 18630 3020 18675 3140
rect 18795 3020 18840 3140
rect 18960 3020 19005 3140
rect 19125 3020 19180 3140
rect 19300 3020 19345 3140
rect 19465 3020 19510 3140
rect 19630 3020 19675 3140
rect 19795 3020 19850 3140
rect 19970 3020 20015 3140
rect 20135 3020 20180 3140
rect 20300 3020 20345 3140
rect 20465 3020 20520 3140
rect 20640 3020 20685 3140
rect 20805 3020 20850 3140
rect 20970 3020 21015 3140
rect 21135 3020 21190 3140
rect 21310 3020 21355 3140
rect 21475 3020 21520 3140
rect 21640 3020 21685 3140
rect 21805 3020 21860 3140
rect 21980 3020 22025 3140
rect 22145 3020 22190 3140
rect 22310 3020 22355 3140
rect 22475 3020 22530 3140
rect 22650 3020 22695 3140
rect 22815 3020 22860 3140
rect 22980 3020 23025 3140
rect 23145 3020 23200 3140
rect 23320 3020 23365 3140
rect 23485 3020 23530 3140
rect 23650 3020 23695 3140
rect 23815 3020 23870 3140
rect 23990 3020 24000 3140
rect 18500 2965 24000 3020
rect 18500 2845 18510 2965
rect 18630 2845 18675 2965
rect 18795 2845 18840 2965
rect 18960 2845 19005 2965
rect 19125 2845 19180 2965
rect 19300 2845 19345 2965
rect 19465 2845 19510 2965
rect 19630 2845 19675 2965
rect 19795 2845 19850 2965
rect 19970 2845 20015 2965
rect 20135 2845 20180 2965
rect 20300 2845 20345 2965
rect 20465 2845 20520 2965
rect 20640 2845 20685 2965
rect 20805 2845 20850 2965
rect 20970 2845 21015 2965
rect 21135 2845 21190 2965
rect 21310 2845 21355 2965
rect 21475 2845 21520 2965
rect 21640 2845 21685 2965
rect 21805 2845 21860 2965
rect 21980 2845 22025 2965
rect 22145 2845 22190 2965
rect 22310 2845 22355 2965
rect 22475 2845 22530 2965
rect 22650 2845 22695 2965
rect 22815 2845 22860 2965
rect 22980 2845 23025 2965
rect 23145 2845 23200 2965
rect 23320 2845 23365 2965
rect 23485 2845 23530 2965
rect 23650 2845 23695 2965
rect 23815 2845 23870 2965
rect 23990 2845 24000 2965
rect 18500 2800 24000 2845
rect 18500 2680 18510 2800
rect 18630 2680 18675 2800
rect 18795 2680 18840 2800
rect 18960 2680 19005 2800
rect 19125 2680 19180 2800
rect 19300 2680 19345 2800
rect 19465 2680 19510 2800
rect 19630 2680 19675 2800
rect 19795 2680 19850 2800
rect 19970 2680 20015 2800
rect 20135 2680 20180 2800
rect 20300 2680 20345 2800
rect 20465 2680 20520 2800
rect 20640 2680 20685 2800
rect 20805 2680 20850 2800
rect 20970 2680 21015 2800
rect 21135 2680 21190 2800
rect 21310 2680 21355 2800
rect 21475 2680 21520 2800
rect 21640 2680 21685 2800
rect 21805 2680 21860 2800
rect 21980 2680 22025 2800
rect 22145 2680 22190 2800
rect 22310 2680 22355 2800
rect 22475 2680 22530 2800
rect 22650 2680 22695 2800
rect 22815 2680 22860 2800
rect 22980 2680 23025 2800
rect 23145 2680 23200 2800
rect 23320 2680 23365 2800
rect 23485 2680 23530 2800
rect 23650 2680 23695 2800
rect 23815 2680 23870 2800
rect 23990 2680 24000 2800
rect 18500 2635 24000 2680
rect 18500 2515 18510 2635
rect 18630 2515 18675 2635
rect 18795 2515 18840 2635
rect 18960 2515 19005 2635
rect 19125 2515 19180 2635
rect 19300 2515 19345 2635
rect 19465 2515 19510 2635
rect 19630 2515 19675 2635
rect 19795 2515 19850 2635
rect 19970 2515 20015 2635
rect 20135 2515 20180 2635
rect 20300 2515 20345 2635
rect 20465 2515 20520 2635
rect 20640 2515 20685 2635
rect 20805 2515 20850 2635
rect 20970 2515 21015 2635
rect 21135 2515 21190 2635
rect 21310 2515 21355 2635
rect 21475 2515 21520 2635
rect 21640 2515 21685 2635
rect 21805 2515 21860 2635
rect 21980 2515 22025 2635
rect 22145 2515 22190 2635
rect 22310 2515 22355 2635
rect 22475 2515 22530 2635
rect 22650 2515 22695 2635
rect 22815 2515 22860 2635
rect 22980 2515 23025 2635
rect 23145 2515 23200 2635
rect 23320 2515 23365 2635
rect 23485 2515 23530 2635
rect 23650 2515 23695 2635
rect 23815 2515 23870 2635
rect 23990 2515 24000 2635
rect 18500 2470 24000 2515
rect 18500 2350 18510 2470
rect 18630 2350 18675 2470
rect 18795 2350 18840 2470
rect 18960 2350 19005 2470
rect 19125 2350 19180 2470
rect 19300 2350 19345 2470
rect 19465 2350 19510 2470
rect 19630 2350 19675 2470
rect 19795 2350 19850 2470
rect 19970 2350 20015 2470
rect 20135 2350 20180 2470
rect 20300 2350 20345 2470
rect 20465 2350 20520 2470
rect 20640 2350 20685 2470
rect 20805 2350 20850 2470
rect 20970 2350 21015 2470
rect 21135 2350 21190 2470
rect 21310 2350 21355 2470
rect 21475 2350 21520 2470
rect 21640 2350 21685 2470
rect 21805 2350 21860 2470
rect 21980 2350 22025 2470
rect 22145 2350 22190 2470
rect 22310 2350 22355 2470
rect 22475 2350 22530 2470
rect 22650 2350 22695 2470
rect 22815 2350 22860 2470
rect 22980 2350 23025 2470
rect 23145 2350 23200 2470
rect 23320 2350 23365 2470
rect 23485 2350 23530 2470
rect 23650 2350 23695 2470
rect 23815 2350 23870 2470
rect 23990 2350 24000 2470
rect 18500 2295 24000 2350
rect 18500 2175 18510 2295
rect 18630 2175 18675 2295
rect 18795 2175 18840 2295
rect 18960 2175 19005 2295
rect 19125 2175 19180 2295
rect 19300 2175 19345 2295
rect 19465 2175 19510 2295
rect 19630 2175 19675 2295
rect 19795 2175 19850 2295
rect 19970 2175 20015 2295
rect 20135 2175 20180 2295
rect 20300 2175 20345 2295
rect 20465 2175 20520 2295
rect 20640 2175 20685 2295
rect 20805 2175 20850 2295
rect 20970 2175 21015 2295
rect 21135 2175 21190 2295
rect 21310 2175 21355 2295
rect 21475 2175 21520 2295
rect 21640 2175 21685 2295
rect 21805 2175 21860 2295
rect 21980 2175 22025 2295
rect 22145 2175 22190 2295
rect 22310 2175 22355 2295
rect 22475 2175 22530 2295
rect 22650 2175 22695 2295
rect 22815 2175 22860 2295
rect 22980 2175 23025 2295
rect 23145 2175 23200 2295
rect 23320 2175 23365 2295
rect 23485 2175 23530 2295
rect 23650 2175 23695 2295
rect 23815 2175 23870 2295
rect 23990 2175 24000 2295
rect 18500 2130 24000 2175
rect 18500 2010 18510 2130
rect 18630 2010 18675 2130
rect 18795 2010 18840 2130
rect 18960 2010 19005 2130
rect 19125 2010 19180 2130
rect 19300 2010 19345 2130
rect 19465 2010 19510 2130
rect 19630 2010 19675 2130
rect 19795 2010 19850 2130
rect 19970 2010 20015 2130
rect 20135 2010 20180 2130
rect 20300 2010 20345 2130
rect 20465 2010 20520 2130
rect 20640 2010 20685 2130
rect 20805 2010 20850 2130
rect 20970 2010 21015 2130
rect 21135 2010 21190 2130
rect 21310 2010 21355 2130
rect 21475 2010 21520 2130
rect 21640 2010 21685 2130
rect 21805 2010 21860 2130
rect 21980 2010 22025 2130
rect 22145 2010 22190 2130
rect 22310 2010 22355 2130
rect 22475 2010 22530 2130
rect 22650 2010 22695 2130
rect 22815 2010 22860 2130
rect 22980 2010 23025 2130
rect 23145 2010 23200 2130
rect 23320 2010 23365 2130
rect 23485 2010 23530 2130
rect 23650 2010 23695 2130
rect 23815 2010 23870 2130
rect 23990 2010 24000 2130
rect 18500 1965 24000 2010
rect 18500 1845 18510 1965
rect 18630 1845 18675 1965
rect 18795 1845 18840 1965
rect 18960 1845 19005 1965
rect 19125 1845 19180 1965
rect 19300 1845 19345 1965
rect 19465 1845 19510 1965
rect 19630 1845 19675 1965
rect 19795 1845 19850 1965
rect 19970 1845 20015 1965
rect 20135 1845 20180 1965
rect 20300 1845 20345 1965
rect 20465 1845 20520 1965
rect 20640 1845 20685 1965
rect 20805 1845 20850 1965
rect 20970 1845 21015 1965
rect 21135 1845 21190 1965
rect 21310 1845 21355 1965
rect 21475 1845 21520 1965
rect 21640 1845 21685 1965
rect 21805 1845 21860 1965
rect 21980 1845 22025 1965
rect 22145 1845 22190 1965
rect 22310 1845 22355 1965
rect 22475 1845 22530 1965
rect 22650 1845 22695 1965
rect 22815 1845 22860 1965
rect 22980 1845 23025 1965
rect 23145 1845 23200 1965
rect 23320 1845 23365 1965
rect 23485 1845 23530 1965
rect 23650 1845 23695 1965
rect 23815 1845 23870 1965
rect 23990 1845 24000 1965
rect 18500 1800 24000 1845
rect 18500 1680 18510 1800
rect 18630 1680 18675 1800
rect 18795 1680 18840 1800
rect 18960 1680 19005 1800
rect 19125 1680 19180 1800
rect 19300 1680 19345 1800
rect 19465 1680 19510 1800
rect 19630 1680 19675 1800
rect 19795 1680 19850 1800
rect 19970 1680 20015 1800
rect 20135 1680 20180 1800
rect 20300 1680 20345 1800
rect 20465 1680 20520 1800
rect 20640 1680 20685 1800
rect 20805 1680 20850 1800
rect 20970 1680 21015 1800
rect 21135 1680 21190 1800
rect 21310 1680 21355 1800
rect 21475 1680 21520 1800
rect 21640 1680 21685 1800
rect 21805 1680 21860 1800
rect 21980 1680 22025 1800
rect 22145 1680 22190 1800
rect 22310 1680 22355 1800
rect 22475 1680 22530 1800
rect 22650 1680 22695 1800
rect 22815 1680 22860 1800
rect 22980 1680 23025 1800
rect 23145 1680 23200 1800
rect 23320 1680 23365 1800
rect 23485 1680 23530 1800
rect 23650 1680 23695 1800
rect 23815 1680 23870 1800
rect 23990 1680 24000 1800
rect 18500 1670 24000 1680
rect 24190 7160 29690 7170
rect 24190 7040 24200 7160
rect 24320 7040 24365 7160
rect 24485 7040 24530 7160
rect 24650 7040 24695 7160
rect 24815 7040 24870 7160
rect 24990 7040 25035 7160
rect 25155 7040 25200 7160
rect 25320 7040 25365 7160
rect 25485 7040 25540 7160
rect 25660 7040 25705 7160
rect 25825 7040 25870 7160
rect 25990 7040 26035 7160
rect 26155 7040 26210 7160
rect 26330 7040 26375 7160
rect 26495 7040 26540 7160
rect 26660 7040 26705 7160
rect 26825 7040 26880 7160
rect 27000 7040 27045 7160
rect 27165 7040 27210 7160
rect 27330 7040 27375 7160
rect 27495 7040 27550 7160
rect 27670 7040 27715 7160
rect 27835 7040 27880 7160
rect 28000 7040 28045 7160
rect 28165 7040 28220 7160
rect 28340 7040 28385 7160
rect 28505 7040 28550 7160
rect 28670 7040 28715 7160
rect 28835 7040 28890 7160
rect 29010 7040 29055 7160
rect 29175 7040 29220 7160
rect 29340 7040 29385 7160
rect 29505 7040 29560 7160
rect 29680 7040 29690 7160
rect 24190 6985 29690 7040
rect 24190 6865 24200 6985
rect 24320 6865 24365 6985
rect 24485 6865 24530 6985
rect 24650 6865 24695 6985
rect 24815 6865 24870 6985
rect 24990 6865 25035 6985
rect 25155 6865 25200 6985
rect 25320 6865 25365 6985
rect 25485 6865 25540 6985
rect 25660 6865 25705 6985
rect 25825 6865 25870 6985
rect 25990 6865 26035 6985
rect 26155 6865 26210 6985
rect 26330 6865 26375 6985
rect 26495 6865 26540 6985
rect 26660 6865 26705 6985
rect 26825 6865 26880 6985
rect 27000 6865 27045 6985
rect 27165 6865 27210 6985
rect 27330 6865 27375 6985
rect 27495 6865 27550 6985
rect 27670 6865 27715 6985
rect 27835 6865 27880 6985
rect 28000 6865 28045 6985
rect 28165 6865 28220 6985
rect 28340 6865 28385 6985
rect 28505 6865 28550 6985
rect 28670 6865 28715 6985
rect 28835 6865 28890 6985
rect 29010 6865 29055 6985
rect 29175 6865 29220 6985
rect 29340 6865 29385 6985
rect 29505 6865 29560 6985
rect 29680 6865 29690 6985
rect 24190 6820 29690 6865
rect 24190 6700 24200 6820
rect 24320 6700 24365 6820
rect 24485 6700 24530 6820
rect 24650 6700 24695 6820
rect 24815 6700 24870 6820
rect 24990 6700 25035 6820
rect 25155 6700 25200 6820
rect 25320 6700 25365 6820
rect 25485 6700 25540 6820
rect 25660 6700 25705 6820
rect 25825 6700 25870 6820
rect 25990 6700 26035 6820
rect 26155 6700 26210 6820
rect 26330 6700 26375 6820
rect 26495 6700 26540 6820
rect 26660 6700 26705 6820
rect 26825 6700 26880 6820
rect 27000 6700 27045 6820
rect 27165 6700 27210 6820
rect 27330 6700 27375 6820
rect 27495 6700 27550 6820
rect 27670 6700 27715 6820
rect 27835 6700 27880 6820
rect 28000 6700 28045 6820
rect 28165 6700 28220 6820
rect 28340 6700 28385 6820
rect 28505 6700 28550 6820
rect 28670 6700 28715 6820
rect 28835 6700 28890 6820
rect 29010 6700 29055 6820
rect 29175 6700 29220 6820
rect 29340 6700 29385 6820
rect 29505 6700 29560 6820
rect 29680 6700 29690 6820
rect 24190 6655 29690 6700
rect 24190 6535 24200 6655
rect 24320 6535 24365 6655
rect 24485 6535 24530 6655
rect 24650 6535 24695 6655
rect 24815 6535 24870 6655
rect 24990 6535 25035 6655
rect 25155 6535 25200 6655
rect 25320 6535 25365 6655
rect 25485 6535 25540 6655
rect 25660 6535 25705 6655
rect 25825 6535 25870 6655
rect 25990 6535 26035 6655
rect 26155 6535 26210 6655
rect 26330 6535 26375 6655
rect 26495 6535 26540 6655
rect 26660 6535 26705 6655
rect 26825 6535 26880 6655
rect 27000 6535 27045 6655
rect 27165 6535 27210 6655
rect 27330 6535 27375 6655
rect 27495 6535 27550 6655
rect 27670 6535 27715 6655
rect 27835 6535 27880 6655
rect 28000 6535 28045 6655
rect 28165 6535 28220 6655
rect 28340 6535 28385 6655
rect 28505 6535 28550 6655
rect 28670 6535 28715 6655
rect 28835 6535 28890 6655
rect 29010 6535 29055 6655
rect 29175 6535 29220 6655
rect 29340 6535 29385 6655
rect 29505 6535 29560 6655
rect 29680 6535 29690 6655
rect 24190 6490 29690 6535
rect 24190 6370 24200 6490
rect 24320 6370 24365 6490
rect 24485 6370 24530 6490
rect 24650 6370 24695 6490
rect 24815 6370 24870 6490
rect 24990 6370 25035 6490
rect 25155 6370 25200 6490
rect 25320 6370 25365 6490
rect 25485 6370 25540 6490
rect 25660 6370 25705 6490
rect 25825 6370 25870 6490
rect 25990 6370 26035 6490
rect 26155 6370 26210 6490
rect 26330 6370 26375 6490
rect 26495 6370 26540 6490
rect 26660 6370 26705 6490
rect 26825 6370 26880 6490
rect 27000 6370 27045 6490
rect 27165 6370 27210 6490
rect 27330 6370 27375 6490
rect 27495 6370 27550 6490
rect 27670 6370 27715 6490
rect 27835 6370 27880 6490
rect 28000 6370 28045 6490
rect 28165 6370 28220 6490
rect 28340 6370 28385 6490
rect 28505 6370 28550 6490
rect 28670 6370 28715 6490
rect 28835 6370 28890 6490
rect 29010 6370 29055 6490
rect 29175 6370 29220 6490
rect 29340 6370 29385 6490
rect 29505 6370 29560 6490
rect 29680 6370 29690 6490
rect 24190 6315 29690 6370
rect 24190 6195 24200 6315
rect 24320 6195 24365 6315
rect 24485 6195 24530 6315
rect 24650 6195 24695 6315
rect 24815 6195 24870 6315
rect 24990 6195 25035 6315
rect 25155 6195 25200 6315
rect 25320 6195 25365 6315
rect 25485 6195 25540 6315
rect 25660 6195 25705 6315
rect 25825 6195 25870 6315
rect 25990 6195 26035 6315
rect 26155 6195 26210 6315
rect 26330 6195 26375 6315
rect 26495 6195 26540 6315
rect 26660 6195 26705 6315
rect 26825 6195 26880 6315
rect 27000 6195 27045 6315
rect 27165 6195 27210 6315
rect 27330 6195 27375 6315
rect 27495 6195 27550 6315
rect 27670 6195 27715 6315
rect 27835 6195 27880 6315
rect 28000 6195 28045 6315
rect 28165 6195 28220 6315
rect 28340 6195 28385 6315
rect 28505 6195 28550 6315
rect 28670 6195 28715 6315
rect 28835 6195 28890 6315
rect 29010 6195 29055 6315
rect 29175 6195 29220 6315
rect 29340 6195 29385 6315
rect 29505 6195 29560 6315
rect 29680 6195 29690 6315
rect 24190 6150 29690 6195
rect 24190 6030 24200 6150
rect 24320 6030 24365 6150
rect 24485 6030 24530 6150
rect 24650 6030 24695 6150
rect 24815 6030 24870 6150
rect 24990 6030 25035 6150
rect 25155 6030 25200 6150
rect 25320 6030 25365 6150
rect 25485 6030 25540 6150
rect 25660 6030 25705 6150
rect 25825 6030 25870 6150
rect 25990 6030 26035 6150
rect 26155 6030 26210 6150
rect 26330 6030 26375 6150
rect 26495 6030 26540 6150
rect 26660 6030 26705 6150
rect 26825 6030 26880 6150
rect 27000 6030 27045 6150
rect 27165 6030 27210 6150
rect 27330 6030 27375 6150
rect 27495 6030 27550 6150
rect 27670 6030 27715 6150
rect 27835 6030 27880 6150
rect 28000 6030 28045 6150
rect 28165 6030 28220 6150
rect 28340 6030 28385 6150
rect 28505 6030 28550 6150
rect 28670 6030 28715 6150
rect 28835 6030 28890 6150
rect 29010 6030 29055 6150
rect 29175 6030 29220 6150
rect 29340 6030 29385 6150
rect 29505 6030 29560 6150
rect 29680 6030 29690 6150
rect 24190 5985 29690 6030
rect 24190 5865 24200 5985
rect 24320 5865 24365 5985
rect 24485 5865 24530 5985
rect 24650 5865 24695 5985
rect 24815 5865 24870 5985
rect 24990 5865 25035 5985
rect 25155 5865 25200 5985
rect 25320 5865 25365 5985
rect 25485 5865 25540 5985
rect 25660 5865 25705 5985
rect 25825 5865 25870 5985
rect 25990 5865 26035 5985
rect 26155 5865 26210 5985
rect 26330 5865 26375 5985
rect 26495 5865 26540 5985
rect 26660 5865 26705 5985
rect 26825 5865 26880 5985
rect 27000 5865 27045 5985
rect 27165 5865 27210 5985
rect 27330 5865 27375 5985
rect 27495 5865 27550 5985
rect 27670 5865 27715 5985
rect 27835 5865 27880 5985
rect 28000 5865 28045 5985
rect 28165 5865 28220 5985
rect 28340 5865 28385 5985
rect 28505 5865 28550 5985
rect 28670 5865 28715 5985
rect 28835 5865 28890 5985
rect 29010 5865 29055 5985
rect 29175 5865 29220 5985
rect 29340 5865 29385 5985
rect 29505 5865 29560 5985
rect 29680 5865 29690 5985
rect 24190 5820 29690 5865
rect 24190 5700 24200 5820
rect 24320 5700 24365 5820
rect 24485 5700 24530 5820
rect 24650 5700 24695 5820
rect 24815 5700 24870 5820
rect 24990 5700 25035 5820
rect 25155 5700 25200 5820
rect 25320 5700 25365 5820
rect 25485 5700 25540 5820
rect 25660 5700 25705 5820
rect 25825 5700 25870 5820
rect 25990 5700 26035 5820
rect 26155 5700 26210 5820
rect 26330 5700 26375 5820
rect 26495 5700 26540 5820
rect 26660 5700 26705 5820
rect 26825 5700 26880 5820
rect 27000 5700 27045 5820
rect 27165 5700 27210 5820
rect 27330 5700 27375 5820
rect 27495 5700 27550 5820
rect 27670 5700 27715 5820
rect 27835 5700 27880 5820
rect 28000 5700 28045 5820
rect 28165 5700 28220 5820
rect 28340 5700 28385 5820
rect 28505 5700 28550 5820
rect 28670 5700 28715 5820
rect 28835 5700 28890 5820
rect 29010 5700 29055 5820
rect 29175 5700 29220 5820
rect 29340 5700 29385 5820
rect 29505 5700 29560 5820
rect 29680 5700 29690 5820
rect 24190 5645 29690 5700
rect 24190 5525 24200 5645
rect 24320 5525 24365 5645
rect 24485 5525 24530 5645
rect 24650 5525 24695 5645
rect 24815 5525 24870 5645
rect 24990 5525 25035 5645
rect 25155 5525 25200 5645
rect 25320 5525 25365 5645
rect 25485 5525 25540 5645
rect 25660 5525 25705 5645
rect 25825 5525 25870 5645
rect 25990 5525 26035 5645
rect 26155 5525 26210 5645
rect 26330 5525 26375 5645
rect 26495 5525 26540 5645
rect 26660 5525 26705 5645
rect 26825 5525 26880 5645
rect 27000 5525 27045 5645
rect 27165 5525 27210 5645
rect 27330 5525 27375 5645
rect 27495 5525 27550 5645
rect 27670 5525 27715 5645
rect 27835 5525 27880 5645
rect 28000 5525 28045 5645
rect 28165 5525 28220 5645
rect 28340 5525 28385 5645
rect 28505 5525 28550 5645
rect 28670 5525 28715 5645
rect 28835 5525 28890 5645
rect 29010 5525 29055 5645
rect 29175 5525 29220 5645
rect 29340 5525 29385 5645
rect 29505 5525 29560 5645
rect 29680 5525 29690 5645
rect 24190 5480 29690 5525
rect 24190 5360 24200 5480
rect 24320 5360 24365 5480
rect 24485 5360 24530 5480
rect 24650 5360 24695 5480
rect 24815 5360 24870 5480
rect 24990 5360 25035 5480
rect 25155 5360 25200 5480
rect 25320 5360 25365 5480
rect 25485 5360 25540 5480
rect 25660 5360 25705 5480
rect 25825 5360 25870 5480
rect 25990 5360 26035 5480
rect 26155 5360 26210 5480
rect 26330 5360 26375 5480
rect 26495 5360 26540 5480
rect 26660 5360 26705 5480
rect 26825 5360 26880 5480
rect 27000 5360 27045 5480
rect 27165 5360 27210 5480
rect 27330 5360 27375 5480
rect 27495 5360 27550 5480
rect 27670 5360 27715 5480
rect 27835 5360 27880 5480
rect 28000 5360 28045 5480
rect 28165 5360 28220 5480
rect 28340 5360 28385 5480
rect 28505 5360 28550 5480
rect 28670 5360 28715 5480
rect 28835 5360 28890 5480
rect 29010 5360 29055 5480
rect 29175 5360 29220 5480
rect 29340 5360 29385 5480
rect 29505 5360 29560 5480
rect 29680 5360 29690 5480
rect 24190 5315 29690 5360
rect 24190 5195 24200 5315
rect 24320 5195 24365 5315
rect 24485 5195 24530 5315
rect 24650 5195 24695 5315
rect 24815 5195 24870 5315
rect 24990 5195 25035 5315
rect 25155 5195 25200 5315
rect 25320 5195 25365 5315
rect 25485 5195 25540 5315
rect 25660 5195 25705 5315
rect 25825 5195 25870 5315
rect 25990 5195 26035 5315
rect 26155 5195 26210 5315
rect 26330 5195 26375 5315
rect 26495 5195 26540 5315
rect 26660 5195 26705 5315
rect 26825 5195 26880 5315
rect 27000 5195 27045 5315
rect 27165 5195 27210 5315
rect 27330 5195 27375 5315
rect 27495 5195 27550 5315
rect 27670 5195 27715 5315
rect 27835 5195 27880 5315
rect 28000 5195 28045 5315
rect 28165 5195 28220 5315
rect 28340 5195 28385 5315
rect 28505 5195 28550 5315
rect 28670 5195 28715 5315
rect 28835 5195 28890 5315
rect 29010 5195 29055 5315
rect 29175 5195 29220 5315
rect 29340 5195 29385 5315
rect 29505 5195 29560 5315
rect 29680 5195 29690 5315
rect 24190 5150 29690 5195
rect 24190 5030 24200 5150
rect 24320 5030 24365 5150
rect 24485 5030 24530 5150
rect 24650 5030 24695 5150
rect 24815 5030 24870 5150
rect 24990 5030 25035 5150
rect 25155 5030 25200 5150
rect 25320 5030 25365 5150
rect 25485 5030 25540 5150
rect 25660 5030 25705 5150
rect 25825 5030 25870 5150
rect 25990 5030 26035 5150
rect 26155 5030 26210 5150
rect 26330 5030 26375 5150
rect 26495 5030 26540 5150
rect 26660 5030 26705 5150
rect 26825 5030 26880 5150
rect 27000 5030 27045 5150
rect 27165 5030 27210 5150
rect 27330 5030 27375 5150
rect 27495 5030 27550 5150
rect 27670 5030 27715 5150
rect 27835 5030 27880 5150
rect 28000 5030 28045 5150
rect 28165 5030 28220 5150
rect 28340 5030 28385 5150
rect 28505 5030 28550 5150
rect 28670 5030 28715 5150
rect 28835 5030 28890 5150
rect 29010 5030 29055 5150
rect 29175 5030 29220 5150
rect 29340 5030 29385 5150
rect 29505 5030 29560 5150
rect 29680 5030 29690 5150
rect 24190 4975 29690 5030
rect 24190 4855 24200 4975
rect 24320 4855 24365 4975
rect 24485 4855 24530 4975
rect 24650 4855 24695 4975
rect 24815 4855 24870 4975
rect 24990 4855 25035 4975
rect 25155 4855 25200 4975
rect 25320 4855 25365 4975
rect 25485 4855 25540 4975
rect 25660 4855 25705 4975
rect 25825 4855 25870 4975
rect 25990 4855 26035 4975
rect 26155 4855 26210 4975
rect 26330 4855 26375 4975
rect 26495 4855 26540 4975
rect 26660 4855 26705 4975
rect 26825 4855 26880 4975
rect 27000 4855 27045 4975
rect 27165 4855 27210 4975
rect 27330 4855 27375 4975
rect 27495 4855 27550 4975
rect 27670 4855 27715 4975
rect 27835 4855 27880 4975
rect 28000 4855 28045 4975
rect 28165 4855 28220 4975
rect 28340 4855 28385 4975
rect 28505 4855 28550 4975
rect 28670 4855 28715 4975
rect 28835 4855 28890 4975
rect 29010 4855 29055 4975
rect 29175 4855 29220 4975
rect 29340 4855 29385 4975
rect 29505 4855 29560 4975
rect 29680 4855 29690 4975
rect 24190 4810 29690 4855
rect 24190 4690 24200 4810
rect 24320 4690 24365 4810
rect 24485 4690 24530 4810
rect 24650 4690 24695 4810
rect 24815 4690 24870 4810
rect 24990 4690 25035 4810
rect 25155 4690 25200 4810
rect 25320 4690 25365 4810
rect 25485 4690 25540 4810
rect 25660 4690 25705 4810
rect 25825 4690 25870 4810
rect 25990 4690 26035 4810
rect 26155 4690 26210 4810
rect 26330 4690 26375 4810
rect 26495 4690 26540 4810
rect 26660 4690 26705 4810
rect 26825 4690 26880 4810
rect 27000 4690 27045 4810
rect 27165 4690 27210 4810
rect 27330 4690 27375 4810
rect 27495 4690 27550 4810
rect 27670 4690 27715 4810
rect 27835 4690 27880 4810
rect 28000 4690 28045 4810
rect 28165 4690 28220 4810
rect 28340 4690 28385 4810
rect 28505 4690 28550 4810
rect 28670 4690 28715 4810
rect 28835 4690 28890 4810
rect 29010 4690 29055 4810
rect 29175 4690 29220 4810
rect 29340 4690 29385 4810
rect 29505 4690 29560 4810
rect 29680 4690 29690 4810
rect 24190 4645 29690 4690
rect 24190 4525 24200 4645
rect 24320 4525 24365 4645
rect 24485 4525 24530 4645
rect 24650 4525 24695 4645
rect 24815 4525 24870 4645
rect 24990 4525 25035 4645
rect 25155 4525 25200 4645
rect 25320 4525 25365 4645
rect 25485 4525 25540 4645
rect 25660 4525 25705 4645
rect 25825 4525 25870 4645
rect 25990 4525 26035 4645
rect 26155 4525 26210 4645
rect 26330 4525 26375 4645
rect 26495 4525 26540 4645
rect 26660 4525 26705 4645
rect 26825 4525 26880 4645
rect 27000 4525 27045 4645
rect 27165 4525 27210 4645
rect 27330 4525 27375 4645
rect 27495 4525 27550 4645
rect 27670 4525 27715 4645
rect 27835 4525 27880 4645
rect 28000 4525 28045 4645
rect 28165 4525 28220 4645
rect 28340 4525 28385 4645
rect 28505 4525 28550 4645
rect 28670 4525 28715 4645
rect 28835 4525 28890 4645
rect 29010 4525 29055 4645
rect 29175 4525 29220 4645
rect 29340 4525 29385 4645
rect 29505 4525 29560 4645
rect 29680 4525 29690 4645
rect 24190 4480 29690 4525
rect 24190 4360 24200 4480
rect 24320 4360 24365 4480
rect 24485 4360 24530 4480
rect 24650 4360 24695 4480
rect 24815 4360 24870 4480
rect 24990 4360 25035 4480
rect 25155 4360 25200 4480
rect 25320 4360 25365 4480
rect 25485 4360 25540 4480
rect 25660 4360 25705 4480
rect 25825 4360 25870 4480
rect 25990 4360 26035 4480
rect 26155 4360 26210 4480
rect 26330 4360 26375 4480
rect 26495 4360 26540 4480
rect 26660 4360 26705 4480
rect 26825 4360 26880 4480
rect 27000 4360 27045 4480
rect 27165 4360 27210 4480
rect 27330 4360 27375 4480
rect 27495 4360 27550 4480
rect 27670 4360 27715 4480
rect 27835 4360 27880 4480
rect 28000 4360 28045 4480
rect 28165 4360 28220 4480
rect 28340 4360 28385 4480
rect 28505 4360 28550 4480
rect 28670 4360 28715 4480
rect 28835 4360 28890 4480
rect 29010 4360 29055 4480
rect 29175 4360 29220 4480
rect 29340 4360 29385 4480
rect 29505 4360 29560 4480
rect 29680 4360 29690 4480
rect 24190 4305 29690 4360
rect 24190 4185 24200 4305
rect 24320 4185 24365 4305
rect 24485 4185 24530 4305
rect 24650 4185 24695 4305
rect 24815 4185 24870 4305
rect 24990 4185 25035 4305
rect 25155 4185 25200 4305
rect 25320 4185 25365 4305
rect 25485 4185 25540 4305
rect 25660 4185 25705 4305
rect 25825 4185 25870 4305
rect 25990 4185 26035 4305
rect 26155 4185 26210 4305
rect 26330 4185 26375 4305
rect 26495 4185 26540 4305
rect 26660 4185 26705 4305
rect 26825 4185 26880 4305
rect 27000 4185 27045 4305
rect 27165 4185 27210 4305
rect 27330 4185 27375 4305
rect 27495 4185 27550 4305
rect 27670 4185 27715 4305
rect 27835 4185 27880 4305
rect 28000 4185 28045 4305
rect 28165 4185 28220 4305
rect 28340 4185 28385 4305
rect 28505 4185 28550 4305
rect 28670 4185 28715 4305
rect 28835 4185 28890 4305
rect 29010 4185 29055 4305
rect 29175 4185 29220 4305
rect 29340 4185 29385 4305
rect 29505 4185 29560 4305
rect 29680 4185 29690 4305
rect 24190 4140 29690 4185
rect 24190 4020 24200 4140
rect 24320 4020 24365 4140
rect 24485 4020 24530 4140
rect 24650 4020 24695 4140
rect 24815 4020 24870 4140
rect 24990 4020 25035 4140
rect 25155 4020 25200 4140
rect 25320 4020 25365 4140
rect 25485 4020 25540 4140
rect 25660 4020 25705 4140
rect 25825 4020 25870 4140
rect 25990 4020 26035 4140
rect 26155 4020 26210 4140
rect 26330 4020 26375 4140
rect 26495 4020 26540 4140
rect 26660 4020 26705 4140
rect 26825 4020 26880 4140
rect 27000 4020 27045 4140
rect 27165 4020 27210 4140
rect 27330 4020 27375 4140
rect 27495 4020 27550 4140
rect 27670 4020 27715 4140
rect 27835 4020 27880 4140
rect 28000 4020 28045 4140
rect 28165 4020 28220 4140
rect 28340 4020 28385 4140
rect 28505 4020 28550 4140
rect 28670 4020 28715 4140
rect 28835 4020 28890 4140
rect 29010 4020 29055 4140
rect 29175 4020 29220 4140
rect 29340 4020 29385 4140
rect 29505 4020 29560 4140
rect 29680 4020 29690 4140
rect 24190 3975 29690 4020
rect 24190 3855 24200 3975
rect 24320 3855 24365 3975
rect 24485 3855 24530 3975
rect 24650 3855 24695 3975
rect 24815 3855 24870 3975
rect 24990 3855 25035 3975
rect 25155 3855 25200 3975
rect 25320 3855 25365 3975
rect 25485 3855 25540 3975
rect 25660 3855 25705 3975
rect 25825 3855 25870 3975
rect 25990 3855 26035 3975
rect 26155 3855 26210 3975
rect 26330 3855 26375 3975
rect 26495 3855 26540 3975
rect 26660 3855 26705 3975
rect 26825 3855 26880 3975
rect 27000 3855 27045 3975
rect 27165 3855 27210 3975
rect 27330 3855 27375 3975
rect 27495 3855 27550 3975
rect 27670 3855 27715 3975
rect 27835 3855 27880 3975
rect 28000 3855 28045 3975
rect 28165 3855 28220 3975
rect 28340 3855 28385 3975
rect 28505 3855 28550 3975
rect 28670 3855 28715 3975
rect 28835 3855 28890 3975
rect 29010 3855 29055 3975
rect 29175 3855 29220 3975
rect 29340 3855 29385 3975
rect 29505 3855 29560 3975
rect 29680 3855 29690 3975
rect 24190 3810 29690 3855
rect 24190 3690 24200 3810
rect 24320 3690 24365 3810
rect 24485 3690 24530 3810
rect 24650 3690 24695 3810
rect 24815 3690 24870 3810
rect 24990 3690 25035 3810
rect 25155 3690 25200 3810
rect 25320 3690 25365 3810
rect 25485 3690 25540 3810
rect 25660 3690 25705 3810
rect 25825 3690 25870 3810
rect 25990 3690 26035 3810
rect 26155 3690 26210 3810
rect 26330 3690 26375 3810
rect 26495 3690 26540 3810
rect 26660 3690 26705 3810
rect 26825 3690 26880 3810
rect 27000 3690 27045 3810
rect 27165 3690 27210 3810
rect 27330 3690 27375 3810
rect 27495 3690 27550 3810
rect 27670 3690 27715 3810
rect 27835 3690 27880 3810
rect 28000 3690 28045 3810
rect 28165 3690 28220 3810
rect 28340 3690 28385 3810
rect 28505 3690 28550 3810
rect 28670 3690 28715 3810
rect 28835 3690 28890 3810
rect 29010 3690 29055 3810
rect 29175 3690 29220 3810
rect 29340 3690 29385 3810
rect 29505 3690 29560 3810
rect 29680 3690 29690 3810
rect 24190 3635 29690 3690
rect 24190 3515 24200 3635
rect 24320 3515 24365 3635
rect 24485 3515 24530 3635
rect 24650 3515 24695 3635
rect 24815 3515 24870 3635
rect 24990 3515 25035 3635
rect 25155 3515 25200 3635
rect 25320 3515 25365 3635
rect 25485 3515 25540 3635
rect 25660 3515 25705 3635
rect 25825 3515 25870 3635
rect 25990 3515 26035 3635
rect 26155 3515 26210 3635
rect 26330 3515 26375 3635
rect 26495 3515 26540 3635
rect 26660 3515 26705 3635
rect 26825 3515 26880 3635
rect 27000 3515 27045 3635
rect 27165 3515 27210 3635
rect 27330 3515 27375 3635
rect 27495 3515 27550 3635
rect 27670 3515 27715 3635
rect 27835 3515 27880 3635
rect 28000 3515 28045 3635
rect 28165 3515 28220 3635
rect 28340 3515 28385 3635
rect 28505 3515 28550 3635
rect 28670 3515 28715 3635
rect 28835 3515 28890 3635
rect 29010 3515 29055 3635
rect 29175 3515 29220 3635
rect 29340 3515 29385 3635
rect 29505 3515 29560 3635
rect 29680 3515 29690 3635
rect 24190 3470 29690 3515
rect 24190 3350 24200 3470
rect 24320 3350 24365 3470
rect 24485 3350 24530 3470
rect 24650 3350 24695 3470
rect 24815 3350 24870 3470
rect 24990 3350 25035 3470
rect 25155 3350 25200 3470
rect 25320 3350 25365 3470
rect 25485 3350 25540 3470
rect 25660 3350 25705 3470
rect 25825 3350 25870 3470
rect 25990 3350 26035 3470
rect 26155 3350 26210 3470
rect 26330 3350 26375 3470
rect 26495 3350 26540 3470
rect 26660 3350 26705 3470
rect 26825 3350 26880 3470
rect 27000 3350 27045 3470
rect 27165 3350 27210 3470
rect 27330 3350 27375 3470
rect 27495 3350 27550 3470
rect 27670 3350 27715 3470
rect 27835 3350 27880 3470
rect 28000 3350 28045 3470
rect 28165 3350 28220 3470
rect 28340 3350 28385 3470
rect 28505 3350 28550 3470
rect 28670 3350 28715 3470
rect 28835 3350 28890 3470
rect 29010 3350 29055 3470
rect 29175 3350 29220 3470
rect 29340 3350 29385 3470
rect 29505 3350 29560 3470
rect 29680 3350 29690 3470
rect 24190 3305 29690 3350
rect 24190 3185 24200 3305
rect 24320 3185 24365 3305
rect 24485 3185 24530 3305
rect 24650 3185 24695 3305
rect 24815 3185 24870 3305
rect 24990 3185 25035 3305
rect 25155 3185 25200 3305
rect 25320 3185 25365 3305
rect 25485 3185 25540 3305
rect 25660 3185 25705 3305
rect 25825 3185 25870 3305
rect 25990 3185 26035 3305
rect 26155 3185 26210 3305
rect 26330 3185 26375 3305
rect 26495 3185 26540 3305
rect 26660 3185 26705 3305
rect 26825 3185 26880 3305
rect 27000 3185 27045 3305
rect 27165 3185 27210 3305
rect 27330 3185 27375 3305
rect 27495 3185 27550 3305
rect 27670 3185 27715 3305
rect 27835 3185 27880 3305
rect 28000 3185 28045 3305
rect 28165 3185 28220 3305
rect 28340 3185 28385 3305
rect 28505 3185 28550 3305
rect 28670 3185 28715 3305
rect 28835 3185 28890 3305
rect 29010 3185 29055 3305
rect 29175 3185 29220 3305
rect 29340 3185 29385 3305
rect 29505 3185 29560 3305
rect 29680 3185 29690 3305
rect 24190 3140 29690 3185
rect 24190 3020 24200 3140
rect 24320 3020 24365 3140
rect 24485 3020 24530 3140
rect 24650 3020 24695 3140
rect 24815 3020 24870 3140
rect 24990 3020 25035 3140
rect 25155 3020 25200 3140
rect 25320 3020 25365 3140
rect 25485 3020 25540 3140
rect 25660 3020 25705 3140
rect 25825 3020 25870 3140
rect 25990 3020 26035 3140
rect 26155 3020 26210 3140
rect 26330 3020 26375 3140
rect 26495 3020 26540 3140
rect 26660 3020 26705 3140
rect 26825 3020 26880 3140
rect 27000 3020 27045 3140
rect 27165 3020 27210 3140
rect 27330 3020 27375 3140
rect 27495 3020 27550 3140
rect 27670 3020 27715 3140
rect 27835 3020 27880 3140
rect 28000 3020 28045 3140
rect 28165 3020 28220 3140
rect 28340 3020 28385 3140
rect 28505 3020 28550 3140
rect 28670 3020 28715 3140
rect 28835 3020 28890 3140
rect 29010 3020 29055 3140
rect 29175 3020 29220 3140
rect 29340 3020 29385 3140
rect 29505 3020 29560 3140
rect 29680 3020 29690 3140
rect 24190 2965 29690 3020
rect 24190 2845 24200 2965
rect 24320 2845 24365 2965
rect 24485 2845 24530 2965
rect 24650 2845 24695 2965
rect 24815 2845 24870 2965
rect 24990 2845 25035 2965
rect 25155 2845 25200 2965
rect 25320 2845 25365 2965
rect 25485 2845 25540 2965
rect 25660 2845 25705 2965
rect 25825 2845 25870 2965
rect 25990 2845 26035 2965
rect 26155 2845 26210 2965
rect 26330 2845 26375 2965
rect 26495 2845 26540 2965
rect 26660 2845 26705 2965
rect 26825 2845 26880 2965
rect 27000 2845 27045 2965
rect 27165 2845 27210 2965
rect 27330 2845 27375 2965
rect 27495 2845 27550 2965
rect 27670 2845 27715 2965
rect 27835 2845 27880 2965
rect 28000 2845 28045 2965
rect 28165 2845 28220 2965
rect 28340 2845 28385 2965
rect 28505 2845 28550 2965
rect 28670 2845 28715 2965
rect 28835 2845 28890 2965
rect 29010 2845 29055 2965
rect 29175 2845 29220 2965
rect 29340 2845 29385 2965
rect 29505 2845 29560 2965
rect 29680 2845 29690 2965
rect 24190 2800 29690 2845
rect 24190 2680 24200 2800
rect 24320 2680 24365 2800
rect 24485 2680 24530 2800
rect 24650 2680 24695 2800
rect 24815 2680 24870 2800
rect 24990 2680 25035 2800
rect 25155 2680 25200 2800
rect 25320 2680 25365 2800
rect 25485 2680 25540 2800
rect 25660 2680 25705 2800
rect 25825 2680 25870 2800
rect 25990 2680 26035 2800
rect 26155 2680 26210 2800
rect 26330 2680 26375 2800
rect 26495 2680 26540 2800
rect 26660 2680 26705 2800
rect 26825 2680 26880 2800
rect 27000 2680 27045 2800
rect 27165 2680 27210 2800
rect 27330 2680 27375 2800
rect 27495 2680 27550 2800
rect 27670 2680 27715 2800
rect 27835 2680 27880 2800
rect 28000 2680 28045 2800
rect 28165 2680 28220 2800
rect 28340 2680 28385 2800
rect 28505 2680 28550 2800
rect 28670 2680 28715 2800
rect 28835 2680 28890 2800
rect 29010 2680 29055 2800
rect 29175 2680 29220 2800
rect 29340 2680 29385 2800
rect 29505 2680 29560 2800
rect 29680 2680 29690 2800
rect 24190 2635 29690 2680
rect 24190 2515 24200 2635
rect 24320 2515 24365 2635
rect 24485 2515 24530 2635
rect 24650 2515 24695 2635
rect 24815 2515 24870 2635
rect 24990 2515 25035 2635
rect 25155 2515 25200 2635
rect 25320 2515 25365 2635
rect 25485 2515 25540 2635
rect 25660 2515 25705 2635
rect 25825 2515 25870 2635
rect 25990 2515 26035 2635
rect 26155 2515 26210 2635
rect 26330 2515 26375 2635
rect 26495 2515 26540 2635
rect 26660 2515 26705 2635
rect 26825 2515 26880 2635
rect 27000 2515 27045 2635
rect 27165 2515 27210 2635
rect 27330 2515 27375 2635
rect 27495 2515 27550 2635
rect 27670 2515 27715 2635
rect 27835 2515 27880 2635
rect 28000 2515 28045 2635
rect 28165 2515 28220 2635
rect 28340 2515 28385 2635
rect 28505 2515 28550 2635
rect 28670 2515 28715 2635
rect 28835 2515 28890 2635
rect 29010 2515 29055 2635
rect 29175 2515 29220 2635
rect 29340 2515 29385 2635
rect 29505 2515 29560 2635
rect 29680 2515 29690 2635
rect 24190 2470 29690 2515
rect 24190 2350 24200 2470
rect 24320 2350 24365 2470
rect 24485 2350 24530 2470
rect 24650 2350 24695 2470
rect 24815 2350 24870 2470
rect 24990 2350 25035 2470
rect 25155 2350 25200 2470
rect 25320 2350 25365 2470
rect 25485 2350 25540 2470
rect 25660 2350 25705 2470
rect 25825 2350 25870 2470
rect 25990 2350 26035 2470
rect 26155 2350 26210 2470
rect 26330 2350 26375 2470
rect 26495 2350 26540 2470
rect 26660 2350 26705 2470
rect 26825 2350 26880 2470
rect 27000 2350 27045 2470
rect 27165 2350 27210 2470
rect 27330 2350 27375 2470
rect 27495 2350 27550 2470
rect 27670 2350 27715 2470
rect 27835 2350 27880 2470
rect 28000 2350 28045 2470
rect 28165 2350 28220 2470
rect 28340 2350 28385 2470
rect 28505 2350 28550 2470
rect 28670 2350 28715 2470
rect 28835 2350 28890 2470
rect 29010 2350 29055 2470
rect 29175 2350 29220 2470
rect 29340 2350 29385 2470
rect 29505 2350 29560 2470
rect 29680 2350 29690 2470
rect 24190 2295 29690 2350
rect 24190 2175 24200 2295
rect 24320 2175 24365 2295
rect 24485 2175 24530 2295
rect 24650 2175 24695 2295
rect 24815 2175 24870 2295
rect 24990 2175 25035 2295
rect 25155 2175 25200 2295
rect 25320 2175 25365 2295
rect 25485 2175 25540 2295
rect 25660 2175 25705 2295
rect 25825 2175 25870 2295
rect 25990 2175 26035 2295
rect 26155 2175 26210 2295
rect 26330 2175 26375 2295
rect 26495 2175 26540 2295
rect 26660 2175 26705 2295
rect 26825 2175 26880 2295
rect 27000 2175 27045 2295
rect 27165 2175 27210 2295
rect 27330 2175 27375 2295
rect 27495 2175 27550 2295
rect 27670 2175 27715 2295
rect 27835 2175 27880 2295
rect 28000 2175 28045 2295
rect 28165 2175 28220 2295
rect 28340 2175 28385 2295
rect 28505 2175 28550 2295
rect 28670 2175 28715 2295
rect 28835 2175 28890 2295
rect 29010 2175 29055 2295
rect 29175 2175 29220 2295
rect 29340 2175 29385 2295
rect 29505 2175 29560 2295
rect 29680 2175 29690 2295
rect 24190 2130 29690 2175
rect 24190 2010 24200 2130
rect 24320 2010 24365 2130
rect 24485 2010 24530 2130
rect 24650 2010 24695 2130
rect 24815 2010 24870 2130
rect 24990 2010 25035 2130
rect 25155 2010 25200 2130
rect 25320 2010 25365 2130
rect 25485 2010 25540 2130
rect 25660 2010 25705 2130
rect 25825 2010 25870 2130
rect 25990 2010 26035 2130
rect 26155 2010 26210 2130
rect 26330 2010 26375 2130
rect 26495 2010 26540 2130
rect 26660 2010 26705 2130
rect 26825 2010 26880 2130
rect 27000 2010 27045 2130
rect 27165 2010 27210 2130
rect 27330 2010 27375 2130
rect 27495 2010 27550 2130
rect 27670 2010 27715 2130
rect 27835 2010 27880 2130
rect 28000 2010 28045 2130
rect 28165 2010 28220 2130
rect 28340 2010 28385 2130
rect 28505 2010 28550 2130
rect 28670 2010 28715 2130
rect 28835 2010 28890 2130
rect 29010 2010 29055 2130
rect 29175 2010 29220 2130
rect 29340 2010 29385 2130
rect 29505 2010 29560 2130
rect 29680 2010 29690 2130
rect 24190 1965 29690 2010
rect 24190 1845 24200 1965
rect 24320 1845 24365 1965
rect 24485 1845 24530 1965
rect 24650 1845 24695 1965
rect 24815 1845 24870 1965
rect 24990 1845 25035 1965
rect 25155 1845 25200 1965
rect 25320 1845 25365 1965
rect 25485 1845 25540 1965
rect 25660 1845 25705 1965
rect 25825 1845 25870 1965
rect 25990 1845 26035 1965
rect 26155 1845 26210 1965
rect 26330 1845 26375 1965
rect 26495 1845 26540 1965
rect 26660 1845 26705 1965
rect 26825 1845 26880 1965
rect 27000 1845 27045 1965
rect 27165 1845 27210 1965
rect 27330 1845 27375 1965
rect 27495 1845 27550 1965
rect 27670 1845 27715 1965
rect 27835 1845 27880 1965
rect 28000 1845 28045 1965
rect 28165 1845 28220 1965
rect 28340 1845 28385 1965
rect 28505 1845 28550 1965
rect 28670 1845 28715 1965
rect 28835 1845 28890 1965
rect 29010 1845 29055 1965
rect 29175 1845 29220 1965
rect 29340 1845 29385 1965
rect 29505 1845 29560 1965
rect 29680 1845 29690 1965
rect 24190 1800 29690 1845
rect 24190 1680 24200 1800
rect 24320 1680 24365 1800
rect 24485 1680 24530 1800
rect 24650 1680 24695 1800
rect 24815 1680 24870 1800
rect 24990 1680 25035 1800
rect 25155 1680 25200 1800
rect 25320 1680 25365 1800
rect 25485 1680 25540 1800
rect 25660 1680 25705 1800
rect 25825 1680 25870 1800
rect 25990 1680 26035 1800
rect 26155 1680 26210 1800
rect 26330 1680 26375 1800
rect 26495 1680 26540 1800
rect 26660 1680 26705 1800
rect 26825 1680 26880 1800
rect 27000 1680 27045 1800
rect 27165 1680 27210 1800
rect 27330 1680 27375 1800
rect 27495 1680 27550 1800
rect 27670 1680 27715 1800
rect 27835 1680 27880 1800
rect 28000 1680 28045 1800
rect 28165 1680 28220 1800
rect 28340 1680 28385 1800
rect 28505 1680 28550 1800
rect 28670 1680 28715 1800
rect 28835 1680 28890 1800
rect 29010 1680 29055 1800
rect 29175 1680 29220 1800
rect 29340 1680 29385 1800
rect 29505 1680 29560 1800
rect 29680 1680 29690 1800
rect 24190 1670 29690 1680
rect 7120 1380 12620 1390
rect 7120 1260 7130 1380
rect 7250 1260 7305 1380
rect 7425 1260 7470 1380
rect 7590 1260 7635 1380
rect 7755 1260 7800 1380
rect 7920 1260 7975 1380
rect 8095 1260 8140 1380
rect 8260 1260 8305 1380
rect 8425 1260 8470 1380
rect 8590 1260 8645 1380
rect 8765 1260 8810 1380
rect 8930 1260 8975 1380
rect 9095 1260 9140 1380
rect 9260 1260 9315 1380
rect 9435 1260 9480 1380
rect 9600 1260 9645 1380
rect 9765 1260 9810 1380
rect 9930 1260 9985 1380
rect 10105 1260 10150 1380
rect 10270 1260 10315 1380
rect 10435 1260 10480 1380
rect 10600 1260 10655 1380
rect 10775 1260 10820 1380
rect 10940 1260 10985 1380
rect 11105 1260 11150 1380
rect 11270 1260 11325 1380
rect 11445 1260 11490 1380
rect 11610 1260 11655 1380
rect 11775 1260 11820 1380
rect 11940 1260 11995 1380
rect 12115 1260 12160 1380
rect 12280 1260 12325 1380
rect 12445 1260 12490 1380
rect 12610 1260 12620 1380
rect 7120 1215 12620 1260
rect 7120 1095 7130 1215
rect 7250 1095 7305 1215
rect 7425 1095 7470 1215
rect 7590 1095 7635 1215
rect 7755 1095 7800 1215
rect 7920 1095 7975 1215
rect 8095 1095 8140 1215
rect 8260 1095 8305 1215
rect 8425 1095 8470 1215
rect 8590 1095 8645 1215
rect 8765 1095 8810 1215
rect 8930 1095 8975 1215
rect 9095 1095 9140 1215
rect 9260 1095 9315 1215
rect 9435 1095 9480 1215
rect 9600 1095 9645 1215
rect 9765 1095 9810 1215
rect 9930 1095 9985 1215
rect 10105 1095 10150 1215
rect 10270 1095 10315 1215
rect 10435 1095 10480 1215
rect 10600 1095 10655 1215
rect 10775 1095 10820 1215
rect 10940 1095 10985 1215
rect 11105 1095 11150 1215
rect 11270 1095 11325 1215
rect 11445 1095 11490 1215
rect 11610 1095 11655 1215
rect 11775 1095 11820 1215
rect 11940 1095 11995 1215
rect 12115 1095 12160 1215
rect 12280 1095 12325 1215
rect 12445 1095 12490 1215
rect 12610 1095 12620 1215
rect 7120 1050 12620 1095
rect 7120 930 7130 1050
rect 7250 930 7305 1050
rect 7425 930 7470 1050
rect 7590 930 7635 1050
rect 7755 930 7800 1050
rect 7920 930 7975 1050
rect 8095 930 8140 1050
rect 8260 930 8305 1050
rect 8425 930 8470 1050
rect 8590 930 8645 1050
rect 8765 930 8810 1050
rect 8930 930 8975 1050
rect 9095 930 9140 1050
rect 9260 930 9315 1050
rect 9435 930 9480 1050
rect 9600 930 9645 1050
rect 9765 930 9810 1050
rect 9930 930 9985 1050
rect 10105 930 10150 1050
rect 10270 930 10315 1050
rect 10435 930 10480 1050
rect 10600 930 10655 1050
rect 10775 930 10820 1050
rect 10940 930 10985 1050
rect 11105 930 11150 1050
rect 11270 930 11325 1050
rect 11445 930 11490 1050
rect 11610 930 11655 1050
rect 11775 930 11820 1050
rect 11940 930 11995 1050
rect 12115 930 12160 1050
rect 12280 930 12325 1050
rect 12445 930 12490 1050
rect 12610 930 12620 1050
rect 7120 885 12620 930
rect 7120 765 7130 885
rect 7250 765 7305 885
rect 7425 765 7470 885
rect 7590 765 7635 885
rect 7755 765 7800 885
rect 7920 765 7975 885
rect 8095 765 8140 885
rect 8260 765 8305 885
rect 8425 765 8470 885
rect 8590 765 8645 885
rect 8765 765 8810 885
rect 8930 765 8975 885
rect 9095 765 9140 885
rect 9260 765 9315 885
rect 9435 765 9480 885
rect 9600 765 9645 885
rect 9765 765 9810 885
rect 9930 765 9985 885
rect 10105 765 10150 885
rect 10270 765 10315 885
rect 10435 765 10480 885
rect 10600 765 10655 885
rect 10775 765 10820 885
rect 10940 765 10985 885
rect 11105 765 11150 885
rect 11270 765 11325 885
rect 11445 765 11490 885
rect 11610 765 11655 885
rect 11775 765 11820 885
rect 11940 765 11995 885
rect 12115 765 12160 885
rect 12280 765 12325 885
rect 12445 765 12490 885
rect 12610 765 12620 885
rect 7120 710 12620 765
rect 7120 590 7130 710
rect 7250 590 7305 710
rect 7425 590 7470 710
rect 7590 590 7635 710
rect 7755 590 7800 710
rect 7920 590 7975 710
rect 8095 590 8140 710
rect 8260 590 8305 710
rect 8425 590 8470 710
rect 8590 590 8645 710
rect 8765 590 8810 710
rect 8930 590 8975 710
rect 9095 590 9140 710
rect 9260 590 9315 710
rect 9435 590 9480 710
rect 9600 590 9645 710
rect 9765 590 9810 710
rect 9930 590 9985 710
rect 10105 590 10150 710
rect 10270 590 10315 710
rect 10435 590 10480 710
rect 10600 590 10655 710
rect 10775 590 10820 710
rect 10940 590 10985 710
rect 11105 590 11150 710
rect 11270 590 11325 710
rect 11445 590 11490 710
rect 11610 590 11655 710
rect 11775 590 11820 710
rect 11940 590 11995 710
rect 12115 590 12160 710
rect 12280 590 12325 710
rect 12445 590 12490 710
rect 12610 590 12620 710
rect 7120 545 12620 590
rect 7120 425 7130 545
rect 7250 425 7305 545
rect 7425 425 7470 545
rect 7590 425 7635 545
rect 7755 425 7800 545
rect 7920 425 7975 545
rect 8095 425 8140 545
rect 8260 425 8305 545
rect 8425 425 8470 545
rect 8590 425 8645 545
rect 8765 425 8810 545
rect 8930 425 8975 545
rect 9095 425 9140 545
rect 9260 425 9315 545
rect 9435 425 9480 545
rect 9600 425 9645 545
rect 9765 425 9810 545
rect 9930 425 9985 545
rect 10105 425 10150 545
rect 10270 425 10315 545
rect 10435 425 10480 545
rect 10600 425 10655 545
rect 10775 425 10820 545
rect 10940 425 10985 545
rect 11105 425 11150 545
rect 11270 425 11325 545
rect 11445 425 11490 545
rect 11610 425 11655 545
rect 11775 425 11820 545
rect 11940 425 11995 545
rect 12115 425 12160 545
rect 12280 425 12325 545
rect 12445 425 12490 545
rect 12610 425 12620 545
rect 7120 380 12620 425
rect 7120 260 7130 380
rect 7250 260 7305 380
rect 7425 260 7470 380
rect 7590 260 7635 380
rect 7755 260 7800 380
rect 7920 260 7975 380
rect 8095 260 8140 380
rect 8260 260 8305 380
rect 8425 260 8470 380
rect 8590 260 8645 380
rect 8765 260 8810 380
rect 8930 260 8975 380
rect 9095 260 9140 380
rect 9260 260 9315 380
rect 9435 260 9480 380
rect 9600 260 9645 380
rect 9765 260 9810 380
rect 9930 260 9985 380
rect 10105 260 10150 380
rect 10270 260 10315 380
rect 10435 260 10480 380
rect 10600 260 10655 380
rect 10775 260 10820 380
rect 10940 260 10985 380
rect 11105 260 11150 380
rect 11270 260 11325 380
rect 11445 260 11490 380
rect 11610 260 11655 380
rect 11775 260 11820 380
rect 11940 260 11995 380
rect 12115 260 12160 380
rect 12280 260 12325 380
rect 12445 260 12490 380
rect 12610 260 12620 380
rect 7120 215 12620 260
rect 7120 95 7130 215
rect 7250 95 7305 215
rect 7425 95 7470 215
rect 7590 95 7635 215
rect 7755 95 7800 215
rect 7920 95 7975 215
rect 8095 95 8140 215
rect 8260 95 8305 215
rect 8425 95 8470 215
rect 8590 95 8645 215
rect 8765 95 8810 215
rect 8930 95 8975 215
rect 9095 95 9140 215
rect 9260 95 9315 215
rect 9435 95 9480 215
rect 9600 95 9645 215
rect 9765 95 9810 215
rect 9930 95 9985 215
rect 10105 95 10150 215
rect 10270 95 10315 215
rect 10435 95 10480 215
rect 10600 95 10655 215
rect 10775 95 10820 215
rect 10940 95 10985 215
rect 11105 95 11150 215
rect 11270 95 11325 215
rect 11445 95 11490 215
rect 11610 95 11655 215
rect 11775 95 11820 215
rect 11940 95 11995 215
rect 12115 95 12160 215
rect 12280 95 12325 215
rect 12445 95 12490 215
rect 12610 95 12620 215
rect 7120 40 12620 95
rect 7120 -80 7130 40
rect 7250 -80 7305 40
rect 7425 -80 7470 40
rect 7590 -80 7635 40
rect 7755 -80 7800 40
rect 7920 -80 7975 40
rect 8095 -80 8140 40
rect 8260 -80 8305 40
rect 8425 -80 8470 40
rect 8590 -80 8645 40
rect 8765 -80 8810 40
rect 8930 -80 8975 40
rect 9095 -80 9140 40
rect 9260 -80 9315 40
rect 9435 -80 9480 40
rect 9600 -80 9645 40
rect 9765 -80 9810 40
rect 9930 -80 9985 40
rect 10105 -80 10150 40
rect 10270 -80 10315 40
rect 10435 -80 10480 40
rect 10600 -80 10655 40
rect 10775 -80 10820 40
rect 10940 -80 10985 40
rect 11105 -80 11150 40
rect 11270 -80 11325 40
rect 11445 -80 11490 40
rect 11610 -80 11655 40
rect 11775 -80 11820 40
rect 11940 -80 11995 40
rect 12115 -80 12160 40
rect 12280 -80 12325 40
rect 12445 -80 12490 40
rect 12610 -80 12620 40
rect 7120 -125 12620 -80
rect 7120 -245 7130 -125
rect 7250 -245 7305 -125
rect 7425 -245 7470 -125
rect 7590 -245 7635 -125
rect 7755 -245 7800 -125
rect 7920 -245 7975 -125
rect 8095 -245 8140 -125
rect 8260 -245 8305 -125
rect 8425 -245 8470 -125
rect 8590 -245 8645 -125
rect 8765 -245 8810 -125
rect 8930 -245 8975 -125
rect 9095 -245 9140 -125
rect 9260 -245 9315 -125
rect 9435 -245 9480 -125
rect 9600 -245 9645 -125
rect 9765 -245 9810 -125
rect 9930 -245 9985 -125
rect 10105 -245 10150 -125
rect 10270 -245 10315 -125
rect 10435 -245 10480 -125
rect 10600 -245 10655 -125
rect 10775 -245 10820 -125
rect 10940 -245 10985 -125
rect 11105 -245 11150 -125
rect 11270 -245 11325 -125
rect 11445 -245 11490 -125
rect 11610 -245 11655 -125
rect 11775 -245 11820 -125
rect 11940 -245 11995 -125
rect 12115 -245 12160 -125
rect 12280 -245 12325 -125
rect 12445 -245 12490 -125
rect 12610 -245 12620 -125
rect 7120 -290 12620 -245
rect 7120 -410 7130 -290
rect 7250 -410 7305 -290
rect 7425 -410 7470 -290
rect 7590 -410 7635 -290
rect 7755 -410 7800 -290
rect 7920 -410 7975 -290
rect 8095 -410 8140 -290
rect 8260 -410 8305 -290
rect 8425 -410 8470 -290
rect 8590 -410 8645 -290
rect 8765 -410 8810 -290
rect 8930 -410 8975 -290
rect 9095 -410 9140 -290
rect 9260 -410 9315 -290
rect 9435 -410 9480 -290
rect 9600 -410 9645 -290
rect 9765 -410 9810 -290
rect 9930 -410 9985 -290
rect 10105 -410 10150 -290
rect 10270 -410 10315 -290
rect 10435 -410 10480 -290
rect 10600 -410 10655 -290
rect 10775 -410 10820 -290
rect 10940 -410 10985 -290
rect 11105 -410 11150 -290
rect 11270 -410 11325 -290
rect 11445 -410 11490 -290
rect 11610 -410 11655 -290
rect 11775 -410 11820 -290
rect 11940 -410 11995 -290
rect 12115 -410 12160 -290
rect 12280 -410 12325 -290
rect 12445 -410 12490 -290
rect 12610 -410 12620 -290
rect 7120 -455 12620 -410
rect 7120 -575 7130 -455
rect 7250 -575 7305 -455
rect 7425 -575 7470 -455
rect 7590 -575 7635 -455
rect 7755 -575 7800 -455
rect 7920 -575 7975 -455
rect 8095 -575 8140 -455
rect 8260 -575 8305 -455
rect 8425 -575 8470 -455
rect 8590 -575 8645 -455
rect 8765 -575 8810 -455
rect 8930 -575 8975 -455
rect 9095 -575 9140 -455
rect 9260 -575 9315 -455
rect 9435 -575 9480 -455
rect 9600 -575 9645 -455
rect 9765 -575 9810 -455
rect 9930 -575 9985 -455
rect 10105 -575 10150 -455
rect 10270 -575 10315 -455
rect 10435 -575 10480 -455
rect 10600 -575 10655 -455
rect 10775 -575 10820 -455
rect 10940 -575 10985 -455
rect 11105 -575 11150 -455
rect 11270 -575 11325 -455
rect 11445 -575 11490 -455
rect 11610 -575 11655 -455
rect 11775 -575 11820 -455
rect 11940 -575 11995 -455
rect 12115 -575 12160 -455
rect 12280 -575 12325 -455
rect 12445 -575 12490 -455
rect 12610 -575 12620 -455
rect 7120 -630 12620 -575
rect 7120 -750 7130 -630
rect 7250 -750 7305 -630
rect 7425 -750 7470 -630
rect 7590 -750 7635 -630
rect 7755 -750 7800 -630
rect 7920 -750 7975 -630
rect 8095 -750 8140 -630
rect 8260 -750 8305 -630
rect 8425 -750 8470 -630
rect 8590 -750 8645 -630
rect 8765 -750 8810 -630
rect 8930 -750 8975 -630
rect 9095 -750 9140 -630
rect 9260 -750 9315 -630
rect 9435 -750 9480 -630
rect 9600 -750 9645 -630
rect 9765 -750 9810 -630
rect 9930 -750 9985 -630
rect 10105 -750 10150 -630
rect 10270 -750 10315 -630
rect 10435 -750 10480 -630
rect 10600 -750 10655 -630
rect 10775 -750 10820 -630
rect 10940 -750 10985 -630
rect 11105 -750 11150 -630
rect 11270 -750 11325 -630
rect 11445 -750 11490 -630
rect 11610 -750 11655 -630
rect 11775 -750 11820 -630
rect 11940 -750 11995 -630
rect 12115 -750 12160 -630
rect 12280 -750 12325 -630
rect 12445 -750 12490 -630
rect 12610 -750 12620 -630
rect 7120 -795 12620 -750
rect 7120 -915 7130 -795
rect 7250 -915 7305 -795
rect 7425 -915 7470 -795
rect 7590 -915 7635 -795
rect 7755 -915 7800 -795
rect 7920 -915 7975 -795
rect 8095 -915 8140 -795
rect 8260 -915 8305 -795
rect 8425 -915 8470 -795
rect 8590 -915 8645 -795
rect 8765 -915 8810 -795
rect 8930 -915 8975 -795
rect 9095 -915 9140 -795
rect 9260 -915 9315 -795
rect 9435 -915 9480 -795
rect 9600 -915 9645 -795
rect 9765 -915 9810 -795
rect 9930 -915 9985 -795
rect 10105 -915 10150 -795
rect 10270 -915 10315 -795
rect 10435 -915 10480 -795
rect 10600 -915 10655 -795
rect 10775 -915 10820 -795
rect 10940 -915 10985 -795
rect 11105 -915 11150 -795
rect 11270 -915 11325 -795
rect 11445 -915 11490 -795
rect 11610 -915 11655 -795
rect 11775 -915 11820 -795
rect 11940 -915 11995 -795
rect 12115 -915 12160 -795
rect 12280 -915 12325 -795
rect 12445 -915 12490 -795
rect 12610 -915 12620 -795
rect 7120 -960 12620 -915
rect 7120 -1080 7130 -960
rect 7250 -1080 7305 -960
rect 7425 -1080 7470 -960
rect 7590 -1080 7635 -960
rect 7755 -1080 7800 -960
rect 7920 -1080 7975 -960
rect 8095 -1080 8140 -960
rect 8260 -1080 8305 -960
rect 8425 -1080 8470 -960
rect 8590 -1080 8645 -960
rect 8765 -1080 8810 -960
rect 8930 -1080 8975 -960
rect 9095 -1080 9140 -960
rect 9260 -1080 9315 -960
rect 9435 -1080 9480 -960
rect 9600 -1080 9645 -960
rect 9765 -1080 9810 -960
rect 9930 -1080 9985 -960
rect 10105 -1080 10150 -960
rect 10270 -1080 10315 -960
rect 10435 -1080 10480 -960
rect 10600 -1080 10655 -960
rect 10775 -1080 10820 -960
rect 10940 -1080 10985 -960
rect 11105 -1080 11150 -960
rect 11270 -1080 11325 -960
rect 11445 -1080 11490 -960
rect 11610 -1080 11655 -960
rect 11775 -1080 11820 -960
rect 11940 -1080 11995 -960
rect 12115 -1080 12160 -960
rect 12280 -1080 12325 -960
rect 12445 -1080 12490 -960
rect 12610 -1080 12620 -960
rect 7120 -1125 12620 -1080
rect 7120 -1245 7130 -1125
rect 7250 -1245 7305 -1125
rect 7425 -1245 7470 -1125
rect 7590 -1245 7635 -1125
rect 7755 -1245 7800 -1125
rect 7920 -1245 7975 -1125
rect 8095 -1245 8140 -1125
rect 8260 -1245 8305 -1125
rect 8425 -1245 8470 -1125
rect 8590 -1245 8645 -1125
rect 8765 -1245 8810 -1125
rect 8930 -1245 8975 -1125
rect 9095 -1245 9140 -1125
rect 9260 -1245 9315 -1125
rect 9435 -1245 9480 -1125
rect 9600 -1245 9645 -1125
rect 9765 -1245 9810 -1125
rect 9930 -1245 9985 -1125
rect 10105 -1245 10150 -1125
rect 10270 -1245 10315 -1125
rect 10435 -1245 10480 -1125
rect 10600 -1245 10655 -1125
rect 10775 -1245 10820 -1125
rect 10940 -1245 10985 -1125
rect 11105 -1245 11150 -1125
rect 11270 -1245 11325 -1125
rect 11445 -1245 11490 -1125
rect 11610 -1245 11655 -1125
rect 11775 -1245 11820 -1125
rect 11940 -1245 11995 -1125
rect 12115 -1245 12160 -1125
rect 12280 -1245 12325 -1125
rect 12445 -1245 12490 -1125
rect 12610 -1245 12620 -1125
rect 7120 -1300 12620 -1245
rect 7120 -1420 7130 -1300
rect 7250 -1420 7305 -1300
rect 7425 -1420 7470 -1300
rect 7590 -1420 7635 -1300
rect 7755 -1420 7800 -1300
rect 7920 -1420 7975 -1300
rect 8095 -1420 8140 -1300
rect 8260 -1420 8305 -1300
rect 8425 -1420 8470 -1300
rect 8590 -1420 8645 -1300
rect 8765 -1420 8810 -1300
rect 8930 -1420 8975 -1300
rect 9095 -1420 9140 -1300
rect 9260 -1420 9315 -1300
rect 9435 -1420 9480 -1300
rect 9600 -1420 9645 -1300
rect 9765 -1420 9810 -1300
rect 9930 -1420 9985 -1300
rect 10105 -1420 10150 -1300
rect 10270 -1420 10315 -1300
rect 10435 -1420 10480 -1300
rect 10600 -1420 10655 -1300
rect 10775 -1420 10820 -1300
rect 10940 -1420 10985 -1300
rect 11105 -1420 11150 -1300
rect 11270 -1420 11325 -1300
rect 11445 -1420 11490 -1300
rect 11610 -1420 11655 -1300
rect 11775 -1420 11820 -1300
rect 11940 -1420 11995 -1300
rect 12115 -1420 12160 -1300
rect 12280 -1420 12325 -1300
rect 12445 -1420 12490 -1300
rect 12610 -1420 12620 -1300
rect 7120 -1465 12620 -1420
rect 7120 -1585 7130 -1465
rect 7250 -1585 7305 -1465
rect 7425 -1585 7470 -1465
rect 7590 -1585 7635 -1465
rect 7755 -1585 7800 -1465
rect 7920 -1585 7975 -1465
rect 8095 -1585 8140 -1465
rect 8260 -1585 8305 -1465
rect 8425 -1585 8470 -1465
rect 8590 -1585 8645 -1465
rect 8765 -1585 8810 -1465
rect 8930 -1585 8975 -1465
rect 9095 -1585 9140 -1465
rect 9260 -1585 9315 -1465
rect 9435 -1585 9480 -1465
rect 9600 -1585 9645 -1465
rect 9765 -1585 9810 -1465
rect 9930 -1585 9985 -1465
rect 10105 -1585 10150 -1465
rect 10270 -1585 10315 -1465
rect 10435 -1585 10480 -1465
rect 10600 -1585 10655 -1465
rect 10775 -1585 10820 -1465
rect 10940 -1585 10985 -1465
rect 11105 -1585 11150 -1465
rect 11270 -1585 11325 -1465
rect 11445 -1585 11490 -1465
rect 11610 -1585 11655 -1465
rect 11775 -1585 11820 -1465
rect 11940 -1585 11995 -1465
rect 12115 -1585 12160 -1465
rect 12280 -1585 12325 -1465
rect 12445 -1585 12490 -1465
rect 12610 -1585 12620 -1465
rect 7120 -1630 12620 -1585
rect 7120 -1750 7130 -1630
rect 7250 -1750 7305 -1630
rect 7425 -1750 7470 -1630
rect 7590 -1750 7635 -1630
rect 7755 -1750 7800 -1630
rect 7920 -1750 7975 -1630
rect 8095 -1750 8140 -1630
rect 8260 -1750 8305 -1630
rect 8425 -1750 8470 -1630
rect 8590 -1750 8645 -1630
rect 8765 -1750 8810 -1630
rect 8930 -1750 8975 -1630
rect 9095 -1750 9140 -1630
rect 9260 -1750 9315 -1630
rect 9435 -1750 9480 -1630
rect 9600 -1750 9645 -1630
rect 9765 -1750 9810 -1630
rect 9930 -1750 9985 -1630
rect 10105 -1750 10150 -1630
rect 10270 -1750 10315 -1630
rect 10435 -1750 10480 -1630
rect 10600 -1750 10655 -1630
rect 10775 -1750 10820 -1630
rect 10940 -1750 10985 -1630
rect 11105 -1750 11150 -1630
rect 11270 -1750 11325 -1630
rect 11445 -1750 11490 -1630
rect 11610 -1750 11655 -1630
rect 11775 -1750 11820 -1630
rect 11940 -1750 11995 -1630
rect 12115 -1750 12160 -1630
rect 12280 -1750 12325 -1630
rect 12445 -1750 12490 -1630
rect 12610 -1750 12620 -1630
rect 7120 -1795 12620 -1750
rect 7120 -1915 7130 -1795
rect 7250 -1915 7305 -1795
rect 7425 -1915 7470 -1795
rect 7590 -1915 7635 -1795
rect 7755 -1915 7800 -1795
rect 7920 -1915 7975 -1795
rect 8095 -1915 8140 -1795
rect 8260 -1915 8305 -1795
rect 8425 -1915 8470 -1795
rect 8590 -1915 8645 -1795
rect 8765 -1915 8810 -1795
rect 8930 -1915 8975 -1795
rect 9095 -1915 9140 -1795
rect 9260 -1915 9315 -1795
rect 9435 -1915 9480 -1795
rect 9600 -1915 9645 -1795
rect 9765 -1915 9810 -1795
rect 9930 -1915 9985 -1795
rect 10105 -1915 10150 -1795
rect 10270 -1915 10315 -1795
rect 10435 -1915 10480 -1795
rect 10600 -1915 10655 -1795
rect 10775 -1915 10820 -1795
rect 10940 -1915 10985 -1795
rect 11105 -1915 11150 -1795
rect 11270 -1915 11325 -1795
rect 11445 -1915 11490 -1795
rect 11610 -1915 11655 -1795
rect 11775 -1915 11820 -1795
rect 11940 -1915 11995 -1795
rect 12115 -1915 12160 -1795
rect 12280 -1915 12325 -1795
rect 12445 -1915 12490 -1795
rect 12610 -1915 12620 -1795
rect 7120 -1970 12620 -1915
rect 7120 -2090 7130 -1970
rect 7250 -2090 7305 -1970
rect 7425 -2090 7470 -1970
rect 7590 -2090 7635 -1970
rect 7755 -2090 7800 -1970
rect 7920 -2090 7975 -1970
rect 8095 -2090 8140 -1970
rect 8260 -2090 8305 -1970
rect 8425 -2090 8470 -1970
rect 8590 -2090 8645 -1970
rect 8765 -2090 8810 -1970
rect 8930 -2090 8975 -1970
rect 9095 -2090 9140 -1970
rect 9260 -2090 9315 -1970
rect 9435 -2090 9480 -1970
rect 9600 -2090 9645 -1970
rect 9765 -2090 9810 -1970
rect 9930 -2090 9985 -1970
rect 10105 -2090 10150 -1970
rect 10270 -2090 10315 -1970
rect 10435 -2090 10480 -1970
rect 10600 -2090 10655 -1970
rect 10775 -2090 10820 -1970
rect 10940 -2090 10985 -1970
rect 11105 -2090 11150 -1970
rect 11270 -2090 11325 -1970
rect 11445 -2090 11490 -1970
rect 11610 -2090 11655 -1970
rect 11775 -2090 11820 -1970
rect 11940 -2090 11995 -1970
rect 12115 -2090 12160 -1970
rect 12280 -2090 12325 -1970
rect 12445 -2090 12490 -1970
rect 12610 -2090 12620 -1970
rect 7120 -2135 12620 -2090
rect 7120 -2255 7130 -2135
rect 7250 -2255 7305 -2135
rect 7425 -2255 7470 -2135
rect 7590 -2255 7635 -2135
rect 7755 -2255 7800 -2135
rect 7920 -2255 7975 -2135
rect 8095 -2255 8140 -2135
rect 8260 -2255 8305 -2135
rect 8425 -2255 8470 -2135
rect 8590 -2255 8645 -2135
rect 8765 -2255 8810 -2135
rect 8930 -2255 8975 -2135
rect 9095 -2255 9140 -2135
rect 9260 -2255 9315 -2135
rect 9435 -2255 9480 -2135
rect 9600 -2255 9645 -2135
rect 9765 -2255 9810 -2135
rect 9930 -2255 9985 -2135
rect 10105 -2255 10150 -2135
rect 10270 -2255 10315 -2135
rect 10435 -2255 10480 -2135
rect 10600 -2255 10655 -2135
rect 10775 -2255 10820 -2135
rect 10940 -2255 10985 -2135
rect 11105 -2255 11150 -2135
rect 11270 -2255 11325 -2135
rect 11445 -2255 11490 -2135
rect 11610 -2255 11655 -2135
rect 11775 -2255 11820 -2135
rect 11940 -2255 11995 -2135
rect 12115 -2255 12160 -2135
rect 12280 -2255 12325 -2135
rect 12445 -2255 12490 -2135
rect 12610 -2255 12620 -2135
rect 7120 -2300 12620 -2255
rect 7120 -2420 7130 -2300
rect 7250 -2420 7305 -2300
rect 7425 -2420 7470 -2300
rect 7590 -2420 7635 -2300
rect 7755 -2420 7800 -2300
rect 7920 -2420 7975 -2300
rect 8095 -2420 8140 -2300
rect 8260 -2420 8305 -2300
rect 8425 -2420 8470 -2300
rect 8590 -2420 8645 -2300
rect 8765 -2420 8810 -2300
rect 8930 -2420 8975 -2300
rect 9095 -2420 9140 -2300
rect 9260 -2420 9315 -2300
rect 9435 -2420 9480 -2300
rect 9600 -2420 9645 -2300
rect 9765 -2420 9810 -2300
rect 9930 -2420 9985 -2300
rect 10105 -2420 10150 -2300
rect 10270 -2420 10315 -2300
rect 10435 -2420 10480 -2300
rect 10600 -2420 10655 -2300
rect 10775 -2420 10820 -2300
rect 10940 -2420 10985 -2300
rect 11105 -2420 11150 -2300
rect 11270 -2420 11325 -2300
rect 11445 -2420 11490 -2300
rect 11610 -2420 11655 -2300
rect 11775 -2420 11820 -2300
rect 11940 -2420 11995 -2300
rect 12115 -2420 12160 -2300
rect 12280 -2420 12325 -2300
rect 12445 -2420 12490 -2300
rect 12610 -2420 12620 -2300
rect 7120 -2465 12620 -2420
rect 7120 -2585 7130 -2465
rect 7250 -2585 7305 -2465
rect 7425 -2585 7470 -2465
rect 7590 -2585 7635 -2465
rect 7755 -2585 7800 -2465
rect 7920 -2585 7975 -2465
rect 8095 -2585 8140 -2465
rect 8260 -2585 8305 -2465
rect 8425 -2585 8470 -2465
rect 8590 -2585 8645 -2465
rect 8765 -2585 8810 -2465
rect 8930 -2585 8975 -2465
rect 9095 -2585 9140 -2465
rect 9260 -2585 9315 -2465
rect 9435 -2585 9480 -2465
rect 9600 -2585 9645 -2465
rect 9765 -2585 9810 -2465
rect 9930 -2585 9985 -2465
rect 10105 -2585 10150 -2465
rect 10270 -2585 10315 -2465
rect 10435 -2585 10480 -2465
rect 10600 -2585 10655 -2465
rect 10775 -2585 10820 -2465
rect 10940 -2585 10985 -2465
rect 11105 -2585 11150 -2465
rect 11270 -2585 11325 -2465
rect 11445 -2585 11490 -2465
rect 11610 -2585 11655 -2465
rect 11775 -2585 11820 -2465
rect 11940 -2585 11995 -2465
rect 12115 -2585 12160 -2465
rect 12280 -2585 12325 -2465
rect 12445 -2585 12490 -2465
rect 12610 -2585 12620 -2465
rect 7120 -2640 12620 -2585
rect 7120 -2760 7130 -2640
rect 7250 -2760 7305 -2640
rect 7425 -2760 7470 -2640
rect 7590 -2760 7635 -2640
rect 7755 -2760 7800 -2640
rect 7920 -2760 7975 -2640
rect 8095 -2760 8140 -2640
rect 8260 -2760 8305 -2640
rect 8425 -2760 8470 -2640
rect 8590 -2760 8645 -2640
rect 8765 -2760 8810 -2640
rect 8930 -2760 8975 -2640
rect 9095 -2760 9140 -2640
rect 9260 -2760 9315 -2640
rect 9435 -2760 9480 -2640
rect 9600 -2760 9645 -2640
rect 9765 -2760 9810 -2640
rect 9930 -2760 9985 -2640
rect 10105 -2760 10150 -2640
rect 10270 -2760 10315 -2640
rect 10435 -2760 10480 -2640
rect 10600 -2760 10655 -2640
rect 10775 -2760 10820 -2640
rect 10940 -2760 10985 -2640
rect 11105 -2760 11150 -2640
rect 11270 -2760 11325 -2640
rect 11445 -2760 11490 -2640
rect 11610 -2760 11655 -2640
rect 11775 -2760 11820 -2640
rect 11940 -2760 11995 -2640
rect 12115 -2760 12160 -2640
rect 12280 -2760 12325 -2640
rect 12445 -2760 12490 -2640
rect 12610 -2760 12620 -2640
rect 7120 -2805 12620 -2760
rect 7120 -2925 7130 -2805
rect 7250 -2925 7305 -2805
rect 7425 -2925 7470 -2805
rect 7590 -2925 7635 -2805
rect 7755 -2925 7800 -2805
rect 7920 -2925 7975 -2805
rect 8095 -2925 8140 -2805
rect 8260 -2925 8305 -2805
rect 8425 -2925 8470 -2805
rect 8590 -2925 8645 -2805
rect 8765 -2925 8810 -2805
rect 8930 -2925 8975 -2805
rect 9095 -2925 9140 -2805
rect 9260 -2925 9315 -2805
rect 9435 -2925 9480 -2805
rect 9600 -2925 9645 -2805
rect 9765 -2925 9810 -2805
rect 9930 -2925 9985 -2805
rect 10105 -2925 10150 -2805
rect 10270 -2925 10315 -2805
rect 10435 -2925 10480 -2805
rect 10600 -2925 10655 -2805
rect 10775 -2925 10820 -2805
rect 10940 -2925 10985 -2805
rect 11105 -2925 11150 -2805
rect 11270 -2925 11325 -2805
rect 11445 -2925 11490 -2805
rect 11610 -2925 11655 -2805
rect 11775 -2925 11820 -2805
rect 11940 -2925 11995 -2805
rect 12115 -2925 12160 -2805
rect 12280 -2925 12325 -2805
rect 12445 -2925 12490 -2805
rect 12610 -2925 12620 -2805
rect 7120 -2970 12620 -2925
rect 7120 -3090 7130 -2970
rect 7250 -3090 7305 -2970
rect 7425 -3090 7470 -2970
rect 7590 -3090 7635 -2970
rect 7755 -3090 7800 -2970
rect 7920 -3090 7975 -2970
rect 8095 -3090 8140 -2970
rect 8260 -3090 8305 -2970
rect 8425 -3090 8470 -2970
rect 8590 -3090 8645 -2970
rect 8765 -3090 8810 -2970
rect 8930 -3090 8975 -2970
rect 9095 -3090 9140 -2970
rect 9260 -3090 9315 -2970
rect 9435 -3090 9480 -2970
rect 9600 -3090 9645 -2970
rect 9765 -3090 9810 -2970
rect 9930 -3090 9985 -2970
rect 10105 -3090 10150 -2970
rect 10270 -3090 10315 -2970
rect 10435 -3090 10480 -2970
rect 10600 -3090 10655 -2970
rect 10775 -3090 10820 -2970
rect 10940 -3090 10985 -2970
rect 11105 -3090 11150 -2970
rect 11270 -3090 11325 -2970
rect 11445 -3090 11490 -2970
rect 11610 -3090 11655 -2970
rect 11775 -3090 11820 -2970
rect 11940 -3090 11995 -2970
rect 12115 -3090 12160 -2970
rect 12280 -3090 12325 -2970
rect 12445 -3090 12490 -2970
rect 12610 -3090 12620 -2970
rect 7120 -3135 12620 -3090
rect 7120 -3255 7130 -3135
rect 7250 -3255 7305 -3135
rect 7425 -3255 7470 -3135
rect 7590 -3255 7635 -3135
rect 7755 -3255 7800 -3135
rect 7920 -3255 7975 -3135
rect 8095 -3255 8140 -3135
rect 8260 -3255 8305 -3135
rect 8425 -3255 8470 -3135
rect 8590 -3255 8645 -3135
rect 8765 -3255 8810 -3135
rect 8930 -3255 8975 -3135
rect 9095 -3255 9140 -3135
rect 9260 -3255 9315 -3135
rect 9435 -3255 9480 -3135
rect 9600 -3255 9645 -3135
rect 9765 -3255 9810 -3135
rect 9930 -3255 9985 -3135
rect 10105 -3255 10150 -3135
rect 10270 -3255 10315 -3135
rect 10435 -3255 10480 -3135
rect 10600 -3255 10655 -3135
rect 10775 -3255 10820 -3135
rect 10940 -3255 10985 -3135
rect 11105 -3255 11150 -3135
rect 11270 -3255 11325 -3135
rect 11445 -3255 11490 -3135
rect 11610 -3255 11655 -3135
rect 11775 -3255 11820 -3135
rect 11940 -3255 11995 -3135
rect 12115 -3255 12160 -3135
rect 12280 -3255 12325 -3135
rect 12445 -3255 12490 -3135
rect 12610 -3255 12620 -3135
rect 7120 -3310 12620 -3255
rect 7120 -3430 7130 -3310
rect 7250 -3430 7305 -3310
rect 7425 -3430 7470 -3310
rect 7590 -3430 7635 -3310
rect 7755 -3430 7800 -3310
rect 7920 -3430 7975 -3310
rect 8095 -3430 8140 -3310
rect 8260 -3430 8305 -3310
rect 8425 -3430 8470 -3310
rect 8590 -3430 8645 -3310
rect 8765 -3430 8810 -3310
rect 8930 -3430 8975 -3310
rect 9095 -3430 9140 -3310
rect 9260 -3430 9315 -3310
rect 9435 -3430 9480 -3310
rect 9600 -3430 9645 -3310
rect 9765 -3430 9810 -3310
rect 9930 -3430 9985 -3310
rect 10105 -3430 10150 -3310
rect 10270 -3430 10315 -3310
rect 10435 -3430 10480 -3310
rect 10600 -3430 10655 -3310
rect 10775 -3430 10820 -3310
rect 10940 -3430 10985 -3310
rect 11105 -3430 11150 -3310
rect 11270 -3430 11325 -3310
rect 11445 -3430 11490 -3310
rect 11610 -3430 11655 -3310
rect 11775 -3430 11820 -3310
rect 11940 -3430 11995 -3310
rect 12115 -3430 12160 -3310
rect 12280 -3430 12325 -3310
rect 12445 -3430 12490 -3310
rect 12610 -3430 12620 -3310
rect 7120 -3475 12620 -3430
rect 7120 -3595 7130 -3475
rect 7250 -3595 7305 -3475
rect 7425 -3595 7470 -3475
rect 7590 -3595 7635 -3475
rect 7755 -3595 7800 -3475
rect 7920 -3595 7975 -3475
rect 8095 -3595 8140 -3475
rect 8260 -3595 8305 -3475
rect 8425 -3595 8470 -3475
rect 8590 -3595 8645 -3475
rect 8765 -3595 8810 -3475
rect 8930 -3595 8975 -3475
rect 9095 -3595 9140 -3475
rect 9260 -3595 9315 -3475
rect 9435 -3595 9480 -3475
rect 9600 -3595 9645 -3475
rect 9765 -3595 9810 -3475
rect 9930 -3595 9985 -3475
rect 10105 -3595 10150 -3475
rect 10270 -3595 10315 -3475
rect 10435 -3595 10480 -3475
rect 10600 -3595 10655 -3475
rect 10775 -3595 10820 -3475
rect 10940 -3595 10985 -3475
rect 11105 -3595 11150 -3475
rect 11270 -3595 11325 -3475
rect 11445 -3595 11490 -3475
rect 11610 -3595 11655 -3475
rect 11775 -3595 11820 -3475
rect 11940 -3595 11995 -3475
rect 12115 -3595 12160 -3475
rect 12280 -3595 12325 -3475
rect 12445 -3595 12490 -3475
rect 12610 -3595 12620 -3475
rect 7120 -3640 12620 -3595
rect 7120 -3760 7130 -3640
rect 7250 -3760 7305 -3640
rect 7425 -3760 7470 -3640
rect 7590 -3760 7635 -3640
rect 7755 -3760 7800 -3640
rect 7920 -3760 7975 -3640
rect 8095 -3760 8140 -3640
rect 8260 -3760 8305 -3640
rect 8425 -3760 8470 -3640
rect 8590 -3760 8645 -3640
rect 8765 -3760 8810 -3640
rect 8930 -3760 8975 -3640
rect 9095 -3760 9140 -3640
rect 9260 -3760 9315 -3640
rect 9435 -3760 9480 -3640
rect 9600 -3760 9645 -3640
rect 9765 -3760 9810 -3640
rect 9930 -3760 9985 -3640
rect 10105 -3760 10150 -3640
rect 10270 -3760 10315 -3640
rect 10435 -3760 10480 -3640
rect 10600 -3760 10655 -3640
rect 10775 -3760 10820 -3640
rect 10940 -3760 10985 -3640
rect 11105 -3760 11150 -3640
rect 11270 -3760 11325 -3640
rect 11445 -3760 11490 -3640
rect 11610 -3760 11655 -3640
rect 11775 -3760 11820 -3640
rect 11940 -3760 11995 -3640
rect 12115 -3760 12160 -3640
rect 12280 -3760 12325 -3640
rect 12445 -3760 12490 -3640
rect 12610 -3760 12620 -3640
rect 7120 -3805 12620 -3760
rect 7120 -3925 7130 -3805
rect 7250 -3925 7305 -3805
rect 7425 -3925 7470 -3805
rect 7590 -3925 7635 -3805
rect 7755 -3925 7800 -3805
rect 7920 -3925 7975 -3805
rect 8095 -3925 8140 -3805
rect 8260 -3925 8305 -3805
rect 8425 -3925 8470 -3805
rect 8590 -3925 8645 -3805
rect 8765 -3925 8810 -3805
rect 8930 -3925 8975 -3805
rect 9095 -3925 9140 -3805
rect 9260 -3925 9315 -3805
rect 9435 -3925 9480 -3805
rect 9600 -3925 9645 -3805
rect 9765 -3925 9810 -3805
rect 9930 -3925 9985 -3805
rect 10105 -3925 10150 -3805
rect 10270 -3925 10315 -3805
rect 10435 -3925 10480 -3805
rect 10600 -3925 10655 -3805
rect 10775 -3925 10820 -3805
rect 10940 -3925 10985 -3805
rect 11105 -3925 11150 -3805
rect 11270 -3925 11325 -3805
rect 11445 -3925 11490 -3805
rect 11610 -3925 11655 -3805
rect 11775 -3925 11820 -3805
rect 11940 -3925 11995 -3805
rect 12115 -3925 12160 -3805
rect 12280 -3925 12325 -3805
rect 12445 -3925 12490 -3805
rect 12610 -3925 12620 -3805
rect 7120 -3980 12620 -3925
rect 7120 -4100 7130 -3980
rect 7250 -4100 7305 -3980
rect 7425 -4100 7470 -3980
rect 7590 -4100 7635 -3980
rect 7755 -4100 7800 -3980
rect 7920 -4100 7975 -3980
rect 8095 -4100 8140 -3980
rect 8260 -4100 8305 -3980
rect 8425 -4100 8470 -3980
rect 8590 -4100 8645 -3980
rect 8765 -4100 8810 -3980
rect 8930 -4100 8975 -3980
rect 9095 -4100 9140 -3980
rect 9260 -4100 9315 -3980
rect 9435 -4100 9480 -3980
rect 9600 -4100 9645 -3980
rect 9765 -4100 9810 -3980
rect 9930 -4100 9985 -3980
rect 10105 -4100 10150 -3980
rect 10270 -4100 10315 -3980
rect 10435 -4100 10480 -3980
rect 10600 -4100 10655 -3980
rect 10775 -4100 10820 -3980
rect 10940 -4100 10985 -3980
rect 11105 -4100 11150 -3980
rect 11270 -4100 11325 -3980
rect 11445 -4100 11490 -3980
rect 11610 -4100 11655 -3980
rect 11775 -4100 11820 -3980
rect 11940 -4100 11995 -3980
rect 12115 -4100 12160 -3980
rect 12280 -4100 12325 -3980
rect 12445 -4100 12490 -3980
rect 12610 -4100 12620 -3980
rect 7120 -4110 12620 -4100
rect 12810 1380 18310 1390
rect 12810 1260 12820 1380
rect 12940 1260 12995 1380
rect 13115 1260 13160 1380
rect 13280 1260 13325 1380
rect 13445 1260 13490 1380
rect 13610 1260 13665 1380
rect 13785 1260 13830 1380
rect 13950 1260 13995 1380
rect 14115 1260 14160 1380
rect 14280 1260 14335 1380
rect 14455 1260 14500 1380
rect 14620 1260 14665 1380
rect 14785 1260 14830 1380
rect 14950 1260 15005 1380
rect 15125 1260 15170 1380
rect 15290 1260 15335 1380
rect 15455 1260 15500 1380
rect 15620 1260 15675 1380
rect 15795 1260 15840 1380
rect 15960 1260 16005 1380
rect 16125 1260 16170 1380
rect 16290 1260 16345 1380
rect 16465 1260 16510 1380
rect 16630 1260 16675 1380
rect 16795 1260 16840 1380
rect 16960 1260 17015 1380
rect 17135 1260 17180 1380
rect 17300 1260 17345 1380
rect 17465 1260 17510 1380
rect 17630 1260 17685 1380
rect 17805 1260 17850 1380
rect 17970 1260 18015 1380
rect 18135 1260 18180 1380
rect 18300 1260 18310 1380
rect 12810 1215 18310 1260
rect 12810 1095 12820 1215
rect 12940 1095 12995 1215
rect 13115 1095 13160 1215
rect 13280 1095 13325 1215
rect 13445 1095 13490 1215
rect 13610 1095 13665 1215
rect 13785 1095 13830 1215
rect 13950 1095 13995 1215
rect 14115 1095 14160 1215
rect 14280 1095 14335 1215
rect 14455 1095 14500 1215
rect 14620 1095 14665 1215
rect 14785 1095 14830 1215
rect 14950 1095 15005 1215
rect 15125 1095 15170 1215
rect 15290 1095 15335 1215
rect 15455 1095 15500 1215
rect 15620 1095 15675 1215
rect 15795 1095 15840 1215
rect 15960 1095 16005 1215
rect 16125 1095 16170 1215
rect 16290 1095 16345 1215
rect 16465 1095 16510 1215
rect 16630 1095 16675 1215
rect 16795 1095 16840 1215
rect 16960 1095 17015 1215
rect 17135 1095 17180 1215
rect 17300 1095 17345 1215
rect 17465 1095 17510 1215
rect 17630 1095 17685 1215
rect 17805 1095 17850 1215
rect 17970 1095 18015 1215
rect 18135 1095 18180 1215
rect 18300 1095 18310 1215
rect 12810 1050 18310 1095
rect 12810 930 12820 1050
rect 12940 930 12995 1050
rect 13115 930 13160 1050
rect 13280 930 13325 1050
rect 13445 930 13490 1050
rect 13610 930 13665 1050
rect 13785 930 13830 1050
rect 13950 930 13995 1050
rect 14115 930 14160 1050
rect 14280 930 14335 1050
rect 14455 930 14500 1050
rect 14620 930 14665 1050
rect 14785 930 14830 1050
rect 14950 930 15005 1050
rect 15125 930 15170 1050
rect 15290 930 15335 1050
rect 15455 930 15500 1050
rect 15620 930 15675 1050
rect 15795 930 15840 1050
rect 15960 930 16005 1050
rect 16125 930 16170 1050
rect 16290 930 16345 1050
rect 16465 930 16510 1050
rect 16630 930 16675 1050
rect 16795 930 16840 1050
rect 16960 930 17015 1050
rect 17135 930 17180 1050
rect 17300 930 17345 1050
rect 17465 930 17510 1050
rect 17630 930 17685 1050
rect 17805 930 17850 1050
rect 17970 930 18015 1050
rect 18135 930 18180 1050
rect 18300 930 18310 1050
rect 12810 885 18310 930
rect 12810 765 12820 885
rect 12940 765 12995 885
rect 13115 765 13160 885
rect 13280 765 13325 885
rect 13445 765 13490 885
rect 13610 765 13665 885
rect 13785 765 13830 885
rect 13950 765 13995 885
rect 14115 765 14160 885
rect 14280 765 14335 885
rect 14455 765 14500 885
rect 14620 765 14665 885
rect 14785 765 14830 885
rect 14950 765 15005 885
rect 15125 765 15170 885
rect 15290 765 15335 885
rect 15455 765 15500 885
rect 15620 765 15675 885
rect 15795 765 15840 885
rect 15960 765 16005 885
rect 16125 765 16170 885
rect 16290 765 16345 885
rect 16465 765 16510 885
rect 16630 765 16675 885
rect 16795 765 16840 885
rect 16960 765 17015 885
rect 17135 765 17180 885
rect 17300 765 17345 885
rect 17465 765 17510 885
rect 17630 765 17685 885
rect 17805 765 17850 885
rect 17970 765 18015 885
rect 18135 765 18180 885
rect 18300 765 18310 885
rect 12810 710 18310 765
rect 12810 590 12820 710
rect 12940 590 12995 710
rect 13115 590 13160 710
rect 13280 590 13325 710
rect 13445 590 13490 710
rect 13610 590 13665 710
rect 13785 590 13830 710
rect 13950 590 13995 710
rect 14115 590 14160 710
rect 14280 590 14335 710
rect 14455 590 14500 710
rect 14620 590 14665 710
rect 14785 590 14830 710
rect 14950 590 15005 710
rect 15125 590 15170 710
rect 15290 590 15335 710
rect 15455 590 15500 710
rect 15620 590 15675 710
rect 15795 590 15840 710
rect 15960 590 16005 710
rect 16125 590 16170 710
rect 16290 590 16345 710
rect 16465 590 16510 710
rect 16630 590 16675 710
rect 16795 590 16840 710
rect 16960 590 17015 710
rect 17135 590 17180 710
rect 17300 590 17345 710
rect 17465 590 17510 710
rect 17630 590 17685 710
rect 17805 590 17850 710
rect 17970 590 18015 710
rect 18135 590 18180 710
rect 18300 590 18310 710
rect 12810 545 18310 590
rect 12810 425 12820 545
rect 12940 425 12995 545
rect 13115 425 13160 545
rect 13280 425 13325 545
rect 13445 425 13490 545
rect 13610 425 13665 545
rect 13785 425 13830 545
rect 13950 425 13995 545
rect 14115 425 14160 545
rect 14280 425 14335 545
rect 14455 425 14500 545
rect 14620 425 14665 545
rect 14785 425 14830 545
rect 14950 425 15005 545
rect 15125 425 15170 545
rect 15290 425 15335 545
rect 15455 425 15500 545
rect 15620 425 15675 545
rect 15795 425 15840 545
rect 15960 425 16005 545
rect 16125 425 16170 545
rect 16290 425 16345 545
rect 16465 425 16510 545
rect 16630 425 16675 545
rect 16795 425 16840 545
rect 16960 425 17015 545
rect 17135 425 17180 545
rect 17300 425 17345 545
rect 17465 425 17510 545
rect 17630 425 17685 545
rect 17805 425 17850 545
rect 17970 425 18015 545
rect 18135 425 18180 545
rect 18300 425 18310 545
rect 12810 380 18310 425
rect 12810 260 12820 380
rect 12940 260 12995 380
rect 13115 260 13160 380
rect 13280 260 13325 380
rect 13445 260 13490 380
rect 13610 260 13665 380
rect 13785 260 13830 380
rect 13950 260 13995 380
rect 14115 260 14160 380
rect 14280 260 14335 380
rect 14455 260 14500 380
rect 14620 260 14665 380
rect 14785 260 14830 380
rect 14950 260 15005 380
rect 15125 260 15170 380
rect 15290 260 15335 380
rect 15455 260 15500 380
rect 15620 260 15675 380
rect 15795 260 15840 380
rect 15960 260 16005 380
rect 16125 260 16170 380
rect 16290 260 16345 380
rect 16465 260 16510 380
rect 16630 260 16675 380
rect 16795 260 16840 380
rect 16960 260 17015 380
rect 17135 260 17180 380
rect 17300 260 17345 380
rect 17465 260 17510 380
rect 17630 260 17685 380
rect 17805 260 17850 380
rect 17970 260 18015 380
rect 18135 260 18180 380
rect 18300 260 18310 380
rect 12810 215 18310 260
rect 12810 95 12820 215
rect 12940 95 12995 215
rect 13115 95 13160 215
rect 13280 95 13325 215
rect 13445 95 13490 215
rect 13610 95 13665 215
rect 13785 95 13830 215
rect 13950 95 13995 215
rect 14115 95 14160 215
rect 14280 95 14335 215
rect 14455 95 14500 215
rect 14620 95 14665 215
rect 14785 95 14830 215
rect 14950 95 15005 215
rect 15125 95 15170 215
rect 15290 95 15335 215
rect 15455 95 15500 215
rect 15620 95 15675 215
rect 15795 95 15840 215
rect 15960 95 16005 215
rect 16125 95 16170 215
rect 16290 95 16345 215
rect 16465 95 16510 215
rect 16630 95 16675 215
rect 16795 95 16840 215
rect 16960 95 17015 215
rect 17135 95 17180 215
rect 17300 95 17345 215
rect 17465 95 17510 215
rect 17630 95 17685 215
rect 17805 95 17850 215
rect 17970 95 18015 215
rect 18135 95 18180 215
rect 18300 95 18310 215
rect 12810 40 18310 95
rect 12810 -80 12820 40
rect 12940 -80 12995 40
rect 13115 -80 13160 40
rect 13280 -80 13325 40
rect 13445 -80 13490 40
rect 13610 -80 13665 40
rect 13785 -80 13830 40
rect 13950 -80 13995 40
rect 14115 -80 14160 40
rect 14280 -80 14335 40
rect 14455 -80 14500 40
rect 14620 -80 14665 40
rect 14785 -80 14830 40
rect 14950 -80 15005 40
rect 15125 -80 15170 40
rect 15290 -80 15335 40
rect 15455 -80 15500 40
rect 15620 -80 15675 40
rect 15795 -80 15840 40
rect 15960 -80 16005 40
rect 16125 -80 16170 40
rect 16290 -80 16345 40
rect 16465 -80 16510 40
rect 16630 -80 16675 40
rect 16795 -80 16840 40
rect 16960 -80 17015 40
rect 17135 -80 17180 40
rect 17300 -80 17345 40
rect 17465 -80 17510 40
rect 17630 -80 17685 40
rect 17805 -80 17850 40
rect 17970 -80 18015 40
rect 18135 -80 18180 40
rect 18300 -80 18310 40
rect 12810 -125 18310 -80
rect 12810 -245 12820 -125
rect 12940 -245 12995 -125
rect 13115 -245 13160 -125
rect 13280 -245 13325 -125
rect 13445 -245 13490 -125
rect 13610 -245 13665 -125
rect 13785 -245 13830 -125
rect 13950 -245 13995 -125
rect 14115 -245 14160 -125
rect 14280 -245 14335 -125
rect 14455 -245 14500 -125
rect 14620 -245 14665 -125
rect 14785 -245 14830 -125
rect 14950 -245 15005 -125
rect 15125 -245 15170 -125
rect 15290 -245 15335 -125
rect 15455 -245 15500 -125
rect 15620 -245 15675 -125
rect 15795 -245 15840 -125
rect 15960 -245 16005 -125
rect 16125 -245 16170 -125
rect 16290 -245 16345 -125
rect 16465 -245 16510 -125
rect 16630 -245 16675 -125
rect 16795 -245 16840 -125
rect 16960 -245 17015 -125
rect 17135 -245 17180 -125
rect 17300 -245 17345 -125
rect 17465 -245 17510 -125
rect 17630 -245 17685 -125
rect 17805 -245 17850 -125
rect 17970 -245 18015 -125
rect 18135 -245 18180 -125
rect 18300 -245 18310 -125
rect 12810 -290 18310 -245
rect 12810 -410 12820 -290
rect 12940 -410 12995 -290
rect 13115 -410 13160 -290
rect 13280 -410 13325 -290
rect 13445 -410 13490 -290
rect 13610 -410 13665 -290
rect 13785 -410 13830 -290
rect 13950 -410 13995 -290
rect 14115 -410 14160 -290
rect 14280 -410 14335 -290
rect 14455 -410 14500 -290
rect 14620 -410 14665 -290
rect 14785 -410 14830 -290
rect 14950 -410 15005 -290
rect 15125 -410 15170 -290
rect 15290 -410 15335 -290
rect 15455 -410 15500 -290
rect 15620 -410 15675 -290
rect 15795 -410 15840 -290
rect 15960 -410 16005 -290
rect 16125 -410 16170 -290
rect 16290 -410 16345 -290
rect 16465 -410 16510 -290
rect 16630 -410 16675 -290
rect 16795 -410 16840 -290
rect 16960 -410 17015 -290
rect 17135 -410 17180 -290
rect 17300 -410 17345 -290
rect 17465 -410 17510 -290
rect 17630 -410 17685 -290
rect 17805 -410 17850 -290
rect 17970 -410 18015 -290
rect 18135 -410 18180 -290
rect 18300 -410 18310 -290
rect 12810 -455 18310 -410
rect 12810 -575 12820 -455
rect 12940 -575 12995 -455
rect 13115 -575 13160 -455
rect 13280 -575 13325 -455
rect 13445 -575 13490 -455
rect 13610 -575 13665 -455
rect 13785 -575 13830 -455
rect 13950 -575 13995 -455
rect 14115 -575 14160 -455
rect 14280 -575 14335 -455
rect 14455 -575 14500 -455
rect 14620 -575 14665 -455
rect 14785 -575 14830 -455
rect 14950 -575 15005 -455
rect 15125 -575 15170 -455
rect 15290 -575 15335 -455
rect 15455 -575 15500 -455
rect 15620 -575 15675 -455
rect 15795 -575 15840 -455
rect 15960 -575 16005 -455
rect 16125 -575 16170 -455
rect 16290 -575 16345 -455
rect 16465 -575 16510 -455
rect 16630 -575 16675 -455
rect 16795 -575 16840 -455
rect 16960 -575 17015 -455
rect 17135 -575 17180 -455
rect 17300 -575 17345 -455
rect 17465 -575 17510 -455
rect 17630 -575 17685 -455
rect 17805 -575 17850 -455
rect 17970 -575 18015 -455
rect 18135 -575 18180 -455
rect 18300 -575 18310 -455
rect 12810 -630 18310 -575
rect 12810 -750 12820 -630
rect 12940 -750 12995 -630
rect 13115 -750 13160 -630
rect 13280 -750 13325 -630
rect 13445 -750 13490 -630
rect 13610 -750 13665 -630
rect 13785 -750 13830 -630
rect 13950 -750 13995 -630
rect 14115 -750 14160 -630
rect 14280 -750 14335 -630
rect 14455 -750 14500 -630
rect 14620 -750 14665 -630
rect 14785 -750 14830 -630
rect 14950 -750 15005 -630
rect 15125 -750 15170 -630
rect 15290 -750 15335 -630
rect 15455 -750 15500 -630
rect 15620 -750 15675 -630
rect 15795 -750 15840 -630
rect 15960 -750 16005 -630
rect 16125 -750 16170 -630
rect 16290 -750 16345 -630
rect 16465 -750 16510 -630
rect 16630 -750 16675 -630
rect 16795 -750 16840 -630
rect 16960 -750 17015 -630
rect 17135 -750 17180 -630
rect 17300 -750 17345 -630
rect 17465 -750 17510 -630
rect 17630 -750 17685 -630
rect 17805 -750 17850 -630
rect 17970 -750 18015 -630
rect 18135 -750 18180 -630
rect 18300 -750 18310 -630
rect 12810 -795 18310 -750
rect 12810 -915 12820 -795
rect 12940 -915 12995 -795
rect 13115 -915 13160 -795
rect 13280 -915 13325 -795
rect 13445 -915 13490 -795
rect 13610 -915 13665 -795
rect 13785 -915 13830 -795
rect 13950 -915 13995 -795
rect 14115 -915 14160 -795
rect 14280 -915 14335 -795
rect 14455 -915 14500 -795
rect 14620 -915 14665 -795
rect 14785 -915 14830 -795
rect 14950 -915 15005 -795
rect 15125 -915 15170 -795
rect 15290 -915 15335 -795
rect 15455 -915 15500 -795
rect 15620 -915 15675 -795
rect 15795 -915 15840 -795
rect 15960 -915 16005 -795
rect 16125 -915 16170 -795
rect 16290 -915 16345 -795
rect 16465 -915 16510 -795
rect 16630 -915 16675 -795
rect 16795 -915 16840 -795
rect 16960 -915 17015 -795
rect 17135 -915 17180 -795
rect 17300 -915 17345 -795
rect 17465 -915 17510 -795
rect 17630 -915 17685 -795
rect 17805 -915 17850 -795
rect 17970 -915 18015 -795
rect 18135 -915 18180 -795
rect 18300 -915 18310 -795
rect 12810 -960 18310 -915
rect 12810 -1080 12820 -960
rect 12940 -1080 12995 -960
rect 13115 -1080 13160 -960
rect 13280 -1080 13325 -960
rect 13445 -1080 13490 -960
rect 13610 -1080 13665 -960
rect 13785 -1080 13830 -960
rect 13950 -1080 13995 -960
rect 14115 -1080 14160 -960
rect 14280 -1080 14335 -960
rect 14455 -1080 14500 -960
rect 14620 -1080 14665 -960
rect 14785 -1080 14830 -960
rect 14950 -1080 15005 -960
rect 15125 -1080 15170 -960
rect 15290 -1080 15335 -960
rect 15455 -1080 15500 -960
rect 15620 -1080 15675 -960
rect 15795 -1080 15840 -960
rect 15960 -1080 16005 -960
rect 16125 -1080 16170 -960
rect 16290 -1080 16345 -960
rect 16465 -1080 16510 -960
rect 16630 -1080 16675 -960
rect 16795 -1080 16840 -960
rect 16960 -1080 17015 -960
rect 17135 -1080 17180 -960
rect 17300 -1080 17345 -960
rect 17465 -1080 17510 -960
rect 17630 -1080 17685 -960
rect 17805 -1080 17850 -960
rect 17970 -1080 18015 -960
rect 18135 -1080 18180 -960
rect 18300 -1080 18310 -960
rect 12810 -1125 18310 -1080
rect 12810 -1245 12820 -1125
rect 12940 -1245 12995 -1125
rect 13115 -1245 13160 -1125
rect 13280 -1245 13325 -1125
rect 13445 -1245 13490 -1125
rect 13610 -1245 13665 -1125
rect 13785 -1245 13830 -1125
rect 13950 -1245 13995 -1125
rect 14115 -1245 14160 -1125
rect 14280 -1245 14335 -1125
rect 14455 -1245 14500 -1125
rect 14620 -1245 14665 -1125
rect 14785 -1245 14830 -1125
rect 14950 -1245 15005 -1125
rect 15125 -1245 15170 -1125
rect 15290 -1245 15335 -1125
rect 15455 -1245 15500 -1125
rect 15620 -1245 15675 -1125
rect 15795 -1245 15840 -1125
rect 15960 -1245 16005 -1125
rect 16125 -1245 16170 -1125
rect 16290 -1245 16345 -1125
rect 16465 -1245 16510 -1125
rect 16630 -1245 16675 -1125
rect 16795 -1245 16840 -1125
rect 16960 -1245 17015 -1125
rect 17135 -1245 17180 -1125
rect 17300 -1245 17345 -1125
rect 17465 -1245 17510 -1125
rect 17630 -1245 17685 -1125
rect 17805 -1245 17850 -1125
rect 17970 -1245 18015 -1125
rect 18135 -1245 18180 -1125
rect 18300 -1245 18310 -1125
rect 12810 -1300 18310 -1245
rect 12810 -1420 12820 -1300
rect 12940 -1420 12995 -1300
rect 13115 -1420 13160 -1300
rect 13280 -1420 13325 -1300
rect 13445 -1420 13490 -1300
rect 13610 -1420 13665 -1300
rect 13785 -1420 13830 -1300
rect 13950 -1420 13995 -1300
rect 14115 -1420 14160 -1300
rect 14280 -1420 14335 -1300
rect 14455 -1420 14500 -1300
rect 14620 -1420 14665 -1300
rect 14785 -1420 14830 -1300
rect 14950 -1420 15005 -1300
rect 15125 -1420 15170 -1300
rect 15290 -1420 15335 -1300
rect 15455 -1420 15500 -1300
rect 15620 -1420 15675 -1300
rect 15795 -1420 15840 -1300
rect 15960 -1420 16005 -1300
rect 16125 -1420 16170 -1300
rect 16290 -1420 16345 -1300
rect 16465 -1420 16510 -1300
rect 16630 -1420 16675 -1300
rect 16795 -1420 16840 -1300
rect 16960 -1420 17015 -1300
rect 17135 -1420 17180 -1300
rect 17300 -1420 17345 -1300
rect 17465 -1420 17510 -1300
rect 17630 -1420 17685 -1300
rect 17805 -1420 17850 -1300
rect 17970 -1420 18015 -1300
rect 18135 -1420 18180 -1300
rect 18300 -1420 18310 -1300
rect 12810 -1465 18310 -1420
rect 12810 -1585 12820 -1465
rect 12940 -1585 12995 -1465
rect 13115 -1585 13160 -1465
rect 13280 -1585 13325 -1465
rect 13445 -1585 13490 -1465
rect 13610 -1585 13665 -1465
rect 13785 -1585 13830 -1465
rect 13950 -1585 13995 -1465
rect 14115 -1585 14160 -1465
rect 14280 -1585 14335 -1465
rect 14455 -1585 14500 -1465
rect 14620 -1585 14665 -1465
rect 14785 -1585 14830 -1465
rect 14950 -1585 15005 -1465
rect 15125 -1585 15170 -1465
rect 15290 -1585 15335 -1465
rect 15455 -1585 15500 -1465
rect 15620 -1585 15675 -1465
rect 15795 -1585 15840 -1465
rect 15960 -1585 16005 -1465
rect 16125 -1585 16170 -1465
rect 16290 -1585 16345 -1465
rect 16465 -1585 16510 -1465
rect 16630 -1585 16675 -1465
rect 16795 -1585 16840 -1465
rect 16960 -1585 17015 -1465
rect 17135 -1585 17180 -1465
rect 17300 -1585 17345 -1465
rect 17465 -1585 17510 -1465
rect 17630 -1585 17685 -1465
rect 17805 -1585 17850 -1465
rect 17970 -1585 18015 -1465
rect 18135 -1585 18180 -1465
rect 18300 -1585 18310 -1465
rect 12810 -1630 18310 -1585
rect 12810 -1750 12820 -1630
rect 12940 -1750 12995 -1630
rect 13115 -1750 13160 -1630
rect 13280 -1750 13325 -1630
rect 13445 -1750 13490 -1630
rect 13610 -1750 13665 -1630
rect 13785 -1750 13830 -1630
rect 13950 -1750 13995 -1630
rect 14115 -1750 14160 -1630
rect 14280 -1750 14335 -1630
rect 14455 -1750 14500 -1630
rect 14620 -1750 14665 -1630
rect 14785 -1750 14830 -1630
rect 14950 -1750 15005 -1630
rect 15125 -1750 15170 -1630
rect 15290 -1750 15335 -1630
rect 15455 -1750 15500 -1630
rect 15620 -1750 15675 -1630
rect 15795 -1750 15840 -1630
rect 15960 -1750 16005 -1630
rect 16125 -1750 16170 -1630
rect 16290 -1750 16345 -1630
rect 16465 -1750 16510 -1630
rect 16630 -1750 16675 -1630
rect 16795 -1750 16840 -1630
rect 16960 -1750 17015 -1630
rect 17135 -1750 17180 -1630
rect 17300 -1750 17345 -1630
rect 17465 -1750 17510 -1630
rect 17630 -1750 17685 -1630
rect 17805 -1750 17850 -1630
rect 17970 -1750 18015 -1630
rect 18135 -1750 18180 -1630
rect 18300 -1750 18310 -1630
rect 12810 -1795 18310 -1750
rect 12810 -1915 12820 -1795
rect 12940 -1915 12995 -1795
rect 13115 -1915 13160 -1795
rect 13280 -1915 13325 -1795
rect 13445 -1915 13490 -1795
rect 13610 -1915 13665 -1795
rect 13785 -1915 13830 -1795
rect 13950 -1915 13995 -1795
rect 14115 -1915 14160 -1795
rect 14280 -1915 14335 -1795
rect 14455 -1915 14500 -1795
rect 14620 -1915 14665 -1795
rect 14785 -1915 14830 -1795
rect 14950 -1915 15005 -1795
rect 15125 -1915 15170 -1795
rect 15290 -1915 15335 -1795
rect 15455 -1915 15500 -1795
rect 15620 -1915 15675 -1795
rect 15795 -1915 15840 -1795
rect 15960 -1915 16005 -1795
rect 16125 -1915 16170 -1795
rect 16290 -1915 16345 -1795
rect 16465 -1915 16510 -1795
rect 16630 -1915 16675 -1795
rect 16795 -1915 16840 -1795
rect 16960 -1915 17015 -1795
rect 17135 -1915 17180 -1795
rect 17300 -1915 17345 -1795
rect 17465 -1915 17510 -1795
rect 17630 -1915 17685 -1795
rect 17805 -1915 17850 -1795
rect 17970 -1915 18015 -1795
rect 18135 -1915 18180 -1795
rect 18300 -1915 18310 -1795
rect 12810 -1970 18310 -1915
rect 12810 -2090 12820 -1970
rect 12940 -2090 12995 -1970
rect 13115 -2090 13160 -1970
rect 13280 -2090 13325 -1970
rect 13445 -2090 13490 -1970
rect 13610 -2090 13665 -1970
rect 13785 -2090 13830 -1970
rect 13950 -2090 13995 -1970
rect 14115 -2090 14160 -1970
rect 14280 -2090 14335 -1970
rect 14455 -2090 14500 -1970
rect 14620 -2090 14665 -1970
rect 14785 -2090 14830 -1970
rect 14950 -2090 15005 -1970
rect 15125 -2090 15170 -1970
rect 15290 -2090 15335 -1970
rect 15455 -2090 15500 -1970
rect 15620 -2090 15675 -1970
rect 15795 -2090 15840 -1970
rect 15960 -2090 16005 -1970
rect 16125 -2090 16170 -1970
rect 16290 -2090 16345 -1970
rect 16465 -2090 16510 -1970
rect 16630 -2090 16675 -1970
rect 16795 -2090 16840 -1970
rect 16960 -2090 17015 -1970
rect 17135 -2090 17180 -1970
rect 17300 -2090 17345 -1970
rect 17465 -2090 17510 -1970
rect 17630 -2090 17685 -1970
rect 17805 -2090 17850 -1970
rect 17970 -2090 18015 -1970
rect 18135 -2090 18180 -1970
rect 18300 -2090 18310 -1970
rect 12810 -2135 18310 -2090
rect 12810 -2255 12820 -2135
rect 12940 -2255 12995 -2135
rect 13115 -2255 13160 -2135
rect 13280 -2255 13325 -2135
rect 13445 -2255 13490 -2135
rect 13610 -2255 13665 -2135
rect 13785 -2255 13830 -2135
rect 13950 -2255 13995 -2135
rect 14115 -2255 14160 -2135
rect 14280 -2255 14335 -2135
rect 14455 -2255 14500 -2135
rect 14620 -2255 14665 -2135
rect 14785 -2255 14830 -2135
rect 14950 -2255 15005 -2135
rect 15125 -2255 15170 -2135
rect 15290 -2255 15335 -2135
rect 15455 -2255 15500 -2135
rect 15620 -2255 15675 -2135
rect 15795 -2255 15840 -2135
rect 15960 -2255 16005 -2135
rect 16125 -2255 16170 -2135
rect 16290 -2255 16345 -2135
rect 16465 -2255 16510 -2135
rect 16630 -2255 16675 -2135
rect 16795 -2255 16840 -2135
rect 16960 -2255 17015 -2135
rect 17135 -2255 17180 -2135
rect 17300 -2255 17345 -2135
rect 17465 -2255 17510 -2135
rect 17630 -2255 17685 -2135
rect 17805 -2255 17850 -2135
rect 17970 -2255 18015 -2135
rect 18135 -2255 18180 -2135
rect 18300 -2255 18310 -2135
rect 12810 -2300 18310 -2255
rect 12810 -2420 12820 -2300
rect 12940 -2420 12995 -2300
rect 13115 -2420 13160 -2300
rect 13280 -2420 13325 -2300
rect 13445 -2420 13490 -2300
rect 13610 -2420 13665 -2300
rect 13785 -2420 13830 -2300
rect 13950 -2420 13995 -2300
rect 14115 -2420 14160 -2300
rect 14280 -2420 14335 -2300
rect 14455 -2420 14500 -2300
rect 14620 -2420 14665 -2300
rect 14785 -2420 14830 -2300
rect 14950 -2420 15005 -2300
rect 15125 -2420 15170 -2300
rect 15290 -2420 15335 -2300
rect 15455 -2420 15500 -2300
rect 15620 -2420 15675 -2300
rect 15795 -2420 15840 -2300
rect 15960 -2420 16005 -2300
rect 16125 -2420 16170 -2300
rect 16290 -2420 16345 -2300
rect 16465 -2420 16510 -2300
rect 16630 -2420 16675 -2300
rect 16795 -2420 16840 -2300
rect 16960 -2420 17015 -2300
rect 17135 -2420 17180 -2300
rect 17300 -2420 17345 -2300
rect 17465 -2420 17510 -2300
rect 17630 -2420 17685 -2300
rect 17805 -2420 17850 -2300
rect 17970 -2420 18015 -2300
rect 18135 -2420 18180 -2300
rect 18300 -2420 18310 -2300
rect 12810 -2465 18310 -2420
rect 12810 -2585 12820 -2465
rect 12940 -2585 12995 -2465
rect 13115 -2585 13160 -2465
rect 13280 -2585 13325 -2465
rect 13445 -2585 13490 -2465
rect 13610 -2585 13665 -2465
rect 13785 -2585 13830 -2465
rect 13950 -2585 13995 -2465
rect 14115 -2585 14160 -2465
rect 14280 -2585 14335 -2465
rect 14455 -2585 14500 -2465
rect 14620 -2585 14665 -2465
rect 14785 -2585 14830 -2465
rect 14950 -2585 15005 -2465
rect 15125 -2585 15170 -2465
rect 15290 -2585 15335 -2465
rect 15455 -2585 15500 -2465
rect 15620 -2585 15675 -2465
rect 15795 -2585 15840 -2465
rect 15960 -2585 16005 -2465
rect 16125 -2585 16170 -2465
rect 16290 -2585 16345 -2465
rect 16465 -2585 16510 -2465
rect 16630 -2585 16675 -2465
rect 16795 -2585 16840 -2465
rect 16960 -2585 17015 -2465
rect 17135 -2585 17180 -2465
rect 17300 -2585 17345 -2465
rect 17465 -2585 17510 -2465
rect 17630 -2585 17685 -2465
rect 17805 -2585 17850 -2465
rect 17970 -2585 18015 -2465
rect 18135 -2585 18180 -2465
rect 18300 -2585 18310 -2465
rect 12810 -2640 18310 -2585
rect 12810 -2760 12820 -2640
rect 12940 -2760 12995 -2640
rect 13115 -2760 13160 -2640
rect 13280 -2760 13325 -2640
rect 13445 -2760 13490 -2640
rect 13610 -2760 13665 -2640
rect 13785 -2760 13830 -2640
rect 13950 -2760 13995 -2640
rect 14115 -2760 14160 -2640
rect 14280 -2760 14335 -2640
rect 14455 -2760 14500 -2640
rect 14620 -2760 14665 -2640
rect 14785 -2760 14830 -2640
rect 14950 -2760 15005 -2640
rect 15125 -2760 15170 -2640
rect 15290 -2760 15335 -2640
rect 15455 -2760 15500 -2640
rect 15620 -2760 15675 -2640
rect 15795 -2760 15840 -2640
rect 15960 -2760 16005 -2640
rect 16125 -2760 16170 -2640
rect 16290 -2760 16345 -2640
rect 16465 -2760 16510 -2640
rect 16630 -2760 16675 -2640
rect 16795 -2760 16840 -2640
rect 16960 -2760 17015 -2640
rect 17135 -2760 17180 -2640
rect 17300 -2760 17345 -2640
rect 17465 -2760 17510 -2640
rect 17630 -2760 17685 -2640
rect 17805 -2760 17850 -2640
rect 17970 -2760 18015 -2640
rect 18135 -2760 18180 -2640
rect 18300 -2760 18310 -2640
rect 12810 -2805 18310 -2760
rect 12810 -2925 12820 -2805
rect 12940 -2925 12995 -2805
rect 13115 -2925 13160 -2805
rect 13280 -2925 13325 -2805
rect 13445 -2925 13490 -2805
rect 13610 -2925 13665 -2805
rect 13785 -2925 13830 -2805
rect 13950 -2925 13995 -2805
rect 14115 -2925 14160 -2805
rect 14280 -2925 14335 -2805
rect 14455 -2925 14500 -2805
rect 14620 -2925 14665 -2805
rect 14785 -2925 14830 -2805
rect 14950 -2925 15005 -2805
rect 15125 -2925 15170 -2805
rect 15290 -2925 15335 -2805
rect 15455 -2925 15500 -2805
rect 15620 -2925 15675 -2805
rect 15795 -2925 15840 -2805
rect 15960 -2925 16005 -2805
rect 16125 -2925 16170 -2805
rect 16290 -2925 16345 -2805
rect 16465 -2925 16510 -2805
rect 16630 -2925 16675 -2805
rect 16795 -2925 16840 -2805
rect 16960 -2925 17015 -2805
rect 17135 -2925 17180 -2805
rect 17300 -2925 17345 -2805
rect 17465 -2925 17510 -2805
rect 17630 -2925 17685 -2805
rect 17805 -2925 17850 -2805
rect 17970 -2925 18015 -2805
rect 18135 -2925 18180 -2805
rect 18300 -2925 18310 -2805
rect 12810 -2970 18310 -2925
rect 12810 -3090 12820 -2970
rect 12940 -3090 12995 -2970
rect 13115 -3090 13160 -2970
rect 13280 -3090 13325 -2970
rect 13445 -3090 13490 -2970
rect 13610 -3090 13665 -2970
rect 13785 -3090 13830 -2970
rect 13950 -3090 13995 -2970
rect 14115 -3090 14160 -2970
rect 14280 -3090 14335 -2970
rect 14455 -3090 14500 -2970
rect 14620 -3090 14665 -2970
rect 14785 -3090 14830 -2970
rect 14950 -3090 15005 -2970
rect 15125 -3090 15170 -2970
rect 15290 -3090 15335 -2970
rect 15455 -3090 15500 -2970
rect 15620 -3090 15675 -2970
rect 15795 -3090 15840 -2970
rect 15960 -3090 16005 -2970
rect 16125 -3090 16170 -2970
rect 16290 -3090 16345 -2970
rect 16465 -3090 16510 -2970
rect 16630 -3090 16675 -2970
rect 16795 -3090 16840 -2970
rect 16960 -3090 17015 -2970
rect 17135 -3090 17180 -2970
rect 17300 -3090 17345 -2970
rect 17465 -3090 17510 -2970
rect 17630 -3090 17685 -2970
rect 17805 -3090 17850 -2970
rect 17970 -3090 18015 -2970
rect 18135 -3090 18180 -2970
rect 18300 -3090 18310 -2970
rect 12810 -3135 18310 -3090
rect 12810 -3255 12820 -3135
rect 12940 -3255 12995 -3135
rect 13115 -3255 13160 -3135
rect 13280 -3255 13325 -3135
rect 13445 -3255 13490 -3135
rect 13610 -3255 13665 -3135
rect 13785 -3255 13830 -3135
rect 13950 -3255 13995 -3135
rect 14115 -3255 14160 -3135
rect 14280 -3255 14335 -3135
rect 14455 -3255 14500 -3135
rect 14620 -3255 14665 -3135
rect 14785 -3255 14830 -3135
rect 14950 -3255 15005 -3135
rect 15125 -3255 15170 -3135
rect 15290 -3255 15335 -3135
rect 15455 -3255 15500 -3135
rect 15620 -3255 15675 -3135
rect 15795 -3255 15840 -3135
rect 15960 -3255 16005 -3135
rect 16125 -3255 16170 -3135
rect 16290 -3255 16345 -3135
rect 16465 -3255 16510 -3135
rect 16630 -3255 16675 -3135
rect 16795 -3255 16840 -3135
rect 16960 -3255 17015 -3135
rect 17135 -3255 17180 -3135
rect 17300 -3255 17345 -3135
rect 17465 -3255 17510 -3135
rect 17630 -3255 17685 -3135
rect 17805 -3255 17850 -3135
rect 17970 -3255 18015 -3135
rect 18135 -3255 18180 -3135
rect 18300 -3255 18310 -3135
rect 12810 -3310 18310 -3255
rect 12810 -3430 12820 -3310
rect 12940 -3430 12995 -3310
rect 13115 -3430 13160 -3310
rect 13280 -3430 13325 -3310
rect 13445 -3430 13490 -3310
rect 13610 -3430 13665 -3310
rect 13785 -3430 13830 -3310
rect 13950 -3430 13995 -3310
rect 14115 -3430 14160 -3310
rect 14280 -3430 14335 -3310
rect 14455 -3430 14500 -3310
rect 14620 -3430 14665 -3310
rect 14785 -3430 14830 -3310
rect 14950 -3430 15005 -3310
rect 15125 -3430 15170 -3310
rect 15290 -3430 15335 -3310
rect 15455 -3430 15500 -3310
rect 15620 -3430 15675 -3310
rect 15795 -3430 15840 -3310
rect 15960 -3430 16005 -3310
rect 16125 -3430 16170 -3310
rect 16290 -3430 16345 -3310
rect 16465 -3430 16510 -3310
rect 16630 -3430 16675 -3310
rect 16795 -3430 16840 -3310
rect 16960 -3430 17015 -3310
rect 17135 -3430 17180 -3310
rect 17300 -3430 17345 -3310
rect 17465 -3430 17510 -3310
rect 17630 -3430 17685 -3310
rect 17805 -3430 17850 -3310
rect 17970 -3430 18015 -3310
rect 18135 -3430 18180 -3310
rect 18300 -3430 18310 -3310
rect 12810 -3475 18310 -3430
rect 12810 -3595 12820 -3475
rect 12940 -3595 12995 -3475
rect 13115 -3595 13160 -3475
rect 13280 -3595 13325 -3475
rect 13445 -3595 13490 -3475
rect 13610 -3595 13665 -3475
rect 13785 -3595 13830 -3475
rect 13950 -3595 13995 -3475
rect 14115 -3595 14160 -3475
rect 14280 -3595 14335 -3475
rect 14455 -3595 14500 -3475
rect 14620 -3595 14665 -3475
rect 14785 -3595 14830 -3475
rect 14950 -3595 15005 -3475
rect 15125 -3595 15170 -3475
rect 15290 -3595 15335 -3475
rect 15455 -3595 15500 -3475
rect 15620 -3595 15675 -3475
rect 15795 -3595 15840 -3475
rect 15960 -3595 16005 -3475
rect 16125 -3595 16170 -3475
rect 16290 -3595 16345 -3475
rect 16465 -3595 16510 -3475
rect 16630 -3595 16675 -3475
rect 16795 -3595 16840 -3475
rect 16960 -3595 17015 -3475
rect 17135 -3595 17180 -3475
rect 17300 -3595 17345 -3475
rect 17465 -3595 17510 -3475
rect 17630 -3595 17685 -3475
rect 17805 -3595 17850 -3475
rect 17970 -3595 18015 -3475
rect 18135 -3595 18180 -3475
rect 18300 -3595 18310 -3475
rect 12810 -3640 18310 -3595
rect 12810 -3760 12820 -3640
rect 12940 -3760 12995 -3640
rect 13115 -3760 13160 -3640
rect 13280 -3760 13325 -3640
rect 13445 -3760 13490 -3640
rect 13610 -3760 13665 -3640
rect 13785 -3760 13830 -3640
rect 13950 -3760 13995 -3640
rect 14115 -3760 14160 -3640
rect 14280 -3760 14335 -3640
rect 14455 -3760 14500 -3640
rect 14620 -3760 14665 -3640
rect 14785 -3760 14830 -3640
rect 14950 -3760 15005 -3640
rect 15125 -3760 15170 -3640
rect 15290 -3760 15335 -3640
rect 15455 -3760 15500 -3640
rect 15620 -3760 15675 -3640
rect 15795 -3760 15840 -3640
rect 15960 -3760 16005 -3640
rect 16125 -3760 16170 -3640
rect 16290 -3760 16345 -3640
rect 16465 -3760 16510 -3640
rect 16630 -3760 16675 -3640
rect 16795 -3760 16840 -3640
rect 16960 -3760 17015 -3640
rect 17135 -3760 17180 -3640
rect 17300 -3760 17345 -3640
rect 17465 -3760 17510 -3640
rect 17630 -3760 17685 -3640
rect 17805 -3760 17850 -3640
rect 17970 -3760 18015 -3640
rect 18135 -3760 18180 -3640
rect 18300 -3760 18310 -3640
rect 12810 -3805 18310 -3760
rect 12810 -3925 12820 -3805
rect 12940 -3925 12995 -3805
rect 13115 -3925 13160 -3805
rect 13280 -3925 13325 -3805
rect 13445 -3925 13490 -3805
rect 13610 -3925 13665 -3805
rect 13785 -3925 13830 -3805
rect 13950 -3925 13995 -3805
rect 14115 -3925 14160 -3805
rect 14280 -3925 14335 -3805
rect 14455 -3925 14500 -3805
rect 14620 -3925 14665 -3805
rect 14785 -3925 14830 -3805
rect 14950 -3925 15005 -3805
rect 15125 -3925 15170 -3805
rect 15290 -3925 15335 -3805
rect 15455 -3925 15500 -3805
rect 15620 -3925 15675 -3805
rect 15795 -3925 15840 -3805
rect 15960 -3925 16005 -3805
rect 16125 -3925 16170 -3805
rect 16290 -3925 16345 -3805
rect 16465 -3925 16510 -3805
rect 16630 -3925 16675 -3805
rect 16795 -3925 16840 -3805
rect 16960 -3925 17015 -3805
rect 17135 -3925 17180 -3805
rect 17300 -3925 17345 -3805
rect 17465 -3925 17510 -3805
rect 17630 -3925 17685 -3805
rect 17805 -3925 17850 -3805
rect 17970 -3925 18015 -3805
rect 18135 -3925 18180 -3805
rect 18300 -3925 18310 -3805
rect 12810 -3980 18310 -3925
rect 12810 -4100 12820 -3980
rect 12940 -4100 12995 -3980
rect 13115 -4100 13160 -3980
rect 13280 -4100 13325 -3980
rect 13445 -4100 13490 -3980
rect 13610 -4100 13665 -3980
rect 13785 -4100 13830 -3980
rect 13950 -4100 13995 -3980
rect 14115 -4100 14160 -3980
rect 14280 -4100 14335 -3980
rect 14455 -4100 14500 -3980
rect 14620 -4100 14665 -3980
rect 14785 -4100 14830 -3980
rect 14950 -4100 15005 -3980
rect 15125 -4100 15170 -3980
rect 15290 -4100 15335 -3980
rect 15455 -4100 15500 -3980
rect 15620 -4100 15675 -3980
rect 15795 -4100 15840 -3980
rect 15960 -4100 16005 -3980
rect 16125 -4100 16170 -3980
rect 16290 -4100 16345 -3980
rect 16465 -4100 16510 -3980
rect 16630 -4100 16675 -3980
rect 16795 -4100 16840 -3980
rect 16960 -4100 17015 -3980
rect 17135 -4100 17180 -3980
rect 17300 -4100 17345 -3980
rect 17465 -4100 17510 -3980
rect 17630 -4100 17685 -3980
rect 17805 -4100 17850 -3980
rect 17970 -4100 18015 -3980
rect 18135 -4100 18180 -3980
rect 18300 -4100 18310 -3980
rect 12810 -4110 18310 -4100
rect 18500 1380 24000 1390
rect 18500 1260 18510 1380
rect 18630 1260 18685 1380
rect 18805 1260 18850 1380
rect 18970 1260 19015 1380
rect 19135 1260 19180 1380
rect 19300 1260 19355 1380
rect 19475 1260 19520 1380
rect 19640 1260 19685 1380
rect 19805 1260 19850 1380
rect 19970 1260 20025 1380
rect 20145 1260 20190 1380
rect 20310 1260 20355 1380
rect 20475 1260 20520 1380
rect 20640 1260 20695 1380
rect 20815 1260 20860 1380
rect 20980 1260 21025 1380
rect 21145 1260 21190 1380
rect 21310 1260 21365 1380
rect 21485 1260 21530 1380
rect 21650 1260 21695 1380
rect 21815 1260 21860 1380
rect 21980 1260 22035 1380
rect 22155 1260 22200 1380
rect 22320 1260 22365 1380
rect 22485 1260 22530 1380
rect 22650 1260 22705 1380
rect 22825 1260 22870 1380
rect 22990 1260 23035 1380
rect 23155 1260 23200 1380
rect 23320 1260 23375 1380
rect 23495 1260 23540 1380
rect 23660 1260 23705 1380
rect 23825 1260 23870 1380
rect 23990 1260 24000 1380
rect 18500 1215 24000 1260
rect 18500 1095 18510 1215
rect 18630 1095 18685 1215
rect 18805 1095 18850 1215
rect 18970 1095 19015 1215
rect 19135 1095 19180 1215
rect 19300 1095 19355 1215
rect 19475 1095 19520 1215
rect 19640 1095 19685 1215
rect 19805 1095 19850 1215
rect 19970 1095 20025 1215
rect 20145 1095 20190 1215
rect 20310 1095 20355 1215
rect 20475 1095 20520 1215
rect 20640 1095 20695 1215
rect 20815 1095 20860 1215
rect 20980 1095 21025 1215
rect 21145 1095 21190 1215
rect 21310 1095 21365 1215
rect 21485 1095 21530 1215
rect 21650 1095 21695 1215
rect 21815 1095 21860 1215
rect 21980 1095 22035 1215
rect 22155 1095 22200 1215
rect 22320 1095 22365 1215
rect 22485 1095 22530 1215
rect 22650 1095 22705 1215
rect 22825 1095 22870 1215
rect 22990 1095 23035 1215
rect 23155 1095 23200 1215
rect 23320 1095 23375 1215
rect 23495 1095 23540 1215
rect 23660 1095 23705 1215
rect 23825 1095 23870 1215
rect 23990 1095 24000 1215
rect 18500 1050 24000 1095
rect 18500 930 18510 1050
rect 18630 930 18685 1050
rect 18805 930 18850 1050
rect 18970 930 19015 1050
rect 19135 930 19180 1050
rect 19300 930 19355 1050
rect 19475 930 19520 1050
rect 19640 930 19685 1050
rect 19805 930 19850 1050
rect 19970 930 20025 1050
rect 20145 930 20190 1050
rect 20310 930 20355 1050
rect 20475 930 20520 1050
rect 20640 930 20695 1050
rect 20815 930 20860 1050
rect 20980 930 21025 1050
rect 21145 930 21190 1050
rect 21310 930 21365 1050
rect 21485 930 21530 1050
rect 21650 930 21695 1050
rect 21815 930 21860 1050
rect 21980 930 22035 1050
rect 22155 930 22200 1050
rect 22320 930 22365 1050
rect 22485 930 22530 1050
rect 22650 930 22705 1050
rect 22825 930 22870 1050
rect 22990 930 23035 1050
rect 23155 930 23200 1050
rect 23320 930 23375 1050
rect 23495 930 23540 1050
rect 23660 930 23705 1050
rect 23825 930 23870 1050
rect 23990 930 24000 1050
rect 18500 885 24000 930
rect 18500 765 18510 885
rect 18630 765 18685 885
rect 18805 765 18850 885
rect 18970 765 19015 885
rect 19135 765 19180 885
rect 19300 765 19355 885
rect 19475 765 19520 885
rect 19640 765 19685 885
rect 19805 765 19850 885
rect 19970 765 20025 885
rect 20145 765 20190 885
rect 20310 765 20355 885
rect 20475 765 20520 885
rect 20640 765 20695 885
rect 20815 765 20860 885
rect 20980 765 21025 885
rect 21145 765 21190 885
rect 21310 765 21365 885
rect 21485 765 21530 885
rect 21650 765 21695 885
rect 21815 765 21860 885
rect 21980 765 22035 885
rect 22155 765 22200 885
rect 22320 765 22365 885
rect 22485 765 22530 885
rect 22650 765 22705 885
rect 22825 765 22870 885
rect 22990 765 23035 885
rect 23155 765 23200 885
rect 23320 765 23375 885
rect 23495 765 23540 885
rect 23660 765 23705 885
rect 23825 765 23870 885
rect 23990 765 24000 885
rect 18500 710 24000 765
rect 18500 590 18510 710
rect 18630 590 18685 710
rect 18805 590 18850 710
rect 18970 590 19015 710
rect 19135 590 19180 710
rect 19300 590 19355 710
rect 19475 590 19520 710
rect 19640 590 19685 710
rect 19805 590 19850 710
rect 19970 590 20025 710
rect 20145 590 20190 710
rect 20310 590 20355 710
rect 20475 590 20520 710
rect 20640 590 20695 710
rect 20815 590 20860 710
rect 20980 590 21025 710
rect 21145 590 21190 710
rect 21310 590 21365 710
rect 21485 590 21530 710
rect 21650 590 21695 710
rect 21815 590 21860 710
rect 21980 590 22035 710
rect 22155 590 22200 710
rect 22320 590 22365 710
rect 22485 590 22530 710
rect 22650 590 22705 710
rect 22825 590 22870 710
rect 22990 590 23035 710
rect 23155 590 23200 710
rect 23320 590 23375 710
rect 23495 590 23540 710
rect 23660 590 23705 710
rect 23825 590 23870 710
rect 23990 590 24000 710
rect 18500 545 24000 590
rect 18500 425 18510 545
rect 18630 425 18685 545
rect 18805 425 18850 545
rect 18970 425 19015 545
rect 19135 425 19180 545
rect 19300 425 19355 545
rect 19475 425 19520 545
rect 19640 425 19685 545
rect 19805 425 19850 545
rect 19970 425 20025 545
rect 20145 425 20190 545
rect 20310 425 20355 545
rect 20475 425 20520 545
rect 20640 425 20695 545
rect 20815 425 20860 545
rect 20980 425 21025 545
rect 21145 425 21190 545
rect 21310 425 21365 545
rect 21485 425 21530 545
rect 21650 425 21695 545
rect 21815 425 21860 545
rect 21980 425 22035 545
rect 22155 425 22200 545
rect 22320 425 22365 545
rect 22485 425 22530 545
rect 22650 425 22705 545
rect 22825 425 22870 545
rect 22990 425 23035 545
rect 23155 425 23200 545
rect 23320 425 23375 545
rect 23495 425 23540 545
rect 23660 425 23705 545
rect 23825 425 23870 545
rect 23990 425 24000 545
rect 18500 380 24000 425
rect 18500 260 18510 380
rect 18630 260 18685 380
rect 18805 260 18850 380
rect 18970 260 19015 380
rect 19135 260 19180 380
rect 19300 260 19355 380
rect 19475 260 19520 380
rect 19640 260 19685 380
rect 19805 260 19850 380
rect 19970 260 20025 380
rect 20145 260 20190 380
rect 20310 260 20355 380
rect 20475 260 20520 380
rect 20640 260 20695 380
rect 20815 260 20860 380
rect 20980 260 21025 380
rect 21145 260 21190 380
rect 21310 260 21365 380
rect 21485 260 21530 380
rect 21650 260 21695 380
rect 21815 260 21860 380
rect 21980 260 22035 380
rect 22155 260 22200 380
rect 22320 260 22365 380
rect 22485 260 22530 380
rect 22650 260 22705 380
rect 22825 260 22870 380
rect 22990 260 23035 380
rect 23155 260 23200 380
rect 23320 260 23375 380
rect 23495 260 23540 380
rect 23660 260 23705 380
rect 23825 260 23870 380
rect 23990 260 24000 380
rect 18500 215 24000 260
rect 18500 95 18510 215
rect 18630 95 18685 215
rect 18805 95 18850 215
rect 18970 95 19015 215
rect 19135 95 19180 215
rect 19300 95 19355 215
rect 19475 95 19520 215
rect 19640 95 19685 215
rect 19805 95 19850 215
rect 19970 95 20025 215
rect 20145 95 20190 215
rect 20310 95 20355 215
rect 20475 95 20520 215
rect 20640 95 20695 215
rect 20815 95 20860 215
rect 20980 95 21025 215
rect 21145 95 21190 215
rect 21310 95 21365 215
rect 21485 95 21530 215
rect 21650 95 21695 215
rect 21815 95 21860 215
rect 21980 95 22035 215
rect 22155 95 22200 215
rect 22320 95 22365 215
rect 22485 95 22530 215
rect 22650 95 22705 215
rect 22825 95 22870 215
rect 22990 95 23035 215
rect 23155 95 23200 215
rect 23320 95 23375 215
rect 23495 95 23540 215
rect 23660 95 23705 215
rect 23825 95 23870 215
rect 23990 95 24000 215
rect 18500 40 24000 95
rect 18500 -80 18510 40
rect 18630 -80 18685 40
rect 18805 -80 18850 40
rect 18970 -80 19015 40
rect 19135 -80 19180 40
rect 19300 -80 19355 40
rect 19475 -80 19520 40
rect 19640 -80 19685 40
rect 19805 -80 19850 40
rect 19970 -80 20025 40
rect 20145 -80 20190 40
rect 20310 -80 20355 40
rect 20475 -80 20520 40
rect 20640 -80 20695 40
rect 20815 -80 20860 40
rect 20980 -80 21025 40
rect 21145 -80 21190 40
rect 21310 -80 21365 40
rect 21485 -80 21530 40
rect 21650 -80 21695 40
rect 21815 -80 21860 40
rect 21980 -80 22035 40
rect 22155 -80 22200 40
rect 22320 -80 22365 40
rect 22485 -80 22530 40
rect 22650 -80 22705 40
rect 22825 -80 22870 40
rect 22990 -80 23035 40
rect 23155 -80 23200 40
rect 23320 -80 23375 40
rect 23495 -80 23540 40
rect 23660 -80 23705 40
rect 23825 -80 23870 40
rect 23990 -80 24000 40
rect 18500 -125 24000 -80
rect 18500 -245 18510 -125
rect 18630 -245 18685 -125
rect 18805 -245 18850 -125
rect 18970 -245 19015 -125
rect 19135 -245 19180 -125
rect 19300 -245 19355 -125
rect 19475 -245 19520 -125
rect 19640 -245 19685 -125
rect 19805 -245 19850 -125
rect 19970 -245 20025 -125
rect 20145 -245 20190 -125
rect 20310 -245 20355 -125
rect 20475 -245 20520 -125
rect 20640 -245 20695 -125
rect 20815 -245 20860 -125
rect 20980 -245 21025 -125
rect 21145 -245 21190 -125
rect 21310 -245 21365 -125
rect 21485 -245 21530 -125
rect 21650 -245 21695 -125
rect 21815 -245 21860 -125
rect 21980 -245 22035 -125
rect 22155 -245 22200 -125
rect 22320 -245 22365 -125
rect 22485 -245 22530 -125
rect 22650 -245 22705 -125
rect 22825 -245 22870 -125
rect 22990 -245 23035 -125
rect 23155 -245 23200 -125
rect 23320 -245 23375 -125
rect 23495 -245 23540 -125
rect 23660 -245 23705 -125
rect 23825 -245 23870 -125
rect 23990 -245 24000 -125
rect 18500 -290 24000 -245
rect 18500 -410 18510 -290
rect 18630 -410 18685 -290
rect 18805 -410 18850 -290
rect 18970 -410 19015 -290
rect 19135 -410 19180 -290
rect 19300 -410 19355 -290
rect 19475 -410 19520 -290
rect 19640 -410 19685 -290
rect 19805 -410 19850 -290
rect 19970 -410 20025 -290
rect 20145 -410 20190 -290
rect 20310 -410 20355 -290
rect 20475 -410 20520 -290
rect 20640 -410 20695 -290
rect 20815 -410 20860 -290
rect 20980 -410 21025 -290
rect 21145 -410 21190 -290
rect 21310 -410 21365 -290
rect 21485 -410 21530 -290
rect 21650 -410 21695 -290
rect 21815 -410 21860 -290
rect 21980 -410 22035 -290
rect 22155 -410 22200 -290
rect 22320 -410 22365 -290
rect 22485 -410 22530 -290
rect 22650 -410 22705 -290
rect 22825 -410 22870 -290
rect 22990 -410 23035 -290
rect 23155 -410 23200 -290
rect 23320 -410 23375 -290
rect 23495 -410 23540 -290
rect 23660 -410 23705 -290
rect 23825 -410 23870 -290
rect 23990 -410 24000 -290
rect 18500 -455 24000 -410
rect 18500 -575 18510 -455
rect 18630 -575 18685 -455
rect 18805 -575 18850 -455
rect 18970 -575 19015 -455
rect 19135 -575 19180 -455
rect 19300 -575 19355 -455
rect 19475 -575 19520 -455
rect 19640 -575 19685 -455
rect 19805 -575 19850 -455
rect 19970 -575 20025 -455
rect 20145 -575 20190 -455
rect 20310 -575 20355 -455
rect 20475 -575 20520 -455
rect 20640 -575 20695 -455
rect 20815 -575 20860 -455
rect 20980 -575 21025 -455
rect 21145 -575 21190 -455
rect 21310 -575 21365 -455
rect 21485 -575 21530 -455
rect 21650 -575 21695 -455
rect 21815 -575 21860 -455
rect 21980 -575 22035 -455
rect 22155 -575 22200 -455
rect 22320 -575 22365 -455
rect 22485 -575 22530 -455
rect 22650 -575 22705 -455
rect 22825 -575 22870 -455
rect 22990 -575 23035 -455
rect 23155 -575 23200 -455
rect 23320 -575 23375 -455
rect 23495 -575 23540 -455
rect 23660 -575 23705 -455
rect 23825 -575 23870 -455
rect 23990 -575 24000 -455
rect 18500 -630 24000 -575
rect 18500 -750 18510 -630
rect 18630 -750 18685 -630
rect 18805 -750 18850 -630
rect 18970 -750 19015 -630
rect 19135 -750 19180 -630
rect 19300 -750 19355 -630
rect 19475 -750 19520 -630
rect 19640 -750 19685 -630
rect 19805 -750 19850 -630
rect 19970 -750 20025 -630
rect 20145 -750 20190 -630
rect 20310 -750 20355 -630
rect 20475 -750 20520 -630
rect 20640 -750 20695 -630
rect 20815 -750 20860 -630
rect 20980 -750 21025 -630
rect 21145 -750 21190 -630
rect 21310 -750 21365 -630
rect 21485 -750 21530 -630
rect 21650 -750 21695 -630
rect 21815 -750 21860 -630
rect 21980 -750 22035 -630
rect 22155 -750 22200 -630
rect 22320 -750 22365 -630
rect 22485 -750 22530 -630
rect 22650 -750 22705 -630
rect 22825 -750 22870 -630
rect 22990 -750 23035 -630
rect 23155 -750 23200 -630
rect 23320 -750 23375 -630
rect 23495 -750 23540 -630
rect 23660 -750 23705 -630
rect 23825 -750 23870 -630
rect 23990 -750 24000 -630
rect 18500 -795 24000 -750
rect 18500 -915 18510 -795
rect 18630 -915 18685 -795
rect 18805 -915 18850 -795
rect 18970 -915 19015 -795
rect 19135 -915 19180 -795
rect 19300 -915 19355 -795
rect 19475 -915 19520 -795
rect 19640 -915 19685 -795
rect 19805 -915 19850 -795
rect 19970 -915 20025 -795
rect 20145 -915 20190 -795
rect 20310 -915 20355 -795
rect 20475 -915 20520 -795
rect 20640 -915 20695 -795
rect 20815 -915 20860 -795
rect 20980 -915 21025 -795
rect 21145 -915 21190 -795
rect 21310 -915 21365 -795
rect 21485 -915 21530 -795
rect 21650 -915 21695 -795
rect 21815 -915 21860 -795
rect 21980 -915 22035 -795
rect 22155 -915 22200 -795
rect 22320 -915 22365 -795
rect 22485 -915 22530 -795
rect 22650 -915 22705 -795
rect 22825 -915 22870 -795
rect 22990 -915 23035 -795
rect 23155 -915 23200 -795
rect 23320 -915 23375 -795
rect 23495 -915 23540 -795
rect 23660 -915 23705 -795
rect 23825 -915 23870 -795
rect 23990 -915 24000 -795
rect 18500 -960 24000 -915
rect 18500 -1080 18510 -960
rect 18630 -1080 18685 -960
rect 18805 -1080 18850 -960
rect 18970 -1080 19015 -960
rect 19135 -1080 19180 -960
rect 19300 -1080 19355 -960
rect 19475 -1080 19520 -960
rect 19640 -1080 19685 -960
rect 19805 -1080 19850 -960
rect 19970 -1080 20025 -960
rect 20145 -1080 20190 -960
rect 20310 -1080 20355 -960
rect 20475 -1080 20520 -960
rect 20640 -1080 20695 -960
rect 20815 -1080 20860 -960
rect 20980 -1080 21025 -960
rect 21145 -1080 21190 -960
rect 21310 -1080 21365 -960
rect 21485 -1080 21530 -960
rect 21650 -1080 21695 -960
rect 21815 -1080 21860 -960
rect 21980 -1080 22035 -960
rect 22155 -1080 22200 -960
rect 22320 -1080 22365 -960
rect 22485 -1080 22530 -960
rect 22650 -1080 22705 -960
rect 22825 -1080 22870 -960
rect 22990 -1080 23035 -960
rect 23155 -1080 23200 -960
rect 23320 -1080 23375 -960
rect 23495 -1080 23540 -960
rect 23660 -1080 23705 -960
rect 23825 -1080 23870 -960
rect 23990 -1080 24000 -960
rect 18500 -1125 24000 -1080
rect 18500 -1245 18510 -1125
rect 18630 -1245 18685 -1125
rect 18805 -1245 18850 -1125
rect 18970 -1245 19015 -1125
rect 19135 -1245 19180 -1125
rect 19300 -1245 19355 -1125
rect 19475 -1245 19520 -1125
rect 19640 -1245 19685 -1125
rect 19805 -1245 19850 -1125
rect 19970 -1245 20025 -1125
rect 20145 -1245 20190 -1125
rect 20310 -1245 20355 -1125
rect 20475 -1245 20520 -1125
rect 20640 -1245 20695 -1125
rect 20815 -1245 20860 -1125
rect 20980 -1245 21025 -1125
rect 21145 -1245 21190 -1125
rect 21310 -1245 21365 -1125
rect 21485 -1245 21530 -1125
rect 21650 -1245 21695 -1125
rect 21815 -1245 21860 -1125
rect 21980 -1245 22035 -1125
rect 22155 -1245 22200 -1125
rect 22320 -1245 22365 -1125
rect 22485 -1245 22530 -1125
rect 22650 -1245 22705 -1125
rect 22825 -1245 22870 -1125
rect 22990 -1245 23035 -1125
rect 23155 -1245 23200 -1125
rect 23320 -1245 23375 -1125
rect 23495 -1245 23540 -1125
rect 23660 -1245 23705 -1125
rect 23825 -1245 23870 -1125
rect 23990 -1245 24000 -1125
rect 18500 -1300 24000 -1245
rect 18500 -1420 18510 -1300
rect 18630 -1420 18685 -1300
rect 18805 -1420 18850 -1300
rect 18970 -1420 19015 -1300
rect 19135 -1420 19180 -1300
rect 19300 -1420 19355 -1300
rect 19475 -1420 19520 -1300
rect 19640 -1420 19685 -1300
rect 19805 -1420 19850 -1300
rect 19970 -1420 20025 -1300
rect 20145 -1420 20190 -1300
rect 20310 -1420 20355 -1300
rect 20475 -1420 20520 -1300
rect 20640 -1420 20695 -1300
rect 20815 -1420 20860 -1300
rect 20980 -1420 21025 -1300
rect 21145 -1420 21190 -1300
rect 21310 -1420 21365 -1300
rect 21485 -1420 21530 -1300
rect 21650 -1420 21695 -1300
rect 21815 -1420 21860 -1300
rect 21980 -1420 22035 -1300
rect 22155 -1420 22200 -1300
rect 22320 -1420 22365 -1300
rect 22485 -1420 22530 -1300
rect 22650 -1420 22705 -1300
rect 22825 -1420 22870 -1300
rect 22990 -1420 23035 -1300
rect 23155 -1420 23200 -1300
rect 23320 -1420 23375 -1300
rect 23495 -1420 23540 -1300
rect 23660 -1420 23705 -1300
rect 23825 -1420 23870 -1300
rect 23990 -1420 24000 -1300
rect 18500 -1465 24000 -1420
rect 18500 -1585 18510 -1465
rect 18630 -1585 18685 -1465
rect 18805 -1585 18850 -1465
rect 18970 -1585 19015 -1465
rect 19135 -1585 19180 -1465
rect 19300 -1585 19355 -1465
rect 19475 -1585 19520 -1465
rect 19640 -1585 19685 -1465
rect 19805 -1585 19850 -1465
rect 19970 -1585 20025 -1465
rect 20145 -1585 20190 -1465
rect 20310 -1585 20355 -1465
rect 20475 -1585 20520 -1465
rect 20640 -1585 20695 -1465
rect 20815 -1585 20860 -1465
rect 20980 -1585 21025 -1465
rect 21145 -1585 21190 -1465
rect 21310 -1585 21365 -1465
rect 21485 -1585 21530 -1465
rect 21650 -1585 21695 -1465
rect 21815 -1585 21860 -1465
rect 21980 -1585 22035 -1465
rect 22155 -1585 22200 -1465
rect 22320 -1585 22365 -1465
rect 22485 -1585 22530 -1465
rect 22650 -1585 22705 -1465
rect 22825 -1585 22870 -1465
rect 22990 -1585 23035 -1465
rect 23155 -1585 23200 -1465
rect 23320 -1585 23375 -1465
rect 23495 -1585 23540 -1465
rect 23660 -1585 23705 -1465
rect 23825 -1585 23870 -1465
rect 23990 -1585 24000 -1465
rect 18500 -1630 24000 -1585
rect 18500 -1750 18510 -1630
rect 18630 -1750 18685 -1630
rect 18805 -1750 18850 -1630
rect 18970 -1750 19015 -1630
rect 19135 -1750 19180 -1630
rect 19300 -1750 19355 -1630
rect 19475 -1750 19520 -1630
rect 19640 -1750 19685 -1630
rect 19805 -1750 19850 -1630
rect 19970 -1750 20025 -1630
rect 20145 -1750 20190 -1630
rect 20310 -1750 20355 -1630
rect 20475 -1750 20520 -1630
rect 20640 -1750 20695 -1630
rect 20815 -1750 20860 -1630
rect 20980 -1750 21025 -1630
rect 21145 -1750 21190 -1630
rect 21310 -1750 21365 -1630
rect 21485 -1750 21530 -1630
rect 21650 -1750 21695 -1630
rect 21815 -1750 21860 -1630
rect 21980 -1750 22035 -1630
rect 22155 -1750 22200 -1630
rect 22320 -1750 22365 -1630
rect 22485 -1750 22530 -1630
rect 22650 -1750 22705 -1630
rect 22825 -1750 22870 -1630
rect 22990 -1750 23035 -1630
rect 23155 -1750 23200 -1630
rect 23320 -1750 23375 -1630
rect 23495 -1750 23540 -1630
rect 23660 -1750 23705 -1630
rect 23825 -1750 23870 -1630
rect 23990 -1750 24000 -1630
rect 18500 -1795 24000 -1750
rect 18500 -1915 18510 -1795
rect 18630 -1915 18685 -1795
rect 18805 -1915 18850 -1795
rect 18970 -1915 19015 -1795
rect 19135 -1915 19180 -1795
rect 19300 -1915 19355 -1795
rect 19475 -1915 19520 -1795
rect 19640 -1915 19685 -1795
rect 19805 -1915 19850 -1795
rect 19970 -1915 20025 -1795
rect 20145 -1915 20190 -1795
rect 20310 -1915 20355 -1795
rect 20475 -1915 20520 -1795
rect 20640 -1915 20695 -1795
rect 20815 -1915 20860 -1795
rect 20980 -1915 21025 -1795
rect 21145 -1915 21190 -1795
rect 21310 -1915 21365 -1795
rect 21485 -1915 21530 -1795
rect 21650 -1915 21695 -1795
rect 21815 -1915 21860 -1795
rect 21980 -1915 22035 -1795
rect 22155 -1915 22200 -1795
rect 22320 -1915 22365 -1795
rect 22485 -1915 22530 -1795
rect 22650 -1915 22705 -1795
rect 22825 -1915 22870 -1795
rect 22990 -1915 23035 -1795
rect 23155 -1915 23200 -1795
rect 23320 -1915 23375 -1795
rect 23495 -1915 23540 -1795
rect 23660 -1915 23705 -1795
rect 23825 -1915 23870 -1795
rect 23990 -1915 24000 -1795
rect 18500 -1970 24000 -1915
rect 18500 -2090 18510 -1970
rect 18630 -2090 18685 -1970
rect 18805 -2090 18850 -1970
rect 18970 -2090 19015 -1970
rect 19135 -2090 19180 -1970
rect 19300 -2090 19355 -1970
rect 19475 -2090 19520 -1970
rect 19640 -2090 19685 -1970
rect 19805 -2090 19850 -1970
rect 19970 -2090 20025 -1970
rect 20145 -2090 20190 -1970
rect 20310 -2090 20355 -1970
rect 20475 -2090 20520 -1970
rect 20640 -2090 20695 -1970
rect 20815 -2090 20860 -1970
rect 20980 -2090 21025 -1970
rect 21145 -2090 21190 -1970
rect 21310 -2090 21365 -1970
rect 21485 -2090 21530 -1970
rect 21650 -2090 21695 -1970
rect 21815 -2090 21860 -1970
rect 21980 -2090 22035 -1970
rect 22155 -2090 22200 -1970
rect 22320 -2090 22365 -1970
rect 22485 -2090 22530 -1970
rect 22650 -2090 22705 -1970
rect 22825 -2090 22870 -1970
rect 22990 -2090 23035 -1970
rect 23155 -2090 23200 -1970
rect 23320 -2090 23375 -1970
rect 23495 -2090 23540 -1970
rect 23660 -2090 23705 -1970
rect 23825 -2090 23870 -1970
rect 23990 -2090 24000 -1970
rect 18500 -2135 24000 -2090
rect 18500 -2255 18510 -2135
rect 18630 -2255 18685 -2135
rect 18805 -2255 18850 -2135
rect 18970 -2255 19015 -2135
rect 19135 -2255 19180 -2135
rect 19300 -2255 19355 -2135
rect 19475 -2255 19520 -2135
rect 19640 -2255 19685 -2135
rect 19805 -2255 19850 -2135
rect 19970 -2255 20025 -2135
rect 20145 -2255 20190 -2135
rect 20310 -2255 20355 -2135
rect 20475 -2255 20520 -2135
rect 20640 -2255 20695 -2135
rect 20815 -2255 20860 -2135
rect 20980 -2255 21025 -2135
rect 21145 -2255 21190 -2135
rect 21310 -2255 21365 -2135
rect 21485 -2255 21530 -2135
rect 21650 -2255 21695 -2135
rect 21815 -2255 21860 -2135
rect 21980 -2255 22035 -2135
rect 22155 -2255 22200 -2135
rect 22320 -2255 22365 -2135
rect 22485 -2255 22530 -2135
rect 22650 -2255 22705 -2135
rect 22825 -2255 22870 -2135
rect 22990 -2255 23035 -2135
rect 23155 -2255 23200 -2135
rect 23320 -2255 23375 -2135
rect 23495 -2255 23540 -2135
rect 23660 -2255 23705 -2135
rect 23825 -2255 23870 -2135
rect 23990 -2255 24000 -2135
rect 18500 -2300 24000 -2255
rect 18500 -2420 18510 -2300
rect 18630 -2420 18685 -2300
rect 18805 -2420 18850 -2300
rect 18970 -2420 19015 -2300
rect 19135 -2420 19180 -2300
rect 19300 -2420 19355 -2300
rect 19475 -2420 19520 -2300
rect 19640 -2420 19685 -2300
rect 19805 -2420 19850 -2300
rect 19970 -2420 20025 -2300
rect 20145 -2420 20190 -2300
rect 20310 -2420 20355 -2300
rect 20475 -2420 20520 -2300
rect 20640 -2420 20695 -2300
rect 20815 -2420 20860 -2300
rect 20980 -2420 21025 -2300
rect 21145 -2420 21190 -2300
rect 21310 -2420 21365 -2300
rect 21485 -2420 21530 -2300
rect 21650 -2420 21695 -2300
rect 21815 -2420 21860 -2300
rect 21980 -2420 22035 -2300
rect 22155 -2420 22200 -2300
rect 22320 -2420 22365 -2300
rect 22485 -2420 22530 -2300
rect 22650 -2420 22705 -2300
rect 22825 -2420 22870 -2300
rect 22990 -2420 23035 -2300
rect 23155 -2420 23200 -2300
rect 23320 -2420 23375 -2300
rect 23495 -2420 23540 -2300
rect 23660 -2420 23705 -2300
rect 23825 -2420 23870 -2300
rect 23990 -2420 24000 -2300
rect 18500 -2465 24000 -2420
rect 18500 -2585 18510 -2465
rect 18630 -2585 18685 -2465
rect 18805 -2585 18850 -2465
rect 18970 -2585 19015 -2465
rect 19135 -2585 19180 -2465
rect 19300 -2585 19355 -2465
rect 19475 -2585 19520 -2465
rect 19640 -2585 19685 -2465
rect 19805 -2585 19850 -2465
rect 19970 -2585 20025 -2465
rect 20145 -2585 20190 -2465
rect 20310 -2585 20355 -2465
rect 20475 -2585 20520 -2465
rect 20640 -2585 20695 -2465
rect 20815 -2585 20860 -2465
rect 20980 -2585 21025 -2465
rect 21145 -2585 21190 -2465
rect 21310 -2585 21365 -2465
rect 21485 -2585 21530 -2465
rect 21650 -2585 21695 -2465
rect 21815 -2585 21860 -2465
rect 21980 -2585 22035 -2465
rect 22155 -2585 22200 -2465
rect 22320 -2585 22365 -2465
rect 22485 -2585 22530 -2465
rect 22650 -2585 22705 -2465
rect 22825 -2585 22870 -2465
rect 22990 -2585 23035 -2465
rect 23155 -2585 23200 -2465
rect 23320 -2585 23375 -2465
rect 23495 -2585 23540 -2465
rect 23660 -2585 23705 -2465
rect 23825 -2585 23870 -2465
rect 23990 -2585 24000 -2465
rect 18500 -2640 24000 -2585
rect 18500 -2760 18510 -2640
rect 18630 -2760 18685 -2640
rect 18805 -2760 18850 -2640
rect 18970 -2760 19015 -2640
rect 19135 -2760 19180 -2640
rect 19300 -2760 19355 -2640
rect 19475 -2760 19520 -2640
rect 19640 -2760 19685 -2640
rect 19805 -2760 19850 -2640
rect 19970 -2760 20025 -2640
rect 20145 -2760 20190 -2640
rect 20310 -2760 20355 -2640
rect 20475 -2760 20520 -2640
rect 20640 -2760 20695 -2640
rect 20815 -2760 20860 -2640
rect 20980 -2760 21025 -2640
rect 21145 -2760 21190 -2640
rect 21310 -2760 21365 -2640
rect 21485 -2760 21530 -2640
rect 21650 -2760 21695 -2640
rect 21815 -2760 21860 -2640
rect 21980 -2760 22035 -2640
rect 22155 -2760 22200 -2640
rect 22320 -2760 22365 -2640
rect 22485 -2760 22530 -2640
rect 22650 -2760 22705 -2640
rect 22825 -2760 22870 -2640
rect 22990 -2760 23035 -2640
rect 23155 -2760 23200 -2640
rect 23320 -2760 23375 -2640
rect 23495 -2760 23540 -2640
rect 23660 -2760 23705 -2640
rect 23825 -2760 23870 -2640
rect 23990 -2760 24000 -2640
rect 18500 -2805 24000 -2760
rect 18500 -2925 18510 -2805
rect 18630 -2925 18685 -2805
rect 18805 -2925 18850 -2805
rect 18970 -2925 19015 -2805
rect 19135 -2925 19180 -2805
rect 19300 -2925 19355 -2805
rect 19475 -2925 19520 -2805
rect 19640 -2925 19685 -2805
rect 19805 -2925 19850 -2805
rect 19970 -2925 20025 -2805
rect 20145 -2925 20190 -2805
rect 20310 -2925 20355 -2805
rect 20475 -2925 20520 -2805
rect 20640 -2925 20695 -2805
rect 20815 -2925 20860 -2805
rect 20980 -2925 21025 -2805
rect 21145 -2925 21190 -2805
rect 21310 -2925 21365 -2805
rect 21485 -2925 21530 -2805
rect 21650 -2925 21695 -2805
rect 21815 -2925 21860 -2805
rect 21980 -2925 22035 -2805
rect 22155 -2925 22200 -2805
rect 22320 -2925 22365 -2805
rect 22485 -2925 22530 -2805
rect 22650 -2925 22705 -2805
rect 22825 -2925 22870 -2805
rect 22990 -2925 23035 -2805
rect 23155 -2925 23200 -2805
rect 23320 -2925 23375 -2805
rect 23495 -2925 23540 -2805
rect 23660 -2925 23705 -2805
rect 23825 -2925 23870 -2805
rect 23990 -2925 24000 -2805
rect 18500 -2970 24000 -2925
rect 18500 -3090 18510 -2970
rect 18630 -3090 18685 -2970
rect 18805 -3090 18850 -2970
rect 18970 -3090 19015 -2970
rect 19135 -3090 19180 -2970
rect 19300 -3090 19355 -2970
rect 19475 -3090 19520 -2970
rect 19640 -3090 19685 -2970
rect 19805 -3090 19850 -2970
rect 19970 -3090 20025 -2970
rect 20145 -3090 20190 -2970
rect 20310 -3090 20355 -2970
rect 20475 -3090 20520 -2970
rect 20640 -3090 20695 -2970
rect 20815 -3090 20860 -2970
rect 20980 -3090 21025 -2970
rect 21145 -3090 21190 -2970
rect 21310 -3090 21365 -2970
rect 21485 -3090 21530 -2970
rect 21650 -3090 21695 -2970
rect 21815 -3090 21860 -2970
rect 21980 -3090 22035 -2970
rect 22155 -3090 22200 -2970
rect 22320 -3090 22365 -2970
rect 22485 -3090 22530 -2970
rect 22650 -3090 22705 -2970
rect 22825 -3090 22870 -2970
rect 22990 -3090 23035 -2970
rect 23155 -3090 23200 -2970
rect 23320 -3090 23375 -2970
rect 23495 -3090 23540 -2970
rect 23660 -3090 23705 -2970
rect 23825 -3090 23870 -2970
rect 23990 -3090 24000 -2970
rect 18500 -3135 24000 -3090
rect 18500 -3255 18510 -3135
rect 18630 -3255 18685 -3135
rect 18805 -3255 18850 -3135
rect 18970 -3255 19015 -3135
rect 19135 -3255 19180 -3135
rect 19300 -3255 19355 -3135
rect 19475 -3255 19520 -3135
rect 19640 -3255 19685 -3135
rect 19805 -3255 19850 -3135
rect 19970 -3255 20025 -3135
rect 20145 -3255 20190 -3135
rect 20310 -3255 20355 -3135
rect 20475 -3255 20520 -3135
rect 20640 -3255 20695 -3135
rect 20815 -3255 20860 -3135
rect 20980 -3255 21025 -3135
rect 21145 -3255 21190 -3135
rect 21310 -3255 21365 -3135
rect 21485 -3255 21530 -3135
rect 21650 -3255 21695 -3135
rect 21815 -3255 21860 -3135
rect 21980 -3255 22035 -3135
rect 22155 -3255 22200 -3135
rect 22320 -3255 22365 -3135
rect 22485 -3255 22530 -3135
rect 22650 -3255 22705 -3135
rect 22825 -3255 22870 -3135
rect 22990 -3255 23035 -3135
rect 23155 -3255 23200 -3135
rect 23320 -3255 23375 -3135
rect 23495 -3255 23540 -3135
rect 23660 -3255 23705 -3135
rect 23825 -3255 23870 -3135
rect 23990 -3255 24000 -3135
rect 18500 -3310 24000 -3255
rect 18500 -3430 18510 -3310
rect 18630 -3430 18685 -3310
rect 18805 -3430 18850 -3310
rect 18970 -3430 19015 -3310
rect 19135 -3430 19180 -3310
rect 19300 -3430 19355 -3310
rect 19475 -3430 19520 -3310
rect 19640 -3430 19685 -3310
rect 19805 -3430 19850 -3310
rect 19970 -3430 20025 -3310
rect 20145 -3430 20190 -3310
rect 20310 -3430 20355 -3310
rect 20475 -3430 20520 -3310
rect 20640 -3430 20695 -3310
rect 20815 -3430 20860 -3310
rect 20980 -3430 21025 -3310
rect 21145 -3430 21190 -3310
rect 21310 -3430 21365 -3310
rect 21485 -3430 21530 -3310
rect 21650 -3430 21695 -3310
rect 21815 -3430 21860 -3310
rect 21980 -3430 22035 -3310
rect 22155 -3430 22200 -3310
rect 22320 -3430 22365 -3310
rect 22485 -3430 22530 -3310
rect 22650 -3430 22705 -3310
rect 22825 -3430 22870 -3310
rect 22990 -3430 23035 -3310
rect 23155 -3430 23200 -3310
rect 23320 -3430 23375 -3310
rect 23495 -3430 23540 -3310
rect 23660 -3430 23705 -3310
rect 23825 -3430 23870 -3310
rect 23990 -3430 24000 -3310
rect 18500 -3475 24000 -3430
rect 18500 -3595 18510 -3475
rect 18630 -3595 18685 -3475
rect 18805 -3595 18850 -3475
rect 18970 -3595 19015 -3475
rect 19135 -3595 19180 -3475
rect 19300 -3595 19355 -3475
rect 19475 -3595 19520 -3475
rect 19640 -3595 19685 -3475
rect 19805 -3595 19850 -3475
rect 19970 -3595 20025 -3475
rect 20145 -3595 20190 -3475
rect 20310 -3595 20355 -3475
rect 20475 -3595 20520 -3475
rect 20640 -3595 20695 -3475
rect 20815 -3595 20860 -3475
rect 20980 -3595 21025 -3475
rect 21145 -3595 21190 -3475
rect 21310 -3595 21365 -3475
rect 21485 -3595 21530 -3475
rect 21650 -3595 21695 -3475
rect 21815 -3595 21860 -3475
rect 21980 -3595 22035 -3475
rect 22155 -3595 22200 -3475
rect 22320 -3595 22365 -3475
rect 22485 -3595 22530 -3475
rect 22650 -3595 22705 -3475
rect 22825 -3595 22870 -3475
rect 22990 -3595 23035 -3475
rect 23155 -3595 23200 -3475
rect 23320 -3595 23375 -3475
rect 23495 -3595 23540 -3475
rect 23660 -3595 23705 -3475
rect 23825 -3595 23870 -3475
rect 23990 -3595 24000 -3475
rect 18500 -3640 24000 -3595
rect 18500 -3760 18510 -3640
rect 18630 -3760 18685 -3640
rect 18805 -3760 18850 -3640
rect 18970 -3760 19015 -3640
rect 19135 -3760 19180 -3640
rect 19300 -3760 19355 -3640
rect 19475 -3760 19520 -3640
rect 19640 -3760 19685 -3640
rect 19805 -3760 19850 -3640
rect 19970 -3760 20025 -3640
rect 20145 -3760 20190 -3640
rect 20310 -3760 20355 -3640
rect 20475 -3760 20520 -3640
rect 20640 -3760 20695 -3640
rect 20815 -3760 20860 -3640
rect 20980 -3760 21025 -3640
rect 21145 -3760 21190 -3640
rect 21310 -3760 21365 -3640
rect 21485 -3760 21530 -3640
rect 21650 -3760 21695 -3640
rect 21815 -3760 21860 -3640
rect 21980 -3760 22035 -3640
rect 22155 -3760 22200 -3640
rect 22320 -3760 22365 -3640
rect 22485 -3760 22530 -3640
rect 22650 -3760 22705 -3640
rect 22825 -3760 22870 -3640
rect 22990 -3760 23035 -3640
rect 23155 -3760 23200 -3640
rect 23320 -3760 23375 -3640
rect 23495 -3760 23540 -3640
rect 23660 -3760 23705 -3640
rect 23825 -3760 23870 -3640
rect 23990 -3760 24000 -3640
rect 18500 -3805 24000 -3760
rect 18500 -3925 18510 -3805
rect 18630 -3925 18685 -3805
rect 18805 -3925 18850 -3805
rect 18970 -3925 19015 -3805
rect 19135 -3925 19180 -3805
rect 19300 -3925 19355 -3805
rect 19475 -3925 19520 -3805
rect 19640 -3925 19685 -3805
rect 19805 -3925 19850 -3805
rect 19970 -3925 20025 -3805
rect 20145 -3925 20190 -3805
rect 20310 -3925 20355 -3805
rect 20475 -3925 20520 -3805
rect 20640 -3925 20695 -3805
rect 20815 -3925 20860 -3805
rect 20980 -3925 21025 -3805
rect 21145 -3925 21190 -3805
rect 21310 -3925 21365 -3805
rect 21485 -3925 21530 -3805
rect 21650 -3925 21695 -3805
rect 21815 -3925 21860 -3805
rect 21980 -3925 22035 -3805
rect 22155 -3925 22200 -3805
rect 22320 -3925 22365 -3805
rect 22485 -3925 22530 -3805
rect 22650 -3925 22705 -3805
rect 22825 -3925 22870 -3805
rect 22990 -3925 23035 -3805
rect 23155 -3925 23200 -3805
rect 23320 -3925 23375 -3805
rect 23495 -3925 23540 -3805
rect 23660 -3925 23705 -3805
rect 23825 -3925 23870 -3805
rect 23990 -3925 24000 -3805
rect 18500 -3980 24000 -3925
rect 18500 -4100 18510 -3980
rect 18630 -4100 18685 -3980
rect 18805 -4100 18850 -3980
rect 18970 -4100 19015 -3980
rect 19135 -4100 19180 -3980
rect 19300 -4100 19355 -3980
rect 19475 -4100 19520 -3980
rect 19640 -4100 19685 -3980
rect 19805 -4100 19850 -3980
rect 19970 -4100 20025 -3980
rect 20145 -4100 20190 -3980
rect 20310 -4100 20355 -3980
rect 20475 -4100 20520 -3980
rect 20640 -4100 20695 -3980
rect 20815 -4100 20860 -3980
rect 20980 -4100 21025 -3980
rect 21145 -4100 21190 -3980
rect 21310 -4100 21365 -3980
rect 21485 -4100 21530 -3980
rect 21650 -4100 21695 -3980
rect 21815 -4100 21860 -3980
rect 21980 -4100 22035 -3980
rect 22155 -4100 22200 -3980
rect 22320 -4100 22365 -3980
rect 22485 -4100 22530 -3980
rect 22650 -4100 22705 -3980
rect 22825 -4100 22870 -3980
rect 22990 -4100 23035 -3980
rect 23155 -4100 23200 -3980
rect 23320 -4100 23375 -3980
rect 23495 -4100 23540 -3980
rect 23660 -4100 23705 -3980
rect 23825 -4100 23870 -3980
rect 23990 -4100 24000 -3980
rect 18500 -4110 24000 -4100
rect 24190 1380 29690 1390
rect 24190 1260 24200 1380
rect 24320 1260 24375 1380
rect 24495 1260 24540 1380
rect 24660 1260 24705 1380
rect 24825 1260 24870 1380
rect 24990 1260 25045 1380
rect 25165 1260 25210 1380
rect 25330 1260 25375 1380
rect 25495 1260 25540 1380
rect 25660 1260 25715 1380
rect 25835 1260 25880 1380
rect 26000 1260 26045 1380
rect 26165 1260 26210 1380
rect 26330 1260 26385 1380
rect 26505 1260 26550 1380
rect 26670 1260 26715 1380
rect 26835 1260 26880 1380
rect 27000 1260 27055 1380
rect 27175 1260 27220 1380
rect 27340 1260 27385 1380
rect 27505 1260 27550 1380
rect 27670 1260 27725 1380
rect 27845 1260 27890 1380
rect 28010 1260 28055 1380
rect 28175 1260 28220 1380
rect 28340 1260 28395 1380
rect 28515 1260 28560 1380
rect 28680 1260 28725 1380
rect 28845 1260 28890 1380
rect 29010 1260 29065 1380
rect 29185 1260 29230 1380
rect 29350 1260 29395 1380
rect 29515 1260 29560 1380
rect 29680 1260 29690 1380
rect 24190 1215 29690 1260
rect 24190 1095 24200 1215
rect 24320 1095 24375 1215
rect 24495 1095 24540 1215
rect 24660 1095 24705 1215
rect 24825 1095 24870 1215
rect 24990 1095 25045 1215
rect 25165 1095 25210 1215
rect 25330 1095 25375 1215
rect 25495 1095 25540 1215
rect 25660 1095 25715 1215
rect 25835 1095 25880 1215
rect 26000 1095 26045 1215
rect 26165 1095 26210 1215
rect 26330 1095 26385 1215
rect 26505 1095 26550 1215
rect 26670 1095 26715 1215
rect 26835 1095 26880 1215
rect 27000 1095 27055 1215
rect 27175 1095 27220 1215
rect 27340 1095 27385 1215
rect 27505 1095 27550 1215
rect 27670 1095 27725 1215
rect 27845 1095 27890 1215
rect 28010 1095 28055 1215
rect 28175 1095 28220 1215
rect 28340 1095 28395 1215
rect 28515 1095 28560 1215
rect 28680 1095 28725 1215
rect 28845 1095 28890 1215
rect 29010 1095 29065 1215
rect 29185 1095 29230 1215
rect 29350 1095 29395 1215
rect 29515 1095 29560 1215
rect 29680 1095 29690 1215
rect 24190 1050 29690 1095
rect 24190 930 24200 1050
rect 24320 930 24375 1050
rect 24495 930 24540 1050
rect 24660 930 24705 1050
rect 24825 930 24870 1050
rect 24990 930 25045 1050
rect 25165 930 25210 1050
rect 25330 930 25375 1050
rect 25495 930 25540 1050
rect 25660 930 25715 1050
rect 25835 930 25880 1050
rect 26000 930 26045 1050
rect 26165 930 26210 1050
rect 26330 930 26385 1050
rect 26505 930 26550 1050
rect 26670 930 26715 1050
rect 26835 930 26880 1050
rect 27000 930 27055 1050
rect 27175 930 27220 1050
rect 27340 930 27385 1050
rect 27505 930 27550 1050
rect 27670 930 27725 1050
rect 27845 930 27890 1050
rect 28010 930 28055 1050
rect 28175 930 28220 1050
rect 28340 930 28395 1050
rect 28515 930 28560 1050
rect 28680 930 28725 1050
rect 28845 930 28890 1050
rect 29010 930 29065 1050
rect 29185 930 29230 1050
rect 29350 930 29395 1050
rect 29515 930 29560 1050
rect 29680 930 29690 1050
rect 24190 885 29690 930
rect 24190 765 24200 885
rect 24320 765 24375 885
rect 24495 765 24540 885
rect 24660 765 24705 885
rect 24825 765 24870 885
rect 24990 765 25045 885
rect 25165 765 25210 885
rect 25330 765 25375 885
rect 25495 765 25540 885
rect 25660 765 25715 885
rect 25835 765 25880 885
rect 26000 765 26045 885
rect 26165 765 26210 885
rect 26330 765 26385 885
rect 26505 765 26550 885
rect 26670 765 26715 885
rect 26835 765 26880 885
rect 27000 765 27055 885
rect 27175 765 27220 885
rect 27340 765 27385 885
rect 27505 765 27550 885
rect 27670 765 27725 885
rect 27845 765 27890 885
rect 28010 765 28055 885
rect 28175 765 28220 885
rect 28340 765 28395 885
rect 28515 765 28560 885
rect 28680 765 28725 885
rect 28845 765 28890 885
rect 29010 765 29065 885
rect 29185 765 29230 885
rect 29350 765 29395 885
rect 29515 765 29560 885
rect 29680 765 29690 885
rect 24190 710 29690 765
rect 24190 590 24200 710
rect 24320 590 24375 710
rect 24495 590 24540 710
rect 24660 590 24705 710
rect 24825 590 24870 710
rect 24990 590 25045 710
rect 25165 590 25210 710
rect 25330 590 25375 710
rect 25495 590 25540 710
rect 25660 590 25715 710
rect 25835 590 25880 710
rect 26000 590 26045 710
rect 26165 590 26210 710
rect 26330 590 26385 710
rect 26505 590 26550 710
rect 26670 590 26715 710
rect 26835 590 26880 710
rect 27000 590 27055 710
rect 27175 590 27220 710
rect 27340 590 27385 710
rect 27505 590 27550 710
rect 27670 590 27725 710
rect 27845 590 27890 710
rect 28010 590 28055 710
rect 28175 590 28220 710
rect 28340 590 28395 710
rect 28515 590 28560 710
rect 28680 590 28725 710
rect 28845 590 28890 710
rect 29010 590 29065 710
rect 29185 590 29230 710
rect 29350 590 29395 710
rect 29515 590 29560 710
rect 29680 590 29690 710
rect 24190 545 29690 590
rect 24190 425 24200 545
rect 24320 425 24375 545
rect 24495 425 24540 545
rect 24660 425 24705 545
rect 24825 425 24870 545
rect 24990 425 25045 545
rect 25165 425 25210 545
rect 25330 425 25375 545
rect 25495 425 25540 545
rect 25660 425 25715 545
rect 25835 425 25880 545
rect 26000 425 26045 545
rect 26165 425 26210 545
rect 26330 425 26385 545
rect 26505 425 26550 545
rect 26670 425 26715 545
rect 26835 425 26880 545
rect 27000 425 27055 545
rect 27175 425 27220 545
rect 27340 425 27385 545
rect 27505 425 27550 545
rect 27670 425 27725 545
rect 27845 425 27890 545
rect 28010 425 28055 545
rect 28175 425 28220 545
rect 28340 425 28395 545
rect 28515 425 28560 545
rect 28680 425 28725 545
rect 28845 425 28890 545
rect 29010 425 29065 545
rect 29185 425 29230 545
rect 29350 425 29395 545
rect 29515 425 29560 545
rect 29680 425 29690 545
rect 24190 380 29690 425
rect 24190 260 24200 380
rect 24320 260 24375 380
rect 24495 260 24540 380
rect 24660 260 24705 380
rect 24825 260 24870 380
rect 24990 260 25045 380
rect 25165 260 25210 380
rect 25330 260 25375 380
rect 25495 260 25540 380
rect 25660 260 25715 380
rect 25835 260 25880 380
rect 26000 260 26045 380
rect 26165 260 26210 380
rect 26330 260 26385 380
rect 26505 260 26550 380
rect 26670 260 26715 380
rect 26835 260 26880 380
rect 27000 260 27055 380
rect 27175 260 27220 380
rect 27340 260 27385 380
rect 27505 260 27550 380
rect 27670 260 27725 380
rect 27845 260 27890 380
rect 28010 260 28055 380
rect 28175 260 28220 380
rect 28340 260 28395 380
rect 28515 260 28560 380
rect 28680 260 28725 380
rect 28845 260 28890 380
rect 29010 260 29065 380
rect 29185 260 29230 380
rect 29350 260 29395 380
rect 29515 260 29560 380
rect 29680 260 29690 380
rect 24190 215 29690 260
rect 24190 95 24200 215
rect 24320 95 24375 215
rect 24495 95 24540 215
rect 24660 95 24705 215
rect 24825 95 24870 215
rect 24990 95 25045 215
rect 25165 95 25210 215
rect 25330 95 25375 215
rect 25495 95 25540 215
rect 25660 95 25715 215
rect 25835 95 25880 215
rect 26000 95 26045 215
rect 26165 95 26210 215
rect 26330 95 26385 215
rect 26505 95 26550 215
rect 26670 95 26715 215
rect 26835 95 26880 215
rect 27000 95 27055 215
rect 27175 95 27220 215
rect 27340 95 27385 215
rect 27505 95 27550 215
rect 27670 95 27725 215
rect 27845 95 27890 215
rect 28010 95 28055 215
rect 28175 95 28220 215
rect 28340 95 28395 215
rect 28515 95 28560 215
rect 28680 95 28725 215
rect 28845 95 28890 215
rect 29010 95 29065 215
rect 29185 95 29230 215
rect 29350 95 29395 215
rect 29515 95 29560 215
rect 29680 95 29690 215
rect 24190 40 29690 95
rect 24190 -80 24200 40
rect 24320 -80 24375 40
rect 24495 -80 24540 40
rect 24660 -80 24705 40
rect 24825 -80 24870 40
rect 24990 -80 25045 40
rect 25165 -80 25210 40
rect 25330 -80 25375 40
rect 25495 -80 25540 40
rect 25660 -80 25715 40
rect 25835 -80 25880 40
rect 26000 -80 26045 40
rect 26165 -80 26210 40
rect 26330 -80 26385 40
rect 26505 -80 26550 40
rect 26670 -80 26715 40
rect 26835 -80 26880 40
rect 27000 -80 27055 40
rect 27175 -80 27220 40
rect 27340 -80 27385 40
rect 27505 -80 27550 40
rect 27670 -80 27725 40
rect 27845 -80 27890 40
rect 28010 -80 28055 40
rect 28175 -80 28220 40
rect 28340 -80 28395 40
rect 28515 -80 28560 40
rect 28680 -80 28725 40
rect 28845 -80 28890 40
rect 29010 -80 29065 40
rect 29185 -80 29230 40
rect 29350 -80 29395 40
rect 29515 -80 29560 40
rect 29680 -80 29690 40
rect 24190 -125 29690 -80
rect 24190 -245 24200 -125
rect 24320 -245 24375 -125
rect 24495 -245 24540 -125
rect 24660 -245 24705 -125
rect 24825 -245 24870 -125
rect 24990 -245 25045 -125
rect 25165 -245 25210 -125
rect 25330 -245 25375 -125
rect 25495 -245 25540 -125
rect 25660 -245 25715 -125
rect 25835 -245 25880 -125
rect 26000 -245 26045 -125
rect 26165 -245 26210 -125
rect 26330 -245 26385 -125
rect 26505 -245 26550 -125
rect 26670 -245 26715 -125
rect 26835 -245 26880 -125
rect 27000 -245 27055 -125
rect 27175 -245 27220 -125
rect 27340 -245 27385 -125
rect 27505 -245 27550 -125
rect 27670 -245 27725 -125
rect 27845 -245 27890 -125
rect 28010 -245 28055 -125
rect 28175 -245 28220 -125
rect 28340 -245 28395 -125
rect 28515 -245 28560 -125
rect 28680 -245 28725 -125
rect 28845 -245 28890 -125
rect 29010 -245 29065 -125
rect 29185 -245 29230 -125
rect 29350 -245 29395 -125
rect 29515 -245 29560 -125
rect 29680 -245 29690 -125
rect 24190 -290 29690 -245
rect 24190 -410 24200 -290
rect 24320 -410 24375 -290
rect 24495 -410 24540 -290
rect 24660 -410 24705 -290
rect 24825 -410 24870 -290
rect 24990 -410 25045 -290
rect 25165 -410 25210 -290
rect 25330 -410 25375 -290
rect 25495 -410 25540 -290
rect 25660 -410 25715 -290
rect 25835 -410 25880 -290
rect 26000 -410 26045 -290
rect 26165 -410 26210 -290
rect 26330 -410 26385 -290
rect 26505 -410 26550 -290
rect 26670 -410 26715 -290
rect 26835 -410 26880 -290
rect 27000 -410 27055 -290
rect 27175 -410 27220 -290
rect 27340 -410 27385 -290
rect 27505 -410 27550 -290
rect 27670 -410 27725 -290
rect 27845 -410 27890 -290
rect 28010 -410 28055 -290
rect 28175 -410 28220 -290
rect 28340 -410 28395 -290
rect 28515 -410 28560 -290
rect 28680 -410 28725 -290
rect 28845 -410 28890 -290
rect 29010 -410 29065 -290
rect 29185 -410 29230 -290
rect 29350 -410 29395 -290
rect 29515 -410 29560 -290
rect 29680 -410 29690 -290
rect 24190 -455 29690 -410
rect 24190 -575 24200 -455
rect 24320 -575 24375 -455
rect 24495 -575 24540 -455
rect 24660 -575 24705 -455
rect 24825 -575 24870 -455
rect 24990 -575 25045 -455
rect 25165 -575 25210 -455
rect 25330 -575 25375 -455
rect 25495 -575 25540 -455
rect 25660 -575 25715 -455
rect 25835 -575 25880 -455
rect 26000 -575 26045 -455
rect 26165 -575 26210 -455
rect 26330 -575 26385 -455
rect 26505 -575 26550 -455
rect 26670 -575 26715 -455
rect 26835 -575 26880 -455
rect 27000 -575 27055 -455
rect 27175 -575 27220 -455
rect 27340 -575 27385 -455
rect 27505 -575 27550 -455
rect 27670 -575 27725 -455
rect 27845 -575 27890 -455
rect 28010 -575 28055 -455
rect 28175 -575 28220 -455
rect 28340 -575 28395 -455
rect 28515 -575 28560 -455
rect 28680 -575 28725 -455
rect 28845 -575 28890 -455
rect 29010 -575 29065 -455
rect 29185 -575 29230 -455
rect 29350 -575 29395 -455
rect 29515 -575 29560 -455
rect 29680 -575 29690 -455
rect 24190 -630 29690 -575
rect 24190 -750 24200 -630
rect 24320 -750 24375 -630
rect 24495 -750 24540 -630
rect 24660 -750 24705 -630
rect 24825 -750 24870 -630
rect 24990 -750 25045 -630
rect 25165 -750 25210 -630
rect 25330 -750 25375 -630
rect 25495 -750 25540 -630
rect 25660 -750 25715 -630
rect 25835 -750 25880 -630
rect 26000 -750 26045 -630
rect 26165 -750 26210 -630
rect 26330 -750 26385 -630
rect 26505 -750 26550 -630
rect 26670 -750 26715 -630
rect 26835 -750 26880 -630
rect 27000 -750 27055 -630
rect 27175 -750 27220 -630
rect 27340 -750 27385 -630
rect 27505 -750 27550 -630
rect 27670 -750 27725 -630
rect 27845 -750 27890 -630
rect 28010 -750 28055 -630
rect 28175 -750 28220 -630
rect 28340 -750 28395 -630
rect 28515 -750 28560 -630
rect 28680 -750 28725 -630
rect 28845 -750 28890 -630
rect 29010 -750 29065 -630
rect 29185 -750 29230 -630
rect 29350 -750 29395 -630
rect 29515 -750 29560 -630
rect 29680 -750 29690 -630
rect 24190 -795 29690 -750
rect 24190 -915 24200 -795
rect 24320 -915 24375 -795
rect 24495 -915 24540 -795
rect 24660 -915 24705 -795
rect 24825 -915 24870 -795
rect 24990 -915 25045 -795
rect 25165 -915 25210 -795
rect 25330 -915 25375 -795
rect 25495 -915 25540 -795
rect 25660 -915 25715 -795
rect 25835 -915 25880 -795
rect 26000 -915 26045 -795
rect 26165 -915 26210 -795
rect 26330 -915 26385 -795
rect 26505 -915 26550 -795
rect 26670 -915 26715 -795
rect 26835 -915 26880 -795
rect 27000 -915 27055 -795
rect 27175 -915 27220 -795
rect 27340 -915 27385 -795
rect 27505 -915 27550 -795
rect 27670 -915 27725 -795
rect 27845 -915 27890 -795
rect 28010 -915 28055 -795
rect 28175 -915 28220 -795
rect 28340 -915 28395 -795
rect 28515 -915 28560 -795
rect 28680 -915 28725 -795
rect 28845 -915 28890 -795
rect 29010 -915 29065 -795
rect 29185 -915 29230 -795
rect 29350 -915 29395 -795
rect 29515 -915 29560 -795
rect 29680 -915 29690 -795
rect 24190 -960 29690 -915
rect 24190 -1080 24200 -960
rect 24320 -1080 24375 -960
rect 24495 -1080 24540 -960
rect 24660 -1080 24705 -960
rect 24825 -1080 24870 -960
rect 24990 -1080 25045 -960
rect 25165 -1080 25210 -960
rect 25330 -1080 25375 -960
rect 25495 -1080 25540 -960
rect 25660 -1080 25715 -960
rect 25835 -1080 25880 -960
rect 26000 -1080 26045 -960
rect 26165 -1080 26210 -960
rect 26330 -1080 26385 -960
rect 26505 -1080 26550 -960
rect 26670 -1080 26715 -960
rect 26835 -1080 26880 -960
rect 27000 -1080 27055 -960
rect 27175 -1080 27220 -960
rect 27340 -1080 27385 -960
rect 27505 -1080 27550 -960
rect 27670 -1080 27725 -960
rect 27845 -1080 27890 -960
rect 28010 -1080 28055 -960
rect 28175 -1080 28220 -960
rect 28340 -1080 28395 -960
rect 28515 -1080 28560 -960
rect 28680 -1080 28725 -960
rect 28845 -1080 28890 -960
rect 29010 -1080 29065 -960
rect 29185 -1080 29230 -960
rect 29350 -1080 29395 -960
rect 29515 -1080 29560 -960
rect 29680 -1080 29690 -960
rect 24190 -1125 29690 -1080
rect 24190 -1245 24200 -1125
rect 24320 -1245 24375 -1125
rect 24495 -1245 24540 -1125
rect 24660 -1245 24705 -1125
rect 24825 -1245 24870 -1125
rect 24990 -1245 25045 -1125
rect 25165 -1245 25210 -1125
rect 25330 -1245 25375 -1125
rect 25495 -1245 25540 -1125
rect 25660 -1245 25715 -1125
rect 25835 -1245 25880 -1125
rect 26000 -1245 26045 -1125
rect 26165 -1245 26210 -1125
rect 26330 -1245 26385 -1125
rect 26505 -1245 26550 -1125
rect 26670 -1245 26715 -1125
rect 26835 -1245 26880 -1125
rect 27000 -1245 27055 -1125
rect 27175 -1245 27220 -1125
rect 27340 -1245 27385 -1125
rect 27505 -1245 27550 -1125
rect 27670 -1245 27725 -1125
rect 27845 -1245 27890 -1125
rect 28010 -1245 28055 -1125
rect 28175 -1245 28220 -1125
rect 28340 -1245 28395 -1125
rect 28515 -1245 28560 -1125
rect 28680 -1245 28725 -1125
rect 28845 -1245 28890 -1125
rect 29010 -1245 29065 -1125
rect 29185 -1245 29230 -1125
rect 29350 -1245 29395 -1125
rect 29515 -1245 29560 -1125
rect 29680 -1245 29690 -1125
rect 24190 -1300 29690 -1245
rect 24190 -1420 24200 -1300
rect 24320 -1420 24375 -1300
rect 24495 -1420 24540 -1300
rect 24660 -1420 24705 -1300
rect 24825 -1420 24870 -1300
rect 24990 -1420 25045 -1300
rect 25165 -1420 25210 -1300
rect 25330 -1420 25375 -1300
rect 25495 -1420 25540 -1300
rect 25660 -1420 25715 -1300
rect 25835 -1420 25880 -1300
rect 26000 -1420 26045 -1300
rect 26165 -1420 26210 -1300
rect 26330 -1420 26385 -1300
rect 26505 -1420 26550 -1300
rect 26670 -1420 26715 -1300
rect 26835 -1420 26880 -1300
rect 27000 -1420 27055 -1300
rect 27175 -1420 27220 -1300
rect 27340 -1420 27385 -1300
rect 27505 -1420 27550 -1300
rect 27670 -1420 27725 -1300
rect 27845 -1420 27890 -1300
rect 28010 -1420 28055 -1300
rect 28175 -1420 28220 -1300
rect 28340 -1420 28395 -1300
rect 28515 -1420 28560 -1300
rect 28680 -1420 28725 -1300
rect 28845 -1420 28890 -1300
rect 29010 -1420 29065 -1300
rect 29185 -1420 29230 -1300
rect 29350 -1420 29395 -1300
rect 29515 -1420 29560 -1300
rect 29680 -1420 29690 -1300
rect 24190 -1465 29690 -1420
rect 24190 -1585 24200 -1465
rect 24320 -1585 24375 -1465
rect 24495 -1585 24540 -1465
rect 24660 -1585 24705 -1465
rect 24825 -1585 24870 -1465
rect 24990 -1585 25045 -1465
rect 25165 -1585 25210 -1465
rect 25330 -1585 25375 -1465
rect 25495 -1585 25540 -1465
rect 25660 -1585 25715 -1465
rect 25835 -1585 25880 -1465
rect 26000 -1585 26045 -1465
rect 26165 -1585 26210 -1465
rect 26330 -1585 26385 -1465
rect 26505 -1585 26550 -1465
rect 26670 -1585 26715 -1465
rect 26835 -1585 26880 -1465
rect 27000 -1585 27055 -1465
rect 27175 -1585 27220 -1465
rect 27340 -1585 27385 -1465
rect 27505 -1585 27550 -1465
rect 27670 -1585 27725 -1465
rect 27845 -1585 27890 -1465
rect 28010 -1585 28055 -1465
rect 28175 -1585 28220 -1465
rect 28340 -1585 28395 -1465
rect 28515 -1585 28560 -1465
rect 28680 -1585 28725 -1465
rect 28845 -1585 28890 -1465
rect 29010 -1585 29065 -1465
rect 29185 -1585 29230 -1465
rect 29350 -1585 29395 -1465
rect 29515 -1585 29560 -1465
rect 29680 -1585 29690 -1465
rect 24190 -1630 29690 -1585
rect 24190 -1750 24200 -1630
rect 24320 -1750 24375 -1630
rect 24495 -1750 24540 -1630
rect 24660 -1750 24705 -1630
rect 24825 -1750 24870 -1630
rect 24990 -1750 25045 -1630
rect 25165 -1750 25210 -1630
rect 25330 -1750 25375 -1630
rect 25495 -1750 25540 -1630
rect 25660 -1750 25715 -1630
rect 25835 -1750 25880 -1630
rect 26000 -1750 26045 -1630
rect 26165 -1750 26210 -1630
rect 26330 -1750 26385 -1630
rect 26505 -1750 26550 -1630
rect 26670 -1750 26715 -1630
rect 26835 -1750 26880 -1630
rect 27000 -1750 27055 -1630
rect 27175 -1750 27220 -1630
rect 27340 -1750 27385 -1630
rect 27505 -1750 27550 -1630
rect 27670 -1750 27725 -1630
rect 27845 -1750 27890 -1630
rect 28010 -1750 28055 -1630
rect 28175 -1750 28220 -1630
rect 28340 -1750 28395 -1630
rect 28515 -1750 28560 -1630
rect 28680 -1750 28725 -1630
rect 28845 -1750 28890 -1630
rect 29010 -1750 29065 -1630
rect 29185 -1750 29230 -1630
rect 29350 -1750 29395 -1630
rect 29515 -1750 29560 -1630
rect 29680 -1750 29690 -1630
rect 24190 -1795 29690 -1750
rect 24190 -1915 24200 -1795
rect 24320 -1915 24375 -1795
rect 24495 -1915 24540 -1795
rect 24660 -1915 24705 -1795
rect 24825 -1915 24870 -1795
rect 24990 -1915 25045 -1795
rect 25165 -1915 25210 -1795
rect 25330 -1915 25375 -1795
rect 25495 -1915 25540 -1795
rect 25660 -1915 25715 -1795
rect 25835 -1915 25880 -1795
rect 26000 -1915 26045 -1795
rect 26165 -1915 26210 -1795
rect 26330 -1915 26385 -1795
rect 26505 -1915 26550 -1795
rect 26670 -1915 26715 -1795
rect 26835 -1915 26880 -1795
rect 27000 -1915 27055 -1795
rect 27175 -1915 27220 -1795
rect 27340 -1915 27385 -1795
rect 27505 -1915 27550 -1795
rect 27670 -1915 27725 -1795
rect 27845 -1915 27890 -1795
rect 28010 -1915 28055 -1795
rect 28175 -1915 28220 -1795
rect 28340 -1915 28395 -1795
rect 28515 -1915 28560 -1795
rect 28680 -1915 28725 -1795
rect 28845 -1915 28890 -1795
rect 29010 -1915 29065 -1795
rect 29185 -1915 29230 -1795
rect 29350 -1915 29395 -1795
rect 29515 -1915 29560 -1795
rect 29680 -1915 29690 -1795
rect 24190 -1970 29690 -1915
rect 24190 -2090 24200 -1970
rect 24320 -2090 24375 -1970
rect 24495 -2090 24540 -1970
rect 24660 -2090 24705 -1970
rect 24825 -2090 24870 -1970
rect 24990 -2090 25045 -1970
rect 25165 -2090 25210 -1970
rect 25330 -2090 25375 -1970
rect 25495 -2090 25540 -1970
rect 25660 -2090 25715 -1970
rect 25835 -2090 25880 -1970
rect 26000 -2090 26045 -1970
rect 26165 -2090 26210 -1970
rect 26330 -2090 26385 -1970
rect 26505 -2090 26550 -1970
rect 26670 -2090 26715 -1970
rect 26835 -2090 26880 -1970
rect 27000 -2090 27055 -1970
rect 27175 -2090 27220 -1970
rect 27340 -2090 27385 -1970
rect 27505 -2090 27550 -1970
rect 27670 -2090 27725 -1970
rect 27845 -2090 27890 -1970
rect 28010 -2090 28055 -1970
rect 28175 -2090 28220 -1970
rect 28340 -2090 28395 -1970
rect 28515 -2090 28560 -1970
rect 28680 -2090 28725 -1970
rect 28845 -2090 28890 -1970
rect 29010 -2090 29065 -1970
rect 29185 -2090 29230 -1970
rect 29350 -2090 29395 -1970
rect 29515 -2090 29560 -1970
rect 29680 -2090 29690 -1970
rect 24190 -2135 29690 -2090
rect 24190 -2255 24200 -2135
rect 24320 -2255 24375 -2135
rect 24495 -2255 24540 -2135
rect 24660 -2255 24705 -2135
rect 24825 -2255 24870 -2135
rect 24990 -2255 25045 -2135
rect 25165 -2255 25210 -2135
rect 25330 -2255 25375 -2135
rect 25495 -2255 25540 -2135
rect 25660 -2255 25715 -2135
rect 25835 -2255 25880 -2135
rect 26000 -2255 26045 -2135
rect 26165 -2255 26210 -2135
rect 26330 -2255 26385 -2135
rect 26505 -2255 26550 -2135
rect 26670 -2255 26715 -2135
rect 26835 -2255 26880 -2135
rect 27000 -2255 27055 -2135
rect 27175 -2255 27220 -2135
rect 27340 -2255 27385 -2135
rect 27505 -2255 27550 -2135
rect 27670 -2255 27725 -2135
rect 27845 -2255 27890 -2135
rect 28010 -2255 28055 -2135
rect 28175 -2255 28220 -2135
rect 28340 -2255 28395 -2135
rect 28515 -2255 28560 -2135
rect 28680 -2255 28725 -2135
rect 28845 -2255 28890 -2135
rect 29010 -2255 29065 -2135
rect 29185 -2255 29230 -2135
rect 29350 -2255 29395 -2135
rect 29515 -2255 29560 -2135
rect 29680 -2255 29690 -2135
rect 24190 -2300 29690 -2255
rect 24190 -2420 24200 -2300
rect 24320 -2420 24375 -2300
rect 24495 -2420 24540 -2300
rect 24660 -2420 24705 -2300
rect 24825 -2420 24870 -2300
rect 24990 -2420 25045 -2300
rect 25165 -2420 25210 -2300
rect 25330 -2420 25375 -2300
rect 25495 -2420 25540 -2300
rect 25660 -2420 25715 -2300
rect 25835 -2420 25880 -2300
rect 26000 -2420 26045 -2300
rect 26165 -2420 26210 -2300
rect 26330 -2420 26385 -2300
rect 26505 -2420 26550 -2300
rect 26670 -2420 26715 -2300
rect 26835 -2420 26880 -2300
rect 27000 -2420 27055 -2300
rect 27175 -2420 27220 -2300
rect 27340 -2420 27385 -2300
rect 27505 -2420 27550 -2300
rect 27670 -2420 27725 -2300
rect 27845 -2420 27890 -2300
rect 28010 -2420 28055 -2300
rect 28175 -2420 28220 -2300
rect 28340 -2420 28395 -2300
rect 28515 -2420 28560 -2300
rect 28680 -2420 28725 -2300
rect 28845 -2420 28890 -2300
rect 29010 -2420 29065 -2300
rect 29185 -2420 29230 -2300
rect 29350 -2420 29395 -2300
rect 29515 -2420 29560 -2300
rect 29680 -2420 29690 -2300
rect 24190 -2465 29690 -2420
rect 24190 -2585 24200 -2465
rect 24320 -2585 24375 -2465
rect 24495 -2585 24540 -2465
rect 24660 -2585 24705 -2465
rect 24825 -2585 24870 -2465
rect 24990 -2585 25045 -2465
rect 25165 -2585 25210 -2465
rect 25330 -2585 25375 -2465
rect 25495 -2585 25540 -2465
rect 25660 -2585 25715 -2465
rect 25835 -2585 25880 -2465
rect 26000 -2585 26045 -2465
rect 26165 -2585 26210 -2465
rect 26330 -2585 26385 -2465
rect 26505 -2585 26550 -2465
rect 26670 -2585 26715 -2465
rect 26835 -2585 26880 -2465
rect 27000 -2585 27055 -2465
rect 27175 -2585 27220 -2465
rect 27340 -2585 27385 -2465
rect 27505 -2585 27550 -2465
rect 27670 -2585 27725 -2465
rect 27845 -2585 27890 -2465
rect 28010 -2585 28055 -2465
rect 28175 -2585 28220 -2465
rect 28340 -2585 28395 -2465
rect 28515 -2585 28560 -2465
rect 28680 -2585 28725 -2465
rect 28845 -2585 28890 -2465
rect 29010 -2585 29065 -2465
rect 29185 -2585 29230 -2465
rect 29350 -2585 29395 -2465
rect 29515 -2585 29560 -2465
rect 29680 -2585 29690 -2465
rect 24190 -2640 29690 -2585
rect 24190 -2760 24200 -2640
rect 24320 -2760 24375 -2640
rect 24495 -2760 24540 -2640
rect 24660 -2760 24705 -2640
rect 24825 -2760 24870 -2640
rect 24990 -2760 25045 -2640
rect 25165 -2760 25210 -2640
rect 25330 -2760 25375 -2640
rect 25495 -2760 25540 -2640
rect 25660 -2760 25715 -2640
rect 25835 -2760 25880 -2640
rect 26000 -2760 26045 -2640
rect 26165 -2760 26210 -2640
rect 26330 -2760 26385 -2640
rect 26505 -2760 26550 -2640
rect 26670 -2760 26715 -2640
rect 26835 -2760 26880 -2640
rect 27000 -2760 27055 -2640
rect 27175 -2760 27220 -2640
rect 27340 -2760 27385 -2640
rect 27505 -2760 27550 -2640
rect 27670 -2760 27725 -2640
rect 27845 -2760 27890 -2640
rect 28010 -2760 28055 -2640
rect 28175 -2760 28220 -2640
rect 28340 -2760 28395 -2640
rect 28515 -2760 28560 -2640
rect 28680 -2760 28725 -2640
rect 28845 -2760 28890 -2640
rect 29010 -2760 29065 -2640
rect 29185 -2760 29230 -2640
rect 29350 -2760 29395 -2640
rect 29515 -2760 29560 -2640
rect 29680 -2760 29690 -2640
rect 24190 -2805 29690 -2760
rect 24190 -2925 24200 -2805
rect 24320 -2925 24375 -2805
rect 24495 -2925 24540 -2805
rect 24660 -2925 24705 -2805
rect 24825 -2925 24870 -2805
rect 24990 -2925 25045 -2805
rect 25165 -2925 25210 -2805
rect 25330 -2925 25375 -2805
rect 25495 -2925 25540 -2805
rect 25660 -2925 25715 -2805
rect 25835 -2925 25880 -2805
rect 26000 -2925 26045 -2805
rect 26165 -2925 26210 -2805
rect 26330 -2925 26385 -2805
rect 26505 -2925 26550 -2805
rect 26670 -2925 26715 -2805
rect 26835 -2925 26880 -2805
rect 27000 -2925 27055 -2805
rect 27175 -2925 27220 -2805
rect 27340 -2925 27385 -2805
rect 27505 -2925 27550 -2805
rect 27670 -2925 27725 -2805
rect 27845 -2925 27890 -2805
rect 28010 -2925 28055 -2805
rect 28175 -2925 28220 -2805
rect 28340 -2925 28395 -2805
rect 28515 -2925 28560 -2805
rect 28680 -2925 28725 -2805
rect 28845 -2925 28890 -2805
rect 29010 -2925 29065 -2805
rect 29185 -2925 29230 -2805
rect 29350 -2925 29395 -2805
rect 29515 -2925 29560 -2805
rect 29680 -2925 29690 -2805
rect 24190 -2970 29690 -2925
rect 24190 -3090 24200 -2970
rect 24320 -3090 24375 -2970
rect 24495 -3090 24540 -2970
rect 24660 -3090 24705 -2970
rect 24825 -3090 24870 -2970
rect 24990 -3090 25045 -2970
rect 25165 -3090 25210 -2970
rect 25330 -3090 25375 -2970
rect 25495 -3090 25540 -2970
rect 25660 -3090 25715 -2970
rect 25835 -3090 25880 -2970
rect 26000 -3090 26045 -2970
rect 26165 -3090 26210 -2970
rect 26330 -3090 26385 -2970
rect 26505 -3090 26550 -2970
rect 26670 -3090 26715 -2970
rect 26835 -3090 26880 -2970
rect 27000 -3090 27055 -2970
rect 27175 -3090 27220 -2970
rect 27340 -3090 27385 -2970
rect 27505 -3090 27550 -2970
rect 27670 -3090 27725 -2970
rect 27845 -3090 27890 -2970
rect 28010 -3090 28055 -2970
rect 28175 -3090 28220 -2970
rect 28340 -3090 28395 -2970
rect 28515 -3090 28560 -2970
rect 28680 -3090 28725 -2970
rect 28845 -3090 28890 -2970
rect 29010 -3090 29065 -2970
rect 29185 -3090 29230 -2970
rect 29350 -3090 29395 -2970
rect 29515 -3090 29560 -2970
rect 29680 -3090 29690 -2970
rect 24190 -3135 29690 -3090
rect 24190 -3255 24200 -3135
rect 24320 -3255 24375 -3135
rect 24495 -3255 24540 -3135
rect 24660 -3255 24705 -3135
rect 24825 -3255 24870 -3135
rect 24990 -3255 25045 -3135
rect 25165 -3255 25210 -3135
rect 25330 -3255 25375 -3135
rect 25495 -3255 25540 -3135
rect 25660 -3255 25715 -3135
rect 25835 -3255 25880 -3135
rect 26000 -3255 26045 -3135
rect 26165 -3255 26210 -3135
rect 26330 -3255 26385 -3135
rect 26505 -3255 26550 -3135
rect 26670 -3255 26715 -3135
rect 26835 -3255 26880 -3135
rect 27000 -3255 27055 -3135
rect 27175 -3255 27220 -3135
rect 27340 -3255 27385 -3135
rect 27505 -3255 27550 -3135
rect 27670 -3255 27725 -3135
rect 27845 -3255 27890 -3135
rect 28010 -3255 28055 -3135
rect 28175 -3255 28220 -3135
rect 28340 -3255 28395 -3135
rect 28515 -3255 28560 -3135
rect 28680 -3255 28725 -3135
rect 28845 -3255 28890 -3135
rect 29010 -3255 29065 -3135
rect 29185 -3255 29230 -3135
rect 29350 -3255 29395 -3135
rect 29515 -3255 29560 -3135
rect 29680 -3255 29690 -3135
rect 24190 -3310 29690 -3255
rect 24190 -3430 24200 -3310
rect 24320 -3430 24375 -3310
rect 24495 -3430 24540 -3310
rect 24660 -3430 24705 -3310
rect 24825 -3430 24870 -3310
rect 24990 -3430 25045 -3310
rect 25165 -3430 25210 -3310
rect 25330 -3430 25375 -3310
rect 25495 -3430 25540 -3310
rect 25660 -3430 25715 -3310
rect 25835 -3430 25880 -3310
rect 26000 -3430 26045 -3310
rect 26165 -3430 26210 -3310
rect 26330 -3430 26385 -3310
rect 26505 -3430 26550 -3310
rect 26670 -3430 26715 -3310
rect 26835 -3430 26880 -3310
rect 27000 -3430 27055 -3310
rect 27175 -3430 27220 -3310
rect 27340 -3430 27385 -3310
rect 27505 -3430 27550 -3310
rect 27670 -3430 27725 -3310
rect 27845 -3430 27890 -3310
rect 28010 -3430 28055 -3310
rect 28175 -3430 28220 -3310
rect 28340 -3430 28395 -3310
rect 28515 -3430 28560 -3310
rect 28680 -3430 28725 -3310
rect 28845 -3430 28890 -3310
rect 29010 -3430 29065 -3310
rect 29185 -3430 29230 -3310
rect 29350 -3430 29395 -3310
rect 29515 -3430 29560 -3310
rect 29680 -3430 29690 -3310
rect 24190 -3475 29690 -3430
rect 24190 -3595 24200 -3475
rect 24320 -3595 24375 -3475
rect 24495 -3595 24540 -3475
rect 24660 -3595 24705 -3475
rect 24825 -3595 24870 -3475
rect 24990 -3595 25045 -3475
rect 25165 -3595 25210 -3475
rect 25330 -3595 25375 -3475
rect 25495 -3595 25540 -3475
rect 25660 -3595 25715 -3475
rect 25835 -3595 25880 -3475
rect 26000 -3595 26045 -3475
rect 26165 -3595 26210 -3475
rect 26330 -3595 26385 -3475
rect 26505 -3595 26550 -3475
rect 26670 -3595 26715 -3475
rect 26835 -3595 26880 -3475
rect 27000 -3595 27055 -3475
rect 27175 -3595 27220 -3475
rect 27340 -3595 27385 -3475
rect 27505 -3595 27550 -3475
rect 27670 -3595 27725 -3475
rect 27845 -3595 27890 -3475
rect 28010 -3595 28055 -3475
rect 28175 -3595 28220 -3475
rect 28340 -3595 28395 -3475
rect 28515 -3595 28560 -3475
rect 28680 -3595 28725 -3475
rect 28845 -3595 28890 -3475
rect 29010 -3595 29065 -3475
rect 29185 -3595 29230 -3475
rect 29350 -3595 29395 -3475
rect 29515 -3595 29560 -3475
rect 29680 -3595 29690 -3475
rect 24190 -3640 29690 -3595
rect 24190 -3760 24200 -3640
rect 24320 -3760 24375 -3640
rect 24495 -3760 24540 -3640
rect 24660 -3760 24705 -3640
rect 24825 -3760 24870 -3640
rect 24990 -3760 25045 -3640
rect 25165 -3760 25210 -3640
rect 25330 -3760 25375 -3640
rect 25495 -3760 25540 -3640
rect 25660 -3760 25715 -3640
rect 25835 -3760 25880 -3640
rect 26000 -3760 26045 -3640
rect 26165 -3760 26210 -3640
rect 26330 -3760 26385 -3640
rect 26505 -3760 26550 -3640
rect 26670 -3760 26715 -3640
rect 26835 -3760 26880 -3640
rect 27000 -3760 27055 -3640
rect 27175 -3760 27220 -3640
rect 27340 -3760 27385 -3640
rect 27505 -3760 27550 -3640
rect 27670 -3760 27725 -3640
rect 27845 -3760 27890 -3640
rect 28010 -3760 28055 -3640
rect 28175 -3760 28220 -3640
rect 28340 -3760 28395 -3640
rect 28515 -3760 28560 -3640
rect 28680 -3760 28725 -3640
rect 28845 -3760 28890 -3640
rect 29010 -3760 29065 -3640
rect 29185 -3760 29230 -3640
rect 29350 -3760 29395 -3640
rect 29515 -3760 29560 -3640
rect 29680 -3760 29690 -3640
rect 24190 -3805 29690 -3760
rect 24190 -3925 24200 -3805
rect 24320 -3925 24375 -3805
rect 24495 -3925 24540 -3805
rect 24660 -3925 24705 -3805
rect 24825 -3925 24870 -3805
rect 24990 -3925 25045 -3805
rect 25165 -3925 25210 -3805
rect 25330 -3925 25375 -3805
rect 25495 -3925 25540 -3805
rect 25660 -3925 25715 -3805
rect 25835 -3925 25880 -3805
rect 26000 -3925 26045 -3805
rect 26165 -3925 26210 -3805
rect 26330 -3925 26385 -3805
rect 26505 -3925 26550 -3805
rect 26670 -3925 26715 -3805
rect 26835 -3925 26880 -3805
rect 27000 -3925 27055 -3805
rect 27175 -3925 27220 -3805
rect 27340 -3925 27385 -3805
rect 27505 -3925 27550 -3805
rect 27670 -3925 27725 -3805
rect 27845 -3925 27890 -3805
rect 28010 -3925 28055 -3805
rect 28175 -3925 28220 -3805
rect 28340 -3925 28395 -3805
rect 28515 -3925 28560 -3805
rect 28680 -3925 28725 -3805
rect 28845 -3925 28890 -3805
rect 29010 -3925 29065 -3805
rect 29185 -3925 29230 -3805
rect 29350 -3925 29395 -3805
rect 29515 -3925 29560 -3805
rect 29680 -3925 29690 -3805
rect 24190 -3980 29690 -3925
rect 24190 -4100 24200 -3980
rect 24320 -4100 24375 -3980
rect 24495 -4100 24540 -3980
rect 24660 -4100 24705 -3980
rect 24825 -4100 24870 -3980
rect 24990 -4100 25045 -3980
rect 25165 -4100 25210 -3980
rect 25330 -4100 25375 -3980
rect 25495 -4100 25540 -3980
rect 25660 -4100 25715 -3980
rect 25835 -4100 25880 -3980
rect 26000 -4100 26045 -3980
rect 26165 -4100 26210 -3980
rect 26330 -4100 26385 -3980
rect 26505 -4100 26550 -3980
rect 26670 -4100 26715 -3980
rect 26835 -4100 26880 -3980
rect 27000 -4100 27055 -3980
rect 27175 -4100 27220 -3980
rect 27340 -4100 27385 -3980
rect 27505 -4100 27550 -3980
rect 27670 -4100 27725 -3980
rect 27845 -4100 27890 -3980
rect 28010 -4100 28055 -3980
rect 28175 -4100 28220 -3980
rect 28340 -4100 28395 -3980
rect 28515 -4100 28560 -3980
rect 28680 -4100 28725 -3980
rect 28845 -4100 28890 -3980
rect 29010 -4100 29065 -3980
rect 29185 -4100 29230 -3980
rect 29350 -4100 29395 -3980
rect 29515 -4100 29560 -3980
rect 29680 -4100 29690 -3980
rect 24190 -4110 29690 -4100
rect 7120 -4310 12620 -4300
rect 7120 -4430 7130 -4310
rect 7250 -4430 7295 -4310
rect 7415 -4430 7460 -4310
rect 7580 -4430 7625 -4310
rect 7745 -4430 7800 -4310
rect 7920 -4430 7965 -4310
rect 8085 -4430 8130 -4310
rect 8250 -4430 8295 -4310
rect 8415 -4430 8470 -4310
rect 8590 -4430 8635 -4310
rect 8755 -4430 8800 -4310
rect 8920 -4430 8965 -4310
rect 9085 -4430 9140 -4310
rect 9260 -4430 9305 -4310
rect 9425 -4430 9470 -4310
rect 9590 -4430 9635 -4310
rect 9755 -4430 9810 -4310
rect 9930 -4430 9975 -4310
rect 10095 -4430 10140 -4310
rect 10260 -4430 10305 -4310
rect 10425 -4430 10480 -4310
rect 10600 -4430 10645 -4310
rect 10765 -4430 10810 -4310
rect 10930 -4430 10975 -4310
rect 11095 -4430 11150 -4310
rect 11270 -4430 11315 -4310
rect 11435 -4430 11480 -4310
rect 11600 -4430 11645 -4310
rect 11765 -4430 11820 -4310
rect 11940 -4430 11985 -4310
rect 12105 -4430 12150 -4310
rect 12270 -4430 12315 -4310
rect 12435 -4430 12490 -4310
rect 12610 -4430 12620 -4310
rect 7120 -4485 12620 -4430
rect 7120 -4605 7130 -4485
rect 7250 -4605 7295 -4485
rect 7415 -4605 7460 -4485
rect 7580 -4605 7625 -4485
rect 7745 -4605 7800 -4485
rect 7920 -4605 7965 -4485
rect 8085 -4605 8130 -4485
rect 8250 -4605 8295 -4485
rect 8415 -4605 8470 -4485
rect 8590 -4605 8635 -4485
rect 8755 -4605 8800 -4485
rect 8920 -4605 8965 -4485
rect 9085 -4605 9140 -4485
rect 9260 -4605 9305 -4485
rect 9425 -4605 9470 -4485
rect 9590 -4605 9635 -4485
rect 9755 -4605 9810 -4485
rect 9930 -4605 9975 -4485
rect 10095 -4605 10140 -4485
rect 10260 -4605 10305 -4485
rect 10425 -4605 10480 -4485
rect 10600 -4605 10645 -4485
rect 10765 -4605 10810 -4485
rect 10930 -4605 10975 -4485
rect 11095 -4605 11150 -4485
rect 11270 -4605 11315 -4485
rect 11435 -4605 11480 -4485
rect 11600 -4605 11645 -4485
rect 11765 -4605 11820 -4485
rect 11940 -4605 11985 -4485
rect 12105 -4605 12150 -4485
rect 12270 -4605 12315 -4485
rect 12435 -4605 12490 -4485
rect 12610 -4605 12620 -4485
rect 7120 -4650 12620 -4605
rect 7120 -4770 7130 -4650
rect 7250 -4770 7295 -4650
rect 7415 -4770 7460 -4650
rect 7580 -4770 7625 -4650
rect 7745 -4770 7800 -4650
rect 7920 -4770 7965 -4650
rect 8085 -4770 8130 -4650
rect 8250 -4770 8295 -4650
rect 8415 -4770 8470 -4650
rect 8590 -4770 8635 -4650
rect 8755 -4770 8800 -4650
rect 8920 -4770 8965 -4650
rect 9085 -4770 9140 -4650
rect 9260 -4770 9305 -4650
rect 9425 -4770 9470 -4650
rect 9590 -4770 9635 -4650
rect 9755 -4770 9810 -4650
rect 9930 -4770 9975 -4650
rect 10095 -4770 10140 -4650
rect 10260 -4770 10305 -4650
rect 10425 -4770 10480 -4650
rect 10600 -4770 10645 -4650
rect 10765 -4770 10810 -4650
rect 10930 -4770 10975 -4650
rect 11095 -4770 11150 -4650
rect 11270 -4770 11315 -4650
rect 11435 -4770 11480 -4650
rect 11600 -4770 11645 -4650
rect 11765 -4770 11820 -4650
rect 11940 -4770 11985 -4650
rect 12105 -4770 12150 -4650
rect 12270 -4770 12315 -4650
rect 12435 -4770 12490 -4650
rect 12610 -4770 12620 -4650
rect 7120 -4815 12620 -4770
rect 7120 -4935 7130 -4815
rect 7250 -4935 7295 -4815
rect 7415 -4935 7460 -4815
rect 7580 -4935 7625 -4815
rect 7745 -4935 7800 -4815
rect 7920 -4935 7965 -4815
rect 8085 -4935 8130 -4815
rect 8250 -4935 8295 -4815
rect 8415 -4935 8470 -4815
rect 8590 -4935 8635 -4815
rect 8755 -4935 8800 -4815
rect 8920 -4935 8965 -4815
rect 9085 -4935 9140 -4815
rect 9260 -4935 9305 -4815
rect 9425 -4935 9470 -4815
rect 9590 -4935 9635 -4815
rect 9755 -4935 9810 -4815
rect 9930 -4935 9975 -4815
rect 10095 -4935 10140 -4815
rect 10260 -4935 10305 -4815
rect 10425 -4935 10480 -4815
rect 10600 -4935 10645 -4815
rect 10765 -4935 10810 -4815
rect 10930 -4935 10975 -4815
rect 11095 -4935 11150 -4815
rect 11270 -4935 11315 -4815
rect 11435 -4935 11480 -4815
rect 11600 -4935 11645 -4815
rect 11765 -4935 11820 -4815
rect 11940 -4935 11985 -4815
rect 12105 -4935 12150 -4815
rect 12270 -4935 12315 -4815
rect 12435 -4935 12490 -4815
rect 12610 -4935 12620 -4815
rect 7120 -4980 12620 -4935
rect 7120 -5100 7130 -4980
rect 7250 -5100 7295 -4980
rect 7415 -5100 7460 -4980
rect 7580 -5100 7625 -4980
rect 7745 -5100 7800 -4980
rect 7920 -5100 7965 -4980
rect 8085 -5100 8130 -4980
rect 8250 -5100 8295 -4980
rect 8415 -5100 8470 -4980
rect 8590 -5100 8635 -4980
rect 8755 -5100 8800 -4980
rect 8920 -5100 8965 -4980
rect 9085 -5100 9140 -4980
rect 9260 -5100 9305 -4980
rect 9425 -5100 9470 -4980
rect 9590 -5100 9635 -4980
rect 9755 -5100 9810 -4980
rect 9930 -5100 9975 -4980
rect 10095 -5100 10140 -4980
rect 10260 -5100 10305 -4980
rect 10425 -5100 10480 -4980
rect 10600 -5100 10645 -4980
rect 10765 -5100 10810 -4980
rect 10930 -5100 10975 -4980
rect 11095 -5100 11150 -4980
rect 11270 -5100 11315 -4980
rect 11435 -5100 11480 -4980
rect 11600 -5100 11645 -4980
rect 11765 -5100 11820 -4980
rect 11940 -5100 11985 -4980
rect 12105 -5100 12150 -4980
rect 12270 -5100 12315 -4980
rect 12435 -5100 12490 -4980
rect 12610 -5100 12620 -4980
rect 7120 -5155 12620 -5100
rect 7120 -5275 7130 -5155
rect 7250 -5275 7295 -5155
rect 7415 -5275 7460 -5155
rect 7580 -5275 7625 -5155
rect 7745 -5275 7800 -5155
rect 7920 -5275 7965 -5155
rect 8085 -5275 8130 -5155
rect 8250 -5275 8295 -5155
rect 8415 -5275 8470 -5155
rect 8590 -5275 8635 -5155
rect 8755 -5275 8800 -5155
rect 8920 -5275 8965 -5155
rect 9085 -5275 9140 -5155
rect 9260 -5275 9305 -5155
rect 9425 -5275 9470 -5155
rect 9590 -5275 9635 -5155
rect 9755 -5275 9810 -5155
rect 9930 -5275 9975 -5155
rect 10095 -5275 10140 -5155
rect 10260 -5275 10305 -5155
rect 10425 -5275 10480 -5155
rect 10600 -5275 10645 -5155
rect 10765 -5275 10810 -5155
rect 10930 -5275 10975 -5155
rect 11095 -5275 11150 -5155
rect 11270 -5275 11315 -5155
rect 11435 -5275 11480 -5155
rect 11600 -5275 11645 -5155
rect 11765 -5275 11820 -5155
rect 11940 -5275 11985 -5155
rect 12105 -5275 12150 -5155
rect 12270 -5275 12315 -5155
rect 12435 -5275 12490 -5155
rect 12610 -5275 12620 -5155
rect 7120 -5320 12620 -5275
rect 7120 -5440 7130 -5320
rect 7250 -5440 7295 -5320
rect 7415 -5440 7460 -5320
rect 7580 -5440 7625 -5320
rect 7745 -5440 7800 -5320
rect 7920 -5440 7965 -5320
rect 8085 -5440 8130 -5320
rect 8250 -5440 8295 -5320
rect 8415 -5440 8470 -5320
rect 8590 -5440 8635 -5320
rect 8755 -5440 8800 -5320
rect 8920 -5440 8965 -5320
rect 9085 -5440 9140 -5320
rect 9260 -5440 9305 -5320
rect 9425 -5440 9470 -5320
rect 9590 -5440 9635 -5320
rect 9755 -5440 9810 -5320
rect 9930 -5440 9975 -5320
rect 10095 -5440 10140 -5320
rect 10260 -5440 10305 -5320
rect 10425 -5440 10480 -5320
rect 10600 -5440 10645 -5320
rect 10765 -5440 10810 -5320
rect 10930 -5440 10975 -5320
rect 11095 -5440 11150 -5320
rect 11270 -5440 11315 -5320
rect 11435 -5440 11480 -5320
rect 11600 -5440 11645 -5320
rect 11765 -5440 11820 -5320
rect 11940 -5440 11985 -5320
rect 12105 -5440 12150 -5320
rect 12270 -5440 12315 -5320
rect 12435 -5440 12490 -5320
rect 12610 -5440 12620 -5320
rect 7120 -5485 12620 -5440
rect 7120 -5605 7130 -5485
rect 7250 -5605 7295 -5485
rect 7415 -5605 7460 -5485
rect 7580 -5605 7625 -5485
rect 7745 -5605 7800 -5485
rect 7920 -5605 7965 -5485
rect 8085 -5605 8130 -5485
rect 8250 -5605 8295 -5485
rect 8415 -5605 8470 -5485
rect 8590 -5605 8635 -5485
rect 8755 -5605 8800 -5485
rect 8920 -5605 8965 -5485
rect 9085 -5605 9140 -5485
rect 9260 -5605 9305 -5485
rect 9425 -5605 9470 -5485
rect 9590 -5605 9635 -5485
rect 9755 -5605 9810 -5485
rect 9930 -5605 9975 -5485
rect 10095 -5605 10140 -5485
rect 10260 -5605 10305 -5485
rect 10425 -5605 10480 -5485
rect 10600 -5605 10645 -5485
rect 10765 -5605 10810 -5485
rect 10930 -5605 10975 -5485
rect 11095 -5605 11150 -5485
rect 11270 -5605 11315 -5485
rect 11435 -5605 11480 -5485
rect 11600 -5605 11645 -5485
rect 11765 -5605 11820 -5485
rect 11940 -5605 11985 -5485
rect 12105 -5605 12150 -5485
rect 12270 -5605 12315 -5485
rect 12435 -5605 12490 -5485
rect 12610 -5605 12620 -5485
rect 7120 -5650 12620 -5605
rect 7120 -5770 7130 -5650
rect 7250 -5770 7295 -5650
rect 7415 -5770 7460 -5650
rect 7580 -5770 7625 -5650
rect 7745 -5770 7800 -5650
rect 7920 -5770 7965 -5650
rect 8085 -5770 8130 -5650
rect 8250 -5770 8295 -5650
rect 8415 -5770 8470 -5650
rect 8590 -5770 8635 -5650
rect 8755 -5770 8800 -5650
rect 8920 -5770 8965 -5650
rect 9085 -5770 9140 -5650
rect 9260 -5770 9305 -5650
rect 9425 -5770 9470 -5650
rect 9590 -5770 9635 -5650
rect 9755 -5770 9810 -5650
rect 9930 -5770 9975 -5650
rect 10095 -5770 10140 -5650
rect 10260 -5770 10305 -5650
rect 10425 -5770 10480 -5650
rect 10600 -5770 10645 -5650
rect 10765 -5770 10810 -5650
rect 10930 -5770 10975 -5650
rect 11095 -5770 11150 -5650
rect 11270 -5770 11315 -5650
rect 11435 -5770 11480 -5650
rect 11600 -5770 11645 -5650
rect 11765 -5770 11820 -5650
rect 11940 -5770 11985 -5650
rect 12105 -5770 12150 -5650
rect 12270 -5770 12315 -5650
rect 12435 -5770 12490 -5650
rect 12610 -5770 12620 -5650
rect 7120 -5825 12620 -5770
rect 7120 -5945 7130 -5825
rect 7250 -5945 7295 -5825
rect 7415 -5945 7460 -5825
rect 7580 -5945 7625 -5825
rect 7745 -5945 7800 -5825
rect 7920 -5945 7965 -5825
rect 8085 -5945 8130 -5825
rect 8250 -5945 8295 -5825
rect 8415 -5945 8470 -5825
rect 8590 -5945 8635 -5825
rect 8755 -5945 8800 -5825
rect 8920 -5945 8965 -5825
rect 9085 -5945 9140 -5825
rect 9260 -5945 9305 -5825
rect 9425 -5945 9470 -5825
rect 9590 -5945 9635 -5825
rect 9755 -5945 9810 -5825
rect 9930 -5945 9975 -5825
rect 10095 -5945 10140 -5825
rect 10260 -5945 10305 -5825
rect 10425 -5945 10480 -5825
rect 10600 -5945 10645 -5825
rect 10765 -5945 10810 -5825
rect 10930 -5945 10975 -5825
rect 11095 -5945 11150 -5825
rect 11270 -5945 11315 -5825
rect 11435 -5945 11480 -5825
rect 11600 -5945 11645 -5825
rect 11765 -5945 11820 -5825
rect 11940 -5945 11985 -5825
rect 12105 -5945 12150 -5825
rect 12270 -5945 12315 -5825
rect 12435 -5945 12490 -5825
rect 12610 -5945 12620 -5825
rect 7120 -5990 12620 -5945
rect 7120 -6110 7130 -5990
rect 7250 -6110 7295 -5990
rect 7415 -6110 7460 -5990
rect 7580 -6110 7625 -5990
rect 7745 -6110 7800 -5990
rect 7920 -6110 7965 -5990
rect 8085 -6110 8130 -5990
rect 8250 -6110 8295 -5990
rect 8415 -6110 8470 -5990
rect 8590 -6110 8635 -5990
rect 8755 -6110 8800 -5990
rect 8920 -6110 8965 -5990
rect 9085 -6110 9140 -5990
rect 9260 -6110 9305 -5990
rect 9425 -6110 9470 -5990
rect 9590 -6110 9635 -5990
rect 9755 -6110 9810 -5990
rect 9930 -6110 9975 -5990
rect 10095 -6110 10140 -5990
rect 10260 -6110 10305 -5990
rect 10425 -6110 10480 -5990
rect 10600 -6110 10645 -5990
rect 10765 -6110 10810 -5990
rect 10930 -6110 10975 -5990
rect 11095 -6110 11150 -5990
rect 11270 -6110 11315 -5990
rect 11435 -6110 11480 -5990
rect 11600 -6110 11645 -5990
rect 11765 -6110 11820 -5990
rect 11940 -6110 11985 -5990
rect 12105 -6110 12150 -5990
rect 12270 -6110 12315 -5990
rect 12435 -6110 12490 -5990
rect 12610 -6110 12620 -5990
rect 7120 -6155 12620 -6110
rect 7120 -6275 7130 -6155
rect 7250 -6275 7295 -6155
rect 7415 -6275 7460 -6155
rect 7580 -6275 7625 -6155
rect 7745 -6275 7800 -6155
rect 7920 -6275 7965 -6155
rect 8085 -6275 8130 -6155
rect 8250 -6275 8295 -6155
rect 8415 -6275 8470 -6155
rect 8590 -6275 8635 -6155
rect 8755 -6275 8800 -6155
rect 8920 -6275 8965 -6155
rect 9085 -6275 9140 -6155
rect 9260 -6275 9305 -6155
rect 9425 -6275 9470 -6155
rect 9590 -6275 9635 -6155
rect 9755 -6275 9810 -6155
rect 9930 -6275 9975 -6155
rect 10095 -6275 10140 -6155
rect 10260 -6275 10305 -6155
rect 10425 -6275 10480 -6155
rect 10600 -6275 10645 -6155
rect 10765 -6275 10810 -6155
rect 10930 -6275 10975 -6155
rect 11095 -6275 11150 -6155
rect 11270 -6275 11315 -6155
rect 11435 -6275 11480 -6155
rect 11600 -6275 11645 -6155
rect 11765 -6275 11820 -6155
rect 11940 -6275 11985 -6155
rect 12105 -6275 12150 -6155
rect 12270 -6275 12315 -6155
rect 12435 -6275 12490 -6155
rect 12610 -6275 12620 -6155
rect 7120 -6320 12620 -6275
rect 7120 -6440 7130 -6320
rect 7250 -6440 7295 -6320
rect 7415 -6440 7460 -6320
rect 7580 -6440 7625 -6320
rect 7745 -6440 7800 -6320
rect 7920 -6440 7965 -6320
rect 8085 -6440 8130 -6320
rect 8250 -6440 8295 -6320
rect 8415 -6440 8470 -6320
rect 8590 -6440 8635 -6320
rect 8755 -6440 8800 -6320
rect 8920 -6440 8965 -6320
rect 9085 -6440 9140 -6320
rect 9260 -6440 9305 -6320
rect 9425 -6440 9470 -6320
rect 9590 -6440 9635 -6320
rect 9755 -6440 9810 -6320
rect 9930 -6440 9975 -6320
rect 10095 -6440 10140 -6320
rect 10260 -6440 10305 -6320
rect 10425 -6440 10480 -6320
rect 10600 -6440 10645 -6320
rect 10765 -6440 10810 -6320
rect 10930 -6440 10975 -6320
rect 11095 -6440 11150 -6320
rect 11270 -6440 11315 -6320
rect 11435 -6440 11480 -6320
rect 11600 -6440 11645 -6320
rect 11765 -6440 11820 -6320
rect 11940 -6440 11985 -6320
rect 12105 -6440 12150 -6320
rect 12270 -6440 12315 -6320
rect 12435 -6440 12490 -6320
rect 12610 -6440 12620 -6320
rect 7120 -6495 12620 -6440
rect 7120 -6615 7130 -6495
rect 7250 -6615 7295 -6495
rect 7415 -6615 7460 -6495
rect 7580 -6615 7625 -6495
rect 7745 -6615 7800 -6495
rect 7920 -6615 7965 -6495
rect 8085 -6615 8130 -6495
rect 8250 -6615 8295 -6495
rect 8415 -6615 8470 -6495
rect 8590 -6615 8635 -6495
rect 8755 -6615 8800 -6495
rect 8920 -6615 8965 -6495
rect 9085 -6615 9140 -6495
rect 9260 -6615 9305 -6495
rect 9425 -6615 9470 -6495
rect 9590 -6615 9635 -6495
rect 9755 -6615 9810 -6495
rect 9930 -6615 9975 -6495
rect 10095 -6615 10140 -6495
rect 10260 -6615 10305 -6495
rect 10425 -6615 10480 -6495
rect 10600 -6615 10645 -6495
rect 10765 -6615 10810 -6495
rect 10930 -6615 10975 -6495
rect 11095 -6615 11150 -6495
rect 11270 -6615 11315 -6495
rect 11435 -6615 11480 -6495
rect 11600 -6615 11645 -6495
rect 11765 -6615 11820 -6495
rect 11940 -6615 11985 -6495
rect 12105 -6615 12150 -6495
rect 12270 -6615 12315 -6495
rect 12435 -6615 12490 -6495
rect 12610 -6615 12620 -6495
rect 7120 -6660 12620 -6615
rect 7120 -6780 7130 -6660
rect 7250 -6780 7295 -6660
rect 7415 -6780 7460 -6660
rect 7580 -6780 7625 -6660
rect 7745 -6780 7800 -6660
rect 7920 -6780 7965 -6660
rect 8085 -6780 8130 -6660
rect 8250 -6780 8295 -6660
rect 8415 -6780 8470 -6660
rect 8590 -6780 8635 -6660
rect 8755 -6780 8800 -6660
rect 8920 -6780 8965 -6660
rect 9085 -6780 9140 -6660
rect 9260 -6780 9305 -6660
rect 9425 -6780 9470 -6660
rect 9590 -6780 9635 -6660
rect 9755 -6780 9810 -6660
rect 9930 -6780 9975 -6660
rect 10095 -6780 10140 -6660
rect 10260 -6780 10305 -6660
rect 10425 -6780 10480 -6660
rect 10600 -6780 10645 -6660
rect 10765 -6780 10810 -6660
rect 10930 -6780 10975 -6660
rect 11095 -6780 11150 -6660
rect 11270 -6780 11315 -6660
rect 11435 -6780 11480 -6660
rect 11600 -6780 11645 -6660
rect 11765 -6780 11820 -6660
rect 11940 -6780 11985 -6660
rect 12105 -6780 12150 -6660
rect 12270 -6780 12315 -6660
rect 12435 -6780 12490 -6660
rect 12610 -6780 12620 -6660
rect 7120 -6825 12620 -6780
rect 7120 -6945 7130 -6825
rect 7250 -6945 7295 -6825
rect 7415 -6945 7460 -6825
rect 7580 -6945 7625 -6825
rect 7745 -6945 7800 -6825
rect 7920 -6945 7965 -6825
rect 8085 -6945 8130 -6825
rect 8250 -6945 8295 -6825
rect 8415 -6945 8470 -6825
rect 8590 -6945 8635 -6825
rect 8755 -6945 8800 -6825
rect 8920 -6945 8965 -6825
rect 9085 -6945 9140 -6825
rect 9260 -6945 9305 -6825
rect 9425 -6945 9470 -6825
rect 9590 -6945 9635 -6825
rect 9755 -6945 9810 -6825
rect 9930 -6945 9975 -6825
rect 10095 -6945 10140 -6825
rect 10260 -6945 10305 -6825
rect 10425 -6945 10480 -6825
rect 10600 -6945 10645 -6825
rect 10765 -6945 10810 -6825
rect 10930 -6945 10975 -6825
rect 11095 -6945 11150 -6825
rect 11270 -6945 11315 -6825
rect 11435 -6945 11480 -6825
rect 11600 -6945 11645 -6825
rect 11765 -6945 11820 -6825
rect 11940 -6945 11985 -6825
rect 12105 -6945 12150 -6825
rect 12270 -6945 12315 -6825
rect 12435 -6945 12490 -6825
rect 12610 -6945 12620 -6825
rect 7120 -6990 12620 -6945
rect 7120 -7110 7130 -6990
rect 7250 -7110 7295 -6990
rect 7415 -7110 7460 -6990
rect 7580 -7110 7625 -6990
rect 7745 -7110 7800 -6990
rect 7920 -7110 7965 -6990
rect 8085 -7110 8130 -6990
rect 8250 -7110 8295 -6990
rect 8415 -7110 8470 -6990
rect 8590 -7110 8635 -6990
rect 8755 -7110 8800 -6990
rect 8920 -7110 8965 -6990
rect 9085 -7110 9140 -6990
rect 9260 -7110 9305 -6990
rect 9425 -7110 9470 -6990
rect 9590 -7110 9635 -6990
rect 9755 -7110 9810 -6990
rect 9930 -7110 9975 -6990
rect 10095 -7110 10140 -6990
rect 10260 -7110 10305 -6990
rect 10425 -7110 10480 -6990
rect 10600 -7110 10645 -6990
rect 10765 -7110 10810 -6990
rect 10930 -7110 10975 -6990
rect 11095 -7110 11150 -6990
rect 11270 -7110 11315 -6990
rect 11435 -7110 11480 -6990
rect 11600 -7110 11645 -6990
rect 11765 -7110 11820 -6990
rect 11940 -7110 11985 -6990
rect 12105 -7110 12150 -6990
rect 12270 -7110 12315 -6990
rect 12435 -7110 12490 -6990
rect 12610 -7110 12620 -6990
rect 7120 -7165 12620 -7110
rect 7120 -7285 7130 -7165
rect 7250 -7285 7295 -7165
rect 7415 -7285 7460 -7165
rect 7580 -7285 7625 -7165
rect 7745 -7285 7800 -7165
rect 7920 -7285 7965 -7165
rect 8085 -7285 8130 -7165
rect 8250 -7285 8295 -7165
rect 8415 -7285 8470 -7165
rect 8590 -7285 8635 -7165
rect 8755 -7285 8800 -7165
rect 8920 -7285 8965 -7165
rect 9085 -7285 9140 -7165
rect 9260 -7285 9305 -7165
rect 9425 -7285 9470 -7165
rect 9590 -7285 9635 -7165
rect 9755 -7285 9810 -7165
rect 9930 -7285 9975 -7165
rect 10095 -7285 10140 -7165
rect 10260 -7285 10305 -7165
rect 10425 -7285 10480 -7165
rect 10600 -7285 10645 -7165
rect 10765 -7285 10810 -7165
rect 10930 -7285 10975 -7165
rect 11095 -7285 11150 -7165
rect 11270 -7285 11315 -7165
rect 11435 -7285 11480 -7165
rect 11600 -7285 11645 -7165
rect 11765 -7285 11820 -7165
rect 11940 -7285 11985 -7165
rect 12105 -7285 12150 -7165
rect 12270 -7285 12315 -7165
rect 12435 -7285 12490 -7165
rect 12610 -7285 12620 -7165
rect 7120 -7330 12620 -7285
rect 7120 -7450 7130 -7330
rect 7250 -7450 7295 -7330
rect 7415 -7450 7460 -7330
rect 7580 -7450 7625 -7330
rect 7745 -7450 7800 -7330
rect 7920 -7450 7965 -7330
rect 8085 -7450 8130 -7330
rect 8250 -7450 8295 -7330
rect 8415 -7450 8470 -7330
rect 8590 -7450 8635 -7330
rect 8755 -7450 8800 -7330
rect 8920 -7450 8965 -7330
rect 9085 -7450 9140 -7330
rect 9260 -7450 9305 -7330
rect 9425 -7450 9470 -7330
rect 9590 -7450 9635 -7330
rect 9755 -7450 9810 -7330
rect 9930 -7450 9975 -7330
rect 10095 -7450 10140 -7330
rect 10260 -7450 10305 -7330
rect 10425 -7450 10480 -7330
rect 10600 -7450 10645 -7330
rect 10765 -7450 10810 -7330
rect 10930 -7450 10975 -7330
rect 11095 -7450 11150 -7330
rect 11270 -7450 11315 -7330
rect 11435 -7450 11480 -7330
rect 11600 -7450 11645 -7330
rect 11765 -7450 11820 -7330
rect 11940 -7450 11985 -7330
rect 12105 -7450 12150 -7330
rect 12270 -7450 12315 -7330
rect 12435 -7450 12490 -7330
rect 12610 -7450 12620 -7330
rect 7120 -7495 12620 -7450
rect 7120 -7615 7130 -7495
rect 7250 -7615 7295 -7495
rect 7415 -7615 7460 -7495
rect 7580 -7615 7625 -7495
rect 7745 -7615 7800 -7495
rect 7920 -7615 7965 -7495
rect 8085 -7615 8130 -7495
rect 8250 -7615 8295 -7495
rect 8415 -7615 8470 -7495
rect 8590 -7615 8635 -7495
rect 8755 -7615 8800 -7495
rect 8920 -7615 8965 -7495
rect 9085 -7615 9140 -7495
rect 9260 -7615 9305 -7495
rect 9425 -7615 9470 -7495
rect 9590 -7615 9635 -7495
rect 9755 -7615 9810 -7495
rect 9930 -7615 9975 -7495
rect 10095 -7615 10140 -7495
rect 10260 -7615 10305 -7495
rect 10425 -7615 10480 -7495
rect 10600 -7615 10645 -7495
rect 10765 -7615 10810 -7495
rect 10930 -7615 10975 -7495
rect 11095 -7615 11150 -7495
rect 11270 -7615 11315 -7495
rect 11435 -7615 11480 -7495
rect 11600 -7615 11645 -7495
rect 11765 -7615 11820 -7495
rect 11940 -7615 11985 -7495
rect 12105 -7615 12150 -7495
rect 12270 -7615 12315 -7495
rect 12435 -7615 12490 -7495
rect 12610 -7615 12620 -7495
rect 7120 -7660 12620 -7615
rect 7120 -7780 7130 -7660
rect 7250 -7780 7295 -7660
rect 7415 -7780 7460 -7660
rect 7580 -7780 7625 -7660
rect 7745 -7780 7800 -7660
rect 7920 -7780 7965 -7660
rect 8085 -7780 8130 -7660
rect 8250 -7780 8295 -7660
rect 8415 -7780 8470 -7660
rect 8590 -7780 8635 -7660
rect 8755 -7780 8800 -7660
rect 8920 -7780 8965 -7660
rect 9085 -7780 9140 -7660
rect 9260 -7780 9305 -7660
rect 9425 -7780 9470 -7660
rect 9590 -7780 9635 -7660
rect 9755 -7780 9810 -7660
rect 9930 -7780 9975 -7660
rect 10095 -7780 10140 -7660
rect 10260 -7780 10305 -7660
rect 10425 -7780 10480 -7660
rect 10600 -7780 10645 -7660
rect 10765 -7780 10810 -7660
rect 10930 -7780 10975 -7660
rect 11095 -7780 11150 -7660
rect 11270 -7780 11315 -7660
rect 11435 -7780 11480 -7660
rect 11600 -7780 11645 -7660
rect 11765 -7780 11820 -7660
rect 11940 -7780 11985 -7660
rect 12105 -7780 12150 -7660
rect 12270 -7780 12315 -7660
rect 12435 -7780 12490 -7660
rect 12610 -7780 12620 -7660
rect 7120 -7835 12620 -7780
rect 7120 -7955 7130 -7835
rect 7250 -7955 7295 -7835
rect 7415 -7955 7460 -7835
rect 7580 -7955 7625 -7835
rect 7745 -7955 7800 -7835
rect 7920 -7955 7965 -7835
rect 8085 -7955 8130 -7835
rect 8250 -7955 8295 -7835
rect 8415 -7955 8470 -7835
rect 8590 -7955 8635 -7835
rect 8755 -7955 8800 -7835
rect 8920 -7955 8965 -7835
rect 9085 -7955 9140 -7835
rect 9260 -7955 9305 -7835
rect 9425 -7955 9470 -7835
rect 9590 -7955 9635 -7835
rect 9755 -7955 9810 -7835
rect 9930 -7955 9975 -7835
rect 10095 -7955 10140 -7835
rect 10260 -7955 10305 -7835
rect 10425 -7955 10480 -7835
rect 10600 -7955 10645 -7835
rect 10765 -7955 10810 -7835
rect 10930 -7955 10975 -7835
rect 11095 -7955 11150 -7835
rect 11270 -7955 11315 -7835
rect 11435 -7955 11480 -7835
rect 11600 -7955 11645 -7835
rect 11765 -7955 11820 -7835
rect 11940 -7955 11985 -7835
rect 12105 -7955 12150 -7835
rect 12270 -7955 12315 -7835
rect 12435 -7955 12490 -7835
rect 12610 -7955 12620 -7835
rect 7120 -8000 12620 -7955
rect 7120 -8120 7130 -8000
rect 7250 -8120 7295 -8000
rect 7415 -8120 7460 -8000
rect 7580 -8120 7625 -8000
rect 7745 -8120 7800 -8000
rect 7920 -8120 7965 -8000
rect 8085 -8120 8130 -8000
rect 8250 -8120 8295 -8000
rect 8415 -8120 8470 -8000
rect 8590 -8120 8635 -8000
rect 8755 -8120 8800 -8000
rect 8920 -8120 8965 -8000
rect 9085 -8120 9140 -8000
rect 9260 -8120 9305 -8000
rect 9425 -8120 9470 -8000
rect 9590 -8120 9635 -8000
rect 9755 -8120 9810 -8000
rect 9930 -8120 9975 -8000
rect 10095 -8120 10140 -8000
rect 10260 -8120 10305 -8000
rect 10425 -8120 10480 -8000
rect 10600 -8120 10645 -8000
rect 10765 -8120 10810 -8000
rect 10930 -8120 10975 -8000
rect 11095 -8120 11150 -8000
rect 11270 -8120 11315 -8000
rect 11435 -8120 11480 -8000
rect 11600 -8120 11645 -8000
rect 11765 -8120 11820 -8000
rect 11940 -8120 11985 -8000
rect 12105 -8120 12150 -8000
rect 12270 -8120 12315 -8000
rect 12435 -8120 12490 -8000
rect 12610 -8120 12620 -8000
rect 7120 -8165 12620 -8120
rect 7120 -8285 7130 -8165
rect 7250 -8285 7295 -8165
rect 7415 -8285 7460 -8165
rect 7580 -8285 7625 -8165
rect 7745 -8285 7800 -8165
rect 7920 -8285 7965 -8165
rect 8085 -8285 8130 -8165
rect 8250 -8285 8295 -8165
rect 8415 -8285 8470 -8165
rect 8590 -8285 8635 -8165
rect 8755 -8285 8800 -8165
rect 8920 -8285 8965 -8165
rect 9085 -8285 9140 -8165
rect 9260 -8285 9305 -8165
rect 9425 -8285 9470 -8165
rect 9590 -8285 9635 -8165
rect 9755 -8285 9810 -8165
rect 9930 -8285 9975 -8165
rect 10095 -8285 10140 -8165
rect 10260 -8285 10305 -8165
rect 10425 -8285 10480 -8165
rect 10600 -8285 10645 -8165
rect 10765 -8285 10810 -8165
rect 10930 -8285 10975 -8165
rect 11095 -8285 11150 -8165
rect 11270 -8285 11315 -8165
rect 11435 -8285 11480 -8165
rect 11600 -8285 11645 -8165
rect 11765 -8285 11820 -8165
rect 11940 -8285 11985 -8165
rect 12105 -8285 12150 -8165
rect 12270 -8285 12315 -8165
rect 12435 -8285 12490 -8165
rect 12610 -8285 12620 -8165
rect 7120 -8330 12620 -8285
rect 7120 -8450 7130 -8330
rect 7250 -8450 7295 -8330
rect 7415 -8450 7460 -8330
rect 7580 -8450 7625 -8330
rect 7745 -8450 7800 -8330
rect 7920 -8450 7965 -8330
rect 8085 -8450 8130 -8330
rect 8250 -8450 8295 -8330
rect 8415 -8450 8470 -8330
rect 8590 -8450 8635 -8330
rect 8755 -8450 8800 -8330
rect 8920 -8450 8965 -8330
rect 9085 -8450 9140 -8330
rect 9260 -8450 9305 -8330
rect 9425 -8450 9470 -8330
rect 9590 -8450 9635 -8330
rect 9755 -8450 9810 -8330
rect 9930 -8450 9975 -8330
rect 10095 -8450 10140 -8330
rect 10260 -8450 10305 -8330
rect 10425 -8450 10480 -8330
rect 10600 -8450 10645 -8330
rect 10765 -8450 10810 -8330
rect 10930 -8450 10975 -8330
rect 11095 -8450 11150 -8330
rect 11270 -8450 11315 -8330
rect 11435 -8450 11480 -8330
rect 11600 -8450 11645 -8330
rect 11765 -8450 11820 -8330
rect 11940 -8450 11985 -8330
rect 12105 -8450 12150 -8330
rect 12270 -8450 12315 -8330
rect 12435 -8450 12490 -8330
rect 12610 -8450 12620 -8330
rect 7120 -8505 12620 -8450
rect 7120 -8625 7130 -8505
rect 7250 -8625 7295 -8505
rect 7415 -8625 7460 -8505
rect 7580 -8625 7625 -8505
rect 7745 -8625 7800 -8505
rect 7920 -8625 7965 -8505
rect 8085 -8625 8130 -8505
rect 8250 -8625 8295 -8505
rect 8415 -8625 8470 -8505
rect 8590 -8625 8635 -8505
rect 8755 -8625 8800 -8505
rect 8920 -8625 8965 -8505
rect 9085 -8625 9140 -8505
rect 9260 -8625 9305 -8505
rect 9425 -8625 9470 -8505
rect 9590 -8625 9635 -8505
rect 9755 -8625 9810 -8505
rect 9930 -8625 9975 -8505
rect 10095 -8625 10140 -8505
rect 10260 -8625 10305 -8505
rect 10425 -8625 10480 -8505
rect 10600 -8625 10645 -8505
rect 10765 -8625 10810 -8505
rect 10930 -8625 10975 -8505
rect 11095 -8625 11150 -8505
rect 11270 -8625 11315 -8505
rect 11435 -8625 11480 -8505
rect 11600 -8625 11645 -8505
rect 11765 -8625 11820 -8505
rect 11940 -8625 11985 -8505
rect 12105 -8625 12150 -8505
rect 12270 -8625 12315 -8505
rect 12435 -8625 12490 -8505
rect 12610 -8625 12620 -8505
rect 7120 -8670 12620 -8625
rect 7120 -8790 7130 -8670
rect 7250 -8790 7295 -8670
rect 7415 -8790 7460 -8670
rect 7580 -8790 7625 -8670
rect 7745 -8790 7800 -8670
rect 7920 -8790 7965 -8670
rect 8085 -8790 8130 -8670
rect 8250 -8790 8295 -8670
rect 8415 -8790 8470 -8670
rect 8590 -8790 8635 -8670
rect 8755 -8790 8800 -8670
rect 8920 -8790 8965 -8670
rect 9085 -8790 9140 -8670
rect 9260 -8790 9305 -8670
rect 9425 -8790 9470 -8670
rect 9590 -8790 9635 -8670
rect 9755 -8790 9810 -8670
rect 9930 -8790 9975 -8670
rect 10095 -8790 10140 -8670
rect 10260 -8790 10305 -8670
rect 10425 -8790 10480 -8670
rect 10600 -8790 10645 -8670
rect 10765 -8790 10810 -8670
rect 10930 -8790 10975 -8670
rect 11095 -8790 11150 -8670
rect 11270 -8790 11315 -8670
rect 11435 -8790 11480 -8670
rect 11600 -8790 11645 -8670
rect 11765 -8790 11820 -8670
rect 11940 -8790 11985 -8670
rect 12105 -8790 12150 -8670
rect 12270 -8790 12315 -8670
rect 12435 -8790 12490 -8670
rect 12610 -8790 12620 -8670
rect 7120 -8835 12620 -8790
rect 7120 -8955 7130 -8835
rect 7250 -8955 7295 -8835
rect 7415 -8955 7460 -8835
rect 7580 -8955 7625 -8835
rect 7745 -8955 7800 -8835
rect 7920 -8955 7965 -8835
rect 8085 -8955 8130 -8835
rect 8250 -8955 8295 -8835
rect 8415 -8955 8470 -8835
rect 8590 -8955 8635 -8835
rect 8755 -8955 8800 -8835
rect 8920 -8955 8965 -8835
rect 9085 -8955 9140 -8835
rect 9260 -8955 9305 -8835
rect 9425 -8955 9470 -8835
rect 9590 -8955 9635 -8835
rect 9755 -8955 9810 -8835
rect 9930 -8955 9975 -8835
rect 10095 -8955 10140 -8835
rect 10260 -8955 10305 -8835
rect 10425 -8955 10480 -8835
rect 10600 -8955 10645 -8835
rect 10765 -8955 10810 -8835
rect 10930 -8955 10975 -8835
rect 11095 -8955 11150 -8835
rect 11270 -8955 11315 -8835
rect 11435 -8955 11480 -8835
rect 11600 -8955 11645 -8835
rect 11765 -8955 11820 -8835
rect 11940 -8955 11985 -8835
rect 12105 -8955 12150 -8835
rect 12270 -8955 12315 -8835
rect 12435 -8955 12490 -8835
rect 12610 -8955 12620 -8835
rect 7120 -9000 12620 -8955
rect 7120 -9120 7130 -9000
rect 7250 -9120 7295 -9000
rect 7415 -9120 7460 -9000
rect 7580 -9120 7625 -9000
rect 7745 -9120 7800 -9000
rect 7920 -9120 7965 -9000
rect 8085 -9120 8130 -9000
rect 8250 -9120 8295 -9000
rect 8415 -9120 8470 -9000
rect 8590 -9120 8635 -9000
rect 8755 -9120 8800 -9000
rect 8920 -9120 8965 -9000
rect 9085 -9120 9140 -9000
rect 9260 -9120 9305 -9000
rect 9425 -9120 9470 -9000
rect 9590 -9120 9635 -9000
rect 9755 -9120 9810 -9000
rect 9930 -9120 9975 -9000
rect 10095 -9120 10140 -9000
rect 10260 -9120 10305 -9000
rect 10425 -9120 10480 -9000
rect 10600 -9120 10645 -9000
rect 10765 -9120 10810 -9000
rect 10930 -9120 10975 -9000
rect 11095 -9120 11150 -9000
rect 11270 -9120 11315 -9000
rect 11435 -9120 11480 -9000
rect 11600 -9120 11645 -9000
rect 11765 -9120 11820 -9000
rect 11940 -9120 11985 -9000
rect 12105 -9120 12150 -9000
rect 12270 -9120 12315 -9000
rect 12435 -9120 12490 -9000
rect 12610 -9120 12620 -9000
rect 7120 -9175 12620 -9120
rect 7120 -9295 7130 -9175
rect 7250 -9295 7295 -9175
rect 7415 -9295 7460 -9175
rect 7580 -9295 7625 -9175
rect 7745 -9295 7800 -9175
rect 7920 -9295 7965 -9175
rect 8085 -9295 8130 -9175
rect 8250 -9295 8295 -9175
rect 8415 -9295 8470 -9175
rect 8590 -9295 8635 -9175
rect 8755 -9295 8800 -9175
rect 8920 -9295 8965 -9175
rect 9085 -9295 9140 -9175
rect 9260 -9295 9305 -9175
rect 9425 -9295 9470 -9175
rect 9590 -9295 9635 -9175
rect 9755 -9295 9810 -9175
rect 9930 -9295 9975 -9175
rect 10095 -9295 10140 -9175
rect 10260 -9295 10305 -9175
rect 10425 -9295 10480 -9175
rect 10600 -9295 10645 -9175
rect 10765 -9295 10810 -9175
rect 10930 -9295 10975 -9175
rect 11095 -9295 11150 -9175
rect 11270 -9295 11315 -9175
rect 11435 -9295 11480 -9175
rect 11600 -9295 11645 -9175
rect 11765 -9295 11820 -9175
rect 11940 -9295 11985 -9175
rect 12105 -9295 12150 -9175
rect 12270 -9295 12315 -9175
rect 12435 -9295 12490 -9175
rect 12610 -9295 12620 -9175
rect 7120 -9340 12620 -9295
rect 7120 -9460 7130 -9340
rect 7250 -9460 7295 -9340
rect 7415 -9460 7460 -9340
rect 7580 -9460 7625 -9340
rect 7745 -9460 7800 -9340
rect 7920 -9460 7965 -9340
rect 8085 -9460 8130 -9340
rect 8250 -9460 8295 -9340
rect 8415 -9460 8470 -9340
rect 8590 -9460 8635 -9340
rect 8755 -9460 8800 -9340
rect 8920 -9460 8965 -9340
rect 9085 -9460 9140 -9340
rect 9260 -9460 9305 -9340
rect 9425 -9460 9470 -9340
rect 9590 -9460 9635 -9340
rect 9755 -9460 9810 -9340
rect 9930 -9460 9975 -9340
rect 10095 -9460 10140 -9340
rect 10260 -9460 10305 -9340
rect 10425 -9460 10480 -9340
rect 10600 -9460 10645 -9340
rect 10765 -9460 10810 -9340
rect 10930 -9460 10975 -9340
rect 11095 -9460 11150 -9340
rect 11270 -9460 11315 -9340
rect 11435 -9460 11480 -9340
rect 11600 -9460 11645 -9340
rect 11765 -9460 11820 -9340
rect 11940 -9460 11985 -9340
rect 12105 -9460 12150 -9340
rect 12270 -9460 12315 -9340
rect 12435 -9460 12490 -9340
rect 12610 -9460 12620 -9340
rect 7120 -9505 12620 -9460
rect 7120 -9625 7130 -9505
rect 7250 -9625 7295 -9505
rect 7415 -9625 7460 -9505
rect 7580 -9625 7625 -9505
rect 7745 -9625 7800 -9505
rect 7920 -9625 7965 -9505
rect 8085 -9625 8130 -9505
rect 8250 -9625 8295 -9505
rect 8415 -9625 8470 -9505
rect 8590 -9625 8635 -9505
rect 8755 -9625 8800 -9505
rect 8920 -9625 8965 -9505
rect 9085 -9625 9140 -9505
rect 9260 -9625 9305 -9505
rect 9425 -9625 9470 -9505
rect 9590 -9625 9635 -9505
rect 9755 -9625 9810 -9505
rect 9930 -9625 9975 -9505
rect 10095 -9625 10140 -9505
rect 10260 -9625 10305 -9505
rect 10425 -9625 10480 -9505
rect 10600 -9625 10645 -9505
rect 10765 -9625 10810 -9505
rect 10930 -9625 10975 -9505
rect 11095 -9625 11150 -9505
rect 11270 -9625 11315 -9505
rect 11435 -9625 11480 -9505
rect 11600 -9625 11645 -9505
rect 11765 -9625 11820 -9505
rect 11940 -9625 11985 -9505
rect 12105 -9625 12150 -9505
rect 12270 -9625 12315 -9505
rect 12435 -9625 12490 -9505
rect 12610 -9625 12620 -9505
rect 7120 -9670 12620 -9625
rect 7120 -9790 7130 -9670
rect 7250 -9790 7295 -9670
rect 7415 -9790 7460 -9670
rect 7580 -9790 7625 -9670
rect 7745 -9790 7800 -9670
rect 7920 -9790 7965 -9670
rect 8085 -9790 8130 -9670
rect 8250 -9790 8295 -9670
rect 8415 -9790 8470 -9670
rect 8590 -9790 8635 -9670
rect 8755 -9790 8800 -9670
rect 8920 -9790 8965 -9670
rect 9085 -9790 9140 -9670
rect 9260 -9790 9305 -9670
rect 9425 -9790 9470 -9670
rect 9590 -9790 9635 -9670
rect 9755 -9790 9810 -9670
rect 9930 -9790 9975 -9670
rect 10095 -9790 10140 -9670
rect 10260 -9790 10305 -9670
rect 10425 -9790 10480 -9670
rect 10600 -9790 10645 -9670
rect 10765 -9790 10810 -9670
rect 10930 -9790 10975 -9670
rect 11095 -9790 11150 -9670
rect 11270 -9790 11315 -9670
rect 11435 -9790 11480 -9670
rect 11600 -9790 11645 -9670
rect 11765 -9790 11820 -9670
rect 11940 -9790 11985 -9670
rect 12105 -9790 12150 -9670
rect 12270 -9790 12315 -9670
rect 12435 -9790 12490 -9670
rect 12610 -9790 12620 -9670
rect 7120 -9800 12620 -9790
rect 12810 -4310 18310 -4300
rect 12810 -4430 12820 -4310
rect 12940 -4430 12985 -4310
rect 13105 -4430 13150 -4310
rect 13270 -4430 13315 -4310
rect 13435 -4430 13490 -4310
rect 13610 -4430 13655 -4310
rect 13775 -4430 13820 -4310
rect 13940 -4430 13985 -4310
rect 14105 -4430 14160 -4310
rect 14280 -4430 14325 -4310
rect 14445 -4430 14490 -4310
rect 14610 -4430 14655 -4310
rect 14775 -4430 14830 -4310
rect 14950 -4430 14995 -4310
rect 15115 -4430 15160 -4310
rect 15280 -4430 15325 -4310
rect 15445 -4430 15500 -4310
rect 15620 -4430 15665 -4310
rect 15785 -4430 15830 -4310
rect 15950 -4430 15995 -4310
rect 16115 -4430 16170 -4310
rect 16290 -4430 16335 -4310
rect 16455 -4430 16500 -4310
rect 16620 -4430 16665 -4310
rect 16785 -4430 16840 -4310
rect 16960 -4430 17005 -4310
rect 17125 -4430 17170 -4310
rect 17290 -4430 17335 -4310
rect 17455 -4430 17510 -4310
rect 17630 -4430 17675 -4310
rect 17795 -4430 17840 -4310
rect 17960 -4430 18005 -4310
rect 18125 -4430 18180 -4310
rect 18300 -4430 18310 -4310
rect 12810 -4485 18310 -4430
rect 12810 -4605 12820 -4485
rect 12940 -4605 12985 -4485
rect 13105 -4605 13150 -4485
rect 13270 -4605 13315 -4485
rect 13435 -4605 13490 -4485
rect 13610 -4605 13655 -4485
rect 13775 -4605 13820 -4485
rect 13940 -4605 13985 -4485
rect 14105 -4605 14160 -4485
rect 14280 -4605 14325 -4485
rect 14445 -4605 14490 -4485
rect 14610 -4605 14655 -4485
rect 14775 -4605 14830 -4485
rect 14950 -4605 14995 -4485
rect 15115 -4605 15160 -4485
rect 15280 -4605 15325 -4485
rect 15445 -4605 15500 -4485
rect 15620 -4605 15665 -4485
rect 15785 -4605 15830 -4485
rect 15950 -4605 15995 -4485
rect 16115 -4605 16170 -4485
rect 16290 -4605 16335 -4485
rect 16455 -4605 16500 -4485
rect 16620 -4605 16665 -4485
rect 16785 -4605 16840 -4485
rect 16960 -4605 17005 -4485
rect 17125 -4605 17170 -4485
rect 17290 -4605 17335 -4485
rect 17455 -4605 17510 -4485
rect 17630 -4605 17675 -4485
rect 17795 -4605 17840 -4485
rect 17960 -4605 18005 -4485
rect 18125 -4605 18180 -4485
rect 18300 -4605 18310 -4485
rect 12810 -4650 18310 -4605
rect 12810 -4770 12820 -4650
rect 12940 -4770 12985 -4650
rect 13105 -4770 13150 -4650
rect 13270 -4770 13315 -4650
rect 13435 -4770 13490 -4650
rect 13610 -4770 13655 -4650
rect 13775 -4770 13820 -4650
rect 13940 -4770 13985 -4650
rect 14105 -4770 14160 -4650
rect 14280 -4770 14325 -4650
rect 14445 -4770 14490 -4650
rect 14610 -4770 14655 -4650
rect 14775 -4770 14830 -4650
rect 14950 -4770 14995 -4650
rect 15115 -4770 15160 -4650
rect 15280 -4770 15325 -4650
rect 15445 -4770 15500 -4650
rect 15620 -4770 15665 -4650
rect 15785 -4770 15830 -4650
rect 15950 -4770 15995 -4650
rect 16115 -4770 16170 -4650
rect 16290 -4770 16335 -4650
rect 16455 -4770 16500 -4650
rect 16620 -4770 16665 -4650
rect 16785 -4770 16840 -4650
rect 16960 -4770 17005 -4650
rect 17125 -4770 17170 -4650
rect 17290 -4770 17335 -4650
rect 17455 -4770 17510 -4650
rect 17630 -4770 17675 -4650
rect 17795 -4770 17840 -4650
rect 17960 -4770 18005 -4650
rect 18125 -4770 18180 -4650
rect 18300 -4770 18310 -4650
rect 12810 -4815 18310 -4770
rect 12810 -4935 12820 -4815
rect 12940 -4935 12985 -4815
rect 13105 -4935 13150 -4815
rect 13270 -4935 13315 -4815
rect 13435 -4935 13490 -4815
rect 13610 -4935 13655 -4815
rect 13775 -4935 13820 -4815
rect 13940 -4935 13985 -4815
rect 14105 -4935 14160 -4815
rect 14280 -4935 14325 -4815
rect 14445 -4935 14490 -4815
rect 14610 -4935 14655 -4815
rect 14775 -4935 14830 -4815
rect 14950 -4935 14995 -4815
rect 15115 -4935 15160 -4815
rect 15280 -4935 15325 -4815
rect 15445 -4935 15500 -4815
rect 15620 -4935 15665 -4815
rect 15785 -4935 15830 -4815
rect 15950 -4935 15995 -4815
rect 16115 -4935 16170 -4815
rect 16290 -4935 16335 -4815
rect 16455 -4935 16500 -4815
rect 16620 -4935 16665 -4815
rect 16785 -4935 16840 -4815
rect 16960 -4935 17005 -4815
rect 17125 -4935 17170 -4815
rect 17290 -4935 17335 -4815
rect 17455 -4935 17510 -4815
rect 17630 -4935 17675 -4815
rect 17795 -4935 17840 -4815
rect 17960 -4935 18005 -4815
rect 18125 -4935 18180 -4815
rect 18300 -4935 18310 -4815
rect 12810 -4980 18310 -4935
rect 12810 -5100 12820 -4980
rect 12940 -5100 12985 -4980
rect 13105 -5100 13150 -4980
rect 13270 -5100 13315 -4980
rect 13435 -5100 13490 -4980
rect 13610 -5100 13655 -4980
rect 13775 -5100 13820 -4980
rect 13940 -5100 13985 -4980
rect 14105 -5100 14160 -4980
rect 14280 -5100 14325 -4980
rect 14445 -5100 14490 -4980
rect 14610 -5100 14655 -4980
rect 14775 -5100 14830 -4980
rect 14950 -5100 14995 -4980
rect 15115 -5100 15160 -4980
rect 15280 -5100 15325 -4980
rect 15445 -5100 15500 -4980
rect 15620 -5100 15665 -4980
rect 15785 -5100 15830 -4980
rect 15950 -5100 15995 -4980
rect 16115 -5100 16170 -4980
rect 16290 -5100 16335 -4980
rect 16455 -5100 16500 -4980
rect 16620 -5100 16665 -4980
rect 16785 -5100 16840 -4980
rect 16960 -5100 17005 -4980
rect 17125 -5100 17170 -4980
rect 17290 -5100 17335 -4980
rect 17455 -5100 17510 -4980
rect 17630 -5100 17675 -4980
rect 17795 -5100 17840 -4980
rect 17960 -5100 18005 -4980
rect 18125 -5100 18180 -4980
rect 18300 -5100 18310 -4980
rect 12810 -5155 18310 -5100
rect 12810 -5275 12820 -5155
rect 12940 -5275 12985 -5155
rect 13105 -5275 13150 -5155
rect 13270 -5275 13315 -5155
rect 13435 -5275 13490 -5155
rect 13610 -5275 13655 -5155
rect 13775 -5275 13820 -5155
rect 13940 -5275 13985 -5155
rect 14105 -5275 14160 -5155
rect 14280 -5275 14325 -5155
rect 14445 -5275 14490 -5155
rect 14610 -5275 14655 -5155
rect 14775 -5275 14830 -5155
rect 14950 -5275 14995 -5155
rect 15115 -5275 15160 -5155
rect 15280 -5275 15325 -5155
rect 15445 -5275 15500 -5155
rect 15620 -5275 15665 -5155
rect 15785 -5275 15830 -5155
rect 15950 -5275 15995 -5155
rect 16115 -5275 16170 -5155
rect 16290 -5275 16335 -5155
rect 16455 -5275 16500 -5155
rect 16620 -5275 16665 -5155
rect 16785 -5275 16840 -5155
rect 16960 -5275 17005 -5155
rect 17125 -5275 17170 -5155
rect 17290 -5275 17335 -5155
rect 17455 -5275 17510 -5155
rect 17630 -5275 17675 -5155
rect 17795 -5275 17840 -5155
rect 17960 -5275 18005 -5155
rect 18125 -5275 18180 -5155
rect 18300 -5275 18310 -5155
rect 12810 -5320 18310 -5275
rect 12810 -5440 12820 -5320
rect 12940 -5440 12985 -5320
rect 13105 -5440 13150 -5320
rect 13270 -5440 13315 -5320
rect 13435 -5440 13490 -5320
rect 13610 -5440 13655 -5320
rect 13775 -5440 13820 -5320
rect 13940 -5440 13985 -5320
rect 14105 -5440 14160 -5320
rect 14280 -5440 14325 -5320
rect 14445 -5440 14490 -5320
rect 14610 -5440 14655 -5320
rect 14775 -5440 14830 -5320
rect 14950 -5440 14995 -5320
rect 15115 -5440 15160 -5320
rect 15280 -5440 15325 -5320
rect 15445 -5440 15500 -5320
rect 15620 -5440 15665 -5320
rect 15785 -5440 15830 -5320
rect 15950 -5440 15995 -5320
rect 16115 -5440 16170 -5320
rect 16290 -5440 16335 -5320
rect 16455 -5440 16500 -5320
rect 16620 -5440 16665 -5320
rect 16785 -5440 16840 -5320
rect 16960 -5440 17005 -5320
rect 17125 -5440 17170 -5320
rect 17290 -5440 17335 -5320
rect 17455 -5440 17510 -5320
rect 17630 -5440 17675 -5320
rect 17795 -5440 17840 -5320
rect 17960 -5440 18005 -5320
rect 18125 -5440 18180 -5320
rect 18300 -5440 18310 -5320
rect 12810 -5485 18310 -5440
rect 12810 -5605 12820 -5485
rect 12940 -5605 12985 -5485
rect 13105 -5605 13150 -5485
rect 13270 -5605 13315 -5485
rect 13435 -5605 13490 -5485
rect 13610 -5605 13655 -5485
rect 13775 -5605 13820 -5485
rect 13940 -5605 13985 -5485
rect 14105 -5605 14160 -5485
rect 14280 -5605 14325 -5485
rect 14445 -5605 14490 -5485
rect 14610 -5605 14655 -5485
rect 14775 -5605 14830 -5485
rect 14950 -5605 14995 -5485
rect 15115 -5605 15160 -5485
rect 15280 -5605 15325 -5485
rect 15445 -5605 15500 -5485
rect 15620 -5605 15665 -5485
rect 15785 -5605 15830 -5485
rect 15950 -5605 15995 -5485
rect 16115 -5605 16170 -5485
rect 16290 -5605 16335 -5485
rect 16455 -5605 16500 -5485
rect 16620 -5605 16665 -5485
rect 16785 -5605 16840 -5485
rect 16960 -5605 17005 -5485
rect 17125 -5605 17170 -5485
rect 17290 -5605 17335 -5485
rect 17455 -5605 17510 -5485
rect 17630 -5605 17675 -5485
rect 17795 -5605 17840 -5485
rect 17960 -5605 18005 -5485
rect 18125 -5605 18180 -5485
rect 18300 -5605 18310 -5485
rect 12810 -5650 18310 -5605
rect 12810 -5770 12820 -5650
rect 12940 -5770 12985 -5650
rect 13105 -5770 13150 -5650
rect 13270 -5770 13315 -5650
rect 13435 -5770 13490 -5650
rect 13610 -5770 13655 -5650
rect 13775 -5770 13820 -5650
rect 13940 -5770 13985 -5650
rect 14105 -5770 14160 -5650
rect 14280 -5770 14325 -5650
rect 14445 -5770 14490 -5650
rect 14610 -5770 14655 -5650
rect 14775 -5770 14830 -5650
rect 14950 -5770 14995 -5650
rect 15115 -5770 15160 -5650
rect 15280 -5770 15325 -5650
rect 15445 -5770 15500 -5650
rect 15620 -5770 15665 -5650
rect 15785 -5770 15830 -5650
rect 15950 -5770 15995 -5650
rect 16115 -5770 16170 -5650
rect 16290 -5770 16335 -5650
rect 16455 -5770 16500 -5650
rect 16620 -5770 16665 -5650
rect 16785 -5770 16840 -5650
rect 16960 -5770 17005 -5650
rect 17125 -5770 17170 -5650
rect 17290 -5770 17335 -5650
rect 17455 -5770 17510 -5650
rect 17630 -5770 17675 -5650
rect 17795 -5770 17840 -5650
rect 17960 -5770 18005 -5650
rect 18125 -5770 18180 -5650
rect 18300 -5770 18310 -5650
rect 12810 -5825 18310 -5770
rect 12810 -5945 12820 -5825
rect 12940 -5945 12985 -5825
rect 13105 -5945 13150 -5825
rect 13270 -5945 13315 -5825
rect 13435 -5945 13490 -5825
rect 13610 -5945 13655 -5825
rect 13775 -5945 13820 -5825
rect 13940 -5945 13985 -5825
rect 14105 -5945 14160 -5825
rect 14280 -5945 14325 -5825
rect 14445 -5945 14490 -5825
rect 14610 -5945 14655 -5825
rect 14775 -5945 14830 -5825
rect 14950 -5945 14995 -5825
rect 15115 -5945 15160 -5825
rect 15280 -5945 15325 -5825
rect 15445 -5945 15500 -5825
rect 15620 -5945 15665 -5825
rect 15785 -5945 15830 -5825
rect 15950 -5945 15995 -5825
rect 16115 -5945 16170 -5825
rect 16290 -5945 16335 -5825
rect 16455 -5945 16500 -5825
rect 16620 -5945 16665 -5825
rect 16785 -5945 16840 -5825
rect 16960 -5945 17005 -5825
rect 17125 -5945 17170 -5825
rect 17290 -5945 17335 -5825
rect 17455 -5945 17510 -5825
rect 17630 -5945 17675 -5825
rect 17795 -5945 17840 -5825
rect 17960 -5945 18005 -5825
rect 18125 -5945 18180 -5825
rect 18300 -5945 18310 -5825
rect 12810 -5990 18310 -5945
rect 12810 -6110 12820 -5990
rect 12940 -6110 12985 -5990
rect 13105 -6110 13150 -5990
rect 13270 -6110 13315 -5990
rect 13435 -6110 13490 -5990
rect 13610 -6110 13655 -5990
rect 13775 -6110 13820 -5990
rect 13940 -6110 13985 -5990
rect 14105 -6110 14160 -5990
rect 14280 -6110 14325 -5990
rect 14445 -6110 14490 -5990
rect 14610 -6110 14655 -5990
rect 14775 -6110 14830 -5990
rect 14950 -6110 14995 -5990
rect 15115 -6110 15160 -5990
rect 15280 -6110 15325 -5990
rect 15445 -6110 15500 -5990
rect 15620 -6110 15665 -5990
rect 15785 -6110 15830 -5990
rect 15950 -6110 15995 -5990
rect 16115 -6110 16170 -5990
rect 16290 -6110 16335 -5990
rect 16455 -6110 16500 -5990
rect 16620 -6110 16665 -5990
rect 16785 -6110 16840 -5990
rect 16960 -6110 17005 -5990
rect 17125 -6110 17170 -5990
rect 17290 -6110 17335 -5990
rect 17455 -6110 17510 -5990
rect 17630 -6110 17675 -5990
rect 17795 -6110 17840 -5990
rect 17960 -6110 18005 -5990
rect 18125 -6110 18180 -5990
rect 18300 -6110 18310 -5990
rect 12810 -6155 18310 -6110
rect 12810 -6275 12820 -6155
rect 12940 -6275 12985 -6155
rect 13105 -6275 13150 -6155
rect 13270 -6275 13315 -6155
rect 13435 -6275 13490 -6155
rect 13610 -6275 13655 -6155
rect 13775 -6275 13820 -6155
rect 13940 -6275 13985 -6155
rect 14105 -6275 14160 -6155
rect 14280 -6275 14325 -6155
rect 14445 -6275 14490 -6155
rect 14610 -6275 14655 -6155
rect 14775 -6275 14830 -6155
rect 14950 -6275 14995 -6155
rect 15115 -6275 15160 -6155
rect 15280 -6275 15325 -6155
rect 15445 -6275 15500 -6155
rect 15620 -6275 15665 -6155
rect 15785 -6275 15830 -6155
rect 15950 -6275 15995 -6155
rect 16115 -6275 16170 -6155
rect 16290 -6275 16335 -6155
rect 16455 -6275 16500 -6155
rect 16620 -6275 16665 -6155
rect 16785 -6275 16840 -6155
rect 16960 -6275 17005 -6155
rect 17125 -6275 17170 -6155
rect 17290 -6275 17335 -6155
rect 17455 -6275 17510 -6155
rect 17630 -6275 17675 -6155
rect 17795 -6275 17840 -6155
rect 17960 -6275 18005 -6155
rect 18125 -6275 18180 -6155
rect 18300 -6275 18310 -6155
rect 12810 -6320 18310 -6275
rect 12810 -6440 12820 -6320
rect 12940 -6440 12985 -6320
rect 13105 -6440 13150 -6320
rect 13270 -6440 13315 -6320
rect 13435 -6440 13490 -6320
rect 13610 -6440 13655 -6320
rect 13775 -6440 13820 -6320
rect 13940 -6440 13985 -6320
rect 14105 -6440 14160 -6320
rect 14280 -6440 14325 -6320
rect 14445 -6440 14490 -6320
rect 14610 -6440 14655 -6320
rect 14775 -6440 14830 -6320
rect 14950 -6440 14995 -6320
rect 15115 -6440 15160 -6320
rect 15280 -6440 15325 -6320
rect 15445 -6440 15500 -6320
rect 15620 -6440 15665 -6320
rect 15785 -6440 15830 -6320
rect 15950 -6440 15995 -6320
rect 16115 -6440 16170 -6320
rect 16290 -6440 16335 -6320
rect 16455 -6440 16500 -6320
rect 16620 -6440 16665 -6320
rect 16785 -6440 16840 -6320
rect 16960 -6440 17005 -6320
rect 17125 -6440 17170 -6320
rect 17290 -6440 17335 -6320
rect 17455 -6440 17510 -6320
rect 17630 -6440 17675 -6320
rect 17795 -6440 17840 -6320
rect 17960 -6440 18005 -6320
rect 18125 -6440 18180 -6320
rect 18300 -6440 18310 -6320
rect 12810 -6495 18310 -6440
rect 12810 -6615 12820 -6495
rect 12940 -6615 12985 -6495
rect 13105 -6615 13150 -6495
rect 13270 -6615 13315 -6495
rect 13435 -6615 13490 -6495
rect 13610 -6615 13655 -6495
rect 13775 -6615 13820 -6495
rect 13940 -6615 13985 -6495
rect 14105 -6615 14160 -6495
rect 14280 -6615 14325 -6495
rect 14445 -6615 14490 -6495
rect 14610 -6615 14655 -6495
rect 14775 -6615 14830 -6495
rect 14950 -6615 14995 -6495
rect 15115 -6615 15160 -6495
rect 15280 -6615 15325 -6495
rect 15445 -6615 15500 -6495
rect 15620 -6615 15665 -6495
rect 15785 -6615 15830 -6495
rect 15950 -6615 15995 -6495
rect 16115 -6615 16170 -6495
rect 16290 -6615 16335 -6495
rect 16455 -6615 16500 -6495
rect 16620 -6615 16665 -6495
rect 16785 -6615 16840 -6495
rect 16960 -6615 17005 -6495
rect 17125 -6615 17170 -6495
rect 17290 -6615 17335 -6495
rect 17455 -6615 17510 -6495
rect 17630 -6615 17675 -6495
rect 17795 -6615 17840 -6495
rect 17960 -6615 18005 -6495
rect 18125 -6615 18180 -6495
rect 18300 -6615 18310 -6495
rect 12810 -6660 18310 -6615
rect 12810 -6780 12820 -6660
rect 12940 -6780 12985 -6660
rect 13105 -6780 13150 -6660
rect 13270 -6780 13315 -6660
rect 13435 -6780 13490 -6660
rect 13610 -6780 13655 -6660
rect 13775 -6780 13820 -6660
rect 13940 -6780 13985 -6660
rect 14105 -6780 14160 -6660
rect 14280 -6780 14325 -6660
rect 14445 -6780 14490 -6660
rect 14610 -6780 14655 -6660
rect 14775 -6780 14830 -6660
rect 14950 -6780 14995 -6660
rect 15115 -6780 15160 -6660
rect 15280 -6780 15325 -6660
rect 15445 -6780 15500 -6660
rect 15620 -6780 15665 -6660
rect 15785 -6780 15830 -6660
rect 15950 -6780 15995 -6660
rect 16115 -6780 16170 -6660
rect 16290 -6780 16335 -6660
rect 16455 -6780 16500 -6660
rect 16620 -6780 16665 -6660
rect 16785 -6780 16840 -6660
rect 16960 -6780 17005 -6660
rect 17125 -6780 17170 -6660
rect 17290 -6780 17335 -6660
rect 17455 -6780 17510 -6660
rect 17630 -6780 17675 -6660
rect 17795 -6780 17840 -6660
rect 17960 -6780 18005 -6660
rect 18125 -6780 18180 -6660
rect 18300 -6780 18310 -6660
rect 12810 -6825 18310 -6780
rect 12810 -6945 12820 -6825
rect 12940 -6945 12985 -6825
rect 13105 -6945 13150 -6825
rect 13270 -6945 13315 -6825
rect 13435 -6945 13490 -6825
rect 13610 -6945 13655 -6825
rect 13775 -6945 13820 -6825
rect 13940 -6945 13985 -6825
rect 14105 -6945 14160 -6825
rect 14280 -6945 14325 -6825
rect 14445 -6945 14490 -6825
rect 14610 -6945 14655 -6825
rect 14775 -6945 14830 -6825
rect 14950 -6945 14995 -6825
rect 15115 -6945 15160 -6825
rect 15280 -6945 15325 -6825
rect 15445 -6945 15500 -6825
rect 15620 -6945 15665 -6825
rect 15785 -6945 15830 -6825
rect 15950 -6945 15995 -6825
rect 16115 -6945 16170 -6825
rect 16290 -6945 16335 -6825
rect 16455 -6945 16500 -6825
rect 16620 -6945 16665 -6825
rect 16785 -6945 16840 -6825
rect 16960 -6945 17005 -6825
rect 17125 -6945 17170 -6825
rect 17290 -6945 17335 -6825
rect 17455 -6945 17510 -6825
rect 17630 -6945 17675 -6825
rect 17795 -6945 17840 -6825
rect 17960 -6945 18005 -6825
rect 18125 -6945 18180 -6825
rect 18300 -6945 18310 -6825
rect 12810 -6990 18310 -6945
rect 12810 -7110 12820 -6990
rect 12940 -7110 12985 -6990
rect 13105 -7110 13150 -6990
rect 13270 -7110 13315 -6990
rect 13435 -7110 13490 -6990
rect 13610 -7110 13655 -6990
rect 13775 -7110 13820 -6990
rect 13940 -7110 13985 -6990
rect 14105 -7110 14160 -6990
rect 14280 -7110 14325 -6990
rect 14445 -7110 14490 -6990
rect 14610 -7110 14655 -6990
rect 14775 -7110 14830 -6990
rect 14950 -7110 14995 -6990
rect 15115 -7110 15160 -6990
rect 15280 -7110 15325 -6990
rect 15445 -7110 15500 -6990
rect 15620 -7110 15665 -6990
rect 15785 -7110 15830 -6990
rect 15950 -7110 15995 -6990
rect 16115 -7110 16170 -6990
rect 16290 -7110 16335 -6990
rect 16455 -7110 16500 -6990
rect 16620 -7110 16665 -6990
rect 16785 -7110 16840 -6990
rect 16960 -7110 17005 -6990
rect 17125 -7110 17170 -6990
rect 17290 -7110 17335 -6990
rect 17455 -7110 17510 -6990
rect 17630 -7110 17675 -6990
rect 17795 -7110 17840 -6990
rect 17960 -7110 18005 -6990
rect 18125 -7110 18180 -6990
rect 18300 -7110 18310 -6990
rect 12810 -7165 18310 -7110
rect 12810 -7285 12820 -7165
rect 12940 -7285 12985 -7165
rect 13105 -7285 13150 -7165
rect 13270 -7285 13315 -7165
rect 13435 -7285 13490 -7165
rect 13610 -7285 13655 -7165
rect 13775 -7285 13820 -7165
rect 13940 -7285 13985 -7165
rect 14105 -7285 14160 -7165
rect 14280 -7285 14325 -7165
rect 14445 -7285 14490 -7165
rect 14610 -7285 14655 -7165
rect 14775 -7285 14830 -7165
rect 14950 -7285 14995 -7165
rect 15115 -7285 15160 -7165
rect 15280 -7285 15325 -7165
rect 15445 -7285 15500 -7165
rect 15620 -7285 15665 -7165
rect 15785 -7285 15830 -7165
rect 15950 -7285 15995 -7165
rect 16115 -7285 16170 -7165
rect 16290 -7285 16335 -7165
rect 16455 -7285 16500 -7165
rect 16620 -7285 16665 -7165
rect 16785 -7285 16840 -7165
rect 16960 -7285 17005 -7165
rect 17125 -7285 17170 -7165
rect 17290 -7285 17335 -7165
rect 17455 -7285 17510 -7165
rect 17630 -7285 17675 -7165
rect 17795 -7285 17840 -7165
rect 17960 -7285 18005 -7165
rect 18125 -7285 18180 -7165
rect 18300 -7285 18310 -7165
rect 12810 -7330 18310 -7285
rect 12810 -7450 12820 -7330
rect 12940 -7450 12985 -7330
rect 13105 -7450 13150 -7330
rect 13270 -7450 13315 -7330
rect 13435 -7450 13490 -7330
rect 13610 -7450 13655 -7330
rect 13775 -7450 13820 -7330
rect 13940 -7450 13985 -7330
rect 14105 -7450 14160 -7330
rect 14280 -7450 14325 -7330
rect 14445 -7450 14490 -7330
rect 14610 -7450 14655 -7330
rect 14775 -7450 14830 -7330
rect 14950 -7450 14995 -7330
rect 15115 -7450 15160 -7330
rect 15280 -7450 15325 -7330
rect 15445 -7450 15500 -7330
rect 15620 -7450 15665 -7330
rect 15785 -7450 15830 -7330
rect 15950 -7450 15995 -7330
rect 16115 -7450 16170 -7330
rect 16290 -7450 16335 -7330
rect 16455 -7450 16500 -7330
rect 16620 -7450 16665 -7330
rect 16785 -7450 16840 -7330
rect 16960 -7450 17005 -7330
rect 17125 -7450 17170 -7330
rect 17290 -7450 17335 -7330
rect 17455 -7450 17510 -7330
rect 17630 -7450 17675 -7330
rect 17795 -7450 17840 -7330
rect 17960 -7450 18005 -7330
rect 18125 -7450 18180 -7330
rect 18300 -7450 18310 -7330
rect 12810 -7495 18310 -7450
rect 12810 -7615 12820 -7495
rect 12940 -7615 12985 -7495
rect 13105 -7615 13150 -7495
rect 13270 -7615 13315 -7495
rect 13435 -7615 13490 -7495
rect 13610 -7615 13655 -7495
rect 13775 -7615 13820 -7495
rect 13940 -7615 13985 -7495
rect 14105 -7615 14160 -7495
rect 14280 -7615 14325 -7495
rect 14445 -7615 14490 -7495
rect 14610 -7615 14655 -7495
rect 14775 -7615 14830 -7495
rect 14950 -7615 14995 -7495
rect 15115 -7615 15160 -7495
rect 15280 -7615 15325 -7495
rect 15445 -7615 15500 -7495
rect 15620 -7615 15665 -7495
rect 15785 -7615 15830 -7495
rect 15950 -7615 15995 -7495
rect 16115 -7615 16170 -7495
rect 16290 -7615 16335 -7495
rect 16455 -7615 16500 -7495
rect 16620 -7615 16665 -7495
rect 16785 -7615 16840 -7495
rect 16960 -7615 17005 -7495
rect 17125 -7615 17170 -7495
rect 17290 -7615 17335 -7495
rect 17455 -7615 17510 -7495
rect 17630 -7615 17675 -7495
rect 17795 -7615 17840 -7495
rect 17960 -7615 18005 -7495
rect 18125 -7615 18180 -7495
rect 18300 -7615 18310 -7495
rect 12810 -7660 18310 -7615
rect 12810 -7780 12820 -7660
rect 12940 -7780 12985 -7660
rect 13105 -7780 13150 -7660
rect 13270 -7780 13315 -7660
rect 13435 -7780 13490 -7660
rect 13610 -7780 13655 -7660
rect 13775 -7780 13820 -7660
rect 13940 -7780 13985 -7660
rect 14105 -7780 14160 -7660
rect 14280 -7780 14325 -7660
rect 14445 -7780 14490 -7660
rect 14610 -7780 14655 -7660
rect 14775 -7780 14830 -7660
rect 14950 -7780 14995 -7660
rect 15115 -7780 15160 -7660
rect 15280 -7780 15325 -7660
rect 15445 -7780 15500 -7660
rect 15620 -7780 15665 -7660
rect 15785 -7780 15830 -7660
rect 15950 -7780 15995 -7660
rect 16115 -7780 16170 -7660
rect 16290 -7780 16335 -7660
rect 16455 -7780 16500 -7660
rect 16620 -7780 16665 -7660
rect 16785 -7780 16840 -7660
rect 16960 -7780 17005 -7660
rect 17125 -7780 17170 -7660
rect 17290 -7780 17335 -7660
rect 17455 -7780 17510 -7660
rect 17630 -7780 17675 -7660
rect 17795 -7780 17840 -7660
rect 17960 -7780 18005 -7660
rect 18125 -7780 18180 -7660
rect 18300 -7780 18310 -7660
rect 12810 -7835 18310 -7780
rect 12810 -7955 12820 -7835
rect 12940 -7955 12985 -7835
rect 13105 -7955 13150 -7835
rect 13270 -7955 13315 -7835
rect 13435 -7955 13490 -7835
rect 13610 -7955 13655 -7835
rect 13775 -7955 13820 -7835
rect 13940 -7955 13985 -7835
rect 14105 -7955 14160 -7835
rect 14280 -7955 14325 -7835
rect 14445 -7955 14490 -7835
rect 14610 -7955 14655 -7835
rect 14775 -7955 14830 -7835
rect 14950 -7955 14995 -7835
rect 15115 -7955 15160 -7835
rect 15280 -7955 15325 -7835
rect 15445 -7955 15500 -7835
rect 15620 -7955 15665 -7835
rect 15785 -7955 15830 -7835
rect 15950 -7955 15995 -7835
rect 16115 -7955 16170 -7835
rect 16290 -7955 16335 -7835
rect 16455 -7955 16500 -7835
rect 16620 -7955 16665 -7835
rect 16785 -7955 16840 -7835
rect 16960 -7955 17005 -7835
rect 17125 -7955 17170 -7835
rect 17290 -7955 17335 -7835
rect 17455 -7955 17510 -7835
rect 17630 -7955 17675 -7835
rect 17795 -7955 17840 -7835
rect 17960 -7955 18005 -7835
rect 18125 -7955 18180 -7835
rect 18300 -7955 18310 -7835
rect 12810 -8000 18310 -7955
rect 12810 -8120 12820 -8000
rect 12940 -8120 12985 -8000
rect 13105 -8120 13150 -8000
rect 13270 -8120 13315 -8000
rect 13435 -8120 13490 -8000
rect 13610 -8120 13655 -8000
rect 13775 -8120 13820 -8000
rect 13940 -8120 13985 -8000
rect 14105 -8120 14160 -8000
rect 14280 -8120 14325 -8000
rect 14445 -8120 14490 -8000
rect 14610 -8120 14655 -8000
rect 14775 -8120 14830 -8000
rect 14950 -8120 14995 -8000
rect 15115 -8120 15160 -8000
rect 15280 -8120 15325 -8000
rect 15445 -8120 15500 -8000
rect 15620 -8120 15665 -8000
rect 15785 -8120 15830 -8000
rect 15950 -8120 15995 -8000
rect 16115 -8120 16170 -8000
rect 16290 -8120 16335 -8000
rect 16455 -8120 16500 -8000
rect 16620 -8120 16665 -8000
rect 16785 -8120 16840 -8000
rect 16960 -8120 17005 -8000
rect 17125 -8120 17170 -8000
rect 17290 -8120 17335 -8000
rect 17455 -8120 17510 -8000
rect 17630 -8120 17675 -8000
rect 17795 -8120 17840 -8000
rect 17960 -8120 18005 -8000
rect 18125 -8120 18180 -8000
rect 18300 -8120 18310 -8000
rect 12810 -8165 18310 -8120
rect 12810 -8285 12820 -8165
rect 12940 -8285 12985 -8165
rect 13105 -8285 13150 -8165
rect 13270 -8285 13315 -8165
rect 13435 -8285 13490 -8165
rect 13610 -8285 13655 -8165
rect 13775 -8285 13820 -8165
rect 13940 -8285 13985 -8165
rect 14105 -8285 14160 -8165
rect 14280 -8285 14325 -8165
rect 14445 -8285 14490 -8165
rect 14610 -8285 14655 -8165
rect 14775 -8285 14830 -8165
rect 14950 -8285 14995 -8165
rect 15115 -8285 15160 -8165
rect 15280 -8285 15325 -8165
rect 15445 -8285 15500 -8165
rect 15620 -8285 15665 -8165
rect 15785 -8285 15830 -8165
rect 15950 -8285 15995 -8165
rect 16115 -8285 16170 -8165
rect 16290 -8285 16335 -8165
rect 16455 -8285 16500 -8165
rect 16620 -8285 16665 -8165
rect 16785 -8285 16840 -8165
rect 16960 -8285 17005 -8165
rect 17125 -8285 17170 -8165
rect 17290 -8285 17335 -8165
rect 17455 -8285 17510 -8165
rect 17630 -8285 17675 -8165
rect 17795 -8285 17840 -8165
rect 17960 -8285 18005 -8165
rect 18125 -8285 18180 -8165
rect 18300 -8285 18310 -8165
rect 12810 -8330 18310 -8285
rect 12810 -8450 12820 -8330
rect 12940 -8450 12985 -8330
rect 13105 -8450 13150 -8330
rect 13270 -8450 13315 -8330
rect 13435 -8450 13490 -8330
rect 13610 -8450 13655 -8330
rect 13775 -8450 13820 -8330
rect 13940 -8450 13985 -8330
rect 14105 -8450 14160 -8330
rect 14280 -8450 14325 -8330
rect 14445 -8450 14490 -8330
rect 14610 -8450 14655 -8330
rect 14775 -8450 14830 -8330
rect 14950 -8450 14995 -8330
rect 15115 -8450 15160 -8330
rect 15280 -8450 15325 -8330
rect 15445 -8450 15500 -8330
rect 15620 -8450 15665 -8330
rect 15785 -8450 15830 -8330
rect 15950 -8450 15995 -8330
rect 16115 -8450 16170 -8330
rect 16290 -8450 16335 -8330
rect 16455 -8450 16500 -8330
rect 16620 -8450 16665 -8330
rect 16785 -8450 16840 -8330
rect 16960 -8450 17005 -8330
rect 17125 -8450 17170 -8330
rect 17290 -8450 17335 -8330
rect 17455 -8450 17510 -8330
rect 17630 -8450 17675 -8330
rect 17795 -8450 17840 -8330
rect 17960 -8450 18005 -8330
rect 18125 -8450 18180 -8330
rect 18300 -8450 18310 -8330
rect 12810 -8505 18310 -8450
rect 12810 -8625 12820 -8505
rect 12940 -8625 12985 -8505
rect 13105 -8625 13150 -8505
rect 13270 -8625 13315 -8505
rect 13435 -8625 13490 -8505
rect 13610 -8625 13655 -8505
rect 13775 -8625 13820 -8505
rect 13940 -8625 13985 -8505
rect 14105 -8625 14160 -8505
rect 14280 -8625 14325 -8505
rect 14445 -8625 14490 -8505
rect 14610 -8625 14655 -8505
rect 14775 -8625 14830 -8505
rect 14950 -8625 14995 -8505
rect 15115 -8625 15160 -8505
rect 15280 -8625 15325 -8505
rect 15445 -8625 15500 -8505
rect 15620 -8625 15665 -8505
rect 15785 -8625 15830 -8505
rect 15950 -8625 15995 -8505
rect 16115 -8625 16170 -8505
rect 16290 -8625 16335 -8505
rect 16455 -8625 16500 -8505
rect 16620 -8625 16665 -8505
rect 16785 -8625 16840 -8505
rect 16960 -8625 17005 -8505
rect 17125 -8625 17170 -8505
rect 17290 -8625 17335 -8505
rect 17455 -8625 17510 -8505
rect 17630 -8625 17675 -8505
rect 17795 -8625 17840 -8505
rect 17960 -8625 18005 -8505
rect 18125 -8625 18180 -8505
rect 18300 -8625 18310 -8505
rect 12810 -8670 18310 -8625
rect 12810 -8790 12820 -8670
rect 12940 -8790 12985 -8670
rect 13105 -8790 13150 -8670
rect 13270 -8790 13315 -8670
rect 13435 -8790 13490 -8670
rect 13610 -8790 13655 -8670
rect 13775 -8790 13820 -8670
rect 13940 -8790 13985 -8670
rect 14105 -8790 14160 -8670
rect 14280 -8790 14325 -8670
rect 14445 -8790 14490 -8670
rect 14610 -8790 14655 -8670
rect 14775 -8790 14830 -8670
rect 14950 -8790 14995 -8670
rect 15115 -8790 15160 -8670
rect 15280 -8790 15325 -8670
rect 15445 -8790 15500 -8670
rect 15620 -8790 15665 -8670
rect 15785 -8790 15830 -8670
rect 15950 -8790 15995 -8670
rect 16115 -8790 16170 -8670
rect 16290 -8790 16335 -8670
rect 16455 -8790 16500 -8670
rect 16620 -8790 16665 -8670
rect 16785 -8790 16840 -8670
rect 16960 -8790 17005 -8670
rect 17125 -8790 17170 -8670
rect 17290 -8790 17335 -8670
rect 17455 -8790 17510 -8670
rect 17630 -8790 17675 -8670
rect 17795 -8790 17840 -8670
rect 17960 -8790 18005 -8670
rect 18125 -8790 18180 -8670
rect 18300 -8790 18310 -8670
rect 12810 -8835 18310 -8790
rect 12810 -8955 12820 -8835
rect 12940 -8955 12985 -8835
rect 13105 -8955 13150 -8835
rect 13270 -8955 13315 -8835
rect 13435 -8955 13490 -8835
rect 13610 -8955 13655 -8835
rect 13775 -8955 13820 -8835
rect 13940 -8955 13985 -8835
rect 14105 -8955 14160 -8835
rect 14280 -8955 14325 -8835
rect 14445 -8955 14490 -8835
rect 14610 -8955 14655 -8835
rect 14775 -8955 14830 -8835
rect 14950 -8955 14995 -8835
rect 15115 -8955 15160 -8835
rect 15280 -8955 15325 -8835
rect 15445 -8955 15500 -8835
rect 15620 -8955 15665 -8835
rect 15785 -8955 15830 -8835
rect 15950 -8955 15995 -8835
rect 16115 -8955 16170 -8835
rect 16290 -8955 16335 -8835
rect 16455 -8955 16500 -8835
rect 16620 -8955 16665 -8835
rect 16785 -8955 16840 -8835
rect 16960 -8955 17005 -8835
rect 17125 -8955 17170 -8835
rect 17290 -8955 17335 -8835
rect 17455 -8955 17510 -8835
rect 17630 -8955 17675 -8835
rect 17795 -8955 17840 -8835
rect 17960 -8955 18005 -8835
rect 18125 -8955 18180 -8835
rect 18300 -8955 18310 -8835
rect 12810 -9000 18310 -8955
rect 12810 -9120 12820 -9000
rect 12940 -9120 12985 -9000
rect 13105 -9120 13150 -9000
rect 13270 -9120 13315 -9000
rect 13435 -9120 13490 -9000
rect 13610 -9120 13655 -9000
rect 13775 -9120 13820 -9000
rect 13940 -9120 13985 -9000
rect 14105 -9120 14160 -9000
rect 14280 -9120 14325 -9000
rect 14445 -9120 14490 -9000
rect 14610 -9120 14655 -9000
rect 14775 -9120 14830 -9000
rect 14950 -9120 14995 -9000
rect 15115 -9120 15160 -9000
rect 15280 -9120 15325 -9000
rect 15445 -9120 15500 -9000
rect 15620 -9120 15665 -9000
rect 15785 -9120 15830 -9000
rect 15950 -9120 15995 -9000
rect 16115 -9120 16170 -9000
rect 16290 -9120 16335 -9000
rect 16455 -9120 16500 -9000
rect 16620 -9120 16665 -9000
rect 16785 -9120 16840 -9000
rect 16960 -9120 17005 -9000
rect 17125 -9120 17170 -9000
rect 17290 -9120 17335 -9000
rect 17455 -9120 17510 -9000
rect 17630 -9120 17675 -9000
rect 17795 -9120 17840 -9000
rect 17960 -9120 18005 -9000
rect 18125 -9120 18180 -9000
rect 18300 -9120 18310 -9000
rect 12810 -9175 18310 -9120
rect 12810 -9295 12820 -9175
rect 12940 -9295 12985 -9175
rect 13105 -9295 13150 -9175
rect 13270 -9295 13315 -9175
rect 13435 -9295 13490 -9175
rect 13610 -9295 13655 -9175
rect 13775 -9295 13820 -9175
rect 13940 -9295 13985 -9175
rect 14105 -9295 14160 -9175
rect 14280 -9295 14325 -9175
rect 14445 -9295 14490 -9175
rect 14610 -9295 14655 -9175
rect 14775 -9295 14830 -9175
rect 14950 -9295 14995 -9175
rect 15115 -9295 15160 -9175
rect 15280 -9295 15325 -9175
rect 15445 -9295 15500 -9175
rect 15620 -9295 15665 -9175
rect 15785 -9295 15830 -9175
rect 15950 -9295 15995 -9175
rect 16115 -9295 16170 -9175
rect 16290 -9295 16335 -9175
rect 16455 -9295 16500 -9175
rect 16620 -9295 16665 -9175
rect 16785 -9295 16840 -9175
rect 16960 -9295 17005 -9175
rect 17125 -9295 17170 -9175
rect 17290 -9295 17335 -9175
rect 17455 -9295 17510 -9175
rect 17630 -9295 17675 -9175
rect 17795 -9295 17840 -9175
rect 17960 -9295 18005 -9175
rect 18125 -9295 18180 -9175
rect 18300 -9295 18310 -9175
rect 12810 -9340 18310 -9295
rect 12810 -9460 12820 -9340
rect 12940 -9460 12985 -9340
rect 13105 -9460 13150 -9340
rect 13270 -9460 13315 -9340
rect 13435 -9460 13490 -9340
rect 13610 -9460 13655 -9340
rect 13775 -9460 13820 -9340
rect 13940 -9460 13985 -9340
rect 14105 -9460 14160 -9340
rect 14280 -9460 14325 -9340
rect 14445 -9460 14490 -9340
rect 14610 -9460 14655 -9340
rect 14775 -9460 14830 -9340
rect 14950 -9460 14995 -9340
rect 15115 -9460 15160 -9340
rect 15280 -9460 15325 -9340
rect 15445 -9460 15500 -9340
rect 15620 -9460 15665 -9340
rect 15785 -9460 15830 -9340
rect 15950 -9460 15995 -9340
rect 16115 -9460 16170 -9340
rect 16290 -9460 16335 -9340
rect 16455 -9460 16500 -9340
rect 16620 -9460 16665 -9340
rect 16785 -9460 16840 -9340
rect 16960 -9460 17005 -9340
rect 17125 -9460 17170 -9340
rect 17290 -9460 17335 -9340
rect 17455 -9460 17510 -9340
rect 17630 -9460 17675 -9340
rect 17795 -9460 17840 -9340
rect 17960 -9460 18005 -9340
rect 18125 -9460 18180 -9340
rect 18300 -9460 18310 -9340
rect 12810 -9505 18310 -9460
rect 12810 -9625 12820 -9505
rect 12940 -9625 12985 -9505
rect 13105 -9625 13150 -9505
rect 13270 -9625 13315 -9505
rect 13435 -9625 13490 -9505
rect 13610 -9625 13655 -9505
rect 13775 -9625 13820 -9505
rect 13940 -9625 13985 -9505
rect 14105 -9625 14160 -9505
rect 14280 -9625 14325 -9505
rect 14445 -9625 14490 -9505
rect 14610 -9625 14655 -9505
rect 14775 -9625 14830 -9505
rect 14950 -9625 14995 -9505
rect 15115 -9625 15160 -9505
rect 15280 -9625 15325 -9505
rect 15445 -9625 15500 -9505
rect 15620 -9625 15665 -9505
rect 15785 -9625 15830 -9505
rect 15950 -9625 15995 -9505
rect 16115 -9625 16170 -9505
rect 16290 -9625 16335 -9505
rect 16455 -9625 16500 -9505
rect 16620 -9625 16665 -9505
rect 16785 -9625 16840 -9505
rect 16960 -9625 17005 -9505
rect 17125 -9625 17170 -9505
rect 17290 -9625 17335 -9505
rect 17455 -9625 17510 -9505
rect 17630 -9625 17675 -9505
rect 17795 -9625 17840 -9505
rect 17960 -9625 18005 -9505
rect 18125 -9625 18180 -9505
rect 18300 -9625 18310 -9505
rect 12810 -9670 18310 -9625
rect 12810 -9790 12820 -9670
rect 12940 -9790 12985 -9670
rect 13105 -9790 13150 -9670
rect 13270 -9790 13315 -9670
rect 13435 -9790 13490 -9670
rect 13610 -9790 13655 -9670
rect 13775 -9790 13820 -9670
rect 13940 -9790 13985 -9670
rect 14105 -9790 14160 -9670
rect 14280 -9790 14325 -9670
rect 14445 -9790 14490 -9670
rect 14610 -9790 14655 -9670
rect 14775 -9790 14830 -9670
rect 14950 -9790 14995 -9670
rect 15115 -9790 15160 -9670
rect 15280 -9790 15325 -9670
rect 15445 -9790 15500 -9670
rect 15620 -9790 15665 -9670
rect 15785 -9790 15830 -9670
rect 15950 -9790 15995 -9670
rect 16115 -9790 16170 -9670
rect 16290 -9790 16335 -9670
rect 16455 -9790 16500 -9670
rect 16620 -9790 16665 -9670
rect 16785 -9790 16840 -9670
rect 16960 -9790 17005 -9670
rect 17125 -9790 17170 -9670
rect 17290 -9790 17335 -9670
rect 17455 -9790 17510 -9670
rect 17630 -9790 17675 -9670
rect 17795 -9790 17840 -9670
rect 17960 -9790 18005 -9670
rect 18125 -9790 18180 -9670
rect 18300 -9790 18310 -9670
rect 12810 -9800 18310 -9790
rect 18500 -4310 24000 -4300
rect 18500 -4430 18510 -4310
rect 18630 -4430 18675 -4310
rect 18795 -4430 18840 -4310
rect 18960 -4430 19005 -4310
rect 19125 -4430 19180 -4310
rect 19300 -4430 19345 -4310
rect 19465 -4430 19510 -4310
rect 19630 -4430 19675 -4310
rect 19795 -4430 19850 -4310
rect 19970 -4430 20015 -4310
rect 20135 -4430 20180 -4310
rect 20300 -4430 20345 -4310
rect 20465 -4430 20520 -4310
rect 20640 -4430 20685 -4310
rect 20805 -4430 20850 -4310
rect 20970 -4430 21015 -4310
rect 21135 -4430 21190 -4310
rect 21310 -4430 21355 -4310
rect 21475 -4430 21520 -4310
rect 21640 -4430 21685 -4310
rect 21805 -4430 21860 -4310
rect 21980 -4430 22025 -4310
rect 22145 -4430 22190 -4310
rect 22310 -4430 22355 -4310
rect 22475 -4430 22530 -4310
rect 22650 -4430 22695 -4310
rect 22815 -4430 22860 -4310
rect 22980 -4430 23025 -4310
rect 23145 -4430 23200 -4310
rect 23320 -4430 23365 -4310
rect 23485 -4430 23530 -4310
rect 23650 -4430 23695 -4310
rect 23815 -4430 23870 -4310
rect 23990 -4430 24000 -4310
rect 18500 -4485 24000 -4430
rect 18500 -4605 18510 -4485
rect 18630 -4605 18675 -4485
rect 18795 -4605 18840 -4485
rect 18960 -4605 19005 -4485
rect 19125 -4605 19180 -4485
rect 19300 -4605 19345 -4485
rect 19465 -4605 19510 -4485
rect 19630 -4605 19675 -4485
rect 19795 -4605 19850 -4485
rect 19970 -4605 20015 -4485
rect 20135 -4605 20180 -4485
rect 20300 -4605 20345 -4485
rect 20465 -4605 20520 -4485
rect 20640 -4605 20685 -4485
rect 20805 -4605 20850 -4485
rect 20970 -4605 21015 -4485
rect 21135 -4605 21190 -4485
rect 21310 -4605 21355 -4485
rect 21475 -4605 21520 -4485
rect 21640 -4605 21685 -4485
rect 21805 -4605 21860 -4485
rect 21980 -4605 22025 -4485
rect 22145 -4605 22190 -4485
rect 22310 -4605 22355 -4485
rect 22475 -4605 22530 -4485
rect 22650 -4605 22695 -4485
rect 22815 -4605 22860 -4485
rect 22980 -4605 23025 -4485
rect 23145 -4605 23200 -4485
rect 23320 -4605 23365 -4485
rect 23485 -4605 23530 -4485
rect 23650 -4605 23695 -4485
rect 23815 -4605 23870 -4485
rect 23990 -4605 24000 -4485
rect 18500 -4650 24000 -4605
rect 18500 -4770 18510 -4650
rect 18630 -4770 18675 -4650
rect 18795 -4770 18840 -4650
rect 18960 -4770 19005 -4650
rect 19125 -4770 19180 -4650
rect 19300 -4770 19345 -4650
rect 19465 -4770 19510 -4650
rect 19630 -4770 19675 -4650
rect 19795 -4770 19850 -4650
rect 19970 -4770 20015 -4650
rect 20135 -4770 20180 -4650
rect 20300 -4770 20345 -4650
rect 20465 -4770 20520 -4650
rect 20640 -4770 20685 -4650
rect 20805 -4770 20850 -4650
rect 20970 -4770 21015 -4650
rect 21135 -4770 21190 -4650
rect 21310 -4770 21355 -4650
rect 21475 -4770 21520 -4650
rect 21640 -4770 21685 -4650
rect 21805 -4770 21860 -4650
rect 21980 -4770 22025 -4650
rect 22145 -4770 22190 -4650
rect 22310 -4770 22355 -4650
rect 22475 -4770 22530 -4650
rect 22650 -4770 22695 -4650
rect 22815 -4770 22860 -4650
rect 22980 -4770 23025 -4650
rect 23145 -4770 23200 -4650
rect 23320 -4770 23365 -4650
rect 23485 -4770 23530 -4650
rect 23650 -4770 23695 -4650
rect 23815 -4770 23870 -4650
rect 23990 -4770 24000 -4650
rect 18500 -4815 24000 -4770
rect 18500 -4935 18510 -4815
rect 18630 -4935 18675 -4815
rect 18795 -4935 18840 -4815
rect 18960 -4935 19005 -4815
rect 19125 -4935 19180 -4815
rect 19300 -4935 19345 -4815
rect 19465 -4935 19510 -4815
rect 19630 -4935 19675 -4815
rect 19795 -4935 19850 -4815
rect 19970 -4935 20015 -4815
rect 20135 -4935 20180 -4815
rect 20300 -4935 20345 -4815
rect 20465 -4935 20520 -4815
rect 20640 -4935 20685 -4815
rect 20805 -4935 20850 -4815
rect 20970 -4935 21015 -4815
rect 21135 -4935 21190 -4815
rect 21310 -4935 21355 -4815
rect 21475 -4935 21520 -4815
rect 21640 -4935 21685 -4815
rect 21805 -4935 21860 -4815
rect 21980 -4935 22025 -4815
rect 22145 -4935 22190 -4815
rect 22310 -4935 22355 -4815
rect 22475 -4935 22530 -4815
rect 22650 -4935 22695 -4815
rect 22815 -4935 22860 -4815
rect 22980 -4935 23025 -4815
rect 23145 -4935 23200 -4815
rect 23320 -4935 23365 -4815
rect 23485 -4935 23530 -4815
rect 23650 -4935 23695 -4815
rect 23815 -4935 23870 -4815
rect 23990 -4935 24000 -4815
rect 18500 -4980 24000 -4935
rect 18500 -5100 18510 -4980
rect 18630 -5100 18675 -4980
rect 18795 -5100 18840 -4980
rect 18960 -5100 19005 -4980
rect 19125 -5100 19180 -4980
rect 19300 -5100 19345 -4980
rect 19465 -5100 19510 -4980
rect 19630 -5100 19675 -4980
rect 19795 -5100 19850 -4980
rect 19970 -5100 20015 -4980
rect 20135 -5100 20180 -4980
rect 20300 -5100 20345 -4980
rect 20465 -5100 20520 -4980
rect 20640 -5100 20685 -4980
rect 20805 -5100 20850 -4980
rect 20970 -5100 21015 -4980
rect 21135 -5100 21190 -4980
rect 21310 -5100 21355 -4980
rect 21475 -5100 21520 -4980
rect 21640 -5100 21685 -4980
rect 21805 -5100 21860 -4980
rect 21980 -5100 22025 -4980
rect 22145 -5100 22190 -4980
rect 22310 -5100 22355 -4980
rect 22475 -5100 22530 -4980
rect 22650 -5100 22695 -4980
rect 22815 -5100 22860 -4980
rect 22980 -5100 23025 -4980
rect 23145 -5100 23200 -4980
rect 23320 -5100 23365 -4980
rect 23485 -5100 23530 -4980
rect 23650 -5100 23695 -4980
rect 23815 -5100 23870 -4980
rect 23990 -5100 24000 -4980
rect 18500 -5155 24000 -5100
rect 18500 -5275 18510 -5155
rect 18630 -5275 18675 -5155
rect 18795 -5275 18840 -5155
rect 18960 -5275 19005 -5155
rect 19125 -5275 19180 -5155
rect 19300 -5275 19345 -5155
rect 19465 -5275 19510 -5155
rect 19630 -5275 19675 -5155
rect 19795 -5275 19850 -5155
rect 19970 -5275 20015 -5155
rect 20135 -5275 20180 -5155
rect 20300 -5275 20345 -5155
rect 20465 -5275 20520 -5155
rect 20640 -5275 20685 -5155
rect 20805 -5275 20850 -5155
rect 20970 -5275 21015 -5155
rect 21135 -5275 21190 -5155
rect 21310 -5275 21355 -5155
rect 21475 -5275 21520 -5155
rect 21640 -5275 21685 -5155
rect 21805 -5275 21860 -5155
rect 21980 -5275 22025 -5155
rect 22145 -5275 22190 -5155
rect 22310 -5275 22355 -5155
rect 22475 -5275 22530 -5155
rect 22650 -5275 22695 -5155
rect 22815 -5275 22860 -5155
rect 22980 -5275 23025 -5155
rect 23145 -5275 23200 -5155
rect 23320 -5275 23365 -5155
rect 23485 -5275 23530 -5155
rect 23650 -5275 23695 -5155
rect 23815 -5275 23870 -5155
rect 23990 -5275 24000 -5155
rect 18500 -5320 24000 -5275
rect 18500 -5440 18510 -5320
rect 18630 -5440 18675 -5320
rect 18795 -5440 18840 -5320
rect 18960 -5440 19005 -5320
rect 19125 -5440 19180 -5320
rect 19300 -5440 19345 -5320
rect 19465 -5440 19510 -5320
rect 19630 -5440 19675 -5320
rect 19795 -5440 19850 -5320
rect 19970 -5440 20015 -5320
rect 20135 -5440 20180 -5320
rect 20300 -5440 20345 -5320
rect 20465 -5440 20520 -5320
rect 20640 -5440 20685 -5320
rect 20805 -5440 20850 -5320
rect 20970 -5440 21015 -5320
rect 21135 -5440 21190 -5320
rect 21310 -5440 21355 -5320
rect 21475 -5440 21520 -5320
rect 21640 -5440 21685 -5320
rect 21805 -5440 21860 -5320
rect 21980 -5440 22025 -5320
rect 22145 -5440 22190 -5320
rect 22310 -5440 22355 -5320
rect 22475 -5440 22530 -5320
rect 22650 -5440 22695 -5320
rect 22815 -5440 22860 -5320
rect 22980 -5440 23025 -5320
rect 23145 -5440 23200 -5320
rect 23320 -5440 23365 -5320
rect 23485 -5440 23530 -5320
rect 23650 -5440 23695 -5320
rect 23815 -5440 23870 -5320
rect 23990 -5440 24000 -5320
rect 18500 -5485 24000 -5440
rect 18500 -5605 18510 -5485
rect 18630 -5605 18675 -5485
rect 18795 -5605 18840 -5485
rect 18960 -5605 19005 -5485
rect 19125 -5605 19180 -5485
rect 19300 -5605 19345 -5485
rect 19465 -5605 19510 -5485
rect 19630 -5605 19675 -5485
rect 19795 -5605 19850 -5485
rect 19970 -5605 20015 -5485
rect 20135 -5605 20180 -5485
rect 20300 -5605 20345 -5485
rect 20465 -5605 20520 -5485
rect 20640 -5605 20685 -5485
rect 20805 -5605 20850 -5485
rect 20970 -5605 21015 -5485
rect 21135 -5605 21190 -5485
rect 21310 -5605 21355 -5485
rect 21475 -5605 21520 -5485
rect 21640 -5605 21685 -5485
rect 21805 -5605 21860 -5485
rect 21980 -5605 22025 -5485
rect 22145 -5605 22190 -5485
rect 22310 -5605 22355 -5485
rect 22475 -5605 22530 -5485
rect 22650 -5605 22695 -5485
rect 22815 -5605 22860 -5485
rect 22980 -5605 23025 -5485
rect 23145 -5605 23200 -5485
rect 23320 -5605 23365 -5485
rect 23485 -5605 23530 -5485
rect 23650 -5605 23695 -5485
rect 23815 -5605 23870 -5485
rect 23990 -5605 24000 -5485
rect 18500 -5650 24000 -5605
rect 18500 -5770 18510 -5650
rect 18630 -5770 18675 -5650
rect 18795 -5770 18840 -5650
rect 18960 -5770 19005 -5650
rect 19125 -5770 19180 -5650
rect 19300 -5770 19345 -5650
rect 19465 -5770 19510 -5650
rect 19630 -5770 19675 -5650
rect 19795 -5770 19850 -5650
rect 19970 -5770 20015 -5650
rect 20135 -5770 20180 -5650
rect 20300 -5770 20345 -5650
rect 20465 -5770 20520 -5650
rect 20640 -5770 20685 -5650
rect 20805 -5770 20850 -5650
rect 20970 -5770 21015 -5650
rect 21135 -5770 21190 -5650
rect 21310 -5770 21355 -5650
rect 21475 -5770 21520 -5650
rect 21640 -5770 21685 -5650
rect 21805 -5770 21860 -5650
rect 21980 -5770 22025 -5650
rect 22145 -5770 22190 -5650
rect 22310 -5770 22355 -5650
rect 22475 -5770 22530 -5650
rect 22650 -5770 22695 -5650
rect 22815 -5770 22860 -5650
rect 22980 -5770 23025 -5650
rect 23145 -5770 23200 -5650
rect 23320 -5770 23365 -5650
rect 23485 -5770 23530 -5650
rect 23650 -5770 23695 -5650
rect 23815 -5770 23870 -5650
rect 23990 -5770 24000 -5650
rect 18500 -5825 24000 -5770
rect 18500 -5945 18510 -5825
rect 18630 -5945 18675 -5825
rect 18795 -5945 18840 -5825
rect 18960 -5945 19005 -5825
rect 19125 -5945 19180 -5825
rect 19300 -5945 19345 -5825
rect 19465 -5945 19510 -5825
rect 19630 -5945 19675 -5825
rect 19795 -5945 19850 -5825
rect 19970 -5945 20015 -5825
rect 20135 -5945 20180 -5825
rect 20300 -5945 20345 -5825
rect 20465 -5945 20520 -5825
rect 20640 -5945 20685 -5825
rect 20805 -5945 20850 -5825
rect 20970 -5945 21015 -5825
rect 21135 -5945 21190 -5825
rect 21310 -5945 21355 -5825
rect 21475 -5945 21520 -5825
rect 21640 -5945 21685 -5825
rect 21805 -5945 21860 -5825
rect 21980 -5945 22025 -5825
rect 22145 -5945 22190 -5825
rect 22310 -5945 22355 -5825
rect 22475 -5945 22530 -5825
rect 22650 -5945 22695 -5825
rect 22815 -5945 22860 -5825
rect 22980 -5945 23025 -5825
rect 23145 -5945 23200 -5825
rect 23320 -5945 23365 -5825
rect 23485 -5945 23530 -5825
rect 23650 -5945 23695 -5825
rect 23815 -5945 23870 -5825
rect 23990 -5945 24000 -5825
rect 18500 -5990 24000 -5945
rect 18500 -6110 18510 -5990
rect 18630 -6110 18675 -5990
rect 18795 -6110 18840 -5990
rect 18960 -6110 19005 -5990
rect 19125 -6110 19180 -5990
rect 19300 -6110 19345 -5990
rect 19465 -6110 19510 -5990
rect 19630 -6110 19675 -5990
rect 19795 -6110 19850 -5990
rect 19970 -6110 20015 -5990
rect 20135 -6110 20180 -5990
rect 20300 -6110 20345 -5990
rect 20465 -6110 20520 -5990
rect 20640 -6110 20685 -5990
rect 20805 -6110 20850 -5990
rect 20970 -6110 21015 -5990
rect 21135 -6110 21190 -5990
rect 21310 -6110 21355 -5990
rect 21475 -6110 21520 -5990
rect 21640 -6110 21685 -5990
rect 21805 -6110 21860 -5990
rect 21980 -6110 22025 -5990
rect 22145 -6110 22190 -5990
rect 22310 -6110 22355 -5990
rect 22475 -6110 22530 -5990
rect 22650 -6110 22695 -5990
rect 22815 -6110 22860 -5990
rect 22980 -6110 23025 -5990
rect 23145 -6110 23200 -5990
rect 23320 -6110 23365 -5990
rect 23485 -6110 23530 -5990
rect 23650 -6110 23695 -5990
rect 23815 -6110 23870 -5990
rect 23990 -6110 24000 -5990
rect 18500 -6155 24000 -6110
rect 18500 -6275 18510 -6155
rect 18630 -6275 18675 -6155
rect 18795 -6275 18840 -6155
rect 18960 -6275 19005 -6155
rect 19125 -6275 19180 -6155
rect 19300 -6275 19345 -6155
rect 19465 -6275 19510 -6155
rect 19630 -6275 19675 -6155
rect 19795 -6275 19850 -6155
rect 19970 -6275 20015 -6155
rect 20135 -6275 20180 -6155
rect 20300 -6275 20345 -6155
rect 20465 -6275 20520 -6155
rect 20640 -6275 20685 -6155
rect 20805 -6275 20850 -6155
rect 20970 -6275 21015 -6155
rect 21135 -6275 21190 -6155
rect 21310 -6275 21355 -6155
rect 21475 -6275 21520 -6155
rect 21640 -6275 21685 -6155
rect 21805 -6275 21860 -6155
rect 21980 -6275 22025 -6155
rect 22145 -6275 22190 -6155
rect 22310 -6275 22355 -6155
rect 22475 -6275 22530 -6155
rect 22650 -6275 22695 -6155
rect 22815 -6275 22860 -6155
rect 22980 -6275 23025 -6155
rect 23145 -6275 23200 -6155
rect 23320 -6275 23365 -6155
rect 23485 -6275 23530 -6155
rect 23650 -6275 23695 -6155
rect 23815 -6275 23870 -6155
rect 23990 -6275 24000 -6155
rect 18500 -6320 24000 -6275
rect 18500 -6440 18510 -6320
rect 18630 -6440 18675 -6320
rect 18795 -6440 18840 -6320
rect 18960 -6440 19005 -6320
rect 19125 -6440 19180 -6320
rect 19300 -6440 19345 -6320
rect 19465 -6440 19510 -6320
rect 19630 -6440 19675 -6320
rect 19795 -6440 19850 -6320
rect 19970 -6440 20015 -6320
rect 20135 -6440 20180 -6320
rect 20300 -6440 20345 -6320
rect 20465 -6440 20520 -6320
rect 20640 -6440 20685 -6320
rect 20805 -6440 20850 -6320
rect 20970 -6440 21015 -6320
rect 21135 -6440 21190 -6320
rect 21310 -6440 21355 -6320
rect 21475 -6440 21520 -6320
rect 21640 -6440 21685 -6320
rect 21805 -6440 21860 -6320
rect 21980 -6440 22025 -6320
rect 22145 -6440 22190 -6320
rect 22310 -6440 22355 -6320
rect 22475 -6440 22530 -6320
rect 22650 -6440 22695 -6320
rect 22815 -6440 22860 -6320
rect 22980 -6440 23025 -6320
rect 23145 -6440 23200 -6320
rect 23320 -6440 23365 -6320
rect 23485 -6440 23530 -6320
rect 23650 -6440 23695 -6320
rect 23815 -6440 23870 -6320
rect 23990 -6440 24000 -6320
rect 18500 -6495 24000 -6440
rect 18500 -6615 18510 -6495
rect 18630 -6615 18675 -6495
rect 18795 -6615 18840 -6495
rect 18960 -6615 19005 -6495
rect 19125 -6615 19180 -6495
rect 19300 -6615 19345 -6495
rect 19465 -6615 19510 -6495
rect 19630 -6615 19675 -6495
rect 19795 -6615 19850 -6495
rect 19970 -6615 20015 -6495
rect 20135 -6615 20180 -6495
rect 20300 -6615 20345 -6495
rect 20465 -6615 20520 -6495
rect 20640 -6615 20685 -6495
rect 20805 -6615 20850 -6495
rect 20970 -6615 21015 -6495
rect 21135 -6615 21190 -6495
rect 21310 -6615 21355 -6495
rect 21475 -6615 21520 -6495
rect 21640 -6615 21685 -6495
rect 21805 -6615 21860 -6495
rect 21980 -6615 22025 -6495
rect 22145 -6615 22190 -6495
rect 22310 -6615 22355 -6495
rect 22475 -6615 22530 -6495
rect 22650 -6615 22695 -6495
rect 22815 -6615 22860 -6495
rect 22980 -6615 23025 -6495
rect 23145 -6615 23200 -6495
rect 23320 -6615 23365 -6495
rect 23485 -6615 23530 -6495
rect 23650 -6615 23695 -6495
rect 23815 -6615 23870 -6495
rect 23990 -6615 24000 -6495
rect 18500 -6660 24000 -6615
rect 18500 -6780 18510 -6660
rect 18630 -6780 18675 -6660
rect 18795 -6780 18840 -6660
rect 18960 -6780 19005 -6660
rect 19125 -6780 19180 -6660
rect 19300 -6780 19345 -6660
rect 19465 -6780 19510 -6660
rect 19630 -6780 19675 -6660
rect 19795 -6780 19850 -6660
rect 19970 -6780 20015 -6660
rect 20135 -6780 20180 -6660
rect 20300 -6780 20345 -6660
rect 20465 -6780 20520 -6660
rect 20640 -6780 20685 -6660
rect 20805 -6780 20850 -6660
rect 20970 -6780 21015 -6660
rect 21135 -6780 21190 -6660
rect 21310 -6780 21355 -6660
rect 21475 -6780 21520 -6660
rect 21640 -6780 21685 -6660
rect 21805 -6780 21860 -6660
rect 21980 -6780 22025 -6660
rect 22145 -6780 22190 -6660
rect 22310 -6780 22355 -6660
rect 22475 -6780 22530 -6660
rect 22650 -6780 22695 -6660
rect 22815 -6780 22860 -6660
rect 22980 -6780 23025 -6660
rect 23145 -6780 23200 -6660
rect 23320 -6780 23365 -6660
rect 23485 -6780 23530 -6660
rect 23650 -6780 23695 -6660
rect 23815 -6780 23870 -6660
rect 23990 -6780 24000 -6660
rect 18500 -6825 24000 -6780
rect 18500 -6945 18510 -6825
rect 18630 -6945 18675 -6825
rect 18795 -6945 18840 -6825
rect 18960 -6945 19005 -6825
rect 19125 -6945 19180 -6825
rect 19300 -6945 19345 -6825
rect 19465 -6945 19510 -6825
rect 19630 -6945 19675 -6825
rect 19795 -6945 19850 -6825
rect 19970 -6945 20015 -6825
rect 20135 -6945 20180 -6825
rect 20300 -6945 20345 -6825
rect 20465 -6945 20520 -6825
rect 20640 -6945 20685 -6825
rect 20805 -6945 20850 -6825
rect 20970 -6945 21015 -6825
rect 21135 -6945 21190 -6825
rect 21310 -6945 21355 -6825
rect 21475 -6945 21520 -6825
rect 21640 -6945 21685 -6825
rect 21805 -6945 21860 -6825
rect 21980 -6945 22025 -6825
rect 22145 -6945 22190 -6825
rect 22310 -6945 22355 -6825
rect 22475 -6945 22530 -6825
rect 22650 -6945 22695 -6825
rect 22815 -6945 22860 -6825
rect 22980 -6945 23025 -6825
rect 23145 -6945 23200 -6825
rect 23320 -6945 23365 -6825
rect 23485 -6945 23530 -6825
rect 23650 -6945 23695 -6825
rect 23815 -6945 23870 -6825
rect 23990 -6945 24000 -6825
rect 18500 -6990 24000 -6945
rect 18500 -7110 18510 -6990
rect 18630 -7110 18675 -6990
rect 18795 -7110 18840 -6990
rect 18960 -7110 19005 -6990
rect 19125 -7110 19180 -6990
rect 19300 -7110 19345 -6990
rect 19465 -7110 19510 -6990
rect 19630 -7110 19675 -6990
rect 19795 -7110 19850 -6990
rect 19970 -7110 20015 -6990
rect 20135 -7110 20180 -6990
rect 20300 -7110 20345 -6990
rect 20465 -7110 20520 -6990
rect 20640 -7110 20685 -6990
rect 20805 -7110 20850 -6990
rect 20970 -7110 21015 -6990
rect 21135 -7110 21190 -6990
rect 21310 -7110 21355 -6990
rect 21475 -7110 21520 -6990
rect 21640 -7110 21685 -6990
rect 21805 -7110 21860 -6990
rect 21980 -7110 22025 -6990
rect 22145 -7110 22190 -6990
rect 22310 -7110 22355 -6990
rect 22475 -7110 22530 -6990
rect 22650 -7110 22695 -6990
rect 22815 -7110 22860 -6990
rect 22980 -7110 23025 -6990
rect 23145 -7110 23200 -6990
rect 23320 -7110 23365 -6990
rect 23485 -7110 23530 -6990
rect 23650 -7110 23695 -6990
rect 23815 -7110 23870 -6990
rect 23990 -7110 24000 -6990
rect 18500 -7165 24000 -7110
rect 18500 -7285 18510 -7165
rect 18630 -7285 18675 -7165
rect 18795 -7285 18840 -7165
rect 18960 -7285 19005 -7165
rect 19125 -7285 19180 -7165
rect 19300 -7285 19345 -7165
rect 19465 -7285 19510 -7165
rect 19630 -7285 19675 -7165
rect 19795 -7285 19850 -7165
rect 19970 -7285 20015 -7165
rect 20135 -7285 20180 -7165
rect 20300 -7285 20345 -7165
rect 20465 -7285 20520 -7165
rect 20640 -7285 20685 -7165
rect 20805 -7285 20850 -7165
rect 20970 -7285 21015 -7165
rect 21135 -7285 21190 -7165
rect 21310 -7285 21355 -7165
rect 21475 -7285 21520 -7165
rect 21640 -7285 21685 -7165
rect 21805 -7285 21860 -7165
rect 21980 -7285 22025 -7165
rect 22145 -7285 22190 -7165
rect 22310 -7285 22355 -7165
rect 22475 -7285 22530 -7165
rect 22650 -7285 22695 -7165
rect 22815 -7285 22860 -7165
rect 22980 -7285 23025 -7165
rect 23145 -7285 23200 -7165
rect 23320 -7285 23365 -7165
rect 23485 -7285 23530 -7165
rect 23650 -7285 23695 -7165
rect 23815 -7285 23870 -7165
rect 23990 -7285 24000 -7165
rect 18500 -7330 24000 -7285
rect 18500 -7450 18510 -7330
rect 18630 -7450 18675 -7330
rect 18795 -7450 18840 -7330
rect 18960 -7450 19005 -7330
rect 19125 -7450 19180 -7330
rect 19300 -7450 19345 -7330
rect 19465 -7450 19510 -7330
rect 19630 -7450 19675 -7330
rect 19795 -7450 19850 -7330
rect 19970 -7450 20015 -7330
rect 20135 -7450 20180 -7330
rect 20300 -7450 20345 -7330
rect 20465 -7450 20520 -7330
rect 20640 -7450 20685 -7330
rect 20805 -7450 20850 -7330
rect 20970 -7450 21015 -7330
rect 21135 -7450 21190 -7330
rect 21310 -7450 21355 -7330
rect 21475 -7450 21520 -7330
rect 21640 -7450 21685 -7330
rect 21805 -7450 21860 -7330
rect 21980 -7450 22025 -7330
rect 22145 -7450 22190 -7330
rect 22310 -7450 22355 -7330
rect 22475 -7450 22530 -7330
rect 22650 -7450 22695 -7330
rect 22815 -7450 22860 -7330
rect 22980 -7450 23025 -7330
rect 23145 -7450 23200 -7330
rect 23320 -7450 23365 -7330
rect 23485 -7450 23530 -7330
rect 23650 -7450 23695 -7330
rect 23815 -7450 23870 -7330
rect 23990 -7450 24000 -7330
rect 18500 -7495 24000 -7450
rect 18500 -7615 18510 -7495
rect 18630 -7615 18675 -7495
rect 18795 -7615 18840 -7495
rect 18960 -7615 19005 -7495
rect 19125 -7615 19180 -7495
rect 19300 -7615 19345 -7495
rect 19465 -7615 19510 -7495
rect 19630 -7615 19675 -7495
rect 19795 -7615 19850 -7495
rect 19970 -7615 20015 -7495
rect 20135 -7615 20180 -7495
rect 20300 -7615 20345 -7495
rect 20465 -7615 20520 -7495
rect 20640 -7615 20685 -7495
rect 20805 -7615 20850 -7495
rect 20970 -7615 21015 -7495
rect 21135 -7615 21190 -7495
rect 21310 -7615 21355 -7495
rect 21475 -7615 21520 -7495
rect 21640 -7615 21685 -7495
rect 21805 -7615 21860 -7495
rect 21980 -7615 22025 -7495
rect 22145 -7615 22190 -7495
rect 22310 -7615 22355 -7495
rect 22475 -7615 22530 -7495
rect 22650 -7615 22695 -7495
rect 22815 -7615 22860 -7495
rect 22980 -7615 23025 -7495
rect 23145 -7615 23200 -7495
rect 23320 -7615 23365 -7495
rect 23485 -7615 23530 -7495
rect 23650 -7615 23695 -7495
rect 23815 -7615 23870 -7495
rect 23990 -7615 24000 -7495
rect 18500 -7660 24000 -7615
rect 18500 -7780 18510 -7660
rect 18630 -7780 18675 -7660
rect 18795 -7780 18840 -7660
rect 18960 -7780 19005 -7660
rect 19125 -7780 19180 -7660
rect 19300 -7780 19345 -7660
rect 19465 -7780 19510 -7660
rect 19630 -7780 19675 -7660
rect 19795 -7780 19850 -7660
rect 19970 -7780 20015 -7660
rect 20135 -7780 20180 -7660
rect 20300 -7780 20345 -7660
rect 20465 -7780 20520 -7660
rect 20640 -7780 20685 -7660
rect 20805 -7780 20850 -7660
rect 20970 -7780 21015 -7660
rect 21135 -7780 21190 -7660
rect 21310 -7780 21355 -7660
rect 21475 -7780 21520 -7660
rect 21640 -7780 21685 -7660
rect 21805 -7780 21860 -7660
rect 21980 -7780 22025 -7660
rect 22145 -7780 22190 -7660
rect 22310 -7780 22355 -7660
rect 22475 -7780 22530 -7660
rect 22650 -7780 22695 -7660
rect 22815 -7780 22860 -7660
rect 22980 -7780 23025 -7660
rect 23145 -7780 23200 -7660
rect 23320 -7780 23365 -7660
rect 23485 -7780 23530 -7660
rect 23650 -7780 23695 -7660
rect 23815 -7780 23870 -7660
rect 23990 -7780 24000 -7660
rect 18500 -7835 24000 -7780
rect 18500 -7955 18510 -7835
rect 18630 -7955 18675 -7835
rect 18795 -7955 18840 -7835
rect 18960 -7955 19005 -7835
rect 19125 -7955 19180 -7835
rect 19300 -7955 19345 -7835
rect 19465 -7955 19510 -7835
rect 19630 -7955 19675 -7835
rect 19795 -7955 19850 -7835
rect 19970 -7955 20015 -7835
rect 20135 -7955 20180 -7835
rect 20300 -7955 20345 -7835
rect 20465 -7955 20520 -7835
rect 20640 -7955 20685 -7835
rect 20805 -7955 20850 -7835
rect 20970 -7955 21015 -7835
rect 21135 -7955 21190 -7835
rect 21310 -7955 21355 -7835
rect 21475 -7955 21520 -7835
rect 21640 -7955 21685 -7835
rect 21805 -7955 21860 -7835
rect 21980 -7955 22025 -7835
rect 22145 -7955 22190 -7835
rect 22310 -7955 22355 -7835
rect 22475 -7955 22530 -7835
rect 22650 -7955 22695 -7835
rect 22815 -7955 22860 -7835
rect 22980 -7955 23025 -7835
rect 23145 -7955 23200 -7835
rect 23320 -7955 23365 -7835
rect 23485 -7955 23530 -7835
rect 23650 -7955 23695 -7835
rect 23815 -7955 23870 -7835
rect 23990 -7955 24000 -7835
rect 18500 -8000 24000 -7955
rect 18500 -8120 18510 -8000
rect 18630 -8120 18675 -8000
rect 18795 -8120 18840 -8000
rect 18960 -8120 19005 -8000
rect 19125 -8120 19180 -8000
rect 19300 -8120 19345 -8000
rect 19465 -8120 19510 -8000
rect 19630 -8120 19675 -8000
rect 19795 -8120 19850 -8000
rect 19970 -8120 20015 -8000
rect 20135 -8120 20180 -8000
rect 20300 -8120 20345 -8000
rect 20465 -8120 20520 -8000
rect 20640 -8120 20685 -8000
rect 20805 -8120 20850 -8000
rect 20970 -8120 21015 -8000
rect 21135 -8120 21190 -8000
rect 21310 -8120 21355 -8000
rect 21475 -8120 21520 -8000
rect 21640 -8120 21685 -8000
rect 21805 -8120 21860 -8000
rect 21980 -8120 22025 -8000
rect 22145 -8120 22190 -8000
rect 22310 -8120 22355 -8000
rect 22475 -8120 22530 -8000
rect 22650 -8120 22695 -8000
rect 22815 -8120 22860 -8000
rect 22980 -8120 23025 -8000
rect 23145 -8120 23200 -8000
rect 23320 -8120 23365 -8000
rect 23485 -8120 23530 -8000
rect 23650 -8120 23695 -8000
rect 23815 -8120 23870 -8000
rect 23990 -8120 24000 -8000
rect 18500 -8165 24000 -8120
rect 18500 -8285 18510 -8165
rect 18630 -8285 18675 -8165
rect 18795 -8285 18840 -8165
rect 18960 -8285 19005 -8165
rect 19125 -8285 19180 -8165
rect 19300 -8285 19345 -8165
rect 19465 -8285 19510 -8165
rect 19630 -8285 19675 -8165
rect 19795 -8285 19850 -8165
rect 19970 -8285 20015 -8165
rect 20135 -8285 20180 -8165
rect 20300 -8285 20345 -8165
rect 20465 -8285 20520 -8165
rect 20640 -8285 20685 -8165
rect 20805 -8285 20850 -8165
rect 20970 -8285 21015 -8165
rect 21135 -8285 21190 -8165
rect 21310 -8285 21355 -8165
rect 21475 -8285 21520 -8165
rect 21640 -8285 21685 -8165
rect 21805 -8285 21860 -8165
rect 21980 -8285 22025 -8165
rect 22145 -8285 22190 -8165
rect 22310 -8285 22355 -8165
rect 22475 -8285 22530 -8165
rect 22650 -8285 22695 -8165
rect 22815 -8285 22860 -8165
rect 22980 -8285 23025 -8165
rect 23145 -8285 23200 -8165
rect 23320 -8285 23365 -8165
rect 23485 -8285 23530 -8165
rect 23650 -8285 23695 -8165
rect 23815 -8285 23870 -8165
rect 23990 -8285 24000 -8165
rect 18500 -8330 24000 -8285
rect 18500 -8450 18510 -8330
rect 18630 -8450 18675 -8330
rect 18795 -8450 18840 -8330
rect 18960 -8450 19005 -8330
rect 19125 -8450 19180 -8330
rect 19300 -8450 19345 -8330
rect 19465 -8450 19510 -8330
rect 19630 -8450 19675 -8330
rect 19795 -8450 19850 -8330
rect 19970 -8450 20015 -8330
rect 20135 -8450 20180 -8330
rect 20300 -8450 20345 -8330
rect 20465 -8450 20520 -8330
rect 20640 -8450 20685 -8330
rect 20805 -8450 20850 -8330
rect 20970 -8450 21015 -8330
rect 21135 -8450 21190 -8330
rect 21310 -8450 21355 -8330
rect 21475 -8450 21520 -8330
rect 21640 -8450 21685 -8330
rect 21805 -8450 21860 -8330
rect 21980 -8450 22025 -8330
rect 22145 -8450 22190 -8330
rect 22310 -8450 22355 -8330
rect 22475 -8450 22530 -8330
rect 22650 -8450 22695 -8330
rect 22815 -8450 22860 -8330
rect 22980 -8450 23025 -8330
rect 23145 -8450 23200 -8330
rect 23320 -8450 23365 -8330
rect 23485 -8450 23530 -8330
rect 23650 -8450 23695 -8330
rect 23815 -8450 23870 -8330
rect 23990 -8450 24000 -8330
rect 18500 -8505 24000 -8450
rect 18500 -8625 18510 -8505
rect 18630 -8625 18675 -8505
rect 18795 -8625 18840 -8505
rect 18960 -8625 19005 -8505
rect 19125 -8625 19180 -8505
rect 19300 -8625 19345 -8505
rect 19465 -8625 19510 -8505
rect 19630 -8625 19675 -8505
rect 19795 -8625 19850 -8505
rect 19970 -8625 20015 -8505
rect 20135 -8625 20180 -8505
rect 20300 -8625 20345 -8505
rect 20465 -8625 20520 -8505
rect 20640 -8625 20685 -8505
rect 20805 -8625 20850 -8505
rect 20970 -8625 21015 -8505
rect 21135 -8625 21190 -8505
rect 21310 -8625 21355 -8505
rect 21475 -8625 21520 -8505
rect 21640 -8625 21685 -8505
rect 21805 -8625 21860 -8505
rect 21980 -8625 22025 -8505
rect 22145 -8625 22190 -8505
rect 22310 -8625 22355 -8505
rect 22475 -8625 22530 -8505
rect 22650 -8625 22695 -8505
rect 22815 -8625 22860 -8505
rect 22980 -8625 23025 -8505
rect 23145 -8625 23200 -8505
rect 23320 -8625 23365 -8505
rect 23485 -8625 23530 -8505
rect 23650 -8625 23695 -8505
rect 23815 -8625 23870 -8505
rect 23990 -8625 24000 -8505
rect 18500 -8670 24000 -8625
rect 18500 -8790 18510 -8670
rect 18630 -8790 18675 -8670
rect 18795 -8790 18840 -8670
rect 18960 -8790 19005 -8670
rect 19125 -8790 19180 -8670
rect 19300 -8790 19345 -8670
rect 19465 -8790 19510 -8670
rect 19630 -8790 19675 -8670
rect 19795 -8790 19850 -8670
rect 19970 -8790 20015 -8670
rect 20135 -8790 20180 -8670
rect 20300 -8790 20345 -8670
rect 20465 -8790 20520 -8670
rect 20640 -8790 20685 -8670
rect 20805 -8790 20850 -8670
rect 20970 -8790 21015 -8670
rect 21135 -8790 21190 -8670
rect 21310 -8790 21355 -8670
rect 21475 -8790 21520 -8670
rect 21640 -8790 21685 -8670
rect 21805 -8790 21860 -8670
rect 21980 -8790 22025 -8670
rect 22145 -8790 22190 -8670
rect 22310 -8790 22355 -8670
rect 22475 -8790 22530 -8670
rect 22650 -8790 22695 -8670
rect 22815 -8790 22860 -8670
rect 22980 -8790 23025 -8670
rect 23145 -8790 23200 -8670
rect 23320 -8790 23365 -8670
rect 23485 -8790 23530 -8670
rect 23650 -8790 23695 -8670
rect 23815 -8790 23870 -8670
rect 23990 -8790 24000 -8670
rect 18500 -8835 24000 -8790
rect 18500 -8955 18510 -8835
rect 18630 -8955 18675 -8835
rect 18795 -8955 18840 -8835
rect 18960 -8955 19005 -8835
rect 19125 -8955 19180 -8835
rect 19300 -8955 19345 -8835
rect 19465 -8955 19510 -8835
rect 19630 -8955 19675 -8835
rect 19795 -8955 19850 -8835
rect 19970 -8955 20015 -8835
rect 20135 -8955 20180 -8835
rect 20300 -8955 20345 -8835
rect 20465 -8955 20520 -8835
rect 20640 -8955 20685 -8835
rect 20805 -8955 20850 -8835
rect 20970 -8955 21015 -8835
rect 21135 -8955 21190 -8835
rect 21310 -8955 21355 -8835
rect 21475 -8955 21520 -8835
rect 21640 -8955 21685 -8835
rect 21805 -8955 21860 -8835
rect 21980 -8955 22025 -8835
rect 22145 -8955 22190 -8835
rect 22310 -8955 22355 -8835
rect 22475 -8955 22530 -8835
rect 22650 -8955 22695 -8835
rect 22815 -8955 22860 -8835
rect 22980 -8955 23025 -8835
rect 23145 -8955 23200 -8835
rect 23320 -8955 23365 -8835
rect 23485 -8955 23530 -8835
rect 23650 -8955 23695 -8835
rect 23815 -8955 23870 -8835
rect 23990 -8955 24000 -8835
rect 18500 -9000 24000 -8955
rect 18500 -9120 18510 -9000
rect 18630 -9120 18675 -9000
rect 18795 -9120 18840 -9000
rect 18960 -9120 19005 -9000
rect 19125 -9120 19180 -9000
rect 19300 -9120 19345 -9000
rect 19465 -9120 19510 -9000
rect 19630 -9120 19675 -9000
rect 19795 -9120 19850 -9000
rect 19970 -9120 20015 -9000
rect 20135 -9120 20180 -9000
rect 20300 -9120 20345 -9000
rect 20465 -9120 20520 -9000
rect 20640 -9120 20685 -9000
rect 20805 -9120 20850 -9000
rect 20970 -9120 21015 -9000
rect 21135 -9120 21190 -9000
rect 21310 -9120 21355 -9000
rect 21475 -9120 21520 -9000
rect 21640 -9120 21685 -9000
rect 21805 -9120 21860 -9000
rect 21980 -9120 22025 -9000
rect 22145 -9120 22190 -9000
rect 22310 -9120 22355 -9000
rect 22475 -9120 22530 -9000
rect 22650 -9120 22695 -9000
rect 22815 -9120 22860 -9000
rect 22980 -9120 23025 -9000
rect 23145 -9120 23200 -9000
rect 23320 -9120 23365 -9000
rect 23485 -9120 23530 -9000
rect 23650 -9120 23695 -9000
rect 23815 -9120 23870 -9000
rect 23990 -9120 24000 -9000
rect 18500 -9175 24000 -9120
rect 18500 -9295 18510 -9175
rect 18630 -9295 18675 -9175
rect 18795 -9295 18840 -9175
rect 18960 -9295 19005 -9175
rect 19125 -9295 19180 -9175
rect 19300 -9295 19345 -9175
rect 19465 -9295 19510 -9175
rect 19630 -9295 19675 -9175
rect 19795 -9295 19850 -9175
rect 19970 -9295 20015 -9175
rect 20135 -9295 20180 -9175
rect 20300 -9295 20345 -9175
rect 20465 -9295 20520 -9175
rect 20640 -9295 20685 -9175
rect 20805 -9295 20850 -9175
rect 20970 -9295 21015 -9175
rect 21135 -9295 21190 -9175
rect 21310 -9295 21355 -9175
rect 21475 -9295 21520 -9175
rect 21640 -9295 21685 -9175
rect 21805 -9295 21860 -9175
rect 21980 -9295 22025 -9175
rect 22145 -9295 22190 -9175
rect 22310 -9295 22355 -9175
rect 22475 -9295 22530 -9175
rect 22650 -9295 22695 -9175
rect 22815 -9295 22860 -9175
rect 22980 -9295 23025 -9175
rect 23145 -9295 23200 -9175
rect 23320 -9295 23365 -9175
rect 23485 -9295 23530 -9175
rect 23650 -9295 23695 -9175
rect 23815 -9295 23870 -9175
rect 23990 -9295 24000 -9175
rect 18500 -9340 24000 -9295
rect 18500 -9460 18510 -9340
rect 18630 -9460 18675 -9340
rect 18795 -9460 18840 -9340
rect 18960 -9460 19005 -9340
rect 19125 -9460 19180 -9340
rect 19300 -9460 19345 -9340
rect 19465 -9460 19510 -9340
rect 19630 -9460 19675 -9340
rect 19795 -9460 19850 -9340
rect 19970 -9460 20015 -9340
rect 20135 -9460 20180 -9340
rect 20300 -9460 20345 -9340
rect 20465 -9460 20520 -9340
rect 20640 -9460 20685 -9340
rect 20805 -9460 20850 -9340
rect 20970 -9460 21015 -9340
rect 21135 -9460 21190 -9340
rect 21310 -9460 21355 -9340
rect 21475 -9460 21520 -9340
rect 21640 -9460 21685 -9340
rect 21805 -9460 21860 -9340
rect 21980 -9460 22025 -9340
rect 22145 -9460 22190 -9340
rect 22310 -9460 22355 -9340
rect 22475 -9460 22530 -9340
rect 22650 -9460 22695 -9340
rect 22815 -9460 22860 -9340
rect 22980 -9460 23025 -9340
rect 23145 -9460 23200 -9340
rect 23320 -9460 23365 -9340
rect 23485 -9460 23530 -9340
rect 23650 -9460 23695 -9340
rect 23815 -9460 23870 -9340
rect 23990 -9460 24000 -9340
rect 18500 -9505 24000 -9460
rect 18500 -9625 18510 -9505
rect 18630 -9625 18675 -9505
rect 18795 -9625 18840 -9505
rect 18960 -9625 19005 -9505
rect 19125 -9625 19180 -9505
rect 19300 -9625 19345 -9505
rect 19465 -9625 19510 -9505
rect 19630 -9625 19675 -9505
rect 19795 -9625 19850 -9505
rect 19970 -9625 20015 -9505
rect 20135 -9625 20180 -9505
rect 20300 -9625 20345 -9505
rect 20465 -9625 20520 -9505
rect 20640 -9625 20685 -9505
rect 20805 -9625 20850 -9505
rect 20970 -9625 21015 -9505
rect 21135 -9625 21190 -9505
rect 21310 -9625 21355 -9505
rect 21475 -9625 21520 -9505
rect 21640 -9625 21685 -9505
rect 21805 -9625 21860 -9505
rect 21980 -9625 22025 -9505
rect 22145 -9625 22190 -9505
rect 22310 -9625 22355 -9505
rect 22475 -9625 22530 -9505
rect 22650 -9625 22695 -9505
rect 22815 -9625 22860 -9505
rect 22980 -9625 23025 -9505
rect 23145 -9625 23200 -9505
rect 23320 -9625 23365 -9505
rect 23485 -9625 23530 -9505
rect 23650 -9625 23695 -9505
rect 23815 -9625 23870 -9505
rect 23990 -9625 24000 -9505
rect 18500 -9670 24000 -9625
rect 18500 -9790 18510 -9670
rect 18630 -9790 18675 -9670
rect 18795 -9790 18840 -9670
rect 18960 -9790 19005 -9670
rect 19125 -9790 19180 -9670
rect 19300 -9790 19345 -9670
rect 19465 -9790 19510 -9670
rect 19630 -9790 19675 -9670
rect 19795 -9790 19850 -9670
rect 19970 -9790 20015 -9670
rect 20135 -9790 20180 -9670
rect 20300 -9790 20345 -9670
rect 20465 -9790 20520 -9670
rect 20640 -9790 20685 -9670
rect 20805 -9790 20850 -9670
rect 20970 -9790 21015 -9670
rect 21135 -9790 21190 -9670
rect 21310 -9790 21355 -9670
rect 21475 -9790 21520 -9670
rect 21640 -9790 21685 -9670
rect 21805 -9790 21860 -9670
rect 21980 -9790 22025 -9670
rect 22145 -9790 22190 -9670
rect 22310 -9790 22355 -9670
rect 22475 -9790 22530 -9670
rect 22650 -9790 22695 -9670
rect 22815 -9790 22860 -9670
rect 22980 -9790 23025 -9670
rect 23145 -9790 23200 -9670
rect 23320 -9790 23365 -9670
rect 23485 -9790 23530 -9670
rect 23650 -9790 23695 -9670
rect 23815 -9790 23870 -9670
rect 23990 -9790 24000 -9670
rect 18500 -9800 24000 -9790
rect 24190 -4310 29690 -4300
rect 24190 -4430 24200 -4310
rect 24320 -4430 24365 -4310
rect 24485 -4430 24530 -4310
rect 24650 -4430 24695 -4310
rect 24815 -4430 24870 -4310
rect 24990 -4430 25035 -4310
rect 25155 -4430 25200 -4310
rect 25320 -4430 25365 -4310
rect 25485 -4430 25540 -4310
rect 25660 -4430 25705 -4310
rect 25825 -4430 25870 -4310
rect 25990 -4430 26035 -4310
rect 26155 -4430 26210 -4310
rect 26330 -4430 26375 -4310
rect 26495 -4430 26540 -4310
rect 26660 -4430 26705 -4310
rect 26825 -4430 26880 -4310
rect 27000 -4430 27045 -4310
rect 27165 -4430 27210 -4310
rect 27330 -4430 27375 -4310
rect 27495 -4430 27550 -4310
rect 27670 -4430 27715 -4310
rect 27835 -4430 27880 -4310
rect 28000 -4430 28045 -4310
rect 28165 -4430 28220 -4310
rect 28340 -4430 28385 -4310
rect 28505 -4430 28550 -4310
rect 28670 -4430 28715 -4310
rect 28835 -4430 28890 -4310
rect 29010 -4430 29055 -4310
rect 29175 -4430 29220 -4310
rect 29340 -4430 29385 -4310
rect 29505 -4430 29560 -4310
rect 29680 -4430 29690 -4310
rect 24190 -4485 29690 -4430
rect 24190 -4605 24200 -4485
rect 24320 -4605 24365 -4485
rect 24485 -4605 24530 -4485
rect 24650 -4605 24695 -4485
rect 24815 -4605 24870 -4485
rect 24990 -4605 25035 -4485
rect 25155 -4605 25200 -4485
rect 25320 -4605 25365 -4485
rect 25485 -4605 25540 -4485
rect 25660 -4605 25705 -4485
rect 25825 -4605 25870 -4485
rect 25990 -4605 26035 -4485
rect 26155 -4605 26210 -4485
rect 26330 -4605 26375 -4485
rect 26495 -4605 26540 -4485
rect 26660 -4605 26705 -4485
rect 26825 -4605 26880 -4485
rect 27000 -4605 27045 -4485
rect 27165 -4605 27210 -4485
rect 27330 -4605 27375 -4485
rect 27495 -4605 27550 -4485
rect 27670 -4605 27715 -4485
rect 27835 -4605 27880 -4485
rect 28000 -4605 28045 -4485
rect 28165 -4605 28220 -4485
rect 28340 -4605 28385 -4485
rect 28505 -4605 28550 -4485
rect 28670 -4605 28715 -4485
rect 28835 -4605 28890 -4485
rect 29010 -4605 29055 -4485
rect 29175 -4605 29220 -4485
rect 29340 -4605 29385 -4485
rect 29505 -4605 29560 -4485
rect 29680 -4605 29690 -4485
rect 24190 -4650 29690 -4605
rect 24190 -4770 24200 -4650
rect 24320 -4770 24365 -4650
rect 24485 -4770 24530 -4650
rect 24650 -4770 24695 -4650
rect 24815 -4770 24870 -4650
rect 24990 -4770 25035 -4650
rect 25155 -4770 25200 -4650
rect 25320 -4770 25365 -4650
rect 25485 -4770 25540 -4650
rect 25660 -4770 25705 -4650
rect 25825 -4770 25870 -4650
rect 25990 -4770 26035 -4650
rect 26155 -4770 26210 -4650
rect 26330 -4770 26375 -4650
rect 26495 -4770 26540 -4650
rect 26660 -4770 26705 -4650
rect 26825 -4770 26880 -4650
rect 27000 -4770 27045 -4650
rect 27165 -4770 27210 -4650
rect 27330 -4770 27375 -4650
rect 27495 -4770 27550 -4650
rect 27670 -4770 27715 -4650
rect 27835 -4770 27880 -4650
rect 28000 -4770 28045 -4650
rect 28165 -4770 28220 -4650
rect 28340 -4770 28385 -4650
rect 28505 -4770 28550 -4650
rect 28670 -4770 28715 -4650
rect 28835 -4770 28890 -4650
rect 29010 -4770 29055 -4650
rect 29175 -4770 29220 -4650
rect 29340 -4770 29385 -4650
rect 29505 -4770 29560 -4650
rect 29680 -4770 29690 -4650
rect 24190 -4815 29690 -4770
rect 24190 -4935 24200 -4815
rect 24320 -4935 24365 -4815
rect 24485 -4935 24530 -4815
rect 24650 -4935 24695 -4815
rect 24815 -4935 24870 -4815
rect 24990 -4935 25035 -4815
rect 25155 -4935 25200 -4815
rect 25320 -4935 25365 -4815
rect 25485 -4935 25540 -4815
rect 25660 -4935 25705 -4815
rect 25825 -4935 25870 -4815
rect 25990 -4935 26035 -4815
rect 26155 -4935 26210 -4815
rect 26330 -4935 26375 -4815
rect 26495 -4935 26540 -4815
rect 26660 -4935 26705 -4815
rect 26825 -4935 26880 -4815
rect 27000 -4935 27045 -4815
rect 27165 -4935 27210 -4815
rect 27330 -4935 27375 -4815
rect 27495 -4935 27550 -4815
rect 27670 -4935 27715 -4815
rect 27835 -4935 27880 -4815
rect 28000 -4935 28045 -4815
rect 28165 -4935 28220 -4815
rect 28340 -4935 28385 -4815
rect 28505 -4935 28550 -4815
rect 28670 -4935 28715 -4815
rect 28835 -4935 28890 -4815
rect 29010 -4935 29055 -4815
rect 29175 -4935 29220 -4815
rect 29340 -4935 29385 -4815
rect 29505 -4935 29560 -4815
rect 29680 -4935 29690 -4815
rect 24190 -4980 29690 -4935
rect 24190 -5100 24200 -4980
rect 24320 -5100 24365 -4980
rect 24485 -5100 24530 -4980
rect 24650 -5100 24695 -4980
rect 24815 -5100 24870 -4980
rect 24990 -5100 25035 -4980
rect 25155 -5100 25200 -4980
rect 25320 -5100 25365 -4980
rect 25485 -5100 25540 -4980
rect 25660 -5100 25705 -4980
rect 25825 -5100 25870 -4980
rect 25990 -5100 26035 -4980
rect 26155 -5100 26210 -4980
rect 26330 -5100 26375 -4980
rect 26495 -5100 26540 -4980
rect 26660 -5100 26705 -4980
rect 26825 -5100 26880 -4980
rect 27000 -5100 27045 -4980
rect 27165 -5100 27210 -4980
rect 27330 -5100 27375 -4980
rect 27495 -5100 27550 -4980
rect 27670 -5100 27715 -4980
rect 27835 -5100 27880 -4980
rect 28000 -5100 28045 -4980
rect 28165 -5100 28220 -4980
rect 28340 -5100 28385 -4980
rect 28505 -5100 28550 -4980
rect 28670 -5100 28715 -4980
rect 28835 -5100 28890 -4980
rect 29010 -5100 29055 -4980
rect 29175 -5100 29220 -4980
rect 29340 -5100 29385 -4980
rect 29505 -5100 29560 -4980
rect 29680 -5100 29690 -4980
rect 24190 -5155 29690 -5100
rect 24190 -5275 24200 -5155
rect 24320 -5275 24365 -5155
rect 24485 -5275 24530 -5155
rect 24650 -5275 24695 -5155
rect 24815 -5275 24870 -5155
rect 24990 -5275 25035 -5155
rect 25155 -5275 25200 -5155
rect 25320 -5275 25365 -5155
rect 25485 -5275 25540 -5155
rect 25660 -5275 25705 -5155
rect 25825 -5275 25870 -5155
rect 25990 -5275 26035 -5155
rect 26155 -5275 26210 -5155
rect 26330 -5275 26375 -5155
rect 26495 -5275 26540 -5155
rect 26660 -5275 26705 -5155
rect 26825 -5275 26880 -5155
rect 27000 -5275 27045 -5155
rect 27165 -5275 27210 -5155
rect 27330 -5275 27375 -5155
rect 27495 -5275 27550 -5155
rect 27670 -5275 27715 -5155
rect 27835 -5275 27880 -5155
rect 28000 -5275 28045 -5155
rect 28165 -5275 28220 -5155
rect 28340 -5275 28385 -5155
rect 28505 -5275 28550 -5155
rect 28670 -5275 28715 -5155
rect 28835 -5275 28890 -5155
rect 29010 -5275 29055 -5155
rect 29175 -5275 29220 -5155
rect 29340 -5275 29385 -5155
rect 29505 -5275 29560 -5155
rect 29680 -5275 29690 -5155
rect 24190 -5320 29690 -5275
rect 24190 -5440 24200 -5320
rect 24320 -5440 24365 -5320
rect 24485 -5440 24530 -5320
rect 24650 -5440 24695 -5320
rect 24815 -5440 24870 -5320
rect 24990 -5440 25035 -5320
rect 25155 -5440 25200 -5320
rect 25320 -5440 25365 -5320
rect 25485 -5440 25540 -5320
rect 25660 -5440 25705 -5320
rect 25825 -5440 25870 -5320
rect 25990 -5440 26035 -5320
rect 26155 -5440 26210 -5320
rect 26330 -5440 26375 -5320
rect 26495 -5440 26540 -5320
rect 26660 -5440 26705 -5320
rect 26825 -5440 26880 -5320
rect 27000 -5440 27045 -5320
rect 27165 -5440 27210 -5320
rect 27330 -5440 27375 -5320
rect 27495 -5440 27550 -5320
rect 27670 -5440 27715 -5320
rect 27835 -5440 27880 -5320
rect 28000 -5440 28045 -5320
rect 28165 -5440 28220 -5320
rect 28340 -5440 28385 -5320
rect 28505 -5440 28550 -5320
rect 28670 -5440 28715 -5320
rect 28835 -5440 28890 -5320
rect 29010 -5440 29055 -5320
rect 29175 -5440 29220 -5320
rect 29340 -5440 29385 -5320
rect 29505 -5440 29560 -5320
rect 29680 -5440 29690 -5320
rect 24190 -5485 29690 -5440
rect 24190 -5605 24200 -5485
rect 24320 -5605 24365 -5485
rect 24485 -5605 24530 -5485
rect 24650 -5605 24695 -5485
rect 24815 -5605 24870 -5485
rect 24990 -5605 25035 -5485
rect 25155 -5605 25200 -5485
rect 25320 -5605 25365 -5485
rect 25485 -5605 25540 -5485
rect 25660 -5605 25705 -5485
rect 25825 -5605 25870 -5485
rect 25990 -5605 26035 -5485
rect 26155 -5605 26210 -5485
rect 26330 -5605 26375 -5485
rect 26495 -5605 26540 -5485
rect 26660 -5605 26705 -5485
rect 26825 -5605 26880 -5485
rect 27000 -5605 27045 -5485
rect 27165 -5605 27210 -5485
rect 27330 -5605 27375 -5485
rect 27495 -5605 27550 -5485
rect 27670 -5605 27715 -5485
rect 27835 -5605 27880 -5485
rect 28000 -5605 28045 -5485
rect 28165 -5605 28220 -5485
rect 28340 -5605 28385 -5485
rect 28505 -5605 28550 -5485
rect 28670 -5605 28715 -5485
rect 28835 -5605 28890 -5485
rect 29010 -5605 29055 -5485
rect 29175 -5605 29220 -5485
rect 29340 -5605 29385 -5485
rect 29505 -5605 29560 -5485
rect 29680 -5605 29690 -5485
rect 24190 -5650 29690 -5605
rect 24190 -5770 24200 -5650
rect 24320 -5770 24365 -5650
rect 24485 -5770 24530 -5650
rect 24650 -5770 24695 -5650
rect 24815 -5770 24870 -5650
rect 24990 -5770 25035 -5650
rect 25155 -5770 25200 -5650
rect 25320 -5770 25365 -5650
rect 25485 -5770 25540 -5650
rect 25660 -5770 25705 -5650
rect 25825 -5770 25870 -5650
rect 25990 -5770 26035 -5650
rect 26155 -5770 26210 -5650
rect 26330 -5770 26375 -5650
rect 26495 -5770 26540 -5650
rect 26660 -5770 26705 -5650
rect 26825 -5770 26880 -5650
rect 27000 -5770 27045 -5650
rect 27165 -5770 27210 -5650
rect 27330 -5770 27375 -5650
rect 27495 -5770 27550 -5650
rect 27670 -5770 27715 -5650
rect 27835 -5770 27880 -5650
rect 28000 -5770 28045 -5650
rect 28165 -5770 28220 -5650
rect 28340 -5770 28385 -5650
rect 28505 -5770 28550 -5650
rect 28670 -5770 28715 -5650
rect 28835 -5770 28890 -5650
rect 29010 -5770 29055 -5650
rect 29175 -5770 29220 -5650
rect 29340 -5770 29385 -5650
rect 29505 -5770 29560 -5650
rect 29680 -5770 29690 -5650
rect 24190 -5825 29690 -5770
rect 24190 -5945 24200 -5825
rect 24320 -5945 24365 -5825
rect 24485 -5945 24530 -5825
rect 24650 -5945 24695 -5825
rect 24815 -5945 24870 -5825
rect 24990 -5945 25035 -5825
rect 25155 -5945 25200 -5825
rect 25320 -5945 25365 -5825
rect 25485 -5945 25540 -5825
rect 25660 -5945 25705 -5825
rect 25825 -5945 25870 -5825
rect 25990 -5945 26035 -5825
rect 26155 -5945 26210 -5825
rect 26330 -5945 26375 -5825
rect 26495 -5945 26540 -5825
rect 26660 -5945 26705 -5825
rect 26825 -5945 26880 -5825
rect 27000 -5945 27045 -5825
rect 27165 -5945 27210 -5825
rect 27330 -5945 27375 -5825
rect 27495 -5945 27550 -5825
rect 27670 -5945 27715 -5825
rect 27835 -5945 27880 -5825
rect 28000 -5945 28045 -5825
rect 28165 -5945 28220 -5825
rect 28340 -5945 28385 -5825
rect 28505 -5945 28550 -5825
rect 28670 -5945 28715 -5825
rect 28835 -5945 28890 -5825
rect 29010 -5945 29055 -5825
rect 29175 -5945 29220 -5825
rect 29340 -5945 29385 -5825
rect 29505 -5945 29560 -5825
rect 29680 -5945 29690 -5825
rect 24190 -5990 29690 -5945
rect 24190 -6110 24200 -5990
rect 24320 -6110 24365 -5990
rect 24485 -6110 24530 -5990
rect 24650 -6110 24695 -5990
rect 24815 -6110 24870 -5990
rect 24990 -6110 25035 -5990
rect 25155 -6110 25200 -5990
rect 25320 -6110 25365 -5990
rect 25485 -6110 25540 -5990
rect 25660 -6110 25705 -5990
rect 25825 -6110 25870 -5990
rect 25990 -6110 26035 -5990
rect 26155 -6110 26210 -5990
rect 26330 -6110 26375 -5990
rect 26495 -6110 26540 -5990
rect 26660 -6110 26705 -5990
rect 26825 -6110 26880 -5990
rect 27000 -6110 27045 -5990
rect 27165 -6110 27210 -5990
rect 27330 -6110 27375 -5990
rect 27495 -6110 27550 -5990
rect 27670 -6110 27715 -5990
rect 27835 -6110 27880 -5990
rect 28000 -6110 28045 -5990
rect 28165 -6110 28220 -5990
rect 28340 -6110 28385 -5990
rect 28505 -6110 28550 -5990
rect 28670 -6110 28715 -5990
rect 28835 -6110 28890 -5990
rect 29010 -6110 29055 -5990
rect 29175 -6110 29220 -5990
rect 29340 -6110 29385 -5990
rect 29505 -6110 29560 -5990
rect 29680 -6110 29690 -5990
rect 24190 -6155 29690 -6110
rect 24190 -6275 24200 -6155
rect 24320 -6275 24365 -6155
rect 24485 -6275 24530 -6155
rect 24650 -6275 24695 -6155
rect 24815 -6275 24870 -6155
rect 24990 -6275 25035 -6155
rect 25155 -6275 25200 -6155
rect 25320 -6275 25365 -6155
rect 25485 -6275 25540 -6155
rect 25660 -6275 25705 -6155
rect 25825 -6275 25870 -6155
rect 25990 -6275 26035 -6155
rect 26155 -6275 26210 -6155
rect 26330 -6275 26375 -6155
rect 26495 -6275 26540 -6155
rect 26660 -6275 26705 -6155
rect 26825 -6275 26880 -6155
rect 27000 -6275 27045 -6155
rect 27165 -6275 27210 -6155
rect 27330 -6275 27375 -6155
rect 27495 -6275 27550 -6155
rect 27670 -6275 27715 -6155
rect 27835 -6275 27880 -6155
rect 28000 -6275 28045 -6155
rect 28165 -6275 28220 -6155
rect 28340 -6275 28385 -6155
rect 28505 -6275 28550 -6155
rect 28670 -6275 28715 -6155
rect 28835 -6275 28890 -6155
rect 29010 -6275 29055 -6155
rect 29175 -6275 29220 -6155
rect 29340 -6275 29385 -6155
rect 29505 -6275 29560 -6155
rect 29680 -6275 29690 -6155
rect 24190 -6320 29690 -6275
rect 24190 -6440 24200 -6320
rect 24320 -6440 24365 -6320
rect 24485 -6440 24530 -6320
rect 24650 -6440 24695 -6320
rect 24815 -6440 24870 -6320
rect 24990 -6440 25035 -6320
rect 25155 -6440 25200 -6320
rect 25320 -6440 25365 -6320
rect 25485 -6440 25540 -6320
rect 25660 -6440 25705 -6320
rect 25825 -6440 25870 -6320
rect 25990 -6440 26035 -6320
rect 26155 -6440 26210 -6320
rect 26330 -6440 26375 -6320
rect 26495 -6440 26540 -6320
rect 26660 -6440 26705 -6320
rect 26825 -6440 26880 -6320
rect 27000 -6440 27045 -6320
rect 27165 -6440 27210 -6320
rect 27330 -6440 27375 -6320
rect 27495 -6440 27550 -6320
rect 27670 -6440 27715 -6320
rect 27835 -6440 27880 -6320
rect 28000 -6440 28045 -6320
rect 28165 -6440 28220 -6320
rect 28340 -6440 28385 -6320
rect 28505 -6440 28550 -6320
rect 28670 -6440 28715 -6320
rect 28835 -6440 28890 -6320
rect 29010 -6440 29055 -6320
rect 29175 -6440 29220 -6320
rect 29340 -6440 29385 -6320
rect 29505 -6440 29560 -6320
rect 29680 -6440 29690 -6320
rect 24190 -6495 29690 -6440
rect 24190 -6615 24200 -6495
rect 24320 -6615 24365 -6495
rect 24485 -6615 24530 -6495
rect 24650 -6615 24695 -6495
rect 24815 -6615 24870 -6495
rect 24990 -6615 25035 -6495
rect 25155 -6615 25200 -6495
rect 25320 -6615 25365 -6495
rect 25485 -6615 25540 -6495
rect 25660 -6615 25705 -6495
rect 25825 -6615 25870 -6495
rect 25990 -6615 26035 -6495
rect 26155 -6615 26210 -6495
rect 26330 -6615 26375 -6495
rect 26495 -6615 26540 -6495
rect 26660 -6615 26705 -6495
rect 26825 -6615 26880 -6495
rect 27000 -6615 27045 -6495
rect 27165 -6615 27210 -6495
rect 27330 -6615 27375 -6495
rect 27495 -6615 27550 -6495
rect 27670 -6615 27715 -6495
rect 27835 -6615 27880 -6495
rect 28000 -6615 28045 -6495
rect 28165 -6615 28220 -6495
rect 28340 -6615 28385 -6495
rect 28505 -6615 28550 -6495
rect 28670 -6615 28715 -6495
rect 28835 -6615 28890 -6495
rect 29010 -6615 29055 -6495
rect 29175 -6615 29220 -6495
rect 29340 -6615 29385 -6495
rect 29505 -6615 29560 -6495
rect 29680 -6615 29690 -6495
rect 24190 -6660 29690 -6615
rect 24190 -6780 24200 -6660
rect 24320 -6780 24365 -6660
rect 24485 -6780 24530 -6660
rect 24650 -6780 24695 -6660
rect 24815 -6780 24870 -6660
rect 24990 -6780 25035 -6660
rect 25155 -6780 25200 -6660
rect 25320 -6780 25365 -6660
rect 25485 -6780 25540 -6660
rect 25660 -6780 25705 -6660
rect 25825 -6780 25870 -6660
rect 25990 -6780 26035 -6660
rect 26155 -6780 26210 -6660
rect 26330 -6780 26375 -6660
rect 26495 -6780 26540 -6660
rect 26660 -6780 26705 -6660
rect 26825 -6780 26880 -6660
rect 27000 -6780 27045 -6660
rect 27165 -6780 27210 -6660
rect 27330 -6780 27375 -6660
rect 27495 -6780 27550 -6660
rect 27670 -6780 27715 -6660
rect 27835 -6780 27880 -6660
rect 28000 -6780 28045 -6660
rect 28165 -6780 28220 -6660
rect 28340 -6780 28385 -6660
rect 28505 -6780 28550 -6660
rect 28670 -6780 28715 -6660
rect 28835 -6780 28890 -6660
rect 29010 -6780 29055 -6660
rect 29175 -6780 29220 -6660
rect 29340 -6780 29385 -6660
rect 29505 -6780 29560 -6660
rect 29680 -6780 29690 -6660
rect 24190 -6825 29690 -6780
rect 24190 -6945 24200 -6825
rect 24320 -6945 24365 -6825
rect 24485 -6945 24530 -6825
rect 24650 -6945 24695 -6825
rect 24815 -6945 24870 -6825
rect 24990 -6945 25035 -6825
rect 25155 -6945 25200 -6825
rect 25320 -6945 25365 -6825
rect 25485 -6945 25540 -6825
rect 25660 -6945 25705 -6825
rect 25825 -6945 25870 -6825
rect 25990 -6945 26035 -6825
rect 26155 -6945 26210 -6825
rect 26330 -6945 26375 -6825
rect 26495 -6945 26540 -6825
rect 26660 -6945 26705 -6825
rect 26825 -6945 26880 -6825
rect 27000 -6945 27045 -6825
rect 27165 -6945 27210 -6825
rect 27330 -6945 27375 -6825
rect 27495 -6945 27550 -6825
rect 27670 -6945 27715 -6825
rect 27835 -6945 27880 -6825
rect 28000 -6945 28045 -6825
rect 28165 -6945 28220 -6825
rect 28340 -6945 28385 -6825
rect 28505 -6945 28550 -6825
rect 28670 -6945 28715 -6825
rect 28835 -6945 28890 -6825
rect 29010 -6945 29055 -6825
rect 29175 -6945 29220 -6825
rect 29340 -6945 29385 -6825
rect 29505 -6945 29560 -6825
rect 29680 -6945 29690 -6825
rect 24190 -6990 29690 -6945
rect 24190 -7110 24200 -6990
rect 24320 -7110 24365 -6990
rect 24485 -7110 24530 -6990
rect 24650 -7110 24695 -6990
rect 24815 -7110 24870 -6990
rect 24990 -7110 25035 -6990
rect 25155 -7110 25200 -6990
rect 25320 -7110 25365 -6990
rect 25485 -7110 25540 -6990
rect 25660 -7110 25705 -6990
rect 25825 -7110 25870 -6990
rect 25990 -7110 26035 -6990
rect 26155 -7110 26210 -6990
rect 26330 -7110 26375 -6990
rect 26495 -7110 26540 -6990
rect 26660 -7110 26705 -6990
rect 26825 -7110 26880 -6990
rect 27000 -7110 27045 -6990
rect 27165 -7110 27210 -6990
rect 27330 -7110 27375 -6990
rect 27495 -7110 27550 -6990
rect 27670 -7110 27715 -6990
rect 27835 -7110 27880 -6990
rect 28000 -7110 28045 -6990
rect 28165 -7110 28220 -6990
rect 28340 -7110 28385 -6990
rect 28505 -7110 28550 -6990
rect 28670 -7110 28715 -6990
rect 28835 -7110 28890 -6990
rect 29010 -7110 29055 -6990
rect 29175 -7110 29220 -6990
rect 29340 -7110 29385 -6990
rect 29505 -7110 29560 -6990
rect 29680 -7110 29690 -6990
rect 24190 -7165 29690 -7110
rect 24190 -7285 24200 -7165
rect 24320 -7285 24365 -7165
rect 24485 -7285 24530 -7165
rect 24650 -7285 24695 -7165
rect 24815 -7285 24870 -7165
rect 24990 -7285 25035 -7165
rect 25155 -7285 25200 -7165
rect 25320 -7285 25365 -7165
rect 25485 -7285 25540 -7165
rect 25660 -7285 25705 -7165
rect 25825 -7285 25870 -7165
rect 25990 -7285 26035 -7165
rect 26155 -7285 26210 -7165
rect 26330 -7285 26375 -7165
rect 26495 -7285 26540 -7165
rect 26660 -7285 26705 -7165
rect 26825 -7285 26880 -7165
rect 27000 -7285 27045 -7165
rect 27165 -7285 27210 -7165
rect 27330 -7285 27375 -7165
rect 27495 -7285 27550 -7165
rect 27670 -7285 27715 -7165
rect 27835 -7285 27880 -7165
rect 28000 -7285 28045 -7165
rect 28165 -7285 28220 -7165
rect 28340 -7285 28385 -7165
rect 28505 -7285 28550 -7165
rect 28670 -7285 28715 -7165
rect 28835 -7285 28890 -7165
rect 29010 -7285 29055 -7165
rect 29175 -7285 29220 -7165
rect 29340 -7285 29385 -7165
rect 29505 -7285 29560 -7165
rect 29680 -7285 29690 -7165
rect 24190 -7330 29690 -7285
rect 24190 -7450 24200 -7330
rect 24320 -7450 24365 -7330
rect 24485 -7450 24530 -7330
rect 24650 -7450 24695 -7330
rect 24815 -7450 24870 -7330
rect 24990 -7450 25035 -7330
rect 25155 -7450 25200 -7330
rect 25320 -7450 25365 -7330
rect 25485 -7450 25540 -7330
rect 25660 -7450 25705 -7330
rect 25825 -7450 25870 -7330
rect 25990 -7450 26035 -7330
rect 26155 -7450 26210 -7330
rect 26330 -7450 26375 -7330
rect 26495 -7450 26540 -7330
rect 26660 -7450 26705 -7330
rect 26825 -7450 26880 -7330
rect 27000 -7450 27045 -7330
rect 27165 -7450 27210 -7330
rect 27330 -7450 27375 -7330
rect 27495 -7450 27550 -7330
rect 27670 -7450 27715 -7330
rect 27835 -7450 27880 -7330
rect 28000 -7450 28045 -7330
rect 28165 -7450 28220 -7330
rect 28340 -7450 28385 -7330
rect 28505 -7450 28550 -7330
rect 28670 -7450 28715 -7330
rect 28835 -7450 28890 -7330
rect 29010 -7450 29055 -7330
rect 29175 -7450 29220 -7330
rect 29340 -7450 29385 -7330
rect 29505 -7450 29560 -7330
rect 29680 -7450 29690 -7330
rect 24190 -7495 29690 -7450
rect 24190 -7615 24200 -7495
rect 24320 -7615 24365 -7495
rect 24485 -7615 24530 -7495
rect 24650 -7615 24695 -7495
rect 24815 -7615 24870 -7495
rect 24990 -7615 25035 -7495
rect 25155 -7615 25200 -7495
rect 25320 -7615 25365 -7495
rect 25485 -7615 25540 -7495
rect 25660 -7615 25705 -7495
rect 25825 -7615 25870 -7495
rect 25990 -7615 26035 -7495
rect 26155 -7615 26210 -7495
rect 26330 -7615 26375 -7495
rect 26495 -7615 26540 -7495
rect 26660 -7615 26705 -7495
rect 26825 -7615 26880 -7495
rect 27000 -7615 27045 -7495
rect 27165 -7615 27210 -7495
rect 27330 -7615 27375 -7495
rect 27495 -7615 27550 -7495
rect 27670 -7615 27715 -7495
rect 27835 -7615 27880 -7495
rect 28000 -7615 28045 -7495
rect 28165 -7615 28220 -7495
rect 28340 -7615 28385 -7495
rect 28505 -7615 28550 -7495
rect 28670 -7615 28715 -7495
rect 28835 -7615 28890 -7495
rect 29010 -7615 29055 -7495
rect 29175 -7615 29220 -7495
rect 29340 -7615 29385 -7495
rect 29505 -7615 29560 -7495
rect 29680 -7615 29690 -7495
rect 24190 -7660 29690 -7615
rect 24190 -7780 24200 -7660
rect 24320 -7780 24365 -7660
rect 24485 -7780 24530 -7660
rect 24650 -7780 24695 -7660
rect 24815 -7780 24870 -7660
rect 24990 -7780 25035 -7660
rect 25155 -7780 25200 -7660
rect 25320 -7780 25365 -7660
rect 25485 -7780 25540 -7660
rect 25660 -7780 25705 -7660
rect 25825 -7780 25870 -7660
rect 25990 -7780 26035 -7660
rect 26155 -7780 26210 -7660
rect 26330 -7780 26375 -7660
rect 26495 -7780 26540 -7660
rect 26660 -7780 26705 -7660
rect 26825 -7780 26880 -7660
rect 27000 -7780 27045 -7660
rect 27165 -7780 27210 -7660
rect 27330 -7780 27375 -7660
rect 27495 -7780 27550 -7660
rect 27670 -7780 27715 -7660
rect 27835 -7780 27880 -7660
rect 28000 -7780 28045 -7660
rect 28165 -7780 28220 -7660
rect 28340 -7780 28385 -7660
rect 28505 -7780 28550 -7660
rect 28670 -7780 28715 -7660
rect 28835 -7780 28890 -7660
rect 29010 -7780 29055 -7660
rect 29175 -7780 29220 -7660
rect 29340 -7780 29385 -7660
rect 29505 -7780 29560 -7660
rect 29680 -7780 29690 -7660
rect 24190 -7835 29690 -7780
rect 24190 -7955 24200 -7835
rect 24320 -7955 24365 -7835
rect 24485 -7955 24530 -7835
rect 24650 -7955 24695 -7835
rect 24815 -7955 24870 -7835
rect 24990 -7955 25035 -7835
rect 25155 -7955 25200 -7835
rect 25320 -7955 25365 -7835
rect 25485 -7955 25540 -7835
rect 25660 -7955 25705 -7835
rect 25825 -7955 25870 -7835
rect 25990 -7955 26035 -7835
rect 26155 -7955 26210 -7835
rect 26330 -7955 26375 -7835
rect 26495 -7955 26540 -7835
rect 26660 -7955 26705 -7835
rect 26825 -7955 26880 -7835
rect 27000 -7955 27045 -7835
rect 27165 -7955 27210 -7835
rect 27330 -7955 27375 -7835
rect 27495 -7955 27550 -7835
rect 27670 -7955 27715 -7835
rect 27835 -7955 27880 -7835
rect 28000 -7955 28045 -7835
rect 28165 -7955 28220 -7835
rect 28340 -7955 28385 -7835
rect 28505 -7955 28550 -7835
rect 28670 -7955 28715 -7835
rect 28835 -7955 28890 -7835
rect 29010 -7955 29055 -7835
rect 29175 -7955 29220 -7835
rect 29340 -7955 29385 -7835
rect 29505 -7955 29560 -7835
rect 29680 -7955 29690 -7835
rect 24190 -8000 29690 -7955
rect 24190 -8120 24200 -8000
rect 24320 -8120 24365 -8000
rect 24485 -8120 24530 -8000
rect 24650 -8120 24695 -8000
rect 24815 -8120 24870 -8000
rect 24990 -8120 25035 -8000
rect 25155 -8120 25200 -8000
rect 25320 -8120 25365 -8000
rect 25485 -8120 25540 -8000
rect 25660 -8120 25705 -8000
rect 25825 -8120 25870 -8000
rect 25990 -8120 26035 -8000
rect 26155 -8120 26210 -8000
rect 26330 -8120 26375 -8000
rect 26495 -8120 26540 -8000
rect 26660 -8120 26705 -8000
rect 26825 -8120 26880 -8000
rect 27000 -8120 27045 -8000
rect 27165 -8120 27210 -8000
rect 27330 -8120 27375 -8000
rect 27495 -8120 27550 -8000
rect 27670 -8120 27715 -8000
rect 27835 -8120 27880 -8000
rect 28000 -8120 28045 -8000
rect 28165 -8120 28220 -8000
rect 28340 -8120 28385 -8000
rect 28505 -8120 28550 -8000
rect 28670 -8120 28715 -8000
rect 28835 -8120 28890 -8000
rect 29010 -8120 29055 -8000
rect 29175 -8120 29220 -8000
rect 29340 -8120 29385 -8000
rect 29505 -8120 29560 -8000
rect 29680 -8120 29690 -8000
rect 24190 -8165 29690 -8120
rect 24190 -8285 24200 -8165
rect 24320 -8285 24365 -8165
rect 24485 -8285 24530 -8165
rect 24650 -8285 24695 -8165
rect 24815 -8285 24870 -8165
rect 24990 -8285 25035 -8165
rect 25155 -8285 25200 -8165
rect 25320 -8285 25365 -8165
rect 25485 -8285 25540 -8165
rect 25660 -8285 25705 -8165
rect 25825 -8285 25870 -8165
rect 25990 -8285 26035 -8165
rect 26155 -8285 26210 -8165
rect 26330 -8285 26375 -8165
rect 26495 -8285 26540 -8165
rect 26660 -8285 26705 -8165
rect 26825 -8285 26880 -8165
rect 27000 -8285 27045 -8165
rect 27165 -8285 27210 -8165
rect 27330 -8285 27375 -8165
rect 27495 -8285 27550 -8165
rect 27670 -8285 27715 -8165
rect 27835 -8285 27880 -8165
rect 28000 -8285 28045 -8165
rect 28165 -8285 28220 -8165
rect 28340 -8285 28385 -8165
rect 28505 -8285 28550 -8165
rect 28670 -8285 28715 -8165
rect 28835 -8285 28890 -8165
rect 29010 -8285 29055 -8165
rect 29175 -8285 29220 -8165
rect 29340 -8285 29385 -8165
rect 29505 -8285 29560 -8165
rect 29680 -8285 29690 -8165
rect 24190 -8330 29690 -8285
rect 24190 -8450 24200 -8330
rect 24320 -8450 24365 -8330
rect 24485 -8450 24530 -8330
rect 24650 -8450 24695 -8330
rect 24815 -8450 24870 -8330
rect 24990 -8450 25035 -8330
rect 25155 -8450 25200 -8330
rect 25320 -8450 25365 -8330
rect 25485 -8450 25540 -8330
rect 25660 -8450 25705 -8330
rect 25825 -8450 25870 -8330
rect 25990 -8450 26035 -8330
rect 26155 -8450 26210 -8330
rect 26330 -8450 26375 -8330
rect 26495 -8450 26540 -8330
rect 26660 -8450 26705 -8330
rect 26825 -8450 26880 -8330
rect 27000 -8450 27045 -8330
rect 27165 -8450 27210 -8330
rect 27330 -8450 27375 -8330
rect 27495 -8450 27550 -8330
rect 27670 -8450 27715 -8330
rect 27835 -8450 27880 -8330
rect 28000 -8450 28045 -8330
rect 28165 -8450 28220 -8330
rect 28340 -8450 28385 -8330
rect 28505 -8450 28550 -8330
rect 28670 -8450 28715 -8330
rect 28835 -8450 28890 -8330
rect 29010 -8450 29055 -8330
rect 29175 -8450 29220 -8330
rect 29340 -8450 29385 -8330
rect 29505 -8450 29560 -8330
rect 29680 -8450 29690 -8330
rect 24190 -8505 29690 -8450
rect 24190 -8625 24200 -8505
rect 24320 -8625 24365 -8505
rect 24485 -8625 24530 -8505
rect 24650 -8625 24695 -8505
rect 24815 -8625 24870 -8505
rect 24990 -8625 25035 -8505
rect 25155 -8625 25200 -8505
rect 25320 -8625 25365 -8505
rect 25485 -8625 25540 -8505
rect 25660 -8625 25705 -8505
rect 25825 -8625 25870 -8505
rect 25990 -8625 26035 -8505
rect 26155 -8625 26210 -8505
rect 26330 -8625 26375 -8505
rect 26495 -8625 26540 -8505
rect 26660 -8625 26705 -8505
rect 26825 -8625 26880 -8505
rect 27000 -8625 27045 -8505
rect 27165 -8625 27210 -8505
rect 27330 -8625 27375 -8505
rect 27495 -8625 27550 -8505
rect 27670 -8625 27715 -8505
rect 27835 -8625 27880 -8505
rect 28000 -8625 28045 -8505
rect 28165 -8625 28220 -8505
rect 28340 -8625 28385 -8505
rect 28505 -8625 28550 -8505
rect 28670 -8625 28715 -8505
rect 28835 -8625 28890 -8505
rect 29010 -8625 29055 -8505
rect 29175 -8625 29220 -8505
rect 29340 -8625 29385 -8505
rect 29505 -8625 29560 -8505
rect 29680 -8625 29690 -8505
rect 24190 -8670 29690 -8625
rect 24190 -8790 24200 -8670
rect 24320 -8790 24365 -8670
rect 24485 -8790 24530 -8670
rect 24650 -8790 24695 -8670
rect 24815 -8790 24870 -8670
rect 24990 -8790 25035 -8670
rect 25155 -8790 25200 -8670
rect 25320 -8790 25365 -8670
rect 25485 -8790 25540 -8670
rect 25660 -8790 25705 -8670
rect 25825 -8790 25870 -8670
rect 25990 -8790 26035 -8670
rect 26155 -8790 26210 -8670
rect 26330 -8790 26375 -8670
rect 26495 -8790 26540 -8670
rect 26660 -8790 26705 -8670
rect 26825 -8790 26880 -8670
rect 27000 -8790 27045 -8670
rect 27165 -8790 27210 -8670
rect 27330 -8790 27375 -8670
rect 27495 -8790 27550 -8670
rect 27670 -8790 27715 -8670
rect 27835 -8790 27880 -8670
rect 28000 -8790 28045 -8670
rect 28165 -8790 28220 -8670
rect 28340 -8790 28385 -8670
rect 28505 -8790 28550 -8670
rect 28670 -8790 28715 -8670
rect 28835 -8790 28890 -8670
rect 29010 -8790 29055 -8670
rect 29175 -8790 29220 -8670
rect 29340 -8790 29385 -8670
rect 29505 -8790 29560 -8670
rect 29680 -8790 29690 -8670
rect 24190 -8835 29690 -8790
rect 24190 -8955 24200 -8835
rect 24320 -8955 24365 -8835
rect 24485 -8955 24530 -8835
rect 24650 -8955 24695 -8835
rect 24815 -8955 24870 -8835
rect 24990 -8955 25035 -8835
rect 25155 -8955 25200 -8835
rect 25320 -8955 25365 -8835
rect 25485 -8955 25540 -8835
rect 25660 -8955 25705 -8835
rect 25825 -8955 25870 -8835
rect 25990 -8955 26035 -8835
rect 26155 -8955 26210 -8835
rect 26330 -8955 26375 -8835
rect 26495 -8955 26540 -8835
rect 26660 -8955 26705 -8835
rect 26825 -8955 26880 -8835
rect 27000 -8955 27045 -8835
rect 27165 -8955 27210 -8835
rect 27330 -8955 27375 -8835
rect 27495 -8955 27550 -8835
rect 27670 -8955 27715 -8835
rect 27835 -8955 27880 -8835
rect 28000 -8955 28045 -8835
rect 28165 -8955 28220 -8835
rect 28340 -8955 28385 -8835
rect 28505 -8955 28550 -8835
rect 28670 -8955 28715 -8835
rect 28835 -8955 28890 -8835
rect 29010 -8955 29055 -8835
rect 29175 -8955 29220 -8835
rect 29340 -8955 29385 -8835
rect 29505 -8955 29560 -8835
rect 29680 -8955 29690 -8835
rect 24190 -9000 29690 -8955
rect 24190 -9120 24200 -9000
rect 24320 -9120 24365 -9000
rect 24485 -9120 24530 -9000
rect 24650 -9120 24695 -9000
rect 24815 -9120 24870 -9000
rect 24990 -9120 25035 -9000
rect 25155 -9120 25200 -9000
rect 25320 -9120 25365 -9000
rect 25485 -9120 25540 -9000
rect 25660 -9120 25705 -9000
rect 25825 -9120 25870 -9000
rect 25990 -9120 26035 -9000
rect 26155 -9120 26210 -9000
rect 26330 -9120 26375 -9000
rect 26495 -9120 26540 -9000
rect 26660 -9120 26705 -9000
rect 26825 -9120 26880 -9000
rect 27000 -9120 27045 -9000
rect 27165 -9120 27210 -9000
rect 27330 -9120 27375 -9000
rect 27495 -9120 27550 -9000
rect 27670 -9120 27715 -9000
rect 27835 -9120 27880 -9000
rect 28000 -9120 28045 -9000
rect 28165 -9120 28220 -9000
rect 28340 -9120 28385 -9000
rect 28505 -9120 28550 -9000
rect 28670 -9120 28715 -9000
rect 28835 -9120 28890 -9000
rect 29010 -9120 29055 -9000
rect 29175 -9120 29220 -9000
rect 29340 -9120 29385 -9000
rect 29505 -9120 29560 -9000
rect 29680 -9120 29690 -9000
rect 24190 -9175 29690 -9120
rect 24190 -9295 24200 -9175
rect 24320 -9295 24365 -9175
rect 24485 -9295 24530 -9175
rect 24650 -9295 24695 -9175
rect 24815 -9295 24870 -9175
rect 24990 -9295 25035 -9175
rect 25155 -9295 25200 -9175
rect 25320 -9295 25365 -9175
rect 25485 -9295 25540 -9175
rect 25660 -9295 25705 -9175
rect 25825 -9295 25870 -9175
rect 25990 -9295 26035 -9175
rect 26155 -9295 26210 -9175
rect 26330 -9295 26375 -9175
rect 26495 -9295 26540 -9175
rect 26660 -9295 26705 -9175
rect 26825 -9295 26880 -9175
rect 27000 -9295 27045 -9175
rect 27165 -9295 27210 -9175
rect 27330 -9295 27375 -9175
rect 27495 -9295 27550 -9175
rect 27670 -9295 27715 -9175
rect 27835 -9295 27880 -9175
rect 28000 -9295 28045 -9175
rect 28165 -9295 28220 -9175
rect 28340 -9295 28385 -9175
rect 28505 -9295 28550 -9175
rect 28670 -9295 28715 -9175
rect 28835 -9295 28890 -9175
rect 29010 -9295 29055 -9175
rect 29175 -9295 29220 -9175
rect 29340 -9295 29385 -9175
rect 29505 -9295 29560 -9175
rect 29680 -9295 29690 -9175
rect 24190 -9340 29690 -9295
rect 24190 -9460 24200 -9340
rect 24320 -9460 24365 -9340
rect 24485 -9460 24530 -9340
rect 24650 -9460 24695 -9340
rect 24815 -9460 24870 -9340
rect 24990 -9460 25035 -9340
rect 25155 -9460 25200 -9340
rect 25320 -9460 25365 -9340
rect 25485 -9460 25540 -9340
rect 25660 -9460 25705 -9340
rect 25825 -9460 25870 -9340
rect 25990 -9460 26035 -9340
rect 26155 -9460 26210 -9340
rect 26330 -9460 26375 -9340
rect 26495 -9460 26540 -9340
rect 26660 -9460 26705 -9340
rect 26825 -9460 26880 -9340
rect 27000 -9460 27045 -9340
rect 27165 -9460 27210 -9340
rect 27330 -9460 27375 -9340
rect 27495 -9460 27550 -9340
rect 27670 -9460 27715 -9340
rect 27835 -9460 27880 -9340
rect 28000 -9460 28045 -9340
rect 28165 -9460 28220 -9340
rect 28340 -9460 28385 -9340
rect 28505 -9460 28550 -9340
rect 28670 -9460 28715 -9340
rect 28835 -9460 28890 -9340
rect 29010 -9460 29055 -9340
rect 29175 -9460 29220 -9340
rect 29340 -9460 29385 -9340
rect 29505 -9460 29560 -9340
rect 29680 -9460 29690 -9340
rect 24190 -9505 29690 -9460
rect 24190 -9625 24200 -9505
rect 24320 -9625 24365 -9505
rect 24485 -9625 24530 -9505
rect 24650 -9625 24695 -9505
rect 24815 -9625 24870 -9505
rect 24990 -9625 25035 -9505
rect 25155 -9625 25200 -9505
rect 25320 -9625 25365 -9505
rect 25485 -9625 25540 -9505
rect 25660 -9625 25705 -9505
rect 25825 -9625 25870 -9505
rect 25990 -9625 26035 -9505
rect 26155 -9625 26210 -9505
rect 26330 -9625 26375 -9505
rect 26495 -9625 26540 -9505
rect 26660 -9625 26705 -9505
rect 26825 -9625 26880 -9505
rect 27000 -9625 27045 -9505
rect 27165 -9625 27210 -9505
rect 27330 -9625 27375 -9505
rect 27495 -9625 27550 -9505
rect 27670 -9625 27715 -9505
rect 27835 -9625 27880 -9505
rect 28000 -9625 28045 -9505
rect 28165 -9625 28220 -9505
rect 28340 -9625 28385 -9505
rect 28505 -9625 28550 -9505
rect 28670 -9625 28715 -9505
rect 28835 -9625 28890 -9505
rect 29010 -9625 29055 -9505
rect 29175 -9625 29220 -9505
rect 29340 -9625 29385 -9505
rect 29505 -9625 29560 -9505
rect 29680 -9625 29690 -9505
rect 24190 -9670 29690 -9625
rect 24190 -9790 24200 -9670
rect 24320 -9790 24365 -9670
rect 24485 -9790 24530 -9670
rect 24650 -9790 24695 -9670
rect 24815 -9790 24870 -9670
rect 24990 -9790 25035 -9670
rect 25155 -9790 25200 -9670
rect 25320 -9790 25365 -9670
rect 25485 -9790 25540 -9670
rect 25660 -9790 25705 -9670
rect 25825 -9790 25870 -9670
rect 25990 -9790 26035 -9670
rect 26155 -9790 26210 -9670
rect 26330 -9790 26375 -9670
rect 26495 -9790 26540 -9670
rect 26660 -9790 26705 -9670
rect 26825 -9790 26880 -9670
rect 27000 -9790 27045 -9670
rect 27165 -9790 27210 -9670
rect 27330 -9790 27375 -9670
rect 27495 -9790 27550 -9670
rect 27670 -9790 27715 -9670
rect 27835 -9790 27880 -9670
rect 28000 -9790 28045 -9670
rect 28165 -9790 28220 -9670
rect 28340 -9790 28385 -9670
rect 28505 -9790 28550 -9670
rect 28670 -9790 28715 -9670
rect 28835 -9790 28890 -9670
rect 29010 -9790 29055 -9670
rect 29175 -9790 29220 -9670
rect 29340 -9790 29385 -9670
rect 29505 -9790 29560 -9670
rect 29680 -9790 29690 -9670
rect 24190 -9800 29690 -9790
rect 7120 -10090 12620 -10080
rect 7120 -10210 7130 -10090
rect 7250 -10210 7305 -10090
rect 7425 -10210 7470 -10090
rect 7590 -10210 7635 -10090
rect 7755 -10210 7800 -10090
rect 7920 -10210 7975 -10090
rect 8095 -10210 8140 -10090
rect 8260 -10210 8305 -10090
rect 8425 -10210 8470 -10090
rect 8590 -10210 8645 -10090
rect 8765 -10210 8810 -10090
rect 8930 -10210 8975 -10090
rect 9095 -10210 9140 -10090
rect 9260 -10210 9315 -10090
rect 9435 -10210 9480 -10090
rect 9600 -10210 9645 -10090
rect 9765 -10210 9810 -10090
rect 9930 -10210 9985 -10090
rect 10105 -10210 10150 -10090
rect 10270 -10210 10315 -10090
rect 10435 -10210 10480 -10090
rect 10600 -10210 10655 -10090
rect 10775 -10210 10820 -10090
rect 10940 -10210 10985 -10090
rect 11105 -10210 11150 -10090
rect 11270 -10210 11325 -10090
rect 11445 -10210 11490 -10090
rect 11610 -10210 11655 -10090
rect 11775 -10210 11820 -10090
rect 11940 -10210 11995 -10090
rect 12115 -10210 12160 -10090
rect 12280 -10210 12325 -10090
rect 12445 -10210 12490 -10090
rect 12610 -10210 12620 -10090
rect 7120 -10255 12620 -10210
rect 7120 -10375 7130 -10255
rect 7250 -10375 7305 -10255
rect 7425 -10375 7470 -10255
rect 7590 -10375 7635 -10255
rect 7755 -10375 7800 -10255
rect 7920 -10375 7975 -10255
rect 8095 -10375 8140 -10255
rect 8260 -10375 8305 -10255
rect 8425 -10375 8470 -10255
rect 8590 -10375 8645 -10255
rect 8765 -10375 8810 -10255
rect 8930 -10375 8975 -10255
rect 9095 -10375 9140 -10255
rect 9260 -10375 9315 -10255
rect 9435 -10375 9480 -10255
rect 9600 -10375 9645 -10255
rect 9765 -10375 9810 -10255
rect 9930 -10375 9985 -10255
rect 10105 -10375 10150 -10255
rect 10270 -10375 10315 -10255
rect 10435 -10375 10480 -10255
rect 10600 -10375 10655 -10255
rect 10775 -10375 10820 -10255
rect 10940 -10375 10985 -10255
rect 11105 -10375 11150 -10255
rect 11270 -10375 11325 -10255
rect 11445 -10375 11490 -10255
rect 11610 -10375 11655 -10255
rect 11775 -10375 11820 -10255
rect 11940 -10375 11995 -10255
rect 12115 -10375 12160 -10255
rect 12280 -10375 12325 -10255
rect 12445 -10375 12490 -10255
rect 12610 -10375 12620 -10255
rect 7120 -10420 12620 -10375
rect 7120 -10540 7130 -10420
rect 7250 -10540 7305 -10420
rect 7425 -10540 7470 -10420
rect 7590 -10540 7635 -10420
rect 7755 -10540 7800 -10420
rect 7920 -10540 7975 -10420
rect 8095 -10540 8140 -10420
rect 8260 -10540 8305 -10420
rect 8425 -10540 8470 -10420
rect 8590 -10540 8645 -10420
rect 8765 -10540 8810 -10420
rect 8930 -10540 8975 -10420
rect 9095 -10540 9140 -10420
rect 9260 -10540 9315 -10420
rect 9435 -10540 9480 -10420
rect 9600 -10540 9645 -10420
rect 9765 -10540 9810 -10420
rect 9930 -10540 9985 -10420
rect 10105 -10540 10150 -10420
rect 10270 -10540 10315 -10420
rect 10435 -10540 10480 -10420
rect 10600 -10540 10655 -10420
rect 10775 -10540 10820 -10420
rect 10940 -10540 10985 -10420
rect 11105 -10540 11150 -10420
rect 11270 -10540 11325 -10420
rect 11445 -10540 11490 -10420
rect 11610 -10540 11655 -10420
rect 11775 -10540 11820 -10420
rect 11940 -10540 11995 -10420
rect 12115 -10540 12160 -10420
rect 12280 -10540 12325 -10420
rect 12445 -10540 12490 -10420
rect 12610 -10540 12620 -10420
rect 7120 -10585 12620 -10540
rect 7120 -10705 7130 -10585
rect 7250 -10705 7305 -10585
rect 7425 -10705 7470 -10585
rect 7590 -10705 7635 -10585
rect 7755 -10705 7800 -10585
rect 7920 -10705 7975 -10585
rect 8095 -10705 8140 -10585
rect 8260 -10705 8305 -10585
rect 8425 -10705 8470 -10585
rect 8590 -10705 8645 -10585
rect 8765 -10705 8810 -10585
rect 8930 -10705 8975 -10585
rect 9095 -10705 9140 -10585
rect 9260 -10705 9315 -10585
rect 9435 -10705 9480 -10585
rect 9600 -10705 9645 -10585
rect 9765 -10705 9810 -10585
rect 9930 -10705 9985 -10585
rect 10105 -10705 10150 -10585
rect 10270 -10705 10315 -10585
rect 10435 -10705 10480 -10585
rect 10600 -10705 10655 -10585
rect 10775 -10705 10820 -10585
rect 10940 -10705 10985 -10585
rect 11105 -10705 11150 -10585
rect 11270 -10705 11325 -10585
rect 11445 -10705 11490 -10585
rect 11610 -10705 11655 -10585
rect 11775 -10705 11820 -10585
rect 11940 -10705 11995 -10585
rect 12115 -10705 12160 -10585
rect 12280 -10705 12325 -10585
rect 12445 -10705 12490 -10585
rect 12610 -10705 12620 -10585
rect 7120 -10760 12620 -10705
rect 7120 -10880 7130 -10760
rect 7250 -10880 7305 -10760
rect 7425 -10880 7470 -10760
rect 7590 -10880 7635 -10760
rect 7755 -10880 7800 -10760
rect 7920 -10880 7975 -10760
rect 8095 -10880 8140 -10760
rect 8260 -10880 8305 -10760
rect 8425 -10880 8470 -10760
rect 8590 -10880 8645 -10760
rect 8765 -10880 8810 -10760
rect 8930 -10880 8975 -10760
rect 9095 -10880 9140 -10760
rect 9260 -10880 9315 -10760
rect 9435 -10880 9480 -10760
rect 9600 -10880 9645 -10760
rect 9765 -10880 9810 -10760
rect 9930 -10880 9985 -10760
rect 10105 -10880 10150 -10760
rect 10270 -10880 10315 -10760
rect 10435 -10880 10480 -10760
rect 10600 -10880 10655 -10760
rect 10775 -10880 10820 -10760
rect 10940 -10880 10985 -10760
rect 11105 -10880 11150 -10760
rect 11270 -10880 11325 -10760
rect 11445 -10880 11490 -10760
rect 11610 -10880 11655 -10760
rect 11775 -10880 11820 -10760
rect 11940 -10880 11995 -10760
rect 12115 -10880 12160 -10760
rect 12280 -10880 12325 -10760
rect 12445 -10880 12490 -10760
rect 12610 -10880 12620 -10760
rect 7120 -10925 12620 -10880
rect 7120 -11045 7130 -10925
rect 7250 -11045 7305 -10925
rect 7425 -11045 7470 -10925
rect 7590 -11045 7635 -10925
rect 7755 -11045 7800 -10925
rect 7920 -11045 7975 -10925
rect 8095 -11045 8140 -10925
rect 8260 -11045 8305 -10925
rect 8425 -11045 8470 -10925
rect 8590 -11045 8645 -10925
rect 8765 -11045 8810 -10925
rect 8930 -11045 8975 -10925
rect 9095 -11045 9140 -10925
rect 9260 -11045 9315 -10925
rect 9435 -11045 9480 -10925
rect 9600 -11045 9645 -10925
rect 9765 -11045 9810 -10925
rect 9930 -11045 9985 -10925
rect 10105 -11045 10150 -10925
rect 10270 -11045 10315 -10925
rect 10435 -11045 10480 -10925
rect 10600 -11045 10655 -10925
rect 10775 -11045 10820 -10925
rect 10940 -11045 10985 -10925
rect 11105 -11045 11150 -10925
rect 11270 -11045 11325 -10925
rect 11445 -11045 11490 -10925
rect 11610 -11045 11655 -10925
rect 11775 -11045 11820 -10925
rect 11940 -11045 11995 -10925
rect 12115 -11045 12160 -10925
rect 12280 -11045 12325 -10925
rect 12445 -11045 12490 -10925
rect 12610 -11045 12620 -10925
rect 7120 -11090 12620 -11045
rect 7120 -11210 7130 -11090
rect 7250 -11210 7305 -11090
rect 7425 -11210 7470 -11090
rect 7590 -11210 7635 -11090
rect 7755 -11210 7800 -11090
rect 7920 -11210 7975 -11090
rect 8095 -11210 8140 -11090
rect 8260 -11210 8305 -11090
rect 8425 -11210 8470 -11090
rect 8590 -11210 8645 -11090
rect 8765 -11210 8810 -11090
rect 8930 -11210 8975 -11090
rect 9095 -11210 9140 -11090
rect 9260 -11210 9315 -11090
rect 9435 -11210 9480 -11090
rect 9600 -11210 9645 -11090
rect 9765 -11210 9810 -11090
rect 9930 -11210 9985 -11090
rect 10105 -11210 10150 -11090
rect 10270 -11210 10315 -11090
rect 10435 -11210 10480 -11090
rect 10600 -11210 10655 -11090
rect 10775 -11210 10820 -11090
rect 10940 -11210 10985 -11090
rect 11105 -11210 11150 -11090
rect 11270 -11210 11325 -11090
rect 11445 -11210 11490 -11090
rect 11610 -11210 11655 -11090
rect 11775 -11210 11820 -11090
rect 11940 -11210 11995 -11090
rect 12115 -11210 12160 -11090
rect 12280 -11210 12325 -11090
rect 12445 -11210 12490 -11090
rect 12610 -11210 12620 -11090
rect 7120 -11255 12620 -11210
rect 7120 -11375 7130 -11255
rect 7250 -11375 7305 -11255
rect 7425 -11375 7470 -11255
rect 7590 -11375 7635 -11255
rect 7755 -11375 7800 -11255
rect 7920 -11375 7975 -11255
rect 8095 -11375 8140 -11255
rect 8260 -11375 8305 -11255
rect 8425 -11375 8470 -11255
rect 8590 -11375 8645 -11255
rect 8765 -11375 8810 -11255
rect 8930 -11375 8975 -11255
rect 9095 -11375 9140 -11255
rect 9260 -11375 9315 -11255
rect 9435 -11375 9480 -11255
rect 9600 -11375 9645 -11255
rect 9765 -11375 9810 -11255
rect 9930 -11375 9985 -11255
rect 10105 -11375 10150 -11255
rect 10270 -11375 10315 -11255
rect 10435 -11375 10480 -11255
rect 10600 -11375 10655 -11255
rect 10775 -11375 10820 -11255
rect 10940 -11375 10985 -11255
rect 11105 -11375 11150 -11255
rect 11270 -11375 11325 -11255
rect 11445 -11375 11490 -11255
rect 11610 -11375 11655 -11255
rect 11775 -11375 11820 -11255
rect 11940 -11375 11995 -11255
rect 12115 -11375 12160 -11255
rect 12280 -11375 12325 -11255
rect 12445 -11375 12490 -11255
rect 12610 -11375 12620 -11255
rect 7120 -11430 12620 -11375
rect 7120 -11550 7130 -11430
rect 7250 -11550 7305 -11430
rect 7425 -11550 7470 -11430
rect 7590 -11550 7635 -11430
rect 7755 -11550 7800 -11430
rect 7920 -11550 7975 -11430
rect 8095 -11550 8140 -11430
rect 8260 -11550 8305 -11430
rect 8425 -11550 8470 -11430
rect 8590 -11550 8645 -11430
rect 8765 -11550 8810 -11430
rect 8930 -11550 8975 -11430
rect 9095 -11550 9140 -11430
rect 9260 -11550 9315 -11430
rect 9435 -11550 9480 -11430
rect 9600 -11550 9645 -11430
rect 9765 -11550 9810 -11430
rect 9930 -11550 9985 -11430
rect 10105 -11550 10150 -11430
rect 10270 -11550 10315 -11430
rect 10435 -11550 10480 -11430
rect 10600 -11550 10655 -11430
rect 10775 -11550 10820 -11430
rect 10940 -11550 10985 -11430
rect 11105 -11550 11150 -11430
rect 11270 -11550 11325 -11430
rect 11445 -11550 11490 -11430
rect 11610 -11550 11655 -11430
rect 11775 -11550 11820 -11430
rect 11940 -11550 11995 -11430
rect 12115 -11550 12160 -11430
rect 12280 -11550 12325 -11430
rect 12445 -11550 12490 -11430
rect 12610 -11550 12620 -11430
rect 7120 -11595 12620 -11550
rect 7120 -11715 7130 -11595
rect 7250 -11715 7305 -11595
rect 7425 -11715 7470 -11595
rect 7590 -11715 7635 -11595
rect 7755 -11715 7800 -11595
rect 7920 -11715 7975 -11595
rect 8095 -11715 8140 -11595
rect 8260 -11715 8305 -11595
rect 8425 -11715 8470 -11595
rect 8590 -11715 8645 -11595
rect 8765 -11715 8810 -11595
rect 8930 -11715 8975 -11595
rect 9095 -11715 9140 -11595
rect 9260 -11715 9315 -11595
rect 9435 -11715 9480 -11595
rect 9600 -11715 9645 -11595
rect 9765 -11715 9810 -11595
rect 9930 -11715 9985 -11595
rect 10105 -11715 10150 -11595
rect 10270 -11715 10315 -11595
rect 10435 -11715 10480 -11595
rect 10600 -11715 10655 -11595
rect 10775 -11715 10820 -11595
rect 10940 -11715 10985 -11595
rect 11105 -11715 11150 -11595
rect 11270 -11715 11325 -11595
rect 11445 -11715 11490 -11595
rect 11610 -11715 11655 -11595
rect 11775 -11715 11820 -11595
rect 11940 -11715 11995 -11595
rect 12115 -11715 12160 -11595
rect 12280 -11715 12325 -11595
rect 12445 -11715 12490 -11595
rect 12610 -11715 12620 -11595
rect 7120 -11760 12620 -11715
rect 7120 -11880 7130 -11760
rect 7250 -11880 7305 -11760
rect 7425 -11880 7470 -11760
rect 7590 -11880 7635 -11760
rect 7755 -11880 7800 -11760
rect 7920 -11880 7975 -11760
rect 8095 -11880 8140 -11760
rect 8260 -11880 8305 -11760
rect 8425 -11880 8470 -11760
rect 8590 -11880 8645 -11760
rect 8765 -11880 8810 -11760
rect 8930 -11880 8975 -11760
rect 9095 -11880 9140 -11760
rect 9260 -11880 9315 -11760
rect 9435 -11880 9480 -11760
rect 9600 -11880 9645 -11760
rect 9765 -11880 9810 -11760
rect 9930 -11880 9985 -11760
rect 10105 -11880 10150 -11760
rect 10270 -11880 10315 -11760
rect 10435 -11880 10480 -11760
rect 10600 -11880 10655 -11760
rect 10775 -11880 10820 -11760
rect 10940 -11880 10985 -11760
rect 11105 -11880 11150 -11760
rect 11270 -11880 11325 -11760
rect 11445 -11880 11490 -11760
rect 11610 -11880 11655 -11760
rect 11775 -11880 11820 -11760
rect 11940 -11880 11995 -11760
rect 12115 -11880 12160 -11760
rect 12280 -11880 12325 -11760
rect 12445 -11880 12490 -11760
rect 12610 -11880 12620 -11760
rect 7120 -11925 12620 -11880
rect 7120 -12045 7130 -11925
rect 7250 -12045 7305 -11925
rect 7425 -12045 7470 -11925
rect 7590 -12045 7635 -11925
rect 7755 -12045 7800 -11925
rect 7920 -12045 7975 -11925
rect 8095 -12045 8140 -11925
rect 8260 -12045 8305 -11925
rect 8425 -12045 8470 -11925
rect 8590 -12045 8645 -11925
rect 8765 -12045 8810 -11925
rect 8930 -12045 8975 -11925
rect 9095 -12045 9140 -11925
rect 9260 -12045 9315 -11925
rect 9435 -12045 9480 -11925
rect 9600 -12045 9645 -11925
rect 9765 -12045 9810 -11925
rect 9930 -12045 9985 -11925
rect 10105 -12045 10150 -11925
rect 10270 -12045 10315 -11925
rect 10435 -12045 10480 -11925
rect 10600 -12045 10655 -11925
rect 10775 -12045 10820 -11925
rect 10940 -12045 10985 -11925
rect 11105 -12045 11150 -11925
rect 11270 -12045 11325 -11925
rect 11445 -12045 11490 -11925
rect 11610 -12045 11655 -11925
rect 11775 -12045 11820 -11925
rect 11940 -12045 11995 -11925
rect 12115 -12045 12160 -11925
rect 12280 -12045 12325 -11925
rect 12445 -12045 12490 -11925
rect 12610 -12045 12620 -11925
rect 7120 -12100 12620 -12045
rect 7120 -12220 7130 -12100
rect 7250 -12220 7305 -12100
rect 7425 -12220 7470 -12100
rect 7590 -12220 7635 -12100
rect 7755 -12220 7800 -12100
rect 7920 -12220 7975 -12100
rect 8095 -12220 8140 -12100
rect 8260 -12220 8305 -12100
rect 8425 -12220 8470 -12100
rect 8590 -12220 8645 -12100
rect 8765 -12220 8810 -12100
rect 8930 -12220 8975 -12100
rect 9095 -12220 9140 -12100
rect 9260 -12220 9315 -12100
rect 9435 -12220 9480 -12100
rect 9600 -12220 9645 -12100
rect 9765 -12220 9810 -12100
rect 9930 -12220 9985 -12100
rect 10105 -12220 10150 -12100
rect 10270 -12220 10315 -12100
rect 10435 -12220 10480 -12100
rect 10600 -12220 10655 -12100
rect 10775 -12220 10820 -12100
rect 10940 -12220 10985 -12100
rect 11105 -12220 11150 -12100
rect 11270 -12220 11325 -12100
rect 11445 -12220 11490 -12100
rect 11610 -12220 11655 -12100
rect 11775 -12220 11820 -12100
rect 11940 -12220 11995 -12100
rect 12115 -12220 12160 -12100
rect 12280 -12220 12325 -12100
rect 12445 -12220 12490 -12100
rect 12610 -12220 12620 -12100
rect 7120 -12265 12620 -12220
rect 7120 -12385 7130 -12265
rect 7250 -12385 7305 -12265
rect 7425 -12385 7470 -12265
rect 7590 -12385 7635 -12265
rect 7755 -12385 7800 -12265
rect 7920 -12385 7975 -12265
rect 8095 -12385 8140 -12265
rect 8260 -12385 8305 -12265
rect 8425 -12385 8470 -12265
rect 8590 -12385 8645 -12265
rect 8765 -12385 8810 -12265
rect 8930 -12385 8975 -12265
rect 9095 -12385 9140 -12265
rect 9260 -12385 9315 -12265
rect 9435 -12385 9480 -12265
rect 9600 -12385 9645 -12265
rect 9765 -12385 9810 -12265
rect 9930 -12385 9985 -12265
rect 10105 -12385 10150 -12265
rect 10270 -12385 10315 -12265
rect 10435 -12385 10480 -12265
rect 10600 -12385 10655 -12265
rect 10775 -12385 10820 -12265
rect 10940 -12385 10985 -12265
rect 11105 -12385 11150 -12265
rect 11270 -12385 11325 -12265
rect 11445 -12385 11490 -12265
rect 11610 -12385 11655 -12265
rect 11775 -12385 11820 -12265
rect 11940 -12385 11995 -12265
rect 12115 -12385 12160 -12265
rect 12280 -12385 12325 -12265
rect 12445 -12385 12490 -12265
rect 12610 -12385 12620 -12265
rect 7120 -12430 12620 -12385
rect 7120 -12550 7130 -12430
rect 7250 -12550 7305 -12430
rect 7425 -12550 7470 -12430
rect 7590 -12550 7635 -12430
rect 7755 -12550 7800 -12430
rect 7920 -12550 7975 -12430
rect 8095 -12550 8140 -12430
rect 8260 -12550 8305 -12430
rect 8425 -12550 8470 -12430
rect 8590 -12550 8645 -12430
rect 8765 -12550 8810 -12430
rect 8930 -12550 8975 -12430
rect 9095 -12550 9140 -12430
rect 9260 -12550 9315 -12430
rect 9435 -12550 9480 -12430
rect 9600 -12550 9645 -12430
rect 9765 -12550 9810 -12430
rect 9930 -12550 9985 -12430
rect 10105 -12550 10150 -12430
rect 10270 -12550 10315 -12430
rect 10435 -12550 10480 -12430
rect 10600 -12550 10655 -12430
rect 10775 -12550 10820 -12430
rect 10940 -12550 10985 -12430
rect 11105 -12550 11150 -12430
rect 11270 -12550 11325 -12430
rect 11445 -12550 11490 -12430
rect 11610 -12550 11655 -12430
rect 11775 -12550 11820 -12430
rect 11940 -12550 11995 -12430
rect 12115 -12550 12160 -12430
rect 12280 -12550 12325 -12430
rect 12445 -12550 12490 -12430
rect 12610 -12550 12620 -12430
rect 7120 -12595 12620 -12550
rect 7120 -12715 7130 -12595
rect 7250 -12715 7305 -12595
rect 7425 -12715 7470 -12595
rect 7590 -12715 7635 -12595
rect 7755 -12715 7800 -12595
rect 7920 -12715 7975 -12595
rect 8095 -12715 8140 -12595
rect 8260 -12715 8305 -12595
rect 8425 -12715 8470 -12595
rect 8590 -12715 8645 -12595
rect 8765 -12715 8810 -12595
rect 8930 -12715 8975 -12595
rect 9095 -12715 9140 -12595
rect 9260 -12715 9315 -12595
rect 9435 -12715 9480 -12595
rect 9600 -12715 9645 -12595
rect 9765 -12715 9810 -12595
rect 9930 -12715 9985 -12595
rect 10105 -12715 10150 -12595
rect 10270 -12715 10315 -12595
rect 10435 -12715 10480 -12595
rect 10600 -12715 10655 -12595
rect 10775 -12715 10820 -12595
rect 10940 -12715 10985 -12595
rect 11105 -12715 11150 -12595
rect 11270 -12715 11325 -12595
rect 11445 -12715 11490 -12595
rect 11610 -12715 11655 -12595
rect 11775 -12715 11820 -12595
rect 11940 -12715 11995 -12595
rect 12115 -12715 12160 -12595
rect 12280 -12715 12325 -12595
rect 12445 -12715 12490 -12595
rect 12610 -12715 12620 -12595
rect 7120 -12770 12620 -12715
rect 7120 -12890 7130 -12770
rect 7250 -12890 7305 -12770
rect 7425 -12890 7470 -12770
rect 7590 -12890 7635 -12770
rect 7755 -12890 7800 -12770
rect 7920 -12890 7975 -12770
rect 8095 -12890 8140 -12770
rect 8260 -12890 8305 -12770
rect 8425 -12890 8470 -12770
rect 8590 -12890 8645 -12770
rect 8765 -12890 8810 -12770
rect 8930 -12890 8975 -12770
rect 9095 -12890 9140 -12770
rect 9260 -12890 9315 -12770
rect 9435 -12890 9480 -12770
rect 9600 -12890 9645 -12770
rect 9765 -12890 9810 -12770
rect 9930 -12890 9985 -12770
rect 10105 -12890 10150 -12770
rect 10270 -12890 10315 -12770
rect 10435 -12890 10480 -12770
rect 10600 -12890 10655 -12770
rect 10775 -12890 10820 -12770
rect 10940 -12890 10985 -12770
rect 11105 -12890 11150 -12770
rect 11270 -12890 11325 -12770
rect 11445 -12890 11490 -12770
rect 11610 -12890 11655 -12770
rect 11775 -12890 11820 -12770
rect 11940 -12890 11995 -12770
rect 12115 -12890 12160 -12770
rect 12280 -12890 12325 -12770
rect 12445 -12890 12490 -12770
rect 12610 -12890 12620 -12770
rect 7120 -12935 12620 -12890
rect 7120 -13055 7130 -12935
rect 7250 -13055 7305 -12935
rect 7425 -13055 7470 -12935
rect 7590 -13055 7635 -12935
rect 7755 -13055 7800 -12935
rect 7920 -13055 7975 -12935
rect 8095 -13055 8140 -12935
rect 8260 -13055 8305 -12935
rect 8425 -13055 8470 -12935
rect 8590 -13055 8645 -12935
rect 8765 -13055 8810 -12935
rect 8930 -13055 8975 -12935
rect 9095 -13055 9140 -12935
rect 9260 -13055 9315 -12935
rect 9435 -13055 9480 -12935
rect 9600 -13055 9645 -12935
rect 9765 -13055 9810 -12935
rect 9930 -13055 9985 -12935
rect 10105 -13055 10150 -12935
rect 10270 -13055 10315 -12935
rect 10435 -13055 10480 -12935
rect 10600 -13055 10655 -12935
rect 10775 -13055 10820 -12935
rect 10940 -13055 10985 -12935
rect 11105 -13055 11150 -12935
rect 11270 -13055 11325 -12935
rect 11445 -13055 11490 -12935
rect 11610 -13055 11655 -12935
rect 11775 -13055 11820 -12935
rect 11940 -13055 11995 -12935
rect 12115 -13055 12160 -12935
rect 12280 -13055 12325 -12935
rect 12445 -13055 12490 -12935
rect 12610 -13055 12620 -12935
rect 7120 -13100 12620 -13055
rect 7120 -13220 7130 -13100
rect 7250 -13220 7305 -13100
rect 7425 -13220 7470 -13100
rect 7590 -13220 7635 -13100
rect 7755 -13220 7800 -13100
rect 7920 -13220 7975 -13100
rect 8095 -13220 8140 -13100
rect 8260 -13220 8305 -13100
rect 8425 -13220 8470 -13100
rect 8590 -13220 8645 -13100
rect 8765 -13220 8810 -13100
rect 8930 -13220 8975 -13100
rect 9095 -13220 9140 -13100
rect 9260 -13220 9315 -13100
rect 9435 -13220 9480 -13100
rect 9600 -13220 9645 -13100
rect 9765 -13220 9810 -13100
rect 9930 -13220 9985 -13100
rect 10105 -13220 10150 -13100
rect 10270 -13220 10315 -13100
rect 10435 -13220 10480 -13100
rect 10600 -13220 10655 -13100
rect 10775 -13220 10820 -13100
rect 10940 -13220 10985 -13100
rect 11105 -13220 11150 -13100
rect 11270 -13220 11325 -13100
rect 11445 -13220 11490 -13100
rect 11610 -13220 11655 -13100
rect 11775 -13220 11820 -13100
rect 11940 -13220 11995 -13100
rect 12115 -13220 12160 -13100
rect 12280 -13220 12325 -13100
rect 12445 -13220 12490 -13100
rect 12610 -13220 12620 -13100
rect 7120 -13265 12620 -13220
rect 7120 -13385 7130 -13265
rect 7250 -13385 7305 -13265
rect 7425 -13385 7470 -13265
rect 7590 -13385 7635 -13265
rect 7755 -13385 7800 -13265
rect 7920 -13385 7975 -13265
rect 8095 -13385 8140 -13265
rect 8260 -13385 8305 -13265
rect 8425 -13385 8470 -13265
rect 8590 -13385 8645 -13265
rect 8765 -13385 8810 -13265
rect 8930 -13385 8975 -13265
rect 9095 -13385 9140 -13265
rect 9260 -13385 9315 -13265
rect 9435 -13385 9480 -13265
rect 9600 -13385 9645 -13265
rect 9765 -13385 9810 -13265
rect 9930 -13385 9985 -13265
rect 10105 -13385 10150 -13265
rect 10270 -13385 10315 -13265
rect 10435 -13385 10480 -13265
rect 10600 -13385 10655 -13265
rect 10775 -13385 10820 -13265
rect 10940 -13385 10985 -13265
rect 11105 -13385 11150 -13265
rect 11270 -13385 11325 -13265
rect 11445 -13385 11490 -13265
rect 11610 -13385 11655 -13265
rect 11775 -13385 11820 -13265
rect 11940 -13385 11995 -13265
rect 12115 -13385 12160 -13265
rect 12280 -13385 12325 -13265
rect 12445 -13385 12490 -13265
rect 12610 -13385 12620 -13265
rect 7120 -13440 12620 -13385
rect 7120 -13560 7130 -13440
rect 7250 -13560 7305 -13440
rect 7425 -13560 7470 -13440
rect 7590 -13560 7635 -13440
rect 7755 -13560 7800 -13440
rect 7920 -13560 7975 -13440
rect 8095 -13560 8140 -13440
rect 8260 -13560 8305 -13440
rect 8425 -13560 8470 -13440
rect 8590 -13560 8645 -13440
rect 8765 -13560 8810 -13440
rect 8930 -13560 8975 -13440
rect 9095 -13560 9140 -13440
rect 9260 -13560 9315 -13440
rect 9435 -13560 9480 -13440
rect 9600 -13560 9645 -13440
rect 9765 -13560 9810 -13440
rect 9930 -13560 9985 -13440
rect 10105 -13560 10150 -13440
rect 10270 -13560 10315 -13440
rect 10435 -13560 10480 -13440
rect 10600 -13560 10655 -13440
rect 10775 -13560 10820 -13440
rect 10940 -13560 10985 -13440
rect 11105 -13560 11150 -13440
rect 11270 -13560 11325 -13440
rect 11445 -13560 11490 -13440
rect 11610 -13560 11655 -13440
rect 11775 -13560 11820 -13440
rect 11940 -13560 11995 -13440
rect 12115 -13560 12160 -13440
rect 12280 -13560 12325 -13440
rect 12445 -13560 12490 -13440
rect 12610 -13560 12620 -13440
rect 7120 -13605 12620 -13560
rect 7120 -13725 7130 -13605
rect 7250 -13725 7305 -13605
rect 7425 -13725 7470 -13605
rect 7590 -13725 7635 -13605
rect 7755 -13725 7800 -13605
rect 7920 -13725 7975 -13605
rect 8095 -13725 8140 -13605
rect 8260 -13725 8305 -13605
rect 8425 -13725 8470 -13605
rect 8590 -13725 8645 -13605
rect 8765 -13725 8810 -13605
rect 8930 -13725 8975 -13605
rect 9095 -13725 9140 -13605
rect 9260 -13725 9315 -13605
rect 9435 -13725 9480 -13605
rect 9600 -13725 9645 -13605
rect 9765 -13725 9810 -13605
rect 9930 -13725 9985 -13605
rect 10105 -13725 10150 -13605
rect 10270 -13725 10315 -13605
rect 10435 -13725 10480 -13605
rect 10600 -13725 10655 -13605
rect 10775 -13725 10820 -13605
rect 10940 -13725 10985 -13605
rect 11105 -13725 11150 -13605
rect 11270 -13725 11325 -13605
rect 11445 -13725 11490 -13605
rect 11610 -13725 11655 -13605
rect 11775 -13725 11820 -13605
rect 11940 -13725 11995 -13605
rect 12115 -13725 12160 -13605
rect 12280 -13725 12325 -13605
rect 12445 -13725 12490 -13605
rect 12610 -13725 12620 -13605
rect 7120 -13770 12620 -13725
rect 7120 -13890 7130 -13770
rect 7250 -13890 7305 -13770
rect 7425 -13890 7470 -13770
rect 7590 -13890 7635 -13770
rect 7755 -13890 7800 -13770
rect 7920 -13890 7975 -13770
rect 8095 -13890 8140 -13770
rect 8260 -13890 8305 -13770
rect 8425 -13890 8470 -13770
rect 8590 -13890 8645 -13770
rect 8765 -13890 8810 -13770
rect 8930 -13890 8975 -13770
rect 9095 -13890 9140 -13770
rect 9260 -13890 9315 -13770
rect 9435 -13890 9480 -13770
rect 9600 -13890 9645 -13770
rect 9765 -13890 9810 -13770
rect 9930 -13890 9985 -13770
rect 10105 -13890 10150 -13770
rect 10270 -13890 10315 -13770
rect 10435 -13890 10480 -13770
rect 10600 -13890 10655 -13770
rect 10775 -13890 10820 -13770
rect 10940 -13890 10985 -13770
rect 11105 -13890 11150 -13770
rect 11270 -13890 11325 -13770
rect 11445 -13890 11490 -13770
rect 11610 -13890 11655 -13770
rect 11775 -13890 11820 -13770
rect 11940 -13890 11995 -13770
rect 12115 -13890 12160 -13770
rect 12280 -13890 12325 -13770
rect 12445 -13890 12490 -13770
rect 12610 -13890 12620 -13770
rect 7120 -13935 12620 -13890
rect 7120 -14055 7130 -13935
rect 7250 -14055 7305 -13935
rect 7425 -14055 7470 -13935
rect 7590 -14055 7635 -13935
rect 7755 -14055 7800 -13935
rect 7920 -14055 7975 -13935
rect 8095 -14055 8140 -13935
rect 8260 -14055 8305 -13935
rect 8425 -14055 8470 -13935
rect 8590 -14055 8645 -13935
rect 8765 -14055 8810 -13935
rect 8930 -14055 8975 -13935
rect 9095 -14055 9140 -13935
rect 9260 -14055 9315 -13935
rect 9435 -14055 9480 -13935
rect 9600 -14055 9645 -13935
rect 9765 -14055 9810 -13935
rect 9930 -14055 9985 -13935
rect 10105 -14055 10150 -13935
rect 10270 -14055 10315 -13935
rect 10435 -14055 10480 -13935
rect 10600 -14055 10655 -13935
rect 10775 -14055 10820 -13935
rect 10940 -14055 10985 -13935
rect 11105 -14055 11150 -13935
rect 11270 -14055 11325 -13935
rect 11445 -14055 11490 -13935
rect 11610 -14055 11655 -13935
rect 11775 -14055 11820 -13935
rect 11940 -14055 11995 -13935
rect 12115 -14055 12160 -13935
rect 12280 -14055 12325 -13935
rect 12445 -14055 12490 -13935
rect 12610 -14055 12620 -13935
rect 7120 -14110 12620 -14055
rect 7120 -14230 7130 -14110
rect 7250 -14230 7305 -14110
rect 7425 -14230 7470 -14110
rect 7590 -14230 7635 -14110
rect 7755 -14230 7800 -14110
rect 7920 -14230 7975 -14110
rect 8095 -14230 8140 -14110
rect 8260 -14230 8305 -14110
rect 8425 -14230 8470 -14110
rect 8590 -14230 8645 -14110
rect 8765 -14230 8810 -14110
rect 8930 -14230 8975 -14110
rect 9095 -14230 9140 -14110
rect 9260 -14230 9315 -14110
rect 9435 -14230 9480 -14110
rect 9600 -14230 9645 -14110
rect 9765 -14230 9810 -14110
rect 9930 -14230 9985 -14110
rect 10105 -14230 10150 -14110
rect 10270 -14230 10315 -14110
rect 10435 -14230 10480 -14110
rect 10600 -14230 10655 -14110
rect 10775 -14230 10820 -14110
rect 10940 -14230 10985 -14110
rect 11105 -14230 11150 -14110
rect 11270 -14230 11325 -14110
rect 11445 -14230 11490 -14110
rect 11610 -14230 11655 -14110
rect 11775 -14230 11820 -14110
rect 11940 -14230 11995 -14110
rect 12115 -14230 12160 -14110
rect 12280 -14230 12325 -14110
rect 12445 -14230 12490 -14110
rect 12610 -14230 12620 -14110
rect 7120 -14275 12620 -14230
rect 7120 -14395 7130 -14275
rect 7250 -14395 7305 -14275
rect 7425 -14395 7470 -14275
rect 7590 -14395 7635 -14275
rect 7755 -14395 7800 -14275
rect 7920 -14395 7975 -14275
rect 8095 -14395 8140 -14275
rect 8260 -14395 8305 -14275
rect 8425 -14395 8470 -14275
rect 8590 -14395 8645 -14275
rect 8765 -14395 8810 -14275
rect 8930 -14395 8975 -14275
rect 9095 -14395 9140 -14275
rect 9260 -14395 9315 -14275
rect 9435 -14395 9480 -14275
rect 9600 -14395 9645 -14275
rect 9765 -14395 9810 -14275
rect 9930 -14395 9985 -14275
rect 10105 -14395 10150 -14275
rect 10270 -14395 10315 -14275
rect 10435 -14395 10480 -14275
rect 10600 -14395 10655 -14275
rect 10775 -14395 10820 -14275
rect 10940 -14395 10985 -14275
rect 11105 -14395 11150 -14275
rect 11270 -14395 11325 -14275
rect 11445 -14395 11490 -14275
rect 11610 -14395 11655 -14275
rect 11775 -14395 11820 -14275
rect 11940 -14395 11995 -14275
rect 12115 -14395 12160 -14275
rect 12280 -14395 12325 -14275
rect 12445 -14395 12490 -14275
rect 12610 -14395 12620 -14275
rect 7120 -14440 12620 -14395
rect 7120 -14560 7130 -14440
rect 7250 -14560 7305 -14440
rect 7425 -14560 7470 -14440
rect 7590 -14560 7635 -14440
rect 7755 -14560 7800 -14440
rect 7920 -14560 7975 -14440
rect 8095 -14560 8140 -14440
rect 8260 -14560 8305 -14440
rect 8425 -14560 8470 -14440
rect 8590 -14560 8645 -14440
rect 8765 -14560 8810 -14440
rect 8930 -14560 8975 -14440
rect 9095 -14560 9140 -14440
rect 9260 -14560 9315 -14440
rect 9435 -14560 9480 -14440
rect 9600 -14560 9645 -14440
rect 9765 -14560 9810 -14440
rect 9930 -14560 9985 -14440
rect 10105 -14560 10150 -14440
rect 10270 -14560 10315 -14440
rect 10435 -14560 10480 -14440
rect 10600 -14560 10655 -14440
rect 10775 -14560 10820 -14440
rect 10940 -14560 10985 -14440
rect 11105 -14560 11150 -14440
rect 11270 -14560 11325 -14440
rect 11445 -14560 11490 -14440
rect 11610 -14560 11655 -14440
rect 11775 -14560 11820 -14440
rect 11940 -14560 11995 -14440
rect 12115 -14560 12160 -14440
rect 12280 -14560 12325 -14440
rect 12445 -14560 12490 -14440
rect 12610 -14560 12620 -14440
rect 7120 -14605 12620 -14560
rect 7120 -14725 7130 -14605
rect 7250 -14725 7305 -14605
rect 7425 -14725 7470 -14605
rect 7590 -14725 7635 -14605
rect 7755 -14725 7800 -14605
rect 7920 -14725 7975 -14605
rect 8095 -14725 8140 -14605
rect 8260 -14725 8305 -14605
rect 8425 -14725 8470 -14605
rect 8590 -14725 8645 -14605
rect 8765 -14725 8810 -14605
rect 8930 -14725 8975 -14605
rect 9095 -14725 9140 -14605
rect 9260 -14725 9315 -14605
rect 9435 -14725 9480 -14605
rect 9600 -14725 9645 -14605
rect 9765 -14725 9810 -14605
rect 9930 -14725 9985 -14605
rect 10105 -14725 10150 -14605
rect 10270 -14725 10315 -14605
rect 10435 -14725 10480 -14605
rect 10600 -14725 10655 -14605
rect 10775 -14725 10820 -14605
rect 10940 -14725 10985 -14605
rect 11105 -14725 11150 -14605
rect 11270 -14725 11325 -14605
rect 11445 -14725 11490 -14605
rect 11610 -14725 11655 -14605
rect 11775 -14725 11820 -14605
rect 11940 -14725 11995 -14605
rect 12115 -14725 12160 -14605
rect 12280 -14725 12325 -14605
rect 12445 -14725 12490 -14605
rect 12610 -14725 12620 -14605
rect 7120 -14780 12620 -14725
rect 7120 -14900 7130 -14780
rect 7250 -14900 7305 -14780
rect 7425 -14900 7470 -14780
rect 7590 -14900 7635 -14780
rect 7755 -14900 7800 -14780
rect 7920 -14900 7975 -14780
rect 8095 -14900 8140 -14780
rect 8260 -14900 8305 -14780
rect 8425 -14900 8470 -14780
rect 8590 -14900 8645 -14780
rect 8765 -14900 8810 -14780
rect 8930 -14900 8975 -14780
rect 9095 -14900 9140 -14780
rect 9260 -14900 9315 -14780
rect 9435 -14900 9480 -14780
rect 9600 -14900 9645 -14780
rect 9765 -14900 9810 -14780
rect 9930 -14900 9985 -14780
rect 10105 -14900 10150 -14780
rect 10270 -14900 10315 -14780
rect 10435 -14900 10480 -14780
rect 10600 -14900 10655 -14780
rect 10775 -14900 10820 -14780
rect 10940 -14900 10985 -14780
rect 11105 -14900 11150 -14780
rect 11270 -14900 11325 -14780
rect 11445 -14900 11490 -14780
rect 11610 -14900 11655 -14780
rect 11775 -14900 11820 -14780
rect 11940 -14900 11995 -14780
rect 12115 -14900 12160 -14780
rect 12280 -14900 12325 -14780
rect 12445 -14900 12490 -14780
rect 12610 -14900 12620 -14780
rect 7120 -14945 12620 -14900
rect 7120 -15065 7130 -14945
rect 7250 -15065 7305 -14945
rect 7425 -15065 7470 -14945
rect 7590 -15065 7635 -14945
rect 7755 -15065 7800 -14945
rect 7920 -15065 7975 -14945
rect 8095 -15065 8140 -14945
rect 8260 -15065 8305 -14945
rect 8425 -15065 8470 -14945
rect 8590 -15065 8645 -14945
rect 8765 -15065 8810 -14945
rect 8930 -15065 8975 -14945
rect 9095 -15065 9140 -14945
rect 9260 -15065 9315 -14945
rect 9435 -15065 9480 -14945
rect 9600 -15065 9645 -14945
rect 9765 -15065 9810 -14945
rect 9930 -15065 9985 -14945
rect 10105 -15065 10150 -14945
rect 10270 -15065 10315 -14945
rect 10435 -15065 10480 -14945
rect 10600 -15065 10655 -14945
rect 10775 -15065 10820 -14945
rect 10940 -15065 10985 -14945
rect 11105 -15065 11150 -14945
rect 11270 -15065 11325 -14945
rect 11445 -15065 11490 -14945
rect 11610 -15065 11655 -14945
rect 11775 -15065 11820 -14945
rect 11940 -15065 11995 -14945
rect 12115 -15065 12160 -14945
rect 12280 -15065 12325 -14945
rect 12445 -15065 12490 -14945
rect 12610 -15065 12620 -14945
rect 7120 -15110 12620 -15065
rect 7120 -15230 7130 -15110
rect 7250 -15230 7305 -15110
rect 7425 -15230 7470 -15110
rect 7590 -15230 7635 -15110
rect 7755 -15230 7800 -15110
rect 7920 -15230 7975 -15110
rect 8095 -15230 8140 -15110
rect 8260 -15230 8305 -15110
rect 8425 -15230 8470 -15110
rect 8590 -15230 8645 -15110
rect 8765 -15230 8810 -15110
rect 8930 -15230 8975 -15110
rect 9095 -15230 9140 -15110
rect 9260 -15230 9315 -15110
rect 9435 -15230 9480 -15110
rect 9600 -15230 9645 -15110
rect 9765 -15230 9810 -15110
rect 9930 -15230 9985 -15110
rect 10105 -15230 10150 -15110
rect 10270 -15230 10315 -15110
rect 10435 -15230 10480 -15110
rect 10600 -15230 10655 -15110
rect 10775 -15230 10820 -15110
rect 10940 -15230 10985 -15110
rect 11105 -15230 11150 -15110
rect 11270 -15230 11325 -15110
rect 11445 -15230 11490 -15110
rect 11610 -15230 11655 -15110
rect 11775 -15230 11820 -15110
rect 11940 -15230 11995 -15110
rect 12115 -15230 12160 -15110
rect 12280 -15230 12325 -15110
rect 12445 -15230 12490 -15110
rect 12610 -15230 12620 -15110
rect 7120 -15275 12620 -15230
rect 7120 -15395 7130 -15275
rect 7250 -15395 7305 -15275
rect 7425 -15395 7470 -15275
rect 7590 -15395 7635 -15275
rect 7755 -15395 7800 -15275
rect 7920 -15395 7975 -15275
rect 8095 -15395 8140 -15275
rect 8260 -15395 8305 -15275
rect 8425 -15395 8470 -15275
rect 8590 -15395 8645 -15275
rect 8765 -15395 8810 -15275
rect 8930 -15395 8975 -15275
rect 9095 -15395 9140 -15275
rect 9260 -15395 9315 -15275
rect 9435 -15395 9480 -15275
rect 9600 -15395 9645 -15275
rect 9765 -15395 9810 -15275
rect 9930 -15395 9985 -15275
rect 10105 -15395 10150 -15275
rect 10270 -15395 10315 -15275
rect 10435 -15395 10480 -15275
rect 10600 -15395 10655 -15275
rect 10775 -15395 10820 -15275
rect 10940 -15395 10985 -15275
rect 11105 -15395 11150 -15275
rect 11270 -15395 11325 -15275
rect 11445 -15395 11490 -15275
rect 11610 -15395 11655 -15275
rect 11775 -15395 11820 -15275
rect 11940 -15395 11995 -15275
rect 12115 -15395 12160 -15275
rect 12280 -15395 12325 -15275
rect 12445 -15395 12490 -15275
rect 12610 -15395 12620 -15275
rect 7120 -15450 12620 -15395
rect 7120 -15570 7130 -15450
rect 7250 -15570 7305 -15450
rect 7425 -15570 7470 -15450
rect 7590 -15570 7635 -15450
rect 7755 -15570 7800 -15450
rect 7920 -15570 7975 -15450
rect 8095 -15570 8140 -15450
rect 8260 -15570 8305 -15450
rect 8425 -15570 8470 -15450
rect 8590 -15570 8645 -15450
rect 8765 -15570 8810 -15450
rect 8930 -15570 8975 -15450
rect 9095 -15570 9140 -15450
rect 9260 -15570 9315 -15450
rect 9435 -15570 9480 -15450
rect 9600 -15570 9645 -15450
rect 9765 -15570 9810 -15450
rect 9930 -15570 9985 -15450
rect 10105 -15570 10150 -15450
rect 10270 -15570 10315 -15450
rect 10435 -15570 10480 -15450
rect 10600 -15570 10655 -15450
rect 10775 -15570 10820 -15450
rect 10940 -15570 10985 -15450
rect 11105 -15570 11150 -15450
rect 11270 -15570 11325 -15450
rect 11445 -15570 11490 -15450
rect 11610 -15570 11655 -15450
rect 11775 -15570 11820 -15450
rect 11940 -15570 11995 -15450
rect 12115 -15570 12160 -15450
rect 12280 -15570 12325 -15450
rect 12445 -15570 12490 -15450
rect 12610 -15570 12620 -15450
rect 7120 -15580 12620 -15570
rect 12810 -10090 18310 -10080
rect 12810 -10210 12820 -10090
rect 12940 -10210 12995 -10090
rect 13115 -10210 13160 -10090
rect 13280 -10210 13325 -10090
rect 13445 -10210 13490 -10090
rect 13610 -10210 13665 -10090
rect 13785 -10210 13830 -10090
rect 13950 -10210 13995 -10090
rect 14115 -10210 14160 -10090
rect 14280 -10210 14335 -10090
rect 14455 -10210 14500 -10090
rect 14620 -10210 14665 -10090
rect 14785 -10210 14830 -10090
rect 14950 -10210 15005 -10090
rect 15125 -10210 15170 -10090
rect 15290 -10210 15335 -10090
rect 15455 -10210 15500 -10090
rect 15620 -10210 15675 -10090
rect 15795 -10210 15840 -10090
rect 15960 -10210 16005 -10090
rect 16125 -10210 16170 -10090
rect 16290 -10210 16345 -10090
rect 16465 -10210 16510 -10090
rect 16630 -10210 16675 -10090
rect 16795 -10210 16840 -10090
rect 16960 -10210 17015 -10090
rect 17135 -10210 17180 -10090
rect 17300 -10210 17345 -10090
rect 17465 -10210 17510 -10090
rect 17630 -10210 17685 -10090
rect 17805 -10210 17850 -10090
rect 17970 -10210 18015 -10090
rect 18135 -10210 18180 -10090
rect 18300 -10210 18310 -10090
rect 12810 -10255 18310 -10210
rect 12810 -10375 12820 -10255
rect 12940 -10375 12995 -10255
rect 13115 -10375 13160 -10255
rect 13280 -10375 13325 -10255
rect 13445 -10375 13490 -10255
rect 13610 -10375 13665 -10255
rect 13785 -10375 13830 -10255
rect 13950 -10375 13995 -10255
rect 14115 -10375 14160 -10255
rect 14280 -10375 14335 -10255
rect 14455 -10375 14500 -10255
rect 14620 -10375 14665 -10255
rect 14785 -10375 14830 -10255
rect 14950 -10375 15005 -10255
rect 15125 -10375 15170 -10255
rect 15290 -10375 15335 -10255
rect 15455 -10375 15500 -10255
rect 15620 -10375 15675 -10255
rect 15795 -10375 15840 -10255
rect 15960 -10375 16005 -10255
rect 16125 -10375 16170 -10255
rect 16290 -10375 16345 -10255
rect 16465 -10375 16510 -10255
rect 16630 -10375 16675 -10255
rect 16795 -10375 16840 -10255
rect 16960 -10375 17015 -10255
rect 17135 -10375 17180 -10255
rect 17300 -10375 17345 -10255
rect 17465 -10375 17510 -10255
rect 17630 -10375 17685 -10255
rect 17805 -10375 17850 -10255
rect 17970 -10375 18015 -10255
rect 18135 -10375 18180 -10255
rect 18300 -10375 18310 -10255
rect 12810 -10420 18310 -10375
rect 12810 -10540 12820 -10420
rect 12940 -10540 12995 -10420
rect 13115 -10540 13160 -10420
rect 13280 -10540 13325 -10420
rect 13445 -10540 13490 -10420
rect 13610 -10540 13665 -10420
rect 13785 -10540 13830 -10420
rect 13950 -10540 13995 -10420
rect 14115 -10540 14160 -10420
rect 14280 -10540 14335 -10420
rect 14455 -10540 14500 -10420
rect 14620 -10540 14665 -10420
rect 14785 -10540 14830 -10420
rect 14950 -10540 15005 -10420
rect 15125 -10540 15170 -10420
rect 15290 -10540 15335 -10420
rect 15455 -10540 15500 -10420
rect 15620 -10540 15675 -10420
rect 15795 -10540 15840 -10420
rect 15960 -10540 16005 -10420
rect 16125 -10540 16170 -10420
rect 16290 -10540 16345 -10420
rect 16465 -10540 16510 -10420
rect 16630 -10540 16675 -10420
rect 16795 -10540 16840 -10420
rect 16960 -10540 17015 -10420
rect 17135 -10540 17180 -10420
rect 17300 -10540 17345 -10420
rect 17465 -10540 17510 -10420
rect 17630 -10540 17685 -10420
rect 17805 -10540 17850 -10420
rect 17970 -10540 18015 -10420
rect 18135 -10540 18180 -10420
rect 18300 -10540 18310 -10420
rect 12810 -10585 18310 -10540
rect 12810 -10705 12820 -10585
rect 12940 -10705 12995 -10585
rect 13115 -10705 13160 -10585
rect 13280 -10705 13325 -10585
rect 13445 -10705 13490 -10585
rect 13610 -10705 13665 -10585
rect 13785 -10705 13830 -10585
rect 13950 -10705 13995 -10585
rect 14115 -10705 14160 -10585
rect 14280 -10705 14335 -10585
rect 14455 -10705 14500 -10585
rect 14620 -10705 14665 -10585
rect 14785 -10705 14830 -10585
rect 14950 -10705 15005 -10585
rect 15125 -10705 15170 -10585
rect 15290 -10705 15335 -10585
rect 15455 -10705 15500 -10585
rect 15620 -10705 15675 -10585
rect 15795 -10705 15840 -10585
rect 15960 -10705 16005 -10585
rect 16125 -10705 16170 -10585
rect 16290 -10705 16345 -10585
rect 16465 -10705 16510 -10585
rect 16630 -10705 16675 -10585
rect 16795 -10705 16840 -10585
rect 16960 -10705 17015 -10585
rect 17135 -10705 17180 -10585
rect 17300 -10705 17345 -10585
rect 17465 -10705 17510 -10585
rect 17630 -10705 17685 -10585
rect 17805 -10705 17850 -10585
rect 17970 -10705 18015 -10585
rect 18135 -10705 18180 -10585
rect 18300 -10705 18310 -10585
rect 12810 -10760 18310 -10705
rect 12810 -10880 12820 -10760
rect 12940 -10880 12995 -10760
rect 13115 -10880 13160 -10760
rect 13280 -10880 13325 -10760
rect 13445 -10880 13490 -10760
rect 13610 -10880 13665 -10760
rect 13785 -10880 13830 -10760
rect 13950 -10880 13995 -10760
rect 14115 -10880 14160 -10760
rect 14280 -10880 14335 -10760
rect 14455 -10880 14500 -10760
rect 14620 -10880 14665 -10760
rect 14785 -10880 14830 -10760
rect 14950 -10880 15005 -10760
rect 15125 -10880 15170 -10760
rect 15290 -10880 15335 -10760
rect 15455 -10880 15500 -10760
rect 15620 -10880 15675 -10760
rect 15795 -10880 15840 -10760
rect 15960 -10880 16005 -10760
rect 16125 -10880 16170 -10760
rect 16290 -10880 16345 -10760
rect 16465 -10880 16510 -10760
rect 16630 -10880 16675 -10760
rect 16795 -10880 16840 -10760
rect 16960 -10880 17015 -10760
rect 17135 -10880 17180 -10760
rect 17300 -10880 17345 -10760
rect 17465 -10880 17510 -10760
rect 17630 -10880 17685 -10760
rect 17805 -10880 17850 -10760
rect 17970 -10880 18015 -10760
rect 18135 -10880 18180 -10760
rect 18300 -10880 18310 -10760
rect 12810 -10925 18310 -10880
rect 12810 -11045 12820 -10925
rect 12940 -11045 12995 -10925
rect 13115 -11045 13160 -10925
rect 13280 -11045 13325 -10925
rect 13445 -11045 13490 -10925
rect 13610 -11045 13665 -10925
rect 13785 -11045 13830 -10925
rect 13950 -11045 13995 -10925
rect 14115 -11045 14160 -10925
rect 14280 -11045 14335 -10925
rect 14455 -11045 14500 -10925
rect 14620 -11045 14665 -10925
rect 14785 -11045 14830 -10925
rect 14950 -11045 15005 -10925
rect 15125 -11045 15170 -10925
rect 15290 -11045 15335 -10925
rect 15455 -11045 15500 -10925
rect 15620 -11045 15675 -10925
rect 15795 -11045 15840 -10925
rect 15960 -11045 16005 -10925
rect 16125 -11045 16170 -10925
rect 16290 -11045 16345 -10925
rect 16465 -11045 16510 -10925
rect 16630 -11045 16675 -10925
rect 16795 -11045 16840 -10925
rect 16960 -11045 17015 -10925
rect 17135 -11045 17180 -10925
rect 17300 -11045 17345 -10925
rect 17465 -11045 17510 -10925
rect 17630 -11045 17685 -10925
rect 17805 -11045 17850 -10925
rect 17970 -11045 18015 -10925
rect 18135 -11045 18180 -10925
rect 18300 -11045 18310 -10925
rect 12810 -11090 18310 -11045
rect 12810 -11210 12820 -11090
rect 12940 -11210 12995 -11090
rect 13115 -11210 13160 -11090
rect 13280 -11210 13325 -11090
rect 13445 -11210 13490 -11090
rect 13610 -11210 13665 -11090
rect 13785 -11210 13830 -11090
rect 13950 -11210 13995 -11090
rect 14115 -11210 14160 -11090
rect 14280 -11210 14335 -11090
rect 14455 -11210 14500 -11090
rect 14620 -11210 14665 -11090
rect 14785 -11210 14830 -11090
rect 14950 -11210 15005 -11090
rect 15125 -11210 15170 -11090
rect 15290 -11210 15335 -11090
rect 15455 -11210 15500 -11090
rect 15620 -11210 15675 -11090
rect 15795 -11210 15840 -11090
rect 15960 -11210 16005 -11090
rect 16125 -11210 16170 -11090
rect 16290 -11210 16345 -11090
rect 16465 -11210 16510 -11090
rect 16630 -11210 16675 -11090
rect 16795 -11210 16840 -11090
rect 16960 -11210 17015 -11090
rect 17135 -11210 17180 -11090
rect 17300 -11210 17345 -11090
rect 17465 -11210 17510 -11090
rect 17630 -11210 17685 -11090
rect 17805 -11210 17850 -11090
rect 17970 -11210 18015 -11090
rect 18135 -11210 18180 -11090
rect 18300 -11210 18310 -11090
rect 12810 -11255 18310 -11210
rect 12810 -11375 12820 -11255
rect 12940 -11375 12995 -11255
rect 13115 -11375 13160 -11255
rect 13280 -11375 13325 -11255
rect 13445 -11375 13490 -11255
rect 13610 -11375 13665 -11255
rect 13785 -11375 13830 -11255
rect 13950 -11375 13995 -11255
rect 14115 -11375 14160 -11255
rect 14280 -11375 14335 -11255
rect 14455 -11375 14500 -11255
rect 14620 -11375 14665 -11255
rect 14785 -11375 14830 -11255
rect 14950 -11375 15005 -11255
rect 15125 -11375 15170 -11255
rect 15290 -11375 15335 -11255
rect 15455 -11375 15500 -11255
rect 15620 -11375 15675 -11255
rect 15795 -11375 15840 -11255
rect 15960 -11375 16005 -11255
rect 16125 -11375 16170 -11255
rect 16290 -11375 16345 -11255
rect 16465 -11375 16510 -11255
rect 16630 -11375 16675 -11255
rect 16795 -11375 16840 -11255
rect 16960 -11375 17015 -11255
rect 17135 -11375 17180 -11255
rect 17300 -11375 17345 -11255
rect 17465 -11375 17510 -11255
rect 17630 -11375 17685 -11255
rect 17805 -11375 17850 -11255
rect 17970 -11375 18015 -11255
rect 18135 -11375 18180 -11255
rect 18300 -11375 18310 -11255
rect 12810 -11430 18310 -11375
rect 12810 -11550 12820 -11430
rect 12940 -11550 12995 -11430
rect 13115 -11550 13160 -11430
rect 13280 -11550 13325 -11430
rect 13445 -11550 13490 -11430
rect 13610 -11550 13665 -11430
rect 13785 -11550 13830 -11430
rect 13950 -11550 13995 -11430
rect 14115 -11550 14160 -11430
rect 14280 -11550 14335 -11430
rect 14455 -11550 14500 -11430
rect 14620 -11550 14665 -11430
rect 14785 -11550 14830 -11430
rect 14950 -11550 15005 -11430
rect 15125 -11550 15170 -11430
rect 15290 -11550 15335 -11430
rect 15455 -11550 15500 -11430
rect 15620 -11550 15675 -11430
rect 15795 -11550 15840 -11430
rect 15960 -11550 16005 -11430
rect 16125 -11550 16170 -11430
rect 16290 -11550 16345 -11430
rect 16465 -11550 16510 -11430
rect 16630 -11550 16675 -11430
rect 16795 -11550 16840 -11430
rect 16960 -11550 17015 -11430
rect 17135 -11550 17180 -11430
rect 17300 -11550 17345 -11430
rect 17465 -11550 17510 -11430
rect 17630 -11550 17685 -11430
rect 17805 -11550 17850 -11430
rect 17970 -11550 18015 -11430
rect 18135 -11550 18180 -11430
rect 18300 -11550 18310 -11430
rect 12810 -11595 18310 -11550
rect 12810 -11715 12820 -11595
rect 12940 -11715 12995 -11595
rect 13115 -11715 13160 -11595
rect 13280 -11715 13325 -11595
rect 13445 -11715 13490 -11595
rect 13610 -11715 13665 -11595
rect 13785 -11715 13830 -11595
rect 13950 -11715 13995 -11595
rect 14115 -11715 14160 -11595
rect 14280 -11715 14335 -11595
rect 14455 -11715 14500 -11595
rect 14620 -11715 14665 -11595
rect 14785 -11715 14830 -11595
rect 14950 -11715 15005 -11595
rect 15125 -11715 15170 -11595
rect 15290 -11715 15335 -11595
rect 15455 -11715 15500 -11595
rect 15620 -11715 15675 -11595
rect 15795 -11715 15840 -11595
rect 15960 -11715 16005 -11595
rect 16125 -11715 16170 -11595
rect 16290 -11715 16345 -11595
rect 16465 -11715 16510 -11595
rect 16630 -11715 16675 -11595
rect 16795 -11715 16840 -11595
rect 16960 -11715 17015 -11595
rect 17135 -11715 17180 -11595
rect 17300 -11715 17345 -11595
rect 17465 -11715 17510 -11595
rect 17630 -11715 17685 -11595
rect 17805 -11715 17850 -11595
rect 17970 -11715 18015 -11595
rect 18135 -11715 18180 -11595
rect 18300 -11715 18310 -11595
rect 12810 -11760 18310 -11715
rect 12810 -11880 12820 -11760
rect 12940 -11880 12995 -11760
rect 13115 -11880 13160 -11760
rect 13280 -11880 13325 -11760
rect 13445 -11880 13490 -11760
rect 13610 -11880 13665 -11760
rect 13785 -11880 13830 -11760
rect 13950 -11880 13995 -11760
rect 14115 -11880 14160 -11760
rect 14280 -11880 14335 -11760
rect 14455 -11880 14500 -11760
rect 14620 -11880 14665 -11760
rect 14785 -11880 14830 -11760
rect 14950 -11880 15005 -11760
rect 15125 -11880 15170 -11760
rect 15290 -11880 15335 -11760
rect 15455 -11880 15500 -11760
rect 15620 -11880 15675 -11760
rect 15795 -11880 15840 -11760
rect 15960 -11880 16005 -11760
rect 16125 -11880 16170 -11760
rect 16290 -11880 16345 -11760
rect 16465 -11880 16510 -11760
rect 16630 -11880 16675 -11760
rect 16795 -11880 16840 -11760
rect 16960 -11880 17015 -11760
rect 17135 -11880 17180 -11760
rect 17300 -11880 17345 -11760
rect 17465 -11880 17510 -11760
rect 17630 -11880 17685 -11760
rect 17805 -11880 17850 -11760
rect 17970 -11880 18015 -11760
rect 18135 -11880 18180 -11760
rect 18300 -11880 18310 -11760
rect 12810 -11925 18310 -11880
rect 12810 -12045 12820 -11925
rect 12940 -12045 12995 -11925
rect 13115 -12045 13160 -11925
rect 13280 -12045 13325 -11925
rect 13445 -12045 13490 -11925
rect 13610 -12045 13665 -11925
rect 13785 -12045 13830 -11925
rect 13950 -12045 13995 -11925
rect 14115 -12045 14160 -11925
rect 14280 -12045 14335 -11925
rect 14455 -12045 14500 -11925
rect 14620 -12045 14665 -11925
rect 14785 -12045 14830 -11925
rect 14950 -12045 15005 -11925
rect 15125 -12045 15170 -11925
rect 15290 -12045 15335 -11925
rect 15455 -12045 15500 -11925
rect 15620 -12045 15675 -11925
rect 15795 -12045 15840 -11925
rect 15960 -12045 16005 -11925
rect 16125 -12045 16170 -11925
rect 16290 -12045 16345 -11925
rect 16465 -12045 16510 -11925
rect 16630 -12045 16675 -11925
rect 16795 -12045 16840 -11925
rect 16960 -12045 17015 -11925
rect 17135 -12045 17180 -11925
rect 17300 -12045 17345 -11925
rect 17465 -12045 17510 -11925
rect 17630 -12045 17685 -11925
rect 17805 -12045 17850 -11925
rect 17970 -12045 18015 -11925
rect 18135 -12045 18180 -11925
rect 18300 -12045 18310 -11925
rect 12810 -12100 18310 -12045
rect 12810 -12220 12820 -12100
rect 12940 -12220 12995 -12100
rect 13115 -12220 13160 -12100
rect 13280 -12220 13325 -12100
rect 13445 -12220 13490 -12100
rect 13610 -12220 13665 -12100
rect 13785 -12220 13830 -12100
rect 13950 -12220 13995 -12100
rect 14115 -12220 14160 -12100
rect 14280 -12220 14335 -12100
rect 14455 -12220 14500 -12100
rect 14620 -12220 14665 -12100
rect 14785 -12220 14830 -12100
rect 14950 -12220 15005 -12100
rect 15125 -12220 15170 -12100
rect 15290 -12220 15335 -12100
rect 15455 -12220 15500 -12100
rect 15620 -12220 15675 -12100
rect 15795 -12220 15840 -12100
rect 15960 -12220 16005 -12100
rect 16125 -12220 16170 -12100
rect 16290 -12220 16345 -12100
rect 16465 -12220 16510 -12100
rect 16630 -12220 16675 -12100
rect 16795 -12220 16840 -12100
rect 16960 -12220 17015 -12100
rect 17135 -12220 17180 -12100
rect 17300 -12220 17345 -12100
rect 17465 -12220 17510 -12100
rect 17630 -12220 17685 -12100
rect 17805 -12220 17850 -12100
rect 17970 -12220 18015 -12100
rect 18135 -12220 18180 -12100
rect 18300 -12220 18310 -12100
rect 12810 -12265 18310 -12220
rect 12810 -12385 12820 -12265
rect 12940 -12385 12995 -12265
rect 13115 -12385 13160 -12265
rect 13280 -12385 13325 -12265
rect 13445 -12385 13490 -12265
rect 13610 -12385 13665 -12265
rect 13785 -12385 13830 -12265
rect 13950 -12385 13995 -12265
rect 14115 -12385 14160 -12265
rect 14280 -12385 14335 -12265
rect 14455 -12385 14500 -12265
rect 14620 -12385 14665 -12265
rect 14785 -12385 14830 -12265
rect 14950 -12385 15005 -12265
rect 15125 -12385 15170 -12265
rect 15290 -12385 15335 -12265
rect 15455 -12385 15500 -12265
rect 15620 -12385 15675 -12265
rect 15795 -12385 15840 -12265
rect 15960 -12385 16005 -12265
rect 16125 -12385 16170 -12265
rect 16290 -12385 16345 -12265
rect 16465 -12385 16510 -12265
rect 16630 -12385 16675 -12265
rect 16795 -12385 16840 -12265
rect 16960 -12385 17015 -12265
rect 17135 -12385 17180 -12265
rect 17300 -12385 17345 -12265
rect 17465 -12385 17510 -12265
rect 17630 -12385 17685 -12265
rect 17805 -12385 17850 -12265
rect 17970 -12385 18015 -12265
rect 18135 -12385 18180 -12265
rect 18300 -12385 18310 -12265
rect 12810 -12430 18310 -12385
rect 12810 -12550 12820 -12430
rect 12940 -12550 12995 -12430
rect 13115 -12550 13160 -12430
rect 13280 -12550 13325 -12430
rect 13445 -12550 13490 -12430
rect 13610 -12550 13665 -12430
rect 13785 -12550 13830 -12430
rect 13950 -12550 13995 -12430
rect 14115 -12550 14160 -12430
rect 14280 -12550 14335 -12430
rect 14455 -12550 14500 -12430
rect 14620 -12550 14665 -12430
rect 14785 -12550 14830 -12430
rect 14950 -12550 15005 -12430
rect 15125 -12550 15170 -12430
rect 15290 -12550 15335 -12430
rect 15455 -12550 15500 -12430
rect 15620 -12550 15675 -12430
rect 15795 -12550 15840 -12430
rect 15960 -12550 16005 -12430
rect 16125 -12550 16170 -12430
rect 16290 -12550 16345 -12430
rect 16465 -12550 16510 -12430
rect 16630 -12550 16675 -12430
rect 16795 -12550 16840 -12430
rect 16960 -12550 17015 -12430
rect 17135 -12550 17180 -12430
rect 17300 -12550 17345 -12430
rect 17465 -12550 17510 -12430
rect 17630 -12550 17685 -12430
rect 17805 -12550 17850 -12430
rect 17970 -12550 18015 -12430
rect 18135 -12550 18180 -12430
rect 18300 -12550 18310 -12430
rect 12810 -12595 18310 -12550
rect 12810 -12715 12820 -12595
rect 12940 -12715 12995 -12595
rect 13115 -12715 13160 -12595
rect 13280 -12715 13325 -12595
rect 13445 -12715 13490 -12595
rect 13610 -12715 13665 -12595
rect 13785 -12715 13830 -12595
rect 13950 -12715 13995 -12595
rect 14115 -12715 14160 -12595
rect 14280 -12715 14335 -12595
rect 14455 -12715 14500 -12595
rect 14620 -12715 14665 -12595
rect 14785 -12715 14830 -12595
rect 14950 -12715 15005 -12595
rect 15125 -12715 15170 -12595
rect 15290 -12715 15335 -12595
rect 15455 -12715 15500 -12595
rect 15620 -12715 15675 -12595
rect 15795 -12715 15840 -12595
rect 15960 -12715 16005 -12595
rect 16125 -12715 16170 -12595
rect 16290 -12715 16345 -12595
rect 16465 -12715 16510 -12595
rect 16630 -12715 16675 -12595
rect 16795 -12715 16840 -12595
rect 16960 -12715 17015 -12595
rect 17135 -12715 17180 -12595
rect 17300 -12715 17345 -12595
rect 17465 -12715 17510 -12595
rect 17630 -12715 17685 -12595
rect 17805 -12715 17850 -12595
rect 17970 -12715 18015 -12595
rect 18135 -12715 18180 -12595
rect 18300 -12715 18310 -12595
rect 12810 -12770 18310 -12715
rect 12810 -12890 12820 -12770
rect 12940 -12890 12995 -12770
rect 13115 -12890 13160 -12770
rect 13280 -12890 13325 -12770
rect 13445 -12890 13490 -12770
rect 13610 -12890 13665 -12770
rect 13785 -12890 13830 -12770
rect 13950 -12890 13995 -12770
rect 14115 -12890 14160 -12770
rect 14280 -12890 14335 -12770
rect 14455 -12890 14500 -12770
rect 14620 -12890 14665 -12770
rect 14785 -12890 14830 -12770
rect 14950 -12890 15005 -12770
rect 15125 -12890 15170 -12770
rect 15290 -12890 15335 -12770
rect 15455 -12890 15500 -12770
rect 15620 -12890 15675 -12770
rect 15795 -12890 15840 -12770
rect 15960 -12890 16005 -12770
rect 16125 -12890 16170 -12770
rect 16290 -12890 16345 -12770
rect 16465 -12890 16510 -12770
rect 16630 -12890 16675 -12770
rect 16795 -12890 16840 -12770
rect 16960 -12890 17015 -12770
rect 17135 -12890 17180 -12770
rect 17300 -12890 17345 -12770
rect 17465 -12890 17510 -12770
rect 17630 -12890 17685 -12770
rect 17805 -12890 17850 -12770
rect 17970 -12890 18015 -12770
rect 18135 -12890 18180 -12770
rect 18300 -12890 18310 -12770
rect 12810 -12935 18310 -12890
rect 12810 -13055 12820 -12935
rect 12940 -13055 12995 -12935
rect 13115 -13055 13160 -12935
rect 13280 -13055 13325 -12935
rect 13445 -13055 13490 -12935
rect 13610 -13055 13665 -12935
rect 13785 -13055 13830 -12935
rect 13950 -13055 13995 -12935
rect 14115 -13055 14160 -12935
rect 14280 -13055 14335 -12935
rect 14455 -13055 14500 -12935
rect 14620 -13055 14665 -12935
rect 14785 -13055 14830 -12935
rect 14950 -13055 15005 -12935
rect 15125 -13055 15170 -12935
rect 15290 -13055 15335 -12935
rect 15455 -13055 15500 -12935
rect 15620 -13055 15675 -12935
rect 15795 -13055 15840 -12935
rect 15960 -13055 16005 -12935
rect 16125 -13055 16170 -12935
rect 16290 -13055 16345 -12935
rect 16465 -13055 16510 -12935
rect 16630 -13055 16675 -12935
rect 16795 -13055 16840 -12935
rect 16960 -13055 17015 -12935
rect 17135 -13055 17180 -12935
rect 17300 -13055 17345 -12935
rect 17465 -13055 17510 -12935
rect 17630 -13055 17685 -12935
rect 17805 -13055 17850 -12935
rect 17970 -13055 18015 -12935
rect 18135 -13055 18180 -12935
rect 18300 -13055 18310 -12935
rect 12810 -13100 18310 -13055
rect 12810 -13220 12820 -13100
rect 12940 -13220 12995 -13100
rect 13115 -13220 13160 -13100
rect 13280 -13220 13325 -13100
rect 13445 -13220 13490 -13100
rect 13610 -13220 13665 -13100
rect 13785 -13220 13830 -13100
rect 13950 -13220 13995 -13100
rect 14115 -13220 14160 -13100
rect 14280 -13220 14335 -13100
rect 14455 -13220 14500 -13100
rect 14620 -13220 14665 -13100
rect 14785 -13220 14830 -13100
rect 14950 -13220 15005 -13100
rect 15125 -13220 15170 -13100
rect 15290 -13220 15335 -13100
rect 15455 -13220 15500 -13100
rect 15620 -13220 15675 -13100
rect 15795 -13220 15840 -13100
rect 15960 -13220 16005 -13100
rect 16125 -13220 16170 -13100
rect 16290 -13220 16345 -13100
rect 16465 -13220 16510 -13100
rect 16630 -13220 16675 -13100
rect 16795 -13220 16840 -13100
rect 16960 -13220 17015 -13100
rect 17135 -13220 17180 -13100
rect 17300 -13220 17345 -13100
rect 17465 -13220 17510 -13100
rect 17630 -13220 17685 -13100
rect 17805 -13220 17850 -13100
rect 17970 -13220 18015 -13100
rect 18135 -13220 18180 -13100
rect 18300 -13220 18310 -13100
rect 12810 -13265 18310 -13220
rect 12810 -13385 12820 -13265
rect 12940 -13385 12995 -13265
rect 13115 -13385 13160 -13265
rect 13280 -13385 13325 -13265
rect 13445 -13385 13490 -13265
rect 13610 -13385 13665 -13265
rect 13785 -13385 13830 -13265
rect 13950 -13385 13995 -13265
rect 14115 -13385 14160 -13265
rect 14280 -13385 14335 -13265
rect 14455 -13385 14500 -13265
rect 14620 -13385 14665 -13265
rect 14785 -13385 14830 -13265
rect 14950 -13385 15005 -13265
rect 15125 -13385 15170 -13265
rect 15290 -13385 15335 -13265
rect 15455 -13385 15500 -13265
rect 15620 -13385 15675 -13265
rect 15795 -13385 15840 -13265
rect 15960 -13385 16005 -13265
rect 16125 -13385 16170 -13265
rect 16290 -13385 16345 -13265
rect 16465 -13385 16510 -13265
rect 16630 -13385 16675 -13265
rect 16795 -13385 16840 -13265
rect 16960 -13385 17015 -13265
rect 17135 -13385 17180 -13265
rect 17300 -13385 17345 -13265
rect 17465 -13385 17510 -13265
rect 17630 -13385 17685 -13265
rect 17805 -13385 17850 -13265
rect 17970 -13385 18015 -13265
rect 18135 -13385 18180 -13265
rect 18300 -13385 18310 -13265
rect 12810 -13440 18310 -13385
rect 12810 -13560 12820 -13440
rect 12940 -13560 12995 -13440
rect 13115 -13560 13160 -13440
rect 13280 -13560 13325 -13440
rect 13445 -13560 13490 -13440
rect 13610 -13560 13665 -13440
rect 13785 -13560 13830 -13440
rect 13950 -13560 13995 -13440
rect 14115 -13560 14160 -13440
rect 14280 -13560 14335 -13440
rect 14455 -13560 14500 -13440
rect 14620 -13560 14665 -13440
rect 14785 -13560 14830 -13440
rect 14950 -13560 15005 -13440
rect 15125 -13560 15170 -13440
rect 15290 -13560 15335 -13440
rect 15455 -13560 15500 -13440
rect 15620 -13560 15675 -13440
rect 15795 -13560 15840 -13440
rect 15960 -13560 16005 -13440
rect 16125 -13560 16170 -13440
rect 16290 -13560 16345 -13440
rect 16465 -13560 16510 -13440
rect 16630 -13560 16675 -13440
rect 16795 -13560 16840 -13440
rect 16960 -13560 17015 -13440
rect 17135 -13560 17180 -13440
rect 17300 -13560 17345 -13440
rect 17465 -13560 17510 -13440
rect 17630 -13560 17685 -13440
rect 17805 -13560 17850 -13440
rect 17970 -13560 18015 -13440
rect 18135 -13560 18180 -13440
rect 18300 -13560 18310 -13440
rect 12810 -13605 18310 -13560
rect 12810 -13725 12820 -13605
rect 12940 -13725 12995 -13605
rect 13115 -13725 13160 -13605
rect 13280 -13725 13325 -13605
rect 13445 -13725 13490 -13605
rect 13610 -13725 13665 -13605
rect 13785 -13725 13830 -13605
rect 13950 -13725 13995 -13605
rect 14115 -13725 14160 -13605
rect 14280 -13725 14335 -13605
rect 14455 -13725 14500 -13605
rect 14620 -13725 14665 -13605
rect 14785 -13725 14830 -13605
rect 14950 -13725 15005 -13605
rect 15125 -13725 15170 -13605
rect 15290 -13725 15335 -13605
rect 15455 -13725 15500 -13605
rect 15620 -13725 15675 -13605
rect 15795 -13725 15840 -13605
rect 15960 -13725 16005 -13605
rect 16125 -13725 16170 -13605
rect 16290 -13725 16345 -13605
rect 16465 -13725 16510 -13605
rect 16630 -13725 16675 -13605
rect 16795 -13725 16840 -13605
rect 16960 -13725 17015 -13605
rect 17135 -13725 17180 -13605
rect 17300 -13725 17345 -13605
rect 17465 -13725 17510 -13605
rect 17630 -13725 17685 -13605
rect 17805 -13725 17850 -13605
rect 17970 -13725 18015 -13605
rect 18135 -13725 18180 -13605
rect 18300 -13725 18310 -13605
rect 12810 -13770 18310 -13725
rect 12810 -13890 12820 -13770
rect 12940 -13890 12995 -13770
rect 13115 -13890 13160 -13770
rect 13280 -13890 13325 -13770
rect 13445 -13890 13490 -13770
rect 13610 -13890 13665 -13770
rect 13785 -13890 13830 -13770
rect 13950 -13890 13995 -13770
rect 14115 -13890 14160 -13770
rect 14280 -13890 14335 -13770
rect 14455 -13890 14500 -13770
rect 14620 -13890 14665 -13770
rect 14785 -13890 14830 -13770
rect 14950 -13890 15005 -13770
rect 15125 -13890 15170 -13770
rect 15290 -13890 15335 -13770
rect 15455 -13890 15500 -13770
rect 15620 -13890 15675 -13770
rect 15795 -13890 15840 -13770
rect 15960 -13890 16005 -13770
rect 16125 -13890 16170 -13770
rect 16290 -13890 16345 -13770
rect 16465 -13890 16510 -13770
rect 16630 -13890 16675 -13770
rect 16795 -13890 16840 -13770
rect 16960 -13890 17015 -13770
rect 17135 -13890 17180 -13770
rect 17300 -13890 17345 -13770
rect 17465 -13890 17510 -13770
rect 17630 -13890 17685 -13770
rect 17805 -13890 17850 -13770
rect 17970 -13890 18015 -13770
rect 18135 -13890 18180 -13770
rect 18300 -13890 18310 -13770
rect 12810 -13935 18310 -13890
rect 12810 -14055 12820 -13935
rect 12940 -14055 12995 -13935
rect 13115 -14055 13160 -13935
rect 13280 -14055 13325 -13935
rect 13445 -14055 13490 -13935
rect 13610 -14055 13665 -13935
rect 13785 -14055 13830 -13935
rect 13950 -14055 13995 -13935
rect 14115 -14055 14160 -13935
rect 14280 -14055 14335 -13935
rect 14455 -14055 14500 -13935
rect 14620 -14055 14665 -13935
rect 14785 -14055 14830 -13935
rect 14950 -14055 15005 -13935
rect 15125 -14055 15170 -13935
rect 15290 -14055 15335 -13935
rect 15455 -14055 15500 -13935
rect 15620 -14055 15675 -13935
rect 15795 -14055 15840 -13935
rect 15960 -14055 16005 -13935
rect 16125 -14055 16170 -13935
rect 16290 -14055 16345 -13935
rect 16465 -14055 16510 -13935
rect 16630 -14055 16675 -13935
rect 16795 -14055 16840 -13935
rect 16960 -14055 17015 -13935
rect 17135 -14055 17180 -13935
rect 17300 -14055 17345 -13935
rect 17465 -14055 17510 -13935
rect 17630 -14055 17685 -13935
rect 17805 -14055 17850 -13935
rect 17970 -14055 18015 -13935
rect 18135 -14055 18180 -13935
rect 18300 -14055 18310 -13935
rect 12810 -14110 18310 -14055
rect 12810 -14230 12820 -14110
rect 12940 -14230 12995 -14110
rect 13115 -14230 13160 -14110
rect 13280 -14230 13325 -14110
rect 13445 -14230 13490 -14110
rect 13610 -14230 13665 -14110
rect 13785 -14230 13830 -14110
rect 13950 -14230 13995 -14110
rect 14115 -14230 14160 -14110
rect 14280 -14230 14335 -14110
rect 14455 -14230 14500 -14110
rect 14620 -14230 14665 -14110
rect 14785 -14230 14830 -14110
rect 14950 -14230 15005 -14110
rect 15125 -14230 15170 -14110
rect 15290 -14230 15335 -14110
rect 15455 -14230 15500 -14110
rect 15620 -14230 15675 -14110
rect 15795 -14230 15840 -14110
rect 15960 -14230 16005 -14110
rect 16125 -14230 16170 -14110
rect 16290 -14230 16345 -14110
rect 16465 -14230 16510 -14110
rect 16630 -14230 16675 -14110
rect 16795 -14230 16840 -14110
rect 16960 -14230 17015 -14110
rect 17135 -14230 17180 -14110
rect 17300 -14230 17345 -14110
rect 17465 -14230 17510 -14110
rect 17630 -14230 17685 -14110
rect 17805 -14230 17850 -14110
rect 17970 -14230 18015 -14110
rect 18135 -14230 18180 -14110
rect 18300 -14230 18310 -14110
rect 12810 -14275 18310 -14230
rect 12810 -14395 12820 -14275
rect 12940 -14395 12995 -14275
rect 13115 -14395 13160 -14275
rect 13280 -14395 13325 -14275
rect 13445 -14395 13490 -14275
rect 13610 -14395 13665 -14275
rect 13785 -14395 13830 -14275
rect 13950 -14395 13995 -14275
rect 14115 -14395 14160 -14275
rect 14280 -14395 14335 -14275
rect 14455 -14395 14500 -14275
rect 14620 -14395 14665 -14275
rect 14785 -14395 14830 -14275
rect 14950 -14395 15005 -14275
rect 15125 -14395 15170 -14275
rect 15290 -14395 15335 -14275
rect 15455 -14395 15500 -14275
rect 15620 -14395 15675 -14275
rect 15795 -14395 15840 -14275
rect 15960 -14395 16005 -14275
rect 16125 -14395 16170 -14275
rect 16290 -14395 16345 -14275
rect 16465 -14395 16510 -14275
rect 16630 -14395 16675 -14275
rect 16795 -14395 16840 -14275
rect 16960 -14395 17015 -14275
rect 17135 -14395 17180 -14275
rect 17300 -14395 17345 -14275
rect 17465 -14395 17510 -14275
rect 17630 -14395 17685 -14275
rect 17805 -14395 17850 -14275
rect 17970 -14395 18015 -14275
rect 18135 -14395 18180 -14275
rect 18300 -14395 18310 -14275
rect 12810 -14440 18310 -14395
rect 12810 -14560 12820 -14440
rect 12940 -14560 12995 -14440
rect 13115 -14560 13160 -14440
rect 13280 -14560 13325 -14440
rect 13445 -14560 13490 -14440
rect 13610 -14560 13665 -14440
rect 13785 -14560 13830 -14440
rect 13950 -14560 13995 -14440
rect 14115 -14560 14160 -14440
rect 14280 -14560 14335 -14440
rect 14455 -14560 14500 -14440
rect 14620 -14560 14665 -14440
rect 14785 -14560 14830 -14440
rect 14950 -14560 15005 -14440
rect 15125 -14560 15170 -14440
rect 15290 -14560 15335 -14440
rect 15455 -14560 15500 -14440
rect 15620 -14560 15675 -14440
rect 15795 -14560 15840 -14440
rect 15960 -14560 16005 -14440
rect 16125 -14560 16170 -14440
rect 16290 -14560 16345 -14440
rect 16465 -14560 16510 -14440
rect 16630 -14560 16675 -14440
rect 16795 -14560 16840 -14440
rect 16960 -14560 17015 -14440
rect 17135 -14560 17180 -14440
rect 17300 -14560 17345 -14440
rect 17465 -14560 17510 -14440
rect 17630 -14560 17685 -14440
rect 17805 -14560 17850 -14440
rect 17970 -14560 18015 -14440
rect 18135 -14560 18180 -14440
rect 18300 -14560 18310 -14440
rect 12810 -14605 18310 -14560
rect 12810 -14725 12820 -14605
rect 12940 -14725 12995 -14605
rect 13115 -14725 13160 -14605
rect 13280 -14725 13325 -14605
rect 13445 -14725 13490 -14605
rect 13610 -14725 13665 -14605
rect 13785 -14725 13830 -14605
rect 13950 -14725 13995 -14605
rect 14115 -14725 14160 -14605
rect 14280 -14725 14335 -14605
rect 14455 -14725 14500 -14605
rect 14620 -14725 14665 -14605
rect 14785 -14725 14830 -14605
rect 14950 -14725 15005 -14605
rect 15125 -14725 15170 -14605
rect 15290 -14725 15335 -14605
rect 15455 -14725 15500 -14605
rect 15620 -14725 15675 -14605
rect 15795 -14725 15840 -14605
rect 15960 -14725 16005 -14605
rect 16125 -14725 16170 -14605
rect 16290 -14725 16345 -14605
rect 16465 -14725 16510 -14605
rect 16630 -14725 16675 -14605
rect 16795 -14725 16840 -14605
rect 16960 -14725 17015 -14605
rect 17135 -14725 17180 -14605
rect 17300 -14725 17345 -14605
rect 17465 -14725 17510 -14605
rect 17630 -14725 17685 -14605
rect 17805 -14725 17850 -14605
rect 17970 -14725 18015 -14605
rect 18135 -14725 18180 -14605
rect 18300 -14725 18310 -14605
rect 12810 -14780 18310 -14725
rect 12810 -14900 12820 -14780
rect 12940 -14900 12995 -14780
rect 13115 -14900 13160 -14780
rect 13280 -14900 13325 -14780
rect 13445 -14900 13490 -14780
rect 13610 -14900 13665 -14780
rect 13785 -14900 13830 -14780
rect 13950 -14900 13995 -14780
rect 14115 -14900 14160 -14780
rect 14280 -14900 14335 -14780
rect 14455 -14900 14500 -14780
rect 14620 -14900 14665 -14780
rect 14785 -14900 14830 -14780
rect 14950 -14900 15005 -14780
rect 15125 -14900 15170 -14780
rect 15290 -14900 15335 -14780
rect 15455 -14900 15500 -14780
rect 15620 -14900 15675 -14780
rect 15795 -14900 15840 -14780
rect 15960 -14900 16005 -14780
rect 16125 -14900 16170 -14780
rect 16290 -14900 16345 -14780
rect 16465 -14900 16510 -14780
rect 16630 -14900 16675 -14780
rect 16795 -14900 16840 -14780
rect 16960 -14900 17015 -14780
rect 17135 -14900 17180 -14780
rect 17300 -14900 17345 -14780
rect 17465 -14900 17510 -14780
rect 17630 -14900 17685 -14780
rect 17805 -14900 17850 -14780
rect 17970 -14900 18015 -14780
rect 18135 -14900 18180 -14780
rect 18300 -14900 18310 -14780
rect 12810 -14945 18310 -14900
rect 12810 -15065 12820 -14945
rect 12940 -15065 12995 -14945
rect 13115 -15065 13160 -14945
rect 13280 -15065 13325 -14945
rect 13445 -15065 13490 -14945
rect 13610 -15065 13665 -14945
rect 13785 -15065 13830 -14945
rect 13950 -15065 13995 -14945
rect 14115 -15065 14160 -14945
rect 14280 -15065 14335 -14945
rect 14455 -15065 14500 -14945
rect 14620 -15065 14665 -14945
rect 14785 -15065 14830 -14945
rect 14950 -15065 15005 -14945
rect 15125 -15065 15170 -14945
rect 15290 -15065 15335 -14945
rect 15455 -15065 15500 -14945
rect 15620 -15065 15675 -14945
rect 15795 -15065 15840 -14945
rect 15960 -15065 16005 -14945
rect 16125 -15065 16170 -14945
rect 16290 -15065 16345 -14945
rect 16465 -15065 16510 -14945
rect 16630 -15065 16675 -14945
rect 16795 -15065 16840 -14945
rect 16960 -15065 17015 -14945
rect 17135 -15065 17180 -14945
rect 17300 -15065 17345 -14945
rect 17465 -15065 17510 -14945
rect 17630 -15065 17685 -14945
rect 17805 -15065 17850 -14945
rect 17970 -15065 18015 -14945
rect 18135 -15065 18180 -14945
rect 18300 -15065 18310 -14945
rect 12810 -15110 18310 -15065
rect 12810 -15230 12820 -15110
rect 12940 -15230 12995 -15110
rect 13115 -15230 13160 -15110
rect 13280 -15230 13325 -15110
rect 13445 -15230 13490 -15110
rect 13610 -15230 13665 -15110
rect 13785 -15230 13830 -15110
rect 13950 -15230 13995 -15110
rect 14115 -15230 14160 -15110
rect 14280 -15230 14335 -15110
rect 14455 -15230 14500 -15110
rect 14620 -15230 14665 -15110
rect 14785 -15230 14830 -15110
rect 14950 -15230 15005 -15110
rect 15125 -15230 15170 -15110
rect 15290 -15230 15335 -15110
rect 15455 -15230 15500 -15110
rect 15620 -15230 15675 -15110
rect 15795 -15230 15840 -15110
rect 15960 -15230 16005 -15110
rect 16125 -15230 16170 -15110
rect 16290 -15230 16345 -15110
rect 16465 -15230 16510 -15110
rect 16630 -15230 16675 -15110
rect 16795 -15230 16840 -15110
rect 16960 -15230 17015 -15110
rect 17135 -15230 17180 -15110
rect 17300 -15230 17345 -15110
rect 17465 -15230 17510 -15110
rect 17630 -15230 17685 -15110
rect 17805 -15230 17850 -15110
rect 17970 -15230 18015 -15110
rect 18135 -15230 18180 -15110
rect 18300 -15230 18310 -15110
rect 12810 -15275 18310 -15230
rect 12810 -15395 12820 -15275
rect 12940 -15395 12995 -15275
rect 13115 -15395 13160 -15275
rect 13280 -15395 13325 -15275
rect 13445 -15395 13490 -15275
rect 13610 -15395 13665 -15275
rect 13785 -15395 13830 -15275
rect 13950 -15395 13995 -15275
rect 14115 -15395 14160 -15275
rect 14280 -15395 14335 -15275
rect 14455 -15395 14500 -15275
rect 14620 -15395 14665 -15275
rect 14785 -15395 14830 -15275
rect 14950 -15395 15005 -15275
rect 15125 -15395 15170 -15275
rect 15290 -15395 15335 -15275
rect 15455 -15395 15500 -15275
rect 15620 -15395 15675 -15275
rect 15795 -15395 15840 -15275
rect 15960 -15395 16005 -15275
rect 16125 -15395 16170 -15275
rect 16290 -15395 16345 -15275
rect 16465 -15395 16510 -15275
rect 16630 -15395 16675 -15275
rect 16795 -15395 16840 -15275
rect 16960 -15395 17015 -15275
rect 17135 -15395 17180 -15275
rect 17300 -15395 17345 -15275
rect 17465 -15395 17510 -15275
rect 17630 -15395 17685 -15275
rect 17805 -15395 17850 -15275
rect 17970 -15395 18015 -15275
rect 18135 -15395 18180 -15275
rect 18300 -15395 18310 -15275
rect 12810 -15450 18310 -15395
rect 12810 -15570 12820 -15450
rect 12940 -15570 12995 -15450
rect 13115 -15570 13160 -15450
rect 13280 -15570 13325 -15450
rect 13445 -15570 13490 -15450
rect 13610 -15570 13665 -15450
rect 13785 -15570 13830 -15450
rect 13950 -15570 13995 -15450
rect 14115 -15570 14160 -15450
rect 14280 -15570 14335 -15450
rect 14455 -15570 14500 -15450
rect 14620 -15570 14665 -15450
rect 14785 -15570 14830 -15450
rect 14950 -15570 15005 -15450
rect 15125 -15570 15170 -15450
rect 15290 -15570 15335 -15450
rect 15455 -15570 15500 -15450
rect 15620 -15570 15675 -15450
rect 15795 -15570 15840 -15450
rect 15960 -15570 16005 -15450
rect 16125 -15570 16170 -15450
rect 16290 -15570 16345 -15450
rect 16465 -15570 16510 -15450
rect 16630 -15570 16675 -15450
rect 16795 -15570 16840 -15450
rect 16960 -15570 17015 -15450
rect 17135 -15570 17180 -15450
rect 17300 -15570 17345 -15450
rect 17465 -15570 17510 -15450
rect 17630 -15570 17685 -15450
rect 17805 -15570 17850 -15450
rect 17970 -15570 18015 -15450
rect 18135 -15570 18180 -15450
rect 18300 -15570 18310 -15450
rect 12810 -15580 18310 -15570
rect 18500 -10090 24000 -10080
rect 18500 -10210 18510 -10090
rect 18630 -10210 18685 -10090
rect 18805 -10210 18850 -10090
rect 18970 -10210 19015 -10090
rect 19135 -10210 19180 -10090
rect 19300 -10210 19355 -10090
rect 19475 -10210 19520 -10090
rect 19640 -10210 19685 -10090
rect 19805 -10210 19850 -10090
rect 19970 -10210 20025 -10090
rect 20145 -10210 20190 -10090
rect 20310 -10210 20355 -10090
rect 20475 -10210 20520 -10090
rect 20640 -10210 20695 -10090
rect 20815 -10210 20860 -10090
rect 20980 -10210 21025 -10090
rect 21145 -10210 21190 -10090
rect 21310 -10210 21365 -10090
rect 21485 -10210 21530 -10090
rect 21650 -10210 21695 -10090
rect 21815 -10210 21860 -10090
rect 21980 -10210 22035 -10090
rect 22155 -10210 22200 -10090
rect 22320 -10210 22365 -10090
rect 22485 -10210 22530 -10090
rect 22650 -10210 22705 -10090
rect 22825 -10210 22870 -10090
rect 22990 -10210 23035 -10090
rect 23155 -10210 23200 -10090
rect 23320 -10210 23375 -10090
rect 23495 -10210 23540 -10090
rect 23660 -10210 23705 -10090
rect 23825 -10210 23870 -10090
rect 23990 -10210 24000 -10090
rect 18500 -10255 24000 -10210
rect 18500 -10375 18510 -10255
rect 18630 -10375 18685 -10255
rect 18805 -10375 18850 -10255
rect 18970 -10375 19015 -10255
rect 19135 -10375 19180 -10255
rect 19300 -10375 19355 -10255
rect 19475 -10375 19520 -10255
rect 19640 -10375 19685 -10255
rect 19805 -10375 19850 -10255
rect 19970 -10375 20025 -10255
rect 20145 -10375 20190 -10255
rect 20310 -10375 20355 -10255
rect 20475 -10375 20520 -10255
rect 20640 -10375 20695 -10255
rect 20815 -10375 20860 -10255
rect 20980 -10375 21025 -10255
rect 21145 -10375 21190 -10255
rect 21310 -10375 21365 -10255
rect 21485 -10375 21530 -10255
rect 21650 -10375 21695 -10255
rect 21815 -10375 21860 -10255
rect 21980 -10375 22035 -10255
rect 22155 -10375 22200 -10255
rect 22320 -10375 22365 -10255
rect 22485 -10375 22530 -10255
rect 22650 -10375 22705 -10255
rect 22825 -10375 22870 -10255
rect 22990 -10375 23035 -10255
rect 23155 -10375 23200 -10255
rect 23320 -10375 23375 -10255
rect 23495 -10375 23540 -10255
rect 23660 -10375 23705 -10255
rect 23825 -10375 23870 -10255
rect 23990 -10375 24000 -10255
rect 18500 -10420 24000 -10375
rect 18500 -10540 18510 -10420
rect 18630 -10540 18685 -10420
rect 18805 -10540 18850 -10420
rect 18970 -10540 19015 -10420
rect 19135 -10540 19180 -10420
rect 19300 -10540 19355 -10420
rect 19475 -10540 19520 -10420
rect 19640 -10540 19685 -10420
rect 19805 -10540 19850 -10420
rect 19970 -10540 20025 -10420
rect 20145 -10540 20190 -10420
rect 20310 -10540 20355 -10420
rect 20475 -10540 20520 -10420
rect 20640 -10540 20695 -10420
rect 20815 -10540 20860 -10420
rect 20980 -10540 21025 -10420
rect 21145 -10540 21190 -10420
rect 21310 -10540 21365 -10420
rect 21485 -10540 21530 -10420
rect 21650 -10540 21695 -10420
rect 21815 -10540 21860 -10420
rect 21980 -10540 22035 -10420
rect 22155 -10540 22200 -10420
rect 22320 -10540 22365 -10420
rect 22485 -10540 22530 -10420
rect 22650 -10540 22705 -10420
rect 22825 -10540 22870 -10420
rect 22990 -10540 23035 -10420
rect 23155 -10540 23200 -10420
rect 23320 -10540 23375 -10420
rect 23495 -10540 23540 -10420
rect 23660 -10540 23705 -10420
rect 23825 -10540 23870 -10420
rect 23990 -10540 24000 -10420
rect 18500 -10585 24000 -10540
rect 18500 -10705 18510 -10585
rect 18630 -10705 18685 -10585
rect 18805 -10705 18850 -10585
rect 18970 -10705 19015 -10585
rect 19135 -10705 19180 -10585
rect 19300 -10705 19355 -10585
rect 19475 -10705 19520 -10585
rect 19640 -10705 19685 -10585
rect 19805 -10705 19850 -10585
rect 19970 -10705 20025 -10585
rect 20145 -10705 20190 -10585
rect 20310 -10705 20355 -10585
rect 20475 -10705 20520 -10585
rect 20640 -10705 20695 -10585
rect 20815 -10705 20860 -10585
rect 20980 -10705 21025 -10585
rect 21145 -10705 21190 -10585
rect 21310 -10705 21365 -10585
rect 21485 -10705 21530 -10585
rect 21650 -10705 21695 -10585
rect 21815 -10705 21860 -10585
rect 21980 -10705 22035 -10585
rect 22155 -10705 22200 -10585
rect 22320 -10705 22365 -10585
rect 22485 -10705 22530 -10585
rect 22650 -10705 22705 -10585
rect 22825 -10705 22870 -10585
rect 22990 -10705 23035 -10585
rect 23155 -10705 23200 -10585
rect 23320 -10705 23375 -10585
rect 23495 -10705 23540 -10585
rect 23660 -10705 23705 -10585
rect 23825 -10705 23870 -10585
rect 23990 -10705 24000 -10585
rect 18500 -10760 24000 -10705
rect 18500 -10880 18510 -10760
rect 18630 -10880 18685 -10760
rect 18805 -10880 18850 -10760
rect 18970 -10880 19015 -10760
rect 19135 -10880 19180 -10760
rect 19300 -10880 19355 -10760
rect 19475 -10880 19520 -10760
rect 19640 -10880 19685 -10760
rect 19805 -10880 19850 -10760
rect 19970 -10880 20025 -10760
rect 20145 -10880 20190 -10760
rect 20310 -10880 20355 -10760
rect 20475 -10880 20520 -10760
rect 20640 -10880 20695 -10760
rect 20815 -10880 20860 -10760
rect 20980 -10880 21025 -10760
rect 21145 -10880 21190 -10760
rect 21310 -10880 21365 -10760
rect 21485 -10880 21530 -10760
rect 21650 -10880 21695 -10760
rect 21815 -10880 21860 -10760
rect 21980 -10880 22035 -10760
rect 22155 -10880 22200 -10760
rect 22320 -10880 22365 -10760
rect 22485 -10880 22530 -10760
rect 22650 -10880 22705 -10760
rect 22825 -10880 22870 -10760
rect 22990 -10880 23035 -10760
rect 23155 -10880 23200 -10760
rect 23320 -10880 23375 -10760
rect 23495 -10880 23540 -10760
rect 23660 -10880 23705 -10760
rect 23825 -10880 23870 -10760
rect 23990 -10880 24000 -10760
rect 18500 -10925 24000 -10880
rect 18500 -11045 18510 -10925
rect 18630 -11045 18685 -10925
rect 18805 -11045 18850 -10925
rect 18970 -11045 19015 -10925
rect 19135 -11045 19180 -10925
rect 19300 -11045 19355 -10925
rect 19475 -11045 19520 -10925
rect 19640 -11045 19685 -10925
rect 19805 -11045 19850 -10925
rect 19970 -11045 20025 -10925
rect 20145 -11045 20190 -10925
rect 20310 -11045 20355 -10925
rect 20475 -11045 20520 -10925
rect 20640 -11045 20695 -10925
rect 20815 -11045 20860 -10925
rect 20980 -11045 21025 -10925
rect 21145 -11045 21190 -10925
rect 21310 -11045 21365 -10925
rect 21485 -11045 21530 -10925
rect 21650 -11045 21695 -10925
rect 21815 -11045 21860 -10925
rect 21980 -11045 22035 -10925
rect 22155 -11045 22200 -10925
rect 22320 -11045 22365 -10925
rect 22485 -11045 22530 -10925
rect 22650 -11045 22705 -10925
rect 22825 -11045 22870 -10925
rect 22990 -11045 23035 -10925
rect 23155 -11045 23200 -10925
rect 23320 -11045 23375 -10925
rect 23495 -11045 23540 -10925
rect 23660 -11045 23705 -10925
rect 23825 -11045 23870 -10925
rect 23990 -11045 24000 -10925
rect 18500 -11090 24000 -11045
rect 18500 -11210 18510 -11090
rect 18630 -11210 18685 -11090
rect 18805 -11210 18850 -11090
rect 18970 -11210 19015 -11090
rect 19135 -11210 19180 -11090
rect 19300 -11210 19355 -11090
rect 19475 -11210 19520 -11090
rect 19640 -11210 19685 -11090
rect 19805 -11210 19850 -11090
rect 19970 -11210 20025 -11090
rect 20145 -11210 20190 -11090
rect 20310 -11210 20355 -11090
rect 20475 -11210 20520 -11090
rect 20640 -11210 20695 -11090
rect 20815 -11210 20860 -11090
rect 20980 -11210 21025 -11090
rect 21145 -11210 21190 -11090
rect 21310 -11210 21365 -11090
rect 21485 -11210 21530 -11090
rect 21650 -11210 21695 -11090
rect 21815 -11210 21860 -11090
rect 21980 -11210 22035 -11090
rect 22155 -11210 22200 -11090
rect 22320 -11210 22365 -11090
rect 22485 -11210 22530 -11090
rect 22650 -11210 22705 -11090
rect 22825 -11210 22870 -11090
rect 22990 -11210 23035 -11090
rect 23155 -11210 23200 -11090
rect 23320 -11210 23375 -11090
rect 23495 -11210 23540 -11090
rect 23660 -11210 23705 -11090
rect 23825 -11210 23870 -11090
rect 23990 -11210 24000 -11090
rect 18500 -11255 24000 -11210
rect 18500 -11375 18510 -11255
rect 18630 -11375 18685 -11255
rect 18805 -11375 18850 -11255
rect 18970 -11375 19015 -11255
rect 19135 -11375 19180 -11255
rect 19300 -11375 19355 -11255
rect 19475 -11375 19520 -11255
rect 19640 -11375 19685 -11255
rect 19805 -11375 19850 -11255
rect 19970 -11375 20025 -11255
rect 20145 -11375 20190 -11255
rect 20310 -11375 20355 -11255
rect 20475 -11375 20520 -11255
rect 20640 -11375 20695 -11255
rect 20815 -11375 20860 -11255
rect 20980 -11375 21025 -11255
rect 21145 -11375 21190 -11255
rect 21310 -11375 21365 -11255
rect 21485 -11375 21530 -11255
rect 21650 -11375 21695 -11255
rect 21815 -11375 21860 -11255
rect 21980 -11375 22035 -11255
rect 22155 -11375 22200 -11255
rect 22320 -11375 22365 -11255
rect 22485 -11375 22530 -11255
rect 22650 -11375 22705 -11255
rect 22825 -11375 22870 -11255
rect 22990 -11375 23035 -11255
rect 23155 -11375 23200 -11255
rect 23320 -11375 23375 -11255
rect 23495 -11375 23540 -11255
rect 23660 -11375 23705 -11255
rect 23825 -11375 23870 -11255
rect 23990 -11375 24000 -11255
rect 18500 -11430 24000 -11375
rect 18500 -11550 18510 -11430
rect 18630 -11550 18685 -11430
rect 18805 -11550 18850 -11430
rect 18970 -11550 19015 -11430
rect 19135 -11550 19180 -11430
rect 19300 -11550 19355 -11430
rect 19475 -11550 19520 -11430
rect 19640 -11550 19685 -11430
rect 19805 -11550 19850 -11430
rect 19970 -11550 20025 -11430
rect 20145 -11550 20190 -11430
rect 20310 -11550 20355 -11430
rect 20475 -11550 20520 -11430
rect 20640 -11550 20695 -11430
rect 20815 -11550 20860 -11430
rect 20980 -11550 21025 -11430
rect 21145 -11550 21190 -11430
rect 21310 -11550 21365 -11430
rect 21485 -11550 21530 -11430
rect 21650 -11550 21695 -11430
rect 21815 -11550 21860 -11430
rect 21980 -11550 22035 -11430
rect 22155 -11550 22200 -11430
rect 22320 -11550 22365 -11430
rect 22485 -11550 22530 -11430
rect 22650 -11550 22705 -11430
rect 22825 -11550 22870 -11430
rect 22990 -11550 23035 -11430
rect 23155 -11550 23200 -11430
rect 23320 -11550 23375 -11430
rect 23495 -11550 23540 -11430
rect 23660 -11550 23705 -11430
rect 23825 -11550 23870 -11430
rect 23990 -11550 24000 -11430
rect 18500 -11595 24000 -11550
rect 18500 -11715 18510 -11595
rect 18630 -11715 18685 -11595
rect 18805 -11715 18850 -11595
rect 18970 -11715 19015 -11595
rect 19135 -11715 19180 -11595
rect 19300 -11715 19355 -11595
rect 19475 -11715 19520 -11595
rect 19640 -11715 19685 -11595
rect 19805 -11715 19850 -11595
rect 19970 -11715 20025 -11595
rect 20145 -11715 20190 -11595
rect 20310 -11715 20355 -11595
rect 20475 -11715 20520 -11595
rect 20640 -11715 20695 -11595
rect 20815 -11715 20860 -11595
rect 20980 -11715 21025 -11595
rect 21145 -11715 21190 -11595
rect 21310 -11715 21365 -11595
rect 21485 -11715 21530 -11595
rect 21650 -11715 21695 -11595
rect 21815 -11715 21860 -11595
rect 21980 -11715 22035 -11595
rect 22155 -11715 22200 -11595
rect 22320 -11715 22365 -11595
rect 22485 -11715 22530 -11595
rect 22650 -11715 22705 -11595
rect 22825 -11715 22870 -11595
rect 22990 -11715 23035 -11595
rect 23155 -11715 23200 -11595
rect 23320 -11715 23375 -11595
rect 23495 -11715 23540 -11595
rect 23660 -11715 23705 -11595
rect 23825 -11715 23870 -11595
rect 23990 -11715 24000 -11595
rect 18500 -11760 24000 -11715
rect 18500 -11880 18510 -11760
rect 18630 -11880 18685 -11760
rect 18805 -11880 18850 -11760
rect 18970 -11880 19015 -11760
rect 19135 -11880 19180 -11760
rect 19300 -11880 19355 -11760
rect 19475 -11880 19520 -11760
rect 19640 -11880 19685 -11760
rect 19805 -11880 19850 -11760
rect 19970 -11880 20025 -11760
rect 20145 -11880 20190 -11760
rect 20310 -11880 20355 -11760
rect 20475 -11880 20520 -11760
rect 20640 -11880 20695 -11760
rect 20815 -11880 20860 -11760
rect 20980 -11880 21025 -11760
rect 21145 -11880 21190 -11760
rect 21310 -11880 21365 -11760
rect 21485 -11880 21530 -11760
rect 21650 -11880 21695 -11760
rect 21815 -11880 21860 -11760
rect 21980 -11880 22035 -11760
rect 22155 -11880 22200 -11760
rect 22320 -11880 22365 -11760
rect 22485 -11880 22530 -11760
rect 22650 -11880 22705 -11760
rect 22825 -11880 22870 -11760
rect 22990 -11880 23035 -11760
rect 23155 -11880 23200 -11760
rect 23320 -11880 23375 -11760
rect 23495 -11880 23540 -11760
rect 23660 -11880 23705 -11760
rect 23825 -11880 23870 -11760
rect 23990 -11880 24000 -11760
rect 18500 -11925 24000 -11880
rect 18500 -12045 18510 -11925
rect 18630 -12045 18685 -11925
rect 18805 -12045 18850 -11925
rect 18970 -12045 19015 -11925
rect 19135 -12045 19180 -11925
rect 19300 -12045 19355 -11925
rect 19475 -12045 19520 -11925
rect 19640 -12045 19685 -11925
rect 19805 -12045 19850 -11925
rect 19970 -12045 20025 -11925
rect 20145 -12045 20190 -11925
rect 20310 -12045 20355 -11925
rect 20475 -12045 20520 -11925
rect 20640 -12045 20695 -11925
rect 20815 -12045 20860 -11925
rect 20980 -12045 21025 -11925
rect 21145 -12045 21190 -11925
rect 21310 -12045 21365 -11925
rect 21485 -12045 21530 -11925
rect 21650 -12045 21695 -11925
rect 21815 -12045 21860 -11925
rect 21980 -12045 22035 -11925
rect 22155 -12045 22200 -11925
rect 22320 -12045 22365 -11925
rect 22485 -12045 22530 -11925
rect 22650 -12045 22705 -11925
rect 22825 -12045 22870 -11925
rect 22990 -12045 23035 -11925
rect 23155 -12045 23200 -11925
rect 23320 -12045 23375 -11925
rect 23495 -12045 23540 -11925
rect 23660 -12045 23705 -11925
rect 23825 -12045 23870 -11925
rect 23990 -12045 24000 -11925
rect 18500 -12100 24000 -12045
rect 18500 -12220 18510 -12100
rect 18630 -12220 18685 -12100
rect 18805 -12220 18850 -12100
rect 18970 -12220 19015 -12100
rect 19135 -12220 19180 -12100
rect 19300 -12220 19355 -12100
rect 19475 -12220 19520 -12100
rect 19640 -12220 19685 -12100
rect 19805 -12220 19850 -12100
rect 19970 -12220 20025 -12100
rect 20145 -12220 20190 -12100
rect 20310 -12220 20355 -12100
rect 20475 -12220 20520 -12100
rect 20640 -12220 20695 -12100
rect 20815 -12220 20860 -12100
rect 20980 -12220 21025 -12100
rect 21145 -12220 21190 -12100
rect 21310 -12220 21365 -12100
rect 21485 -12220 21530 -12100
rect 21650 -12220 21695 -12100
rect 21815 -12220 21860 -12100
rect 21980 -12220 22035 -12100
rect 22155 -12220 22200 -12100
rect 22320 -12220 22365 -12100
rect 22485 -12220 22530 -12100
rect 22650 -12220 22705 -12100
rect 22825 -12220 22870 -12100
rect 22990 -12220 23035 -12100
rect 23155 -12220 23200 -12100
rect 23320 -12220 23375 -12100
rect 23495 -12220 23540 -12100
rect 23660 -12220 23705 -12100
rect 23825 -12220 23870 -12100
rect 23990 -12220 24000 -12100
rect 18500 -12265 24000 -12220
rect 18500 -12385 18510 -12265
rect 18630 -12385 18685 -12265
rect 18805 -12385 18850 -12265
rect 18970 -12385 19015 -12265
rect 19135 -12385 19180 -12265
rect 19300 -12385 19355 -12265
rect 19475 -12385 19520 -12265
rect 19640 -12385 19685 -12265
rect 19805 -12385 19850 -12265
rect 19970 -12385 20025 -12265
rect 20145 -12385 20190 -12265
rect 20310 -12385 20355 -12265
rect 20475 -12385 20520 -12265
rect 20640 -12385 20695 -12265
rect 20815 -12385 20860 -12265
rect 20980 -12385 21025 -12265
rect 21145 -12385 21190 -12265
rect 21310 -12385 21365 -12265
rect 21485 -12385 21530 -12265
rect 21650 -12385 21695 -12265
rect 21815 -12385 21860 -12265
rect 21980 -12385 22035 -12265
rect 22155 -12385 22200 -12265
rect 22320 -12385 22365 -12265
rect 22485 -12385 22530 -12265
rect 22650 -12385 22705 -12265
rect 22825 -12385 22870 -12265
rect 22990 -12385 23035 -12265
rect 23155 -12385 23200 -12265
rect 23320 -12385 23375 -12265
rect 23495 -12385 23540 -12265
rect 23660 -12385 23705 -12265
rect 23825 -12385 23870 -12265
rect 23990 -12385 24000 -12265
rect 18500 -12430 24000 -12385
rect 18500 -12550 18510 -12430
rect 18630 -12550 18685 -12430
rect 18805 -12550 18850 -12430
rect 18970 -12550 19015 -12430
rect 19135 -12550 19180 -12430
rect 19300 -12550 19355 -12430
rect 19475 -12550 19520 -12430
rect 19640 -12550 19685 -12430
rect 19805 -12550 19850 -12430
rect 19970 -12550 20025 -12430
rect 20145 -12550 20190 -12430
rect 20310 -12550 20355 -12430
rect 20475 -12550 20520 -12430
rect 20640 -12550 20695 -12430
rect 20815 -12550 20860 -12430
rect 20980 -12550 21025 -12430
rect 21145 -12550 21190 -12430
rect 21310 -12550 21365 -12430
rect 21485 -12550 21530 -12430
rect 21650 -12550 21695 -12430
rect 21815 -12550 21860 -12430
rect 21980 -12550 22035 -12430
rect 22155 -12550 22200 -12430
rect 22320 -12550 22365 -12430
rect 22485 -12550 22530 -12430
rect 22650 -12550 22705 -12430
rect 22825 -12550 22870 -12430
rect 22990 -12550 23035 -12430
rect 23155 -12550 23200 -12430
rect 23320 -12550 23375 -12430
rect 23495 -12550 23540 -12430
rect 23660 -12550 23705 -12430
rect 23825 -12550 23870 -12430
rect 23990 -12550 24000 -12430
rect 18500 -12595 24000 -12550
rect 18500 -12715 18510 -12595
rect 18630 -12715 18685 -12595
rect 18805 -12715 18850 -12595
rect 18970 -12715 19015 -12595
rect 19135 -12715 19180 -12595
rect 19300 -12715 19355 -12595
rect 19475 -12715 19520 -12595
rect 19640 -12715 19685 -12595
rect 19805 -12715 19850 -12595
rect 19970 -12715 20025 -12595
rect 20145 -12715 20190 -12595
rect 20310 -12715 20355 -12595
rect 20475 -12715 20520 -12595
rect 20640 -12715 20695 -12595
rect 20815 -12715 20860 -12595
rect 20980 -12715 21025 -12595
rect 21145 -12715 21190 -12595
rect 21310 -12715 21365 -12595
rect 21485 -12715 21530 -12595
rect 21650 -12715 21695 -12595
rect 21815 -12715 21860 -12595
rect 21980 -12715 22035 -12595
rect 22155 -12715 22200 -12595
rect 22320 -12715 22365 -12595
rect 22485 -12715 22530 -12595
rect 22650 -12715 22705 -12595
rect 22825 -12715 22870 -12595
rect 22990 -12715 23035 -12595
rect 23155 -12715 23200 -12595
rect 23320 -12715 23375 -12595
rect 23495 -12715 23540 -12595
rect 23660 -12715 23705 -12595
rect 23825 -12715 23870 -12595
rect 23990 -12715 24000 -12595
rect 18500 -12770 24000 -12715
rect 18500 -12890 18510 -12770
rect 18630 -12890 18685 -12770
rect 18805 -12890 18850 -12770
rect 18970 -12890 19015 -12770
rect 19135 -12890 19180 -12770
rect 19300 -12890 19355 -12770
rect 19475 -12890 19520 -12770
rect 19640 -12890 19685 -12770
rect 19805 -12890 19850 -12770
rect 19970 -12890 20025 -12770
rect 20145 -12890 20190 -12770
rect 20310 -12890 20355 -12770
rect 20475 -12890 20520 -12770
rect 20640 -12890 20695 -12770
rect 20815 -12890 20860 -12770
rect 20980 -12890 21025 -12770
rect 21145 -12890 21190 -12770
rect 21310 -12890 21365 -12770
rect 21485 -12890 21530 -12770
rect 21650 -12890 21695 -12770
rect 21815 -12890 21860 -12770
rect 21980 -12890 22035 -12770
rect 22155 -12890 22200 -12770
rect 22320 -12890 22365 -12770
rect 22485 -12890 22530 -12770
rect 22650 -12890 22705 -12770
rect 22825 -12890 22870 -12770
rect 22990 -12890 23035 -12770
rect 23155 -12890 23200 -12770
rect 23320 -12890 23375 -12770
rect 23495 -12890 23540 -12770
rect 23660 -12890 23705 -12770
rect 23825 -12890 23870 -12770
rect 23990 -12890 24000 -12770
rect 18500 -12935 24000 -12890
rect 18500 -13055 18510 -12935
rect 18630 -13055 18685 -12935
rect 18805 -13055 18850 -12935
rect 18970 -13055 19015 -12935
rect 19135 -13055 19180 -12935
rect 19300 -13055 19355 -12935
rect 19475 -13055 19520 -12935
rect 19640 -13055 19685 -12935
rect 19805 -13055 19850 -12935
rect 19970 -13055 20025 -12935
rect 20145 -13055 20190 -12935
rect 20310 -13055 20355 -12935
rect 20475 -13055 20520 -12935
rect 20640 -13055 20695 -12935
rect 20815 -13055 20860 -12935
rect 20980 -13055 21025 -12935
rect 21145 -13055 21190 -12935
rect 21310 -13055 21365 -12935
rect 21485 -13055 21530 -12935
rect 21650 -13055 21695 -12935
rect 21815 -13055 21860 -12935
rect 21980 -13055 22035 -12935
rect 22155 -13055 22200 -12935
rect 22320 -13055 22365 -12935
rect 22485 -13055 22530 -12935
rect 22650 -13055 22705 -12935
rect 22825 -13055 22870 -12935
rect 22990 -13055 23035 -12935
rect 23155 -13055 23200 -12935
rect 23320 -13055 23375 -12935
rect 23495 -13055 23540 -12935
rect 23660 -13055 23705 -12935
rect 23825 -13055 23870 -12935
rect 23990 -13055 24000 -12935
rect 18500 -13100 24000 -13055
rect 18500 -13220 18510 -13100
rect 18630 -13220 18685 -13100
rect 18805 -13220 18850 -13100
rect 18970 -13220 19015 -13100
rect 19135 -13220 19180 -13100
rect 19300 -13220 19355 -13100
rect 19475 -13220 19520 -13100
rect 19640 -13220 19685 -13100
rect 19805 -13220 19850 -13100
rect 19970 -13220 20025 -13100
rect 20145 -13220 20190 -13100
rect 20310 -13220 20355 -13100
rect 20475 -13220 20520 -13100
rect 20640 -13220 20695 -13100
rect 20815 -13220 20860 -13100
rect 20980 -13220 21025 -13100
rect 21145 -13220 21190 -13100
rect 21310 -13220 21365 -13100
rect 21485 -13220 21530 -13100
rect 21650 -13220 21695 -13100
rect 21815 -13220 21860 -13100
rect 21980 -13220 22035 -13100
rect 22155 -13220 22200 -13100
rect 22320 -13220 22365 -13100
rect 22485 -13220 22530 -13100
rect 22650 -13220 22705 -13100
rect 22825 -13220 22870 -13100
rect 22990 -13220 23035 -13100
rect 23155 -13220 23200 -13100
rect 23320 -13220 23375 -13100
rect 23495 -13220 23540 -13100
rect 23660 -13220 23705 -13100
rect 23825 -13220 23870 -13100
rect 23990 -13220 24000 -13100
rect 18500 -13265 24000 -13220
rect 18500 -13385 18510 -13265
rect 18630 -13385 18685 -13265
rect 18805 -13385 18850 -13265
rect 18970 -13385 19015 -13265
rect 19135 -13385 19180 -13265
rect 19300 -13385 19355 -13265
rect 19475 -13385 19520 -13265
rect 19640 -13385 19685 -13265
rect 19805 -13385 19850 -13265
rect 19970 -13385 20025 -13265
rect 20145 -13385 20190 -13265
rect 20310 -13385 20355 -13265
rect 20475 -13385 20520 -13265
rect 20640 -13385 20695 -13265
rect 20815 -13385 20860 -13265
rect 20980 -13385 21025 -13265
rect 21145 -13385 21190 -13265
rect 21310 -13385 21365 -13265
rect 21485 -13385 21530 -13265
rect 21650 -13385 21695 -13265
rect 21815 -13385 21860 -13265
rect 21980 -13385 22035 -13265
rect 22155 -13385 22200 -13265
rect 22320 -13385 22365 -13265
rect 22485 -13385 22530 -13265
rect 22650 -13385 22705 -13265
rect 22825 -13385 22870 -13265
rect 22990 -13385 23035 -13265
rect 23155 -13385 23200 -13265
rect 23320 -13385 23375 -13265
rect 23495 -13385 23540 -13265
rect 23660 -13385 23705 -13265
rect 23825 -13385 23870 -13265
rect 23990 -13385 24000 -13265
rect 18500 -13440 24000 -13385
rect 18500 -13560 18510 -13440
rect 18630 -13560 18685 -13440
rect 18805 -13560 18850 -13440
rect 18970 -13560 19015 -13440
rect 19135 -13560 19180 -13440
rect 19300 -13560 19355 -13440
rect 19475 -13560 19520 -13440
rect 19640 -13560 19685 -13440
rect 19805 -13560 19850 -13440
rect 19970 -13560 20025 -13440
rect 20145 -13560 20190 -13440
rect 20310 -13560 20355 -13440
rect 20475 -13560 20520 -13440
rect 20640 -13560 20695 -13440
rect 20815 -13560 20860 -13440
rect 20980 -13560 21025 -13440
rect 21145 -13560 21190 -13440
rect 21310 -13560 21365 -13440
rect 21485 -13560 21530 -13440
rect 21650 -13560 21695 -13440
rect 21815 -13560 21860 -13440
rect 21980 -13560 22035 -13440
rect 22155 -13560 22200 -13440
rect 22320 -13560 22365 -13440
rect 22485 -13560 22530 -13440
rect 22650 -13560 22705 -13440
rect 22825 -13560 22870 -13440
rect 22990 -13560 23035 -13440
rect 23155 -13560 23200 -13440
rect 23320 -13560 23375 -13440
rect 23495 -13560 23540 -13440
rect 23660 -13560 23705 -13440
rect 23825 -13560 23870 -13440
rect 23990 -13560 24000 -13440
rect 18500 -13605 24000 -13560
rect 18500 -13725 18510 -13605
rect 18630 -13725 18685 -13605
rect 18805 -13725 18850 -13605
rect 18970 -13725 19015 -13605
rect 19135 -13725 19180 -13605
rect 19300 -13725 19355 -13605
rect 19475 -13725 19520 -13605
rect 19640 -13725 19685 -13605
rect 19805 -13725 19850 -13605
rect 19970 -13725 20025 -13605
rect 20145 -13725 20190 -13605
rect 20310 -13725 20355 -13605
rect 20475 -13725 20520 -13605
rect 20640 -13725 20695 -13605
rect 20815 -13725 20860 -13605
rect 20980 -13725 21025 -13605
rect 21145 -13725 21190 -13605
rect 21310 -13725 21365 -13605
rect 21485 -13725 21530 -13605
rect 21650 -13725 21695 -13605
rect 21815 -13725 21860 -13605
rect 21980 -13725 22035 -13605
rect 22155 -13725 22200 -13605
rect 22320 -13725 22365 -13605
rect 22485 -13725 22530 -13605
rect 22650 -13725 22705 -13605
rect 22825 -13725 22870 -13605
rect 22990 -13725 23035 -13605
rect 23155 -13725 23200 -13605
rect 23320 -13725 23375 -13605
rect 23495 -13725 23540 -13605
rect 23660 -13725 23705 -13605
rect 23825 -13725 23870 -13605
rect 23990 -13725 24000 -13605
rect 18500 -13770 24000 -13725
rect 18500 -13890 18510 -13770
rect 18630 -13890 18685 -13770
rect 18805 -13890 18850 -13770
rect 18970 -13890 19015 -13770
rect 19135 -13890 19180 -13770
rect 19300 -13890 19355 -13770
rect 19475 -13890 19520 -13770
rect 19640 -13890 19685 -13770
rect 19805 -13890 19850 -13770
rect 19970 -13890 20025 -13770
rect 20145 -13890 20190 -13770
rect 20310 -13890 20355 -13770
rect 20475 -13890 20520 -13770
rect 20640 -13890 20695 -13770
rect 20815 -13890 20860 -13770
rect 20980 -13890 21025 -13770
rect 21145 -13890 21190 -13770
rect 21310 -13890 21365 -13770
rect 21485 -13890 21530 -13770
rect 21650 -13890 21695 -13770
rect 21815 -13890 21860 -13770
rect 21980 -13890 22035 -13770
rect 22155 -13890 22200 -13770
rect 22320 -13890 22365 -13770
rect 22485 -13890 22530 -13770
rect 22650 -13890 22705 -13770
rect 22825 -13890 22870 -13770
rect 22990 -13890 23035 -13770
rect 23155 -13890 23200 -13770
rect 23320 -13890 23375 -13770
rect 23495 -13890 23540 -13770
rect 23660 -13890 23705 -13770
rect 23825 -13890 23870 -13770
rect 23990 -13890 24000 -13770
rect 18500 -13935 24000 -13890
rect 18500 -14055 18510 -13935
rect 18630 -14055 18685 -13935
rect 18805 -14055 18850 -13935
rect 18970 -14055 19015 -13935
rect 19135 -14055 19180 -13935
rect 19300 -14055 19355 -13935
rect 19475 -14055 19520 -13935
rect 19640 -14055 19685 -13935
rect 19805 -14055 19850 -13935
rect 19970 -14055 20025 -13935
rect 20145 -14055 20190 -13935
rect 20310 -14055 20355 -13935
rect 20475 -14055 20520 -13935
rect 20640 -14055 20695 -13935
rect 20815 -14055 20860 -13935
rect 20980 -14055 21025 -13935
rect 21145 -14055 21190 -13935
rect 21310 -14055 21365 -13935
rect 21485 -14055 21530 -13935
rect 21650 -14055 21695 -13935
rect 21815 -14055 21860 -13935
rect 21980 -14055 22035 -13935
rect 22155 -14055 22200 -13935
rect 22320 -14055 22365 -13935
rect 22485 -14055 22530 -13935
rect 22650 -14055 22705 -13935
rect 22825 -14055 22870 -13935
rect 22990 -14055 23035 -13935
rect 23155 -14055 23200 -13935
rect 23320 -14055 23375 -13935
rect 23495 -14055 23540 -13935
rect 23660 -14055 23705 -13935
rect 23825 -14055 23870 -13935
rect 23990 -14055 24000 -13935
rect 18500 -14110 24000 -14055
rect 18500 -14230 18510 -14110
rect 18630 -14230 18685 -14110
rect 18805 -14230 18850 -14110
rect 18970 -14230 19015 -14110
rect 19135 -14230 19180 -14110
rect 19300 -14230 19355 -14110
rect 19475 -14230 19520 -14110
rect 19640 -14230 19685 -14110
rect 19805 -14230 19850 -14110
rect 19970 -14230 20025 -14110
rect 20145 -14230 20190 -14110
rect 20310 -14230 20355 -14110
rect 20475 -14230 20520 -14110
rect 20640 -14230 20695 -14110
rect 20815 -14230 20860 -14110
rect 20980 -14230 21025 -14110
rect 21145 -14230 21190 -14110
rect 21310 -14230 21365 -14110
rect 21485 -14230 21530 -14110
rect 21650 -14230 21695 -14110
rect 21815 -14230 21860 -14110
rect 21980 -14230 22035 -14110
rect 22155 -14230 22200 -14110
rect 22320 -14230 22365 -14110
rect 22485 -14230 22530 -14110
rect 22650 -14230 22705 -14110
rect 22825 -14230 22870 -14110
rect 22990 -14230 23035 -14110
rect 23155 -14230 23200 -14110
rect 23320 -14230 23375 -14110
rect 23495 -14230 23540 -14110
rect 23660 -14230 23705 -14110
rect 23825 -14230 23870 -14110
rect 23990 -14230 24000 -14110
rect 18500 -14275 24000 -14230
rect 18500 -14395 18510 -14275
rect 18630 -14395 18685 -14275
rect 18805 -14395 18850 -14275
rect 18970 -14395 19015 -14275
rect 19135 -14395 19180 -14275
rect 19300 -14395 19355 -14275
rect 19475 -14395 19520 -14275
rect 19640 -14395 19685 -14275
rect 19805 -14395 19850 -14275
rect 19970 -14395 20025 -14275
rect 20145 -14395 20190 -14275
rect 20310 -14395 20355 -14275
rect 20475 -14395 20520 -14275
rect 20640 -14395 20695 -14275
rect 20815 -14395 20860 -14275
rect 20980 -14395 21025 -14275
rect 21145 -14395 21190 -14275
rect 21310 -14395 21365 -14275
rect 21485 -14395 21530 -14275
rect 21650 -14395 21695 -14275
rect 21815 -14395 21860 -14275
rect 21980 -14395 22035 -14275
rect 22155 -14395 22200 -14275
rect 22320 -14395 22365 -14275
rect 22485 -14395 22530 -14275
rect 22650 -14395 22705 -14275
rect 22825 -14395 22870 -14275
rect 22990 -14395 23035 -14275
rect 23155 -14395 23200 -14275
rect 23320 -14395 23375 -14275
rect 23495 -14395 23540 -14275
rect 23660 -14395 23705 -14275
rect 23825 -14395 23870 -14275
rect 23990 -14395 24000 -14275
rect 18500 -14440 24000 -14395
rect 18500 -14560 18510 -14440
rect 18630 -14560 18685 -14440
rect 18805 -14560 18850 -14440
rect 18970 -14560 19015 -14440
rect 19135 -14560 19180 -14440
rect 19300 -14560 19355 -14440
rect 19475 -14560 19520 -14440
rect 19640 -14560 19685 -14440
rect 19805 -14560 19850 -14440
rect 19970 -14560 20025 -14440
rect 20145 -14560 20190 -14440
rect 20310 -14560 20355 -14440
rect 20475 -14560 20520 -14440
rect 20640 -14560 20695 -14440
rect 20815 -14560 20860 -14440
rect 20980 -14560 21025 -14440
rect 21145 -14560 21190 -14440
rect 21310 -14560 21365 -14440
rect 21485 -14560 21530 -14440
rect 21650 -14560 21695 -14440
rect 21815 -14560 21860 -14440
rect 21980 -14560 22035 -14440
rect 22155 -14560 22200 -14440
rect 22320 -14560 22365 -14440
rect 22485 -14560 22530 -14440
rect 22650 -14560 22705 -14440
rect 22825 -14560 22870 -14440
rect 22990 -14560 23035 -14440
rect 23155 -14560 23200 -14440
rect 23320 -14560 23375 -14440
rect 23495 -14560 23540 -14440
rect 23660 -14560 23705 -14440
rect 23825 -14560 23870 -14440
rect 23990 -14560 24000 -14440
rect 18500 -14605 24000 -14560
rect 18500 -14725 18510 -14605
rect 18630 -14725 18685 -14605
rect 18805 -14725 18850 -14605
rect 18970 -14725 19015 -14605
rect 19135 -14725 19180 -14605
rect 19300 -14725 19355 -14605
rect 19475 -14725 19520 -14605
rect 19640 -14725 19685 -14605
rect 19805 -14725 19850 -14605
rect 19970 -14725 20025 -14605
rect 20145 -14725 20190 -14605
rect 20310 -14725 20355 -14605
rect 20475 -14725 20520 -14605
rect 20640 -14725 20695 -14605
rect 20815 -14725 20860 -14605
rect 20980 -14725 21025 -14605
rect 21145 -14725 21190 -14605
rect 21310 -14725 21365 -14605
rect 21485 -14725 21530 -14605
rect 21650 -14725 21695 -14605
rect 21815 -14725 21860 -14605
rect 21980 -14725 22035 -14605
rect 22155 -14725 22200 -14605
rect 22320 -14725 22365 -14605
rect 22485 -14725 22530 -14605
rect 22650 -14725 22705 -14605
rect 22825 -14725 22870 -14605
rect 22990 -14725 23035 -14605
rect 23155 -14725 23200 -14605
rect 23320 -14725 23375 -14605
rect 23495 -14725 23540 -14605
rect 23660 -14725 23705 -14605
rect 23825 -14725 23870 -14605
rect 23990 -14725 24000 -14605
rect 18500 -14780 24000 -14725
rect 18500 -14900 18510 -14780
rect 18630 -14900 18685 -14780
rect 18805 -14900 18850 -14780
rect 18970 -14900 19015 -14780
rect 19135 -14900 19180 -14780
rect 19300 -14900 19355 -14780
rect 19475 -14900 19520 -14780
rect 19640 -14900 19685 -14780
rect 19805 -14900 19850 -14780
rect 19970 -14900 20025 -14780
rect 20145 -14900 20190 -14780
rect 20310 -14900 20355 -14780
rect 20475 -14900 20520 -14780
rect 20640 -14900 20695 -14780
rect 20815 -14900 20860 -14780
rect 20980 -14900 21025 -14780
rect 21145 -14900 21190 -14780
rect 21310 -14900 21365 -14780
rect 21485 -14900 21530 -14780
rect 21650 -14900 21695 -14780
rect 21815 -14900 21860 -14780
rect 21980 -14900 22035 -14780
rect 22155 -14900 22200 -14780
rect 22320 -14900 22365 -14780
rect 22485 -14900 22530 -14780
rect 22650 -14900 22705 -14780
rect 22825 -14900 22870 -14780
rect 22990 -14900 23035 -14780
rect 23155 -14900 23200 -14780
rect 23320 -14900 23375 -14780
rect 23495 -14900 23540 -14780
rect 23660 -14900 23705 -14780
rect 23825 -14900 23870 -14780
rect 23990 -14900 24000 -14780
rect 18500 -14945 24000 -14900
rect 18500 -15065 18510 -14945
rect 18630 -15065 18685 -14945
rect 18805 -15065 18850 -14945
rect 18970 -15065 19015 -14945
rect 19135 -15065 19180 -14945
rect 19300 -15065 19355 -14945
rect 19475 -15065 19520 -14945
rect 19640 -15065 19685 -14945
rect 19805 -15065 19850 -14945
rect 19970 -15065 20025 -14945
rect 20145 -15065 20190 -14945
rect 20310 -15065 20355 -14945
rect 20475 -15065 20520 -14945
rect 20640 -15065 20695 -14945
rect 20815 -15065 20860 -14945
rect 20980 -15065 21025 -14945
rect 21145 -15065 21190 -14945
rect 21310 -15065 21365 -14945
rect 21485 -15065 21530 -14945
rect 21650 -15065 21695 -14945
rect 21815 -15065 21860 -14945
rect 21980 -15065 22035 -14945
rect 22155 -15065 22200 -14945
rect 22320 -15065 22365 -14945
rect 22485 -15065 22530 -14945
rect 22650 -15065 22705 -14945
rect 22825 -15065 22870 -14945
rect 22990 -15065 23035 -14945
rect 23155 -15065 23200 -14945
rect 23320 -15065 23375 -14945
rect 23495 -15065 23540 -14945
rect 23660 -15065 23705 -14945
rect 23825 -15065 23870 -14945
rect 23990 -15065 24000 -14945
rect 18500 -15110 24000 -15065
rect 18500 -15230 18510 -15110
rect 18630 -15230 18685 -15110
rect 18805 -15230 18850 -15110
rect 18970 -15230 19015 -15110
rect 19135 -15230 19180 -15110
rect 19300 -15230 19355 -15110
rect 19475 -15230 19520 -15110
rect 19640 -15230 19685 -15110
rect 19805 -15230 19850 -15110
rect 19970 -15230 20025 -15110
rect 20145 -15230 20190 -15110
rect 20310 -15230 20355 -15110
rect 20475 -15230 20520 -15110
rect 20640 -15230 20695 -15110
rect 20815 -15230 20860 -15110
rect 20980 -15230 21025 -15110
rect 21145 -15230 21190 -15110
rect 21310 -15230 21365 -15110
rect 21485 -15230 21530 -15110
rect 21650 -15230 21695 -15110
rect 21815 -15230 21860 -15110
rect 21980 -15230 22035 -15110
rect 22155 -15230 22200 -15110
rect 22320 -15230 22365 -15110
rect 22485 -15230 22530 -15110
rect 22650 -15230 22705 -15110
rect 22825 -15230 22870 -15110
rect 22990 -15230 23035 -15110
rect 23155 -15230 23200 -15110
rect 23320 -15230 23375 -15110
rect 23495 -15230 23540 -15110
rect 23660 -15230 23705 -15110
rect 23825 -15230 23870 -15110
rect 23990 -15230 24000 -15110
rect 18500 -15275 24000 -15230
rect 18500 -15395 18510 -15275
rect 18630 -15395 18685 -15275
rect 18805 -15395 18850 -15275
rect 18970 -15395 19015 -15275
rect 19135 -15395 19180 -15275
rect 19300 -15395 19355 -15275
rect 19475 -15395 19520 -15275
rect 19640 -15395 19685 -15275
rect 19805 -15395 19850 -15275
rect 19970 -15395 20025 -15275
rect 20145 -15395 20190 -15275
rect 20310 -15395 20355 -15275
rect 20475 -15395 20520 -15275
rect 20640 -15395 20695 -15275
rect 20815 -15395 20860 -15275
rect 20980 -15395 21025 -15275
rect 21145 -15395 21190 -15275
rect 21310 -15395 21365 -15275
rect 21485 -15395 21530 -15275
rect 21650 -15395 21695 -15275
rect 21815 -15395 21860 -15275
rect 21980 -15395 22035 -15275
rect 22155 -15395 22200 -15275
rect 22320 -15395 22365 -15275
rect 22485 -15395 22530 -15275
rect 22650 -15395 22705 -15275
rect 22825 -15395 22870 -15275
rect 22990 -15395 23035 -15275
rect 23155 -15395 23200 -15275
rect 23320 -15395 23375 -15275
rect 23495 -15395 23540 -15275
rect 23660 -15395 23705 -15275
rect 23825 -15395 23870 -15275
rect 23990 -15395 24000 -15275
rect 18500 -15450 24000 -15395
rect 18500 -15570 18510 -15450
rect 18630 -15570 18685 -15450
rect 18805 -15570 18850 -15450
rect 18970 -15570 19015 -15450
rect 19135 -15570 19180 -15450
rect 19300 -15570 19355 -15450
rect 19475 -15570 19520 -15450
rect 19640 -15570 19685 -15450
rect 19805 -15570 19850 -15450
rect 19970 -15570 20025 -15450
rect 20145 -15570 20190 -15450
rect 20310 -15570 20355 -15450
rect 20475 -15570 20520 -15450
rect 20640 -15570 20695 -15450
rect 20815 -15570 20860 -15450
rect 20980 -15570 21025 -15450
rect 21145 -15570 21190 -15450
rect 21310 -15570 21365 -15450
rect 21485 -15570 21530 -15450
rect 21650 -15570 21695 -15450
rect 21815 -15570 21860 -15450
rect 21980 -15570 22035 -15450
rect 22155 -15570 22200 -15450
rect 22320 -15570 22365 -15450
rect 22485 -15570 22530 -15450
rect 22650 -15570 22705 -15450
rect 22825 -15570 22870 -15450
rect 22990 -15570 23035 -15450
rect 23155 -15570 23200 -15450
rect 23320 -15570 23375 -15450
rect 23495 -15570 23540 -15450
rect 23660 -15570 23705 -15450
rect 23825 -15570 23870 -15450
rect 23990 -15570 24000 -15450
rect 18500 -15580 24000 -15570
rect 24190 -10090 29690 -10080
rect 24190 -10210 24200 -10090
rect 24320 -10210 24375 -10090
rect 24495 -10210 24540 -10090
rect 24660 -10210 24705 -10090
rect 24825 -10210 24870 -10090
rect 24990 -10210 25045 -10090
rect 25165 -10210 25210 -10090
rect 25330 -10210 25375 -10090
rect 25495 -10210 25540 -10090
rect 25660 -10210 25715 -10090
rect 25835 -10210 25880 -10090
rect 26000 -10210 26045 -10090
rect 26165 -10210 26210 -10090
rect 26330 -10210 26385 -10090
rect 26505 -10210 26550 -10090
rect 26670 -10210 26715 -10090
rect 26835 -10210 26880 -10090
rect 27000 -10210 27055 -10090
rect 27175 -10210 27220 -10090
rect 27340 -10210 27385 -10090
rect 27505 -10210 27550 -10090
rect 27670 -10210 27725 -10090
rect 27845 -10210 27890 -10090
rect 28010 -10210 28055 -10090
rect 28175 -10210 28220 -10090
rect 28340 -10210 28395 -10090
rect 28515 -10210 28560 -10090
rect 28680 -10210 28725 -10090
rect 28845 -10210 28890 -10090
rect 29010 -10210 29065 -10090
rect 29185 -10210 29230 -10090
rect 29350 -10210 29395 -10090
rect 29515 -10210 29560 -10090
rect 29680 -10210 29690 -10090
rect 24190 -10255 29690 -10210
rect 24190 -10375 24200 -10255
rect 24320 -10375 24375 -10255
rect 24495 -10375 24540 -10255
rect 24660 -10375 24705 -10255
rect 24825 -10375 24870 -10255
rect 24990 -10375 25045 -10255
rect 25165 -10375 25210 -10255
rect 25330 -10375 25375 -10255
rect 25495 -10375 25540 -10255
rect 25660 -10375 25715 -10255
rect 25835 -10375 25880 -10255
rect 26000 -10375 26045 -10255
rect 26165 -10375 26210 -10255
rect 26330 -10375 26385 -10255
rect 26505 -10375 26550 -10255
rect 26670 -10375 26715 -10255
rect 26835 -10375 26880 -10255
rect 27000 -10375 27055 -10255
rect 27175 -10375 27220 -10255
rect 27340 -10375 27385 -10255
rect 27505 -10375 27550 -10255
rect 27670 -10375 27725 -10255
rect 27845 -10375 27890 -10255
rect 28010 -10375 28055 -10255
rect 28175 -10375 28220 -10255
rect 28340 -10375 28395 -10255
rect 28515 -10375 28560 -10255
rect 28680 -10375 28725 -10255
rect 28845 -10375 28890 -10255
rect 29010 -10375 29065 -10255
rect 29185 -10375 29230 -10255
rect 29350 -10375 29395 -10255
rect 29515 -10375 29560 -10255
rect 29680 -10375 29690 -10255
rect 24190 -10420 29690 -10375
rect 24190 -10540 24200 -10420
rect 24320 -10540 24375 -10420
rect 24495 -10540 24540 -10420
rect 24660 -10540 24705 -10420
rect 24825 -10540 24870 -10420
rect 24990 -10540 25045 -10420
rect 25165 -10540 25210 -10420
rect 25330 -10540 25375 -10420
rect 25495 -10540 25540 -10420
rect 25660 -10540 25715 -10420
rect 25835 -10540 25880 -10420
rect 26000 -10540 26045 -10420
rect 26165 -10540 26210 -10420
rect 26330 -10540 26385 -10420
rect 26505 -10540 26550 -10420
rect 26670 -10540 26715 -10420
rect 26835 -10540 26880 -10420
rect 27000 -10540 27055 -10420
rect 27175 -10540 27220 -10420
rect 27340 -10540 27385 -10420
rect 27505 -10540 27550 -10420
rect 27670 -10540 27725 -10420
rect 27845 -10540 27890 -10420
rect 28010 -10540 28055 -10420
rect 28175 -10540 28220 -10420
rect 28340 -10540 28395 -10420
rect 28515 -10540 28560 -10420
rect 28680 -10540 28725 -10420
rect 28845 -10540 28890 -10420
rect 29010 -10540 29065 -10420
rect 29185 -10540 29230 -10420
rect 29350 -10540 29395 -10420
rect 29515 -10540 29560 -10420
rect 29680 -10540 29690 -10420
rect 24190 -10585 29690 -10540
rect 24190 -10705 24200 -10585
rect 24320 -10705 24375 -10585
rect 24495 -10705 24540 -10585
rect 24660 -10705 24705 -10585
rect 24825 -10705 24870 -10585
rect 24990 -10705 25045 -10585
rect 25165 -10705 25210 -10585
rect 25330 -10705 25375 -10585
rect 25495 -10705 25540 -10585
rect 25660 -10705 25715 -10585
rect 25835 -10705 25880 -10585
rect 26000 -10705 26045 -10585
rect 26165 -10705 26210 -10585
rect 26330 -10705 26385 -10585
rect 26505 -10705 26550 -10585
rect 26670 -10705 26715 -10585
rect 26835 -10705 26880 -10585
rect 27000 -10705 27055 -10585
rect 27175 -10705 27220 -10585
rect 27340 -10705 27385 -10585
rect 27505 -10705 27550 -10585
rect 27670 -10705 27725 -10585
rect 27845 -10705 27890 -10585
rect 28010 -10705 28055 -10585
rect 28175 -10705 28220 -10585
rect 28340 -10705 28395 -10585
rect 28515 -10705 28560 -10585
rect 28680 -10705 28725 -10585
rect 28845 -10705 28890 -10585
rect 29010 -10705 29065 -10585
rect 29185 -10705 29230 -10585
rect 29350 -10705 29395 -10585
rect 29515 -10705 29560 -10585
rect 29680 -10705 29690 -10585
rect 24190 -10760 29690 -10705
rect 24190 -10880 24200 -10760
rect 24320 -10880 24375 -10760
rect 24495 -10880 24540 -10760
rect 24660 -10880 24705 -10760
rect 24825 -10880 24870 -10760
rect 24990 -10880 25045 -10760
rect 25165 -10880 25210 -10760
rect 25330 -10880 25375 -10760
rect 25495 -10880 25540 -10760
rect 25660 -10880 25715 -10760
rect 25835 -10880 25880 -10760
rect 26000 -10880 26045 -10760
rect 26165 -10880 26210 -10760
rect 26330 -10880 26385 -10760
rect 26505 -10880 26550 -10760
rect 26670 -10880 26715 -10760
rect 26835 -10880 26880 -10760
rect 27000 -10880 27055 -10760
rect 27175 -10880 27220 -10760
rect 27340 -10880 27385 -10760
rect 27505 -10880 27550 -10760
rect 27670 -10880 27725 -10760
rect 27845 -10880 27890 -10760
rect 28010 -10880 28055 -10760
rect 28175 -10880 28220 -10760
rect 28340 -10880 28395 -10760
rect 28515 -10880 28560 -10760
rect 28680 -10880 28725 -10760
rect 28845 -10880 28890 -10760
rect 29010 -10880 29065 -10760
rect 29185 -10880 29230 -10760
rect 29350 -10880 29395 -10760
rect 29515 -10880 29560 -10760
rect 29680 -10880 29690 -10760
rect 24190 -10925 29690 -10880
rect 24190 -11045 24200 -10925
rect 24320 -11045 24375 -10925
rect 24495 -11045 24540 -10925
rect 24660 -11045 24705 -10925
rect 24825 -11045 24870 -10925
rect 24990 -11045 25045 -10925
rect 25165 -11045 25210 -10925
rect 25330 -11045 25375 -10925
rect 25495 -11045 25540 -10925
rect 25660 -11045 25715 -10925
rect 25835 -11045 25880 -10925
rect 26000 -11045 26045 -10925
rect 26165 -11045 26210 -10925
rect 26330 -11045 26385 -10925
rect 26505 -11045 26550 -10925
rect 26670 -11045 26715 -10925
rect 26835 -11045 26880 -10925
rect 27000 -11045 27055 -10925
rect 27175 -11045 27220 -10925
rect 27340 -11045 27385 -10925
rect 27505 -11045 27550 -10925
rect 27670 -11045 27725 -10925
rect 27845 -11045 27890 -10925
rect 28010 -11045 28055 -10925
rect 28175 -11045 28220 -10925
rect 28340 -11045 28395 -10925
rect 28515 -11045 28560 -10925
rect 28680 -11045 28725 -10925
rect 28845 -11045 28890 -10925
rect 29010 -11045 29065 -10925
rect 29185 -11045 29230 -10925
rect 29350 -11045 29395 -10925
rect 29515 -11045 29560 -10925
rect 29680 -11045 29690 -10925
rect 24190 -11090 29690 -11045
rect 24190 -11210 24200 -11090
rect 24320 -11210 24375 -11090
rect 24495 -11210 24540 -11090
rect 24660 -11210 24705 -11090
rect 24825 -11210 24870 -11090
rect 24990 -11210 25045 -11090
rect 25165 -11210 25210 -11090
rect 25330 -11210 25375 -11090
rect 25495 -11210 25540 -11090
rect 25660 -11210 25715 -11090
rect 25835 -11210 25880 -11090
rect 26000 -11210 26045 -11090
rect 26165 -11210 26210 -11090
rect 26330 -11210 26385 -11090
rect 26505 -11210 26550 -11090
rect 26670 -11210 26715 -11090
rect 26835 -11210 26880 -11090
rect 27000 -11210 27055 -11090
rect 27175 -11210 27220 -11090
rect 27340 -11210 27385 -11090
rect 27505 -11210 27550 -11090
rect 27670 -11210 27725 -11090
rect 27845 -11210 27890 -11090
rect 28010 -11210 28055 -11090
rect 28175 -11210 28220 -11090
rect 28340 -11210 28395 -11090
rect 28515 -11210 28560 -11090
rect 28680 -11210 28725 -11090
rect 28845 -11210 28890 -11090
rect 29010 -11210 29065 -11090
rect 29185 -11210 29230 -11090
rect 29350 -11210 29395 -11090
rect 29515 -11210 29560 -11090
rect 29680 -11210 29690 -11090
rect 24190 -11255 29690 -11210
rect 24190 -11375 24200 -11255
rect 24320 -11375 24375 -11255
rect 24495 -11375 24540 -11255
rect 24660 -11375 24705 -11255
rect 24825 -11375 24870 -11255
rect 24990 -11375 25045 -11255
rect 25165 -11375 25210 -11255
rect 25330 -11375 25375 -11255
rect 25495 -11375 25540 -11255
rect 25660 -11375 25715 -11255
rect 25835 -11375 25880 -11255
rect 26000 -11375 26045 -11255
rect 26165 -11375 26210 -11255
rect 26330 -11375 26385 -11255
rect 26505 -11375 26550 -11255
rect 26670 -11375 26715 -11255
rect 26835 -11375 26880 -11255
rect 27000 -11375 27055 -11255
rect 27175 -11375 27220 -11255
rect 27340 -11375 27385 -11255
rect 27505 -11375 27550 -11255
rect 27670 -11375 27725 -11255
rect 27845 -11375 27890 -11255
rect 28010 -11375 28055 -11255
rect 28175 -11375 28220 -11255
rect 28340 -11375 28395 -11255
rect 28515 -11375 28560 -11255
rect 28680 -11375 28725 -11255
rect 28845 -11375 28890 -11255
rect 29010 -11375 29065 -11255
rect 29185 -11375 29230 -11255
rect 29350 -11375 29395 -11255
rect 29515 -11375 29560 -11255
rect 29680 -11375 29690 -11255
rect 24190 -11430 29690 -11375
rect 24190 -11550 24200 -11430
rect 24320 -11550 24375 -11430
rect 24495 -11550 24540 -11430
rect 24660 -11550 24705 -11430
rect 24825 -11550 24870 -11430
rect 24990 -11550 25045 -11430
rect 25165 -11550 25210 -11430
rect 25330 -11550 25375 -11430
rect 25495 -11550 25540 -11430
rect 25660 -11550 25715 -11430
rect 25835 -11550 25880 -11430
rect 26000 -11550 26045 -11430
rect 26165 -11550 26210 -11430
rect 26330 -11550 26385 -11430
rect 26505 -11550 26550 -11430
rect 26670 -11550 26715 -11430
rect 26835 -11550 26880 -11430
rect 27000 -11550 27055 -11430
rect 27175 -11550 27220 -11430
rect 27340 -11550 27385 -11430
rect 27505 -11550 27550 -11430
rect 27670 -11550 27725 -11430
rect 27845 -11550 27890 -11430
rect 28010 -11550 28055 -11430
rect 28175 -11550 28220 -11430
rect 28340 -11550 28395 -11430
rect 28515 -11550 28560 -11430
rect 28680 -11550 28725 -11430
rect 28845 -11550 28890 -11430
rect 29010 -11550 29065 -11430
rect 29185 -11550 29230 -11430
rect 29350 -11550 29395 -11430
rect 29515 -11550 29560 -11430
rect 29680 -11550 29690 -11430
rect 24190 -11595 29690 -11550
rect 24190 -11715 24200 -11595
rect 24320 -11715 24375 -11595
rect 24495 -11715 24540 -11595
rect 24660 -11715 24705 -11595
rect 24825 -11715 24870 -11595
rect 24990 -11715 25045 -11595
rect 25165 -11715 25210 -11595
rect 25330 -11715 25375 -11595
rect 25495 -11715 25540 -11595
rect 25660 -11715 25715 -11595
rect 25835 -11715 25880 -11595
rect 26000 -11715 26045 -11595
rect 26165 -11715 26210 -11595
rect 26330 -11715 26385 -11595
rect 26505 -11715 26550 -11595
rect 26670 -11715 26715 -11595
rect 26835 -11715 26880 -11595
rect 27000 -11715 27055 -11595
rect 27175 -11715 27220 -11595
rect 27340 -11715 27385 -11595
rect 27505 -11715 27550 -11595
rect 27670 -11715 27725 -11595
rect 27845 -11715 27890 -11595
rect 28010 -11715 28055 -11595
rect 28175 -11715 28220 -11595
rect 28340 -11715 28395 -11595
rect 28515 -11715 28560 -11595
rect 28680 -11715 28725 -11595
rect 28845 -11715 28890 -11595
rect 29010 -11715 29065 -11595
rect 29185 -11715 29230 -11595
rect 29350 -11715 29395 -11595
rect 29515 -11715 29560 -11595
rect 29680 -11715 29690 -11595
rect 24190 -11760 29690 -11715
rect 24190 -11880 24200 -11760
rect 24320 -11880 24375 -11760
rect 24495 -11880 24540 -11760
rect 24660 -11880 24705 -11760
rect 24825 -11880 24870 -11760
rect 24990 -11880 25045 -11760
rect 25165 -11880 25210 -11760
rect 25330 -11880 25375 -11760
rect 25495 -11880 25540 -11760
rect 25660 -11880 25715 -11760
rect 25835 -11880 25880 -11760
rect 26000 -11880 26045 -11760
rect 26165 -11880 26210 -11760
rect 26330 -11880 26385 -11760
rect 26505 -11880 26550 -11760
rect 26670 -11880 26715 -11760
rect 26835 -11880 26880 -11760
rect 27000 -11880 27055 -11760
rect 27175 -11880 27220 -11760
rect 27340 -11880 27385 -11760
rect 27505 -11880 27550 -11760
rect 27670 -11880 27725 -11760
rect 27845 -11880 27890 -11760
rect 28010 -11880 28055 -11760
rect 28175 -11880 28220 -11760
rect 28340 -11880 28395 -11760
rect 28515 -11880 28560 -11760
rect 28680 -11880 28725 -11760
rect 28845 -11880 28890 -11760
rect 29010 -11880 29065 -11760
rect 29185 -11880 29230 -11760
rect 29350 -11880 29395 -11760
rect 29515 -11880 29560 -11760
rect 29680 -11880 29690 -11760
rect 24190 -11925 29690 -11880
rect 24190 -12045 24200 -11925
rect 24320 -12045 24375 -11925
rect 24495 -12045 24540 -11925
rect 24660 -12045 24705 -11925
rect 24825 -12045 24870 -11925
rect 24990 -12045 25045 -11925
rect 25165 -12045 25210 -11925
rect 25330 -12045 25375 -11925
rect 25495 -12045 25540 -11925
rect 25660 -12045 25715 -11925
rect 25835 -12045 25880 -11925
rect 26000 -12045 26045 -11925
rect 26165 -12045 26210 -11925
rect 26330 -12045 26385 -11925
rect 26505 -12045 26550 -11925
rect 26670 -12045 26715 -11925
rect 26835 -12045 26880 -11925
rect 27000 -12045 27055 -11925
rect 27175 -12045 27220 -11925
rect 27340 -12045 27385 -11925
rect 27505 -12045 27550 -11925
rect 27670 -12045 27725 -11925
rect 27845 -12045 27890 -11925
rect 28010 -12045 28055 -11925
rect 28175 -12045 28220 -11925
rect 28340 -12045 28395 -11925
rect 28515 -12045 28560 -11925
rect 28680 -12045 28725 -11925
rect 28845 -12045 28890 -11925
rect 29010 -12045 29065 -11925
rect 29185 -12045 29230 -11925
rect 29350 -12045 29395 -11925
rect 29515 -12045 29560 -11925
rect 29680 -12045 29690 -11925
rect 24190 -12100 29690 -12045
rect 24190 -12220 24200 -12100
rect 24320 -12220 24375 -12100
rect 24495 -12220 24540 -12100
rect 24660 -12220 24705 -12100
rect 24825 -12220 24870 -12100
rect 24990 -12220 25045 -12100
rect 25165 -12220 25210 -12100
rect 25330 -12220 25375 -12100
rect 25495 -12220 25540 -12100
rect 25660 -12220 25715 -12100
rect 25835 -12220 25880 -12100
rect 26000 -12220 26045 -12100
rect 26165 -12220 26210 -12100
rect 26330 -12220 26385 -12100
rect 26505 -12220 26550 -12100
rect 26670 -12220 26715 -12100
rect 26835 -12220 26880 -12100
rect 27000 -12220 27055 -12100
rect 27175 -12220 27220 -12100
rect 27340 -12220 27385 -12100
rect 27505 -12220 27550 -12100
rect 27670 -12220 27725 -12100
rect 27845 -12220 27890 -12100
rect 28010 -12220 28055 -12100
rect 28175 -12220 28220 -12100
rect 28340 -12220 28395 -12100
rect 28515 -12220 28560 -12100
rect 28680 -12220 28725 -12100
rect 28845 -12220 28890 -12100
rect 29010 -12220 29065 -12100
rect 29185 -12220 29230 -12100
rect 29350 -12220 29395 -12100
rect 29515 -12220 29560 -12100
rect 29680 -12220 29690 -12100
rect 24190 -12265 29690 -12220
rect 24190 -12385 24200 -12265
rect 24320 -12385 24375 -12265
rect 24495 -12385 24540 -12265
rect 24660 -12385 24705 -12265
rect 24825 -12385 24870 -12265
rect 24990 -12385 25045 -12265
rect 25165 -12385 25210 -12265
rect 25330 -12385 25375 -12265
rect 25495 -12385 25540 -12265
rect 25660 -12385 25715 -12265
rect 25835 -12385 25880 -12265
rect 26000 -12385 26045 -12265
rect 26165 -12385 26210 -12265
rect 26330 -12385 26385 -12265
rect 26505 -12385 26550 -12265
rect 26670 -12385 26715 -12265
rect 26835 -12385 26880 -12265
rect 27000 -12385 27055 -12265
rect 27175 -12385 27220 -12265
rect 27340 -12385 27385 -12265
rect 27505 -12385 27550 -12265
rect 27670 -12385 27725 -12265
rect 27845 -12385 27890 -12265
rect 28010 -12385 28055 -12265
rect 28175 -12385 28220 -12265
rect 28340 -12385 28395 -12265
rect 28515 -12385 28560 -12265
rect 28680 -12385 28725 -12265
rect 28845 -12385 28890 -12265
rect 29010 -12385 29065 -12265
rect 29185 -12385 29230 -12265
rect 29350 -12385 29395 -12265
rect 29515 -12385 29560 -12265
rect 29680 -12385 29690 -12265
rect 24190 -12430 29690 -12385
rect 24190 -12550 24200 -12430
rect 24320 -12550 24375 -12430
rect 24495 -12550 24540 -12430
rect 24660 -12550 24705 -12430
rect 24825 -12550 24870 -12430
rect 24990 -12550 25045 -12430
rect 25165 -12550 25210 -12430
rect 25330 -12550 25375 -12430
rect 25495 -12550 25540 -12430
rect 25660 -12550 25715 -12430
rect 25835 -12550 25880 -12430
rect 26000 -12550 26045 -12430
rect 26165 -12550 26210 -12430
rect 26330 -12550 26385 -12430
rect 26505 -12550 26550 -12430
rect 26670 -12550 26715 -12430
rect 26835 -12550 26880 -12430
rect 27000 -12550 27055 -12430
rect 27175 -12550 27220 -12430
rect 27340 -12550 27385 -12430
rect 27505 -12550 27550 -12430
rect 27670 -12550 27725 -12430
rect 27845 -12550 27890 -12430
rect 28010 -12550 28055 -12430
rect 28175 -12550 28220 -12430
rect 28340 -12550 28395 -12430
rect 28515 -12550 28560 -12430
rect 28680 -12550 28725 -12430
rect 28845 -12550 28890 -12430
rect 29010 -12550 29065 -12430
rect 29185 -12550 29230 -12430
rect 29350 -12550 29395 -12430
rect 29515 -12550 29560 -12430
rect 29680 -12550 29690 -12430
rect 24190 -12595 29690 -12550
rect 24190 -12715 24200 -12595
rect 24320 -12715 24375 -12595
rect 24495 -12715 24540 -12595
rect 24660 -12715 24705 -12595
rect 24825 -12715 24870 -12595
rect 24990 -12715 25045 -12595
rect 25165 -12715 25210 -12595
rect 25330 -12715 25375 -12595
rect 25495 -12715 25540 -12595
rect 25660 -12715 25715 -12595
rect 25835 -12715 25880 -12595
rect 26000 -12715 26045 -12595
rect 26165 -12715 26210 -12595
rect 26330 -12715 26385 -12595
rect 26505 -12715 26550 -12595
rect 26670 -12715 26715 -12595
rect 26835 -12715 26880 -12595
rect 27000 -12715 27055 -12595
rect 27175 -12715 27220 -12595
rect 27340 -12715 27385 -12595
rect 27505 -12715 27550 -12595
rect 27670 -12715 27725 -12595
rect 27845 -12715 27890 -12595
rect 28010 -12715 28055 -12595
rect 28175 -12715 28220 -12595
rect 28340 -12715 28395 -12595
rect 28515 -12715 28560 -12595
rect 28680 -12715 28725 -12595
rect 28845 -12715 28890 -12595
rect 29010 -12715 29065 -12595
rect 29185 -12715 29230 -12595
rect 29350 -12715 29395 -12595
rect 29515 -12715 29560 -12595
rect 29680 -12715 29690 -12595
rect 24190 -12770 29690 -12715
rect 24190 -12890 24200 -12770
rect 24320 -12890 24375 -12770
rect 24495 -12890 24540 -12770
rect 24660 -12890 24705 -12770
rect 24825 -12890 24870 -12770
rect 24990 -12890 25045 -12770
rect 25165 -12890 25210 -12770
rect 25330 -12890 25375 -12770
rect 25495 -12890 25540 -12770
rect 25660 -12890 25715 -12770
rect 25835 -12890 25880 -12770
rect 26000 -12890 26045 -12770
rect 26165 -12890 26210 -12770
rect 26330 -12890 26385 -12770
rect 26505 -12890 26550 -12770
rect 26670 -12890 26715 -12770
rect 26835 -12890 26880 -12770
rect 27000 -12890 27055 -12770
rect 27175 -12890 27220 -12770
rect 27340 -12890 27385 -12770
rect 27505 -12890 27550 -12770
rect 27670 -12890 27725 -12770
rect 27845 -12890 27890 -12770
rect 28010 -12890 28055 -12770
rect 28175 -12890 28220 -12770
rect 28340 -12890 28395 -12770
rect 28515 -12890 28560 -12770
rect 28680 -12890 28725 -12770
rect 28845 -12890 28890 -12770
rect 29010 -12890 29065 -12770
rect 29185 -12890 29230 -12770
rect 29350 -12890 29395 -12770
rect 29515 -12890 29560 -12770
rect 29680 -12890 29690 -12770
rect 24190 -12935 29690 -12890
rect 24190 -13055 24200 -12935
rect 24320 -13055 24375 -12935
rect 24495 -13055 24540 -12935
rect 24660 -13055 24705 -12935
rect 24825 -13055 24870 -12935
rect 24990 -13055 25045 -12935
rect 25165 -13055 25210 -12935
rect 25330 -13055 25375 -12935
rect 25495 -13055 25540 -12935
rect 25660 -13055 25715 -12935
rect 25835 -13055 25880 -12935
rect 26000 -13055 26045 -12935
rect 26165 -13055 26210 -12935
rect 26330 -13055 26385 -12935
rect 26505 -13055 26550 -12935
rect 26670 -13055 26715 -12935
rect 26835 -13055 26880 -12935
rect 27000 -13055 27055 -12935
rect 27175 -13055 27220 -12935
rect 27340 -13055 27385 -12935
rect 27505 -13055 27550 -12935
rect 27670 -13055 27725 -12935
rect 27845 -13055 27890 -12935
rect 28010 -13055 28055 -12935
rect 28175 -13055 28220 -12935
rect 28340 -13055 28395 -12935
rect 28515 -13055 28560 -12935
rect 28680 -13055 28725 -12935
rect 28845 -13055 28890 -12935
rect 29010 -13055 29065 -12935
rect 29185 -13055 29230 -12935
rect 29350 -13055 29395 -12935
rect 29515 -13055 29560 -12935
rect 29680 -13055 29690 -12935
rect 24190 -13100 29690 -13055
rect 24190 -13220 24200 -13100
rect 24320 -13220 24375 -13100
rect 24495 -13220 24540 -13100
rect 24660 -13220 24705 -13100
rect 24825 -13220 24870 -13100
rect 24990 -13220 25045 -13100
rect 25165 -13220 25210 -13100
rect 25330 -13220 25375 -13100
rect 25495 -13220 25540 -13100
rect 25660 -13220 25715 -13100
rect 25835 -13220 25880 -13100
rect 26000 -13220 26045 -13100
rect 26165 -13220 26210 -13100
rect 26330 -13220 26385 -13100
rect 26505 -13220 26550 -13100
rect 26670 -13220 26715 -13100
rect 26835 -13220 26880 -13100
rect 27000 -13220 27055 -13100
rect 27175 -13220 27220 -13100
rect 27340 -13220 27385 -13100
rect 27505 -13220 27550 -13100
rect 27670 -13220 27725 -13100
rect 27845 -13220 27890 -13100
rect 28010 -13220 28055 -13100
rect 28175 -13220 28220 -13100
rect 28340 -13220 28395 -13100
rect 28515 -13220 28560 -13100
rect 28680 -13220 28725 -13100
rect 28845 -13220 28890 -13100
rect 29010 -13220 29065 -13100
rect 29185 -13220 29230 -13100
rect 29350 -13220 29395 -13100
rect 29515 -13220 29560 -13100
rect 29680 -13220 29690 -13100
rect 24190 -13265 29690 -13220
rect 24190 -13385 24200 -13265
rect 24320 -13385 24375 -13265
rect 24495 -13385 24540 -13265
rect 24660 -13385 24705 -13265
rect 24825 -13385 24870 -13265
rect 24990 -13385 25045 -13265
rect 25165 -13385 25210 -13265
rect 25330 -13385 25375 -13265
rect 25495 -13385 25540 -13265
rect 25660 -13385 25715 -13265
rect 25835 -13385 25880 -13265
rect 26000 -13385 26045 -13265
rect 26165 -13385 26210 -13265
rect 26330 -13385 26385 -13265
rect 26505 -13385 26550 -13265
rect 26670 -13385 26715 -13265
rect 26835 -13385 26880 -13265
rect 27000 -13385 27055 -13265
rect 27175 -13385 27220 -13265
rect 27340 -13385 27385 -13265
rect 27505 -13385 27550 -13265
rect 27670 -13385 27725 -13265
rect 27845 -13385 27890 -13265
rect 28010 -13385 28055 -13265
rect 28175 -13385 28220 -13265
rect 28340 -13385 28395 -13265
rect 28515 -13385 28560 -13265
rect 28680 -13385 28725 -13265
rect 28845 -13385 28890 -13265
rect 29010 -13385 29065 -13265
rect 29185 -13385 29230 -13265
rect 29350 -13385 29395 -13265
rect 29515 -13385 29560 -13265
rect 29680 -13385 29690 -13265
rect 24190 -13440 29690 -13385
rect 24190 -13560 24200 -13440
rect 24320 -13560 24375 -13440
rect 24495 -13560 24540 -13440
rect 24660 -13560 24705 -13440
rect 24825 -13560 24870 -13440
rect 24990 -13560 25045 -13440
rect 25165 -13560 25210 -13440
rect 25330 -13560 25375 -13440
rect 25495 -13560 25540 -13440
rect 25660 -13560 25715 -13440
rect 25835 -13560 25880 -13440
rect 26000 -13560 26045 -13440
rect 26165 -13560 26210 -13440
rect 26330 -13560 26385 -13440
rect 26505 -13560 26550 -13440
rect 26670 -13560 26715 -13440
rect 26835 -13560 26880 -13440
rect 27000 -13560 27055 -13440
rect 27175 -13560 27220 -13440
rect 27340 -13560 27385 -13440
rect 27505 -13560 27550 -13440
rect 27670 -13560 27725 -13440
rect 27845 -13560 27890 -13440
rect 28010 -13560 28055 -13440
rect 28175 -13560 28220 -13440
rect 28340 -13560 28395 -13440
rect 28515 -13560 28560 -13440
rect 28680 -13560 28725 -13440
rect 28845 -13560 28890 -13440
rect 29010 -13560 29065 -13440
rect 29185 -13560 29230 -13440
rect 29350 -13560 29395 -13440
rect 29515 -13560 29560 -13440
rect 29680 -13560 29690 -13440
rect 24190 -13605 29690 -13560
rect 24190 -13725 24200 -13605
rect 24320 -13725 24375 -13605
rect 24495 -13725 24540 -13605
rect 24660 -13725 24705 -13605
rect 24825 -13725 24870 -13605
rect 24990 -13725 25045 -13605
rect 25165 -13725 25210 -13605
rect 25330 -13725 25375 -13605
rect 25495 -13725 25540 -13605
rect 25660 -13725 25715 -13605
rect 25835 -13725 25880 -13605
rect 26000 -13725 26045 -13605
rect 26165 -13725 26210 -13605
rect 26330 -13725 26385 -13605
rect 26505 -13725 26550 -13605
rect 26670 -13725 26715 -13605
rect 26835 -13725 26880 -13605
rect 27000 -13725 27055 -13605
rect 27175 -13725 27220 -13605
rect 27340 -13725 27385 -13605
rect 27505 -13725 27550 -13605
rect 27670 -13725 27725 -13605
rect 27845 -13725 27890 -13605
rect 28010 -13725 28055 -13605
rect 28175 -13725 28220 -13605
rect 28340 -13725 28395 -13605
rect 28515 -13725 28560 -13605
rect 28680 -13725 28725 -13605
rect 28845 -13725 28890 -13605
rect 29010 -13725 29065 -13605
rect 29185 -13725 29230 -13605
rect 29350 -13725 29395 -13605
rect 29515 -13725 29560 -13605
rect 29680 -13725 29690 -13605
rect 24190 -13770 29690 -13725
rect 24190 -13890 24200 -13770
rect 24320 -13890 24375 -13770
rect 24495 -13890 24540 -13770
rect 24660 -13890 24705 -13770
rect 24825 -13890 24870 -13770
rect 24990 -13890 25045 -13770
rect 25165 -13890 25210 -13770
rect 25330 -13890 25375 -13770
rect 25495 -13890 25540 -13770
rect 25660 -13890 25715 -13770
rect 25835 -13890 25880 -13770
rect 26000 -13890 26045 -13770
rect 26165 -13890 26210 -13770
rect 26330 -13890 26385 -13770
rect 26505 -13890 26550 -13770
rect 26670 -13890 26715 -13770
rect 26835 -13890 26880 -13770
rect 27000 -13890 27055 -13770
rect 27175 -13890 27220 -13770
rect 27340 -13890 27385 -13770
rect 27505 -13890 27550 -13770
rect 27670 -13890 27725 -13770
rect 27845 -13890 27890 -13770
rect 28010 -13890 28055 -13770
rect 28175 -13890 28220 -13770
rect 28340 -13890 28395 -13770
rect 28515 -13890 28560 -13770
rect 28680 -13890 28725 -13770
rect 28845 -13890 28890 -13770
rect 29010 -13890 29065 -13770
rect 29185 -13890 29230 -13770
rect 29350 -13890 29395 -13770
rect 29515 -13890 29560 -13770
rect 29680 -13890 29690 -13770
rect 24190 -13935 29690 -13890
rect 24190 -14055 24200 -13935
rect 24320 -14055 24375 -13935
rect 24495 -14055 24540 -13935
rect 24660 -14055 24705 -13935
rect 24825 -14055 24870 -13935
rect 24990 -14055 25045 -13935
rect 25165 -14055 25210 -13935
rect 25330 -14055 25375 -13935
rect 25495 -14055 25540 -13935
rect 25660 -14055 25715 -13935
rect 25835 -14055 25880 -13935
rect 26000 -14055 26045 -13935
rect 26165 -14055 26210 -13935
rect 26330 -14055 26385 -13935
rect 26505 -14055 26550 -13935
rect 26670 -14055 26715 -13935
rect 26835 -14055 26880 -13935
rect 27000 -14055 27055 -13935
rect 27175 -14055 27220 -13935
rect 27340 -14055 27385 -13935
rect 27505 -14055 27550 -13935
rect 27670 -14055 27725 -13935
rect 27845 -14055 27890 -13935
rect 28010 -14055 28055 -13935
rect 28175 -14055 28220 -13935
rect 28340 -14055 28395 -13935
rect 28515 -14055 28560 -13935
rect 28680 -14055 28725 -13935
rect 28845 -14055 28890 -13935
rect 29010 -14055 29065 -13935
rect 29185 -14055 29230 -13935
rect 29350 -14055 29395 -13935
rect 29515 -14055 29560 -13935
rect 29680 -14055 29690 -13935
rect 24190 -14110 29690 -14055
rect 24190 -14230 24200 -14110
rect 24320 -14230 24375 -14110
rect 24495 -14230 24540 -14110
rect 24660 -14230 24705 -14110
rect 24825 -14230 24870 -14110
rect 24990 -14230 25045 -14110
rect 25165 -14230 25210 -14110
rect 25330 -14230 25375 -14110
rect 25495 -14230 25540 -14110
rect 25660 -14230 25715 -14110
rect 25835 -14230 25880 -14110
rect 26000 -14230 26045 -14110
rect 26165 -14230 26210 -14110
rect 26330 -14230 26385 -14110
rect 26505 -14230 26550 -14110
rect 26670 -14230 26715 -14110
rect 26835 -14230 26880 -14110
rect 27000 -14230 27055 -14110
rect 27175 -14230 27220 -14110
rect 27340 -14230 27385 -14110
rect 27505 -14230 27550 -14110
rect 27670 -14230 27725 -14110
rect 27845 -14230 27890 -14110
rect 28010 -14230 28055 -14110
rect 28175 -14230 28220 -14110
rect 28340 -14230 28395 -14110
rect 28515 -14230 28560 -14110
rect 28680 -14230 28725 -14110
rect 28845 -14230 28890 -14110
rect 29010 -14230 29065 -14110
rect 29185 -14230 29230 -14110
rect 29350 -14230 29395 -14110
rect 29515 -14230 29560 -14110
rect 29680 -14230 29690 -14110
rect 24190 -14275 29690 -14230
rect 24190 -14395 24200 -14275
rect 24320 -14395 24375 -14275
rect 24495 -14395 24540 -14275
rect 24660 -14395 24705 -14275
rect 24825 -14395 24870 -14275
rect 24990 -14395 25045 -14275
rect 25165 -14395 25210 -14275
rect 25330 -14395 25375 -14275
rect 25495 -14395 25540 -14275
rect 25660 -14395 25715 -14275
rect 25835 -14395 25880 -14275
rect 26000 -14395 26045 -14275
rect 26165 -14395 26210 -14275
rect 26330 -14395 26385 -14275
rect 26505 -14395 26550 -14275
rect 26670 -14395 26715 -14275
rect 26835 -14395 26880 -14275
rect 27000 -14395 27055 -14275
rect 27175 -14395 27220 -14275
rect 27340 -14395 27385 -14275
rect 27505 -14395 27550 -14275
rect 27670 -14395 27725 -14275
rect 27845 -14395 27890 -14275
rect 28010 -14395 28055 -14275
rect 28175 -14395 28220 -14275
rect 28340 -14395 28395 -14275
rect 28515 -14395 28560 -14275
rect 28680 -14395 28725 -14275
rect 28845 -14395 28890 -14275
rect 29010 -14395 29065 -14275
rect 29185 -14395 29230 -14275
rect 29350 -14395 29395 -14275
rect 29515 -14395 29560 -14275
rect 29680 -14395 29690 -14275
rect 24190 -14440 29690 -14395
rect 24190 -14560 24200 -14440
rect 24320 -14560 24375 -14440
rect 24495 -14560 24540 -14440
rect 24660 -14560 24705 -14440
rect 24825 -14560 24870 -14440
rect 24990 -14560 25045 -14440
rect 25165 -14560 25210 -14440
rect 25330 -14560 25375 -14440
rect 25495 -14560 25540 -14440
rect 25660 -14560 25715 -14440
rect 25835 -14560 25880 -14440
rect 26000 -14560 26045 -14440
rect 26165 -14560 26210 -14440
rect 26330 -14560 26385 -14440
rect 26505 -14560 26550 -14440
rect 26670 -14560 26715 -14440
rect 26835 -14560 26880 -14440
rect 27000 -14560 27055 -14440
rect 27175 -14560 27220 -14440
rect 27340 -14560 27385 -14440
rect 27505 -14560 27550 -14440
rect 27670 -14560 27725 -14440
rect 27845 -14560 27890 -14440
rect 28010 -14560 28055 -14440
rect 28175 -14560 28220 -14440
rect 28340 -14560 28395 -14440
rect 28515 -14560 28560 -14440
rect 28680 -14560 28725 -14440
rect 28845 -14560 28890 -14440
rect 29010 -14560 29065 -14440
rect 29185 -14560 29230 -14440
rect 29350 -14560 29395 -14440
rect 29515 -14560 29560 -14440
rect 29680 -14560 29690 -14440
rect 24190 -14605 29690 -14560
rect 24190 -14725 24200 -14605
rect 24320 -14725 24375 -14605
rect 24495 -14725 24540 -14605
rect 24660 -14725 24705 -14605
rect 24825 -14725 24870 -14605
rect 24990 -14725 25045 -14605
rect 25165 -14725 25210 -14605
rect 25330 -14725 25375 -14605
rect 25495 -14725 25540 -14605
rect 25660 -14725 25715 -14605
rect 25835 -14725 25880 -14605
rect 26000 -14725 26045 -14605
rect 26165 -14725 26210 -14605
rect 26330 -14725 26385 -14605
rect 26505 -14725 26550 -14605
rect 26670 -14725 26715 -14605
rect 26835 -14725 26880 -14605
rect 27000 -14725 27055 -14605
rect 27175 -14725 27220 -14605
rect 27340 -14725 27385 -14605
rect 27505 -14725 27550 -14605
rect 27670 -14725 27725 -14605
rect 27845 -14725 27890 -14605
rect 28010 -14725 28055 -14605
rect 28175 -14725 28220 -14605
rect 28340 -14725 28395 -14605
rect 28515 -14725 28560 -14605
rect 28680 -14725 28725 -14605
rect 28845 -14725 28890 -14605
rect 29010 -14725 29065 -14605
rect 29185 -14725 29230 -14605
rect 29350 -14725 29395 -14605
rect 29515 -14725 29560 -14605
rect 29680 -14725 29690 -14605
rect 24190 -14780 29690 -14725
rect 24190 -14900 24200 -14780
rect 24320 -14900 24375 -14780
rect 24495 -14900 24540 -14780
rect 24660 -14900 24705 -14780
rect 24825 -14900 24870 -14780
rect 24990 -14900 25045 -14780
rect 25165 -14900 25210 -14780
rect 25330 -14900 25375 -14780
rect 25495 -14900 25540 -14780
rect 25660 -14900 25715 -14780
rect 25835 -14900 25880 -14780
rect 26000 -14900 26045 -14780
rect 26165 -14900 26210 -14780
rect 26330 -14900 26385 -14780
rect 26505 -14900 26550 -14780
rect 26670 -14900 26715 -14780
rect 26835 -14900 26880 -14780
rect 27000 -14900 27055 -14780
rect 27175 -14900 27220 -14780
rect 27340 -14900 27385 -14780
rect 27505 -14900 27550 -14780
rect 27670 -14900 27725 -14780
rect 27845 -14900 27890 -14780
rect 28010 -14900 28055 -14780
rect 28175 -14900 28220 -14780
rect 28340 -14900 28395 -14780
rect 28515 -14900 28560 -14780
rect 28680 -14900 28725 -14780
rect 28845 -14900 28890 -14780
rect 29010 -14900 29065 -14780
rect 29185 -14900 29230 -14780
rect 29350 -14900 29395 -14780
rect 29515 -14900 29560 -14780
rect 29680 -14900 29690 -14780
rect 24190 -14945 29690 -14900
rect 24190 -15065 24200 -14945
rect 24320 -15065 24375 -14945
rect 24495 -15065 24540 -14945
rect 24660 -15065 24705 -14945
rect 24825 -15065 24870 -14945
rect 24990 -15065 25045 -14945
rect 25165 -15065 25210 -14945
rect 25330 -15065 25375 -14945
rect 25495 -15065 25540 -14945
rect 25660 -15065 25715 -14945
rect 25835 -15065 25880 -14945
rect 26000 -15065 26045 -14945
rect 26165 -15065 26210 -14945
rect 26330 -15065 26385 -14945
rect 26505 -15065 26550 -14945
rect 26670 -15065 26715 -14945
rect 26835 -15065 26880 -14945
rect 27000 -15065 27055 -14945
rect 27175 -15065 27220 -14945
rect 27340 -15065 27385 -14945
rect 27505 -15065 27550 -14945
rect 27670 -15065 27725 -14945
rect 27845 -15065 27890 -14945
rect 28010 -15065 28055 -14945
rect 28175 -15065 28220 -14945
rect 28340 -15065 28395 -14945
rect 28515 -15065 28560 -14945
rect 28680 -15065 28725 -14945
rect 28845 -15065 28890 -14945
rect 29010 -15065 29065 -14945
rect 29185 -15065 29230 -14945
rect 29350 -15065 29395 -14945
rect 29515 -15065 29560 -14945
rect 29680 -15065 29690 -14945
rect 24190 -15110 29690 -15065
rect 24190 -15230 24200 -15110
rect 24320 -15230 24375 -15110
rect 24495 -15230 24540 -15110
rect 24660 -15230 24705 -15110
rect 24825 -15230 24870 -15110
rect 24990 -15230 25045 -15110
rect 25165 -15230 25210 -15110
rect 25330 -15230 25375 -15110
rect 25495 -15230 25540 -15110
rect 25660 -15230 25715 -15110
rect 25835 -15230 25880 -15110
rect 26000 -15230 26045 -15110
rect 26165 -15230 26210 -15110
rect 26330 -15230 26385 -15110
rect 26505 -15230 26550 -15110
rect 26670 -15230 26715 -15110
rect 26835 -15230 26880 -15110
rect 27000 -15230 27055 -15110
rect 27175 -15230 27220 -15110
rect 27340 -15230 27385 -15110
rect 27505 -15230 27550 -15110
rect 27670 -15230 27725 -15110
rect 27845 -15230 27890 -15110
rect 28010 -15230 28055 -15110
rect 28175 -15230 28220 -15110
rect 28340 -15230 28395 -15110
rect 28515 -15230 28560 -15110
rect 28680 -15230 28725 -15110
rect 28845 -15230 28890 -15110
rect 29010 -15230 29065 -15110
rect 29185 -15230 29230 -15110
rect 29350 -15230 29395 -15110
rect 29515 -15230 29560 -15110
rect 29680 -15230 29690 -15110
rect 24190 -15275 29690 -15230
rect 24190 -15395 24200 -15275
rect 24320 -15395 24375 -15275
rect 24495 -15395 24540 -15275
rect 24660 -15395 24705 -15275
rect 24825 -15395 24870 -15275
rect 24990 -15395 25045 -15275
rect 25165 -15395 25210 -15275
rect 25330 -15395 25375 -15275
rect 25495 -15395 25540 -15275
rect 25660 -15395 25715 -15275
rect 25835 -15395 25880 -15275
rect 26000 -15395 26045 -15275
rect 26165 -15395 26210 -15275
rect 26330 -15395 26385 -15275
rect 26505 -15395 26550 -15275
rect 26670 -15395 26715 -15275
rect 26835 -15395 26880 -15275
rect 27000 -15395 27055 -15275
rect 27175 -15395 27220 -15275
rect 27340 -15395 27385 -15275
rect 27505 -15395 27550 -15275
rect 27670 -15395 27725 -15275
rect 27845 -15395 27890 -15275
rect 28010 -15395 28055 -15275
rect 28175 -15395 28220 -15275
rect 28340 -15395 28395 -15275
rect 28515 -15395 28560 -15275
rect 28680 -15395 28725 -15275
rect 28845 -15395 28890 -15275
rect 29010 -15395 29065 -15275
rect 29185 -15395 29230 -15275
rect 29350 -15395 29395 -15275
rect 29515 -15395 29560 -15275
rect 29680 -15395 29690 -15275
rect 24190 -15450 29690 -15395
rect 24190 -15570 24200 -15450
rect 24320 -15570 24375 -15450
rect 24495 -15570 24540 -15450
rect 24660 -15570 24705 -15450
rect 24825 -15570 24870 -15450
rect 24990 -15570 25045 -15450
rect 25165 -15570 25210 -15450
rect 25330 -15570 25375 -15450
rect 25495 -15570 25540 -15450
rect 25660 -15570 25715 -15450
rect 25835 -15570 25880 -15450
rect 26000 -15570 26045 -15450
rect 26165 -15570 26210 -15450
rect 26330 -15570 26385 -15450
rect 26505 -15570 26550 -15450
rect 26670 -15570 26715 -15450
rect 26835 -15570 26880 -15450
rect 27000 -15570 27055 -15450
rect 27175 -15570 27220 -15450
rect 27340 -15570 27385 -15450
rect 27505 -15570 27550 -15450
rect 27670 -15570 27725 -15450
rect 27845 -15570 27890 -15450
rect 28010 -15570 28055 -15450
rect 28175 -15570 28220 -15450
rect 28340 -15570 28395 -15450
rect 28515 -15570 28560 -15450
rect 28680 -15570 28725 -15450
rect 28845 -15570 28890 -15450
rect 29010 -15570 29065 -15450
rect 29185 -15570 29230 -15450
rect 29350 -15570 29395 -15450
rect 29515 -15570 29560 -15450
rect 29680 -15570 29690 -15450
rect 24190 -15580 29690 -15570
<< mimcap2contact >>
rect 7130 7040 7250 7160
rect 7295 7040 7415 7160
rect 7460 7040 7580 7160
rect 7625 7040 7745 7160
rect 7800 7040 7920 7160
rect 7965 7040 8085 7160
rect 8130 7040 8250 7160
rect 8295 7040 8415 7160
rect 8470 7040 8590 7160
rect 8635 7040 8755 7160
rect 8800 7040 8920 7160
rect 8965 7040 9085 7160
rect 9140 7040 9260 7160
rect 9305 7040 9425 7160
rect 9470 7040 9590 7160
rect 9635 7040 9755 7160
rect 9810 7040 9930 7160
rect 9975 7040 10095 7160
rect 10140 7040 10260 7160
rect 10305 7040 10425 7160
rect 10480 7040 10600 7160
rect 10645 7040 10765 7160
rect 10810 7040 10930 7160
rect 10975 7040 11095 7160
rect 11150 7040 11270 7160
rect 11315 7040 11435 7160
rect 11480 7040 11600 7160
rect 11645 7040 11765 7160
rect 11820 7040 11940 7160
rect 11985 7040 12105 7160
rect 12150 7040 12270 7160
rect 12315 7040 12435 7160
rect 12490 7040 12610 7160
rect 7130 6865 7250 6985
rect 7295 6865 7415 6985
rect 7460 6865 7580 6985
rect 7625 6865 7745 6985
rect 7800 6865 7920 6985
rect 7965 6865 8085 6985
rect 8130 6865 8250 6985
rect 8295 6865 8415 6985
rect 8470 6865 8590 6985
rect 8635 6865 8755 6985
rect 8800 6865 8920 6985
rect 8965 6865 9085 6985
rect 9140 6865 9260 6985
rect 9305 6865 9425 6985
rect 9470 6865 9590 6985
rect 9635 6865 9755 6985
rect 9810 6865 9930 6985
rect 9975 6865 10095 6985
rect 10140 6865 10260 6985
rect 10305 6865 10425 6985
rect 10480 6865 10600 6985
rect 10645 6865 10765 6985
rect 10810 6865 10930 6985
rect 10975 6865 11095 6985
rect 11150 6865 11270 6985
rect 11315 6865 11435 6985
rect 11480 6865 11600 6985
rect 11645 6865 11765 6985
rect 11820 6865 11940 6985
rect 11985 6865 12105 6985
rect 12150 6865 12270 6985
rect 12315 6865 12435 6985
rect 12490 6865 12610 6985
rect 7130 6700 7250 6820
rect 7295 6700 7415 6820
rect 7460 6700 7580 6820
rect 7625 6700 7745 6820
rect 7800 6700 7920 6820
rect 7965 6700 8085 6820
rect 8130 6700 8250 6820
rect 8295 6700 8415 6820
rect 8470 6700 8590 6820
rect 8635 6700 8755 6820
rect 8800 6700 8920 6820
rect 8965 6700 9085 6820
rect 9140 6700 9260 6820
rect 9305 6700 9425 6820
rect 9470 6700 9590 6820
rect 9635 6700 9755 6820
rect 9810 6700 9930 6820
rect 9975 6700 10095 6820
rect 10140 6700 10260 6820
rect 10305 6700 10425 6820
rect 10480 6700 10600 6820
rect 10645 6700 10765 6820
rect 10810 6700 10930 6820
rect 10975 6700 11095 6820
rect 11150 6700 11270 6820
rect 11315 6700 11435 6820
rect 11480 6700 11600 6820
rect 11645 6700 11765 6820
rect 11820 6700 11940 6820
rect 11985 6700 12105 6820
rect 12150 6700 12270 6820
rect 12315 6700 12435 6820
rect 12490 6700 12610 6820
rect 7130 6535 7250 6655
rect 7295 6535 7415 6655
rect 7460 6535 7580 6655
rect 7625 6535 7745 6655
rect 7800 6535 7920 6655
rect 7965 6535 8085 6655
rect 8130 6535 8250 6655
rect 8295 6535 8415 6655
rect 8470 6535 8590 6655
rect 8635 6535 8755 6655
rect 8800 6535 8920 6655
rect 8965 6535 9085 6655
rect 9140 6535 9260 6655
rect 9305 6535 9425 6655
rect 9470 6535 9590 6655
rect 9635 6535 9755 6655
rect 9810 6535 9930 6655
rect 9975 6535 10095 6655
rect 10140 6535 10260 6655
rect 10305 6535 10425 6655
rect 10480 6535 10600 6655
rect 10645 6535 10765 6655
rect 10810 6535 10930 6655
rect 10975 6535 11095 6655
rect 11150 6535 11270 6655
rect 11315 6535 11435 6655
rect 11480 6535 11600 6655
rect 11645 6535 11765 6655
rect 11820 6535 11940 6655
rect 11985 6535 12105 6655
rect 12150 6535 12270 6655
rect 12315 6535 12435 6655
rect 12490 6535 12610 6655
rect 7130 6370 7250 6490
rect 7295 6370 7415 6490
rect 7460 6370 7580 6490
rect 7625 6370 7745 6490
rect 7800 6370 7920 6490
rect 7965 6370 8085 6490
rect 8130 6370 8250 6490
rect 8295 6370 8415 6490
rect 8470 6370 8590 6490
rect 8635 6370 8755 6490
rect 8800 6370 8920 6490
rect 8965 6370 9085 6490
rect 9140 6370 9260 6490
rect 9305 6370 9425 6490
rect 9470 6370 9590 6490
rect 9635 6370 9755 6490
rect 9810 6370 9930 6490
rect 9975 6370 10095 6490
rect 10140 6370 10260 6490
rect 10305 6370 10425 6490
rect 10480 6370 10600 6490
rect 10645 6370 10765 6490
rect 10810 6370 10930 6490
rect 10975 6370 11095 6490
rect 11150 6370 11270 6490
rect 11315 6370 11435 6490
rect 11480 6370 11600 6490
rect 11645 6370 11765 6490
rect 11820 6370 11940 6490
rect 11985 6370 12105 6490
rect 12150 6370 12270 6490
rect 12315 6370 12435 6490
rect 12490 6370 12610 6490
rect 7130 6195 7250 6315
rect 7295 6195 7415 6315
rect 7460 6195 7580 6315
rect 7625 6195 7745 6315
rect 7800 6195 7920 6315
rect 7965 6195 8085 6315
rect 8130 6195 8250 6315
rect 8295 6195 8415 6315
rect 8470 6195 8590 6315
rect 8635 6195 8755 6315
rect 8800 6195 8920 6315
rect 8965 6195 9085 6315
rect 9140 6195 9260 6315
rect 9305 6195 9425 6315
rect 9470 6195 9590 6315
rect 9635 6195 9755 6315
rect 9810 6195 9930 6315
rect 9975 6195 10095 6315
rect 10140 6195 10260 6315
rect 10305 6195 10425 6315
rect 10480 6195 10600 6315
rect 10645 6195 10765 6315
rect 10810 6195 10930 6315
rect 10975 6195 11095 6315
rect 11150 6195 11270 6315
rect 11315 6195 11435 6315
rect 11480 6195 11600 6315
rect 11645 6195 11765 6315
rect 11820 6195 11940 6315
rect 11985 6195 12105 6315
rect 12150 6195 12270 6315
rect 12315 6195 12435 6315
rect 12490 6195 12610 6315
rect 7130 6030 7250 6150
rect 7295 6030 7415 6150
rect 7460 6030 7580 6150
rect 7625 6030 7745 6150
rect 7800 6030 7920 6150
rect 7965 6030 8085 6150
rect 8130 6030 8250 6150
rect 8295 6030 8415 6150
rect 8470 6030 8590 6150
rect 8635 6030 8755 6150
rect 8800 6030 8920 6150
rect 8965 6030 9085 6150
rect 9140 6030 9260 6150
rect 9305 6030 9425 6150
rect 9470 6030 9590 6150
rect 9635 6030 9755 6150
rect 9810 6030 9930 6150
rect 9975 6030 10095 6150
rect 10140 6030 10260 6150
rect 10305 6030 10425 6150
rect 10480 6030 10600 6150
rect 10645 6030 10765 6150
rect 10810 6030 10930 6150
rect 10975 6030 11095 6150
rect 11150 6030 11270 6150
rect 11315 6030 11435 6150
rect 11480 6030 11600 6150
rect 11645 6030 11765 6150
rect 11820 6030 11940 6150
rect 11985 6030 12105 6150
rect 12150 6030 12270 6150
rect 12315 6030 12435 6150
rect 12490 6030 12610 6150
rect 7130 5865 7250 5985
rect 7295 5865 7415 5985
rect 7460 5865 7580 5985
rect 7625 5865 7745 5985
rect 7800 5865 7920 5985
rect 7965 5865 8085 5985
rect 8130 5865 8250 5985
rect 8295 5865 8415 5985
rect 8470 5865 8590 5985
rect 8635 5865 8755 5985
rect 8800 5865 8920 5985
rect 8965 5865 9085 5985
rect 9140 5865 9260 5985
rect 9305 5865 9425 5985
rect 9470 5865 9590 5985
rect 9635 5865 9755 5985
rect 9810 5865 9930 5985
rect 9975 5865 10095 5985
rect 10140 5865 10260 5985
rect 10305 5865 10425 5985
rect 10480 5865 10600 5985
rect 10645 5865 10765 5985
rect 10810 5865 10930 5985
rect 10975 5865 11095 5985
rect 11150 5865 11270 5985
rect 11315 5865 11435 5985
rect 11480 5865 11600 5985
rect 11645 5865 11765 5985
rect 11820 5865 11940 5985
rect 11985 5865 12105 5985
rect 12150 5865 12270 5985
rect 12315 5865 12435 5985
rect 12490 5865 12610 5985
rect 7130 5700 7250 5820
rect 7295 5700 7415 5820
rect 7460 5700 7580 5820
rect 7625 5700 7745 5820
rect 7800 5700 7920 5820
rect 7965 5700 8085 5820
rect 8130 5700 8250 5820
rect 8295 5700 8415 5820
rect 8470 5700 8590 5820
rect 8635 5700 8755 5820
rect 8800 5700 8920 5820
rect 8965 5700 9085 5820
rect 9140 5700 9260 5820
rect 9305 5700 9425 5820
rect 9470 5700 9590 5820
rect 9635 5700 9755 5820
rect 9810 5700 9930 5820
rect 9975 5700 10095 5820
rect 10140 5700 10260 5820
rect 10305 5700 10425 5820
rect 10480 5700 10600 5820
rect 10645 5700 10765 5820
rect 10810 5700 10930 5820
rect 10975 5700 11095 5820
rect 11150 5700 11270 5820
rect 11315 5700 11435 5820
rect 11480 5700 11600 5820
rect 11645 5700 11765 5820
rect 11820 5700 11940 5820
rect 11985 5700 12105 5820
rect 12150 5700 12270 5820
rect 12315 5700 12435 5820
rect 12490 5700 12610 5820
rect 7130 5525 7250 5645
rect 7295 5525 7415 5645
rect 7460 5525 7580 5645
rect 7625 5525 7745 5645
rect 7800 5525 7920 5645
rect 7965 5525 8085 5645
rect 8130 5525 8250 5645
rect 8295 5525 8415 5645
rect 8470 5525 8590 5645
rect 8635 5525 8755 5645
rect 8800 5525 8920 5645
rect 8965 5525 9085 5645
rect 9140 5525 9260 5645
rect 9305 5525 9425 5645
rect 9470 5525 9590 5645
rect 9635 5525 9755 5645
rect 9810 5525 9930 5645
rect 9975 5525 10095 5645
rect 10140 5525 10260 5645
rect 10305 5525 10425 5645
rect 10480 5525 10600 5645
rect 10645 5525 10765 5645
rect 10810 5525 10930 5645
rect 10975 5525 11095 5645
rect 11150 5525 11270 5645
rect 11315 5525 11435 5645
rect 11480 5525 11600 5645
rect 11645 5525 11765 5645
rect 11820 5525 11940 5645
rect 11985 5525 12105 5645
rect 12150 5525 12270 5645
rect 12315 5525 12435 5645
rect 12490 5525 12610 5645
rect 7130 5360 7250 5480
rect 7295 5360 7415 5480
rect 7460 5360 7580 5480
rect 7625 5360 7745 5480
rect 7800 5360 7920 5480
rect 7965 5360 8085 5480
rect 8130 5360 8250 5480
rect 8295 5360 8415 5480
rect 8470 5360 8590 5480
rect 8635 5360 8755 5480
rect 8800 5360 8920 5480
rect 8965 5360 9085 5480
rect 9140 5360 9260 5480
rect 9305 5360 9425 5480
rect 9470 5360 9590 5480
rect 9635 5360 9755 5480
rect 9810 5360 9930 5480
rect 9975 5360 10095 5480
rect 10140 5360 10260 5480
rect 10305 5360 10425 5480
rect 10480 5360 10600 5480
rect 10645 5360 10765 5480
rect 10810 5360 10930 5480
rect 10975 5360 11095 5480
rect 11150 5360 11270 5480
rect 11315 5360 11435 5480
rect 11480 5360 11600 5480
rect 11645 5360 11765 5480
rect 11820 5360 11940 5480
rect 11985 5360 12105 5480
rect 12150 5360 12270 5480
rect 12315 5360 12435 5480
rect 12490 5360 12610 5480
rect 7130 5195 7250 5315
rect 7295 5195 7415 5315
rect 7460 5195 7580 5315
rect 7625 5195 7745 5315
rect 7800 5195 7920 5315
rect 7965 5195 8085 5315
rect 8130 5195 8250 5315
rect 8295 5195 8415 5315
rect 8470 5195 8590 5315
rect 8635 5195 8755 5315
rect 8800 5195 8920 5315
rect 8965 5195 9085 5315
rect 9140 5195 9260 5315
rect 9305 5195 9425 5315
rect 9470 5195 9590 5315
rect 9635 5195 9755 5315
rect 9810 5195 9930 5315
rect 9975 5195 10095 5315
rect 10140 5195 10260 5315
rect 10305 5195 10425 5315
rect 10480 5195 10600 5315
rect 10645 5195 10765 5315
rect 10810 5195 10930 5315
rect 10975 5195 11095 5315
rect 11150 5195 11270 5315
rect 11315 5195 11435 5315
rect 11480 5195 11600 5315
rect 11645 5195 11765 5315
rect 11820 5195 11940 5315
rect 11985 5195 12105 5315
rect 12150 5195 12270 5315
rect 12315 5195 12435 5315
rect 12490 5195 12610 5315
rect 7130 5030 7250 5150
rect 7295 5030 7415 5150
rect 7460 5030 7580 5150
rect 7625 5030 7745 5150
rect 7800 5030 7920 5150
rect 7965 5030 8085 5150
rect 8130 5030 8250 5150
rect 8295 5030 8415 5150
rect 8470 5030 8590 5150
rect 8635 5030 8755 5150
rect 8800 5030 8920 5150
rect 8965 5030 9085 5150
rect 9140 5030 9260 5150
rect 9305 5030 9425 5150
rect 9470 5030 9590 5150
rect 9635 5030 9755 5150
rect 9810 5030 9930 5150
rect 9975 5030 10095 5150
rect 10140 5030 10260 5150
rect 10305 5030 10425 5150
rect 10480 5030 10600 5150
rect 10645 5030 10765 5150
rect 10810 5030 10930 5150
rect 10975 5030 11095 5150
rect 11150 5030 11270 5150
rect 11315 5030 11435 5150
rect 11480 5030 11600 5150
rect 11645 5030 11765 5150
rect 11820 5030 11940 5150
rect 11985 5030 12105 5150
rect 12150 5030 12270 5150
rect 12315 5030 12435 5150
rect 12490 5030 12610 5150
rect 7130 4855 7250 4975
rect 7295 4855 7415 4975
rect 7460 4855 7580 4975
rect 7625 4855 7745 4975
rect 7800 4855 7920 4975
rect 7965 4855 8085 4975
rect 8130 4855 8250 4975
rect 8295 4855 8415 4975
rect 8470 4855 8590 4975
rect 8635 4855 8755 4975
rect 8800 4855 8920 4975
rect 8965 4855 9085 4975
rect 9140 4855 9260 4975
rect 9305 4855 9425 4975
rect 9470 4855 9590 4975
rect 9635 4855 9755 4975
rect 9810 4855 9930 4975
rect 9975 4855 10095 4975
rect 10140 4855 10260 4975
rect 10305 4855 10425 4975
rect 10480 4855 10600 4975
rect 10645 4855 10765 4975
rect 10810 4855 10930 4975
rect 10975 4855 11095 4975
rect 11150 4855 11270 4975
rect 11315 4855 11435 4975
rect 11480 4855 11600 4975
rect 11645 4855 11765 4975
rect 11820 4855 11940 4975
rect 11985 4855 12105 4975
rect 12150 4855 12270 4975
rect 12315 4855 12435 4975
rect 12490 4855 12610 4975
rect 7130 4690 7250 4810
rect 7295 4690 7415 4810
rect 7460 4690 7580 4810
rect 7625 4690 7745 4810
rect 7800 4690 7920 4810
rect 7965 4690 8085 4810
rect 8130 4690 8250 4810
rect 8295 4690 8415 4810
rect 8470 4690 8590 4810
rect 8635 4690 8755 4810
rect 8800 4690 8920 4810
rect 8965 4690 9085 4810
rect 9140 4690 9260 4810
rect 9305 4690 9425 4810
rect 9470 4690 9590 4810
rect 9635 4690 9755 4810
rect 9810 4690 9930 4810
rect 9975 4690 10095 4810
rect 10140 4690 10260 4810
rect 10305 4690 10425 4810
rect 10480 4690 10600 4810
rect 10645 4690 10765 4810
rect 10810 4690 10930 4810
rect 10975 4690 11095 4810
rect 11150 4690 11270 4810
rect 11315 4690 11435 4810
rect 11480 4690 11600 4810
rect 11645 4690 11765 4810
rect 11820 4690 11940 4810
rect 11985 4690 12105 4810
rect 12150 4690 12270 4810
rect 12315 4690 12435 4810
rect 12490 4690 12610 4810
rect 7130 4525 7250 4645
rect 7295 4525 7415 4645
rect 7460 4525 7580 4645
rect 7625 4525 7745 4645
rect 7800 4525 7920 4645
rect 7965 4525 8085 4645
rect 8130 4525 8250 4645
rect 8295 4525 8415 4645
rect 8470 4525 8590 4645
rect 8635 4525 8755 4645
rect 8800 4525 8920 4645
rect 8965 4525 9085 4645
rect 9140 4525 9260 4645
rect 9305 4525 9425 4645
rect 9470 4525 9590 4645
rect 9635 4525 9755 4645
rect 9810 4525 9930 4645
rect 9975 4525 10095 4645
rect 10140 4525 10260 4645
rect 10305 4525 10425 4645
rect 10480 4525 10600 4645
rect 10645 4525 10765 4645
rect 10810 4525 10930 4645
rect 10975 4525 11095 4645
rect 11150 4525 11270 4645
rect 11315 4525 11435 4645
rect 11480 4525 11600 4645
rect 11645 4525 11765 4645
rect 11820 4525 11940 4645
rect 11985 4525 12105 4645
rect 12150 4525 12270 4645
rect 12315 4525 12435 4645
rect 12490 4525 12610 4645
rect 7130 4360 7250 4480
rect 7295 4360 7415 4480
rect 7460 4360 7580 4480
rect 7625 4360 7745 4480
rect 7800 4360 7920 4480
rect 7965 4360 8085 4480
rect 8130 4360 8250 4480
rect 8295 4360 8415 4480
rect 8470 4360 8590 4480
rect 8635 4360 8755 4480
rect 8800 4360 8920 4480
rect 8965 4360 9085 4480
rect 9140 4360 9260 4480
rect 9305 4360 9425 4480
rect 9470 4360 9590 4480
rect 9635 4360 9755 4480
rect 9810 4360 9930 4480
rect 9975 4360 10095 4480
rect 10140 4360 10260 4480
rect 10305 4360 10425 4480
rect 10480 4360 10600 4480
rect 10645 4360 10765 4480
rect 10810 4360 10930 4480
rect 10975 4360 11095 4480
rect 11150 4360 11270 4480
rect 11315 4360 11435 4480
rect 11480 4360 11600 4480
rect 11645 4360 11765 4480
rect 11820 4360 11940 4480
rect 11985 4360 12105 4480
rect 12150 4360 12270 4480
rect 12315 4360 12435 4480
rect 12490 4360 12610 4480
rect 7130 4185 7250 4305
rect 7295 4185 7415 4305
rect 7460 4185 7580 4305
rect 7625 4185 7745 4305
rect 7800 4185 7920 4305
rect 7965 4185 8085 4305
rect 8130 4185 8250 4305
rect 8295 4185 8415 4305
rect 8470 4185 8590 4305
rect 8635 4185 8755 4305
rect 8800 4185 8920 4305
rect 8965 4185 9085 4305
rect 9140 4185 9260 4305
rect 9305 4185 9425 4305
rect 9470 4185 9590 4305
rect 9635 4185 9755 4305
rect 9810 4185 9930 4305
rect 9975 4185 10095 4305
rect 10140 4185 10260 4305
rect 10305 4185 10425 4305
rect 10480 4185 10600 4305
rect 10645 4185 10765 4305
rect 10810 4185 10930 4305
rect 10975 4185 11095 4305
rect 11150 4185 11270 4305
rect 11315 4185 11435 4305
rect 11480 4185 11600 4305
rect 11645 4185 11765 4305
rect 11820 4185 11940 4305
rect 11985 4185 12105 4305
rect 12150 4185 12270 4305
rect 12315 4185 12435 4305
rect 12490 4185 12610 4305
rect 7130 4020 7250 4140
rect 7295 4020 7415 4140
rect 7460 4020 7580 4140
rect 7625 4020 7745 4140
rect 7800 4020 7920 4140
rect 7965 4020 8085 4140
rect 8130 4020 8250 4140
rect 8295 4020 8415 4140
rect 8470 4020 8590 4140
rect 8635 4020 8755 4140
rect 8800 4020 8920 4140
rect 8965 4020 9085 4140
rect 9140 4020 9260 4140
rect 9305 4020 9425 4140
rect 9470 4020 9590 4140
rect 9635 4020 9755 4140
rect 9810 4020 9930 4140
rect 9975 4020 10095 4140
rect 10140 4020 10260 4140
rect 10305 4020 10425 4140
rect 10480 4020 10600 4140
rect 10645 4020 10765 4140
rect 10810 4020 10930 4140
rect 10975 4020 11095 4140
rect 11150 4020 11270 4140
rect 11315 4020 11435 4140
rect 11480 4020 11600 4140
rect 11645 4020 11765 4140
rect 11820 4020 11940 4140
rect 11985 4020 12105 4140
rect 12150 4020 12270 4140
rect 12315 4020 12435 4140
rect 12490 4020 12610 4140
rect 7130 3855 7250 3975
rect 7295 3855 7415 3975
rect 7460 3855 7580 3975
rect 7625 3855 7745 3975
rect 7800 3855 7920 3975
rect 7965 3855 8085 3975
rect 8130 3855 8250 3975
rect 8295 3855 8415 3975
rect 8470 3855 8590 3975
rect 8635 3855 8755 3975
rect 8800 3855 8920 3975
rect 8965 3855 9085 3975
rect 9140 3855 9260 3975
rect 9305 3855 9425 3975
rect 9470 3855 9590 3975
rect 9635 3855 9755 3975
rect 9810 3855 9930 3975
rect 9975 3855 10095 3975
rect 10140 3855 10260 3975
rect 10305 3855 10425 3975
rect 10480 3855 10600 3975
rect 10645 3855 10765 3975
rect 10810 3855 10930 3975
rect 10975 3855 11095 3975
rect 11150 3855 11270 3975
rect 11315 3855 11435 3975
rect 11480 3855 11600 3975
rect 11645 3855 11765 3975
rect 11820 3855 11940 3975
rect 11985 3855 12105 3975
rect 12150 3855 12270 3975
rect 12315 3855 12435 3975
rect 12490 3855 12610 3975
rect 7130 3690 7250 3810
rect 7295 3690 7415 3810
rect 7460 3690 7580 3810
rect 7625 3690 7745 3810
rect 7800 3690 7920 3810
rect 7965 3690 8085 3810
rect 8130 3690 8250 3810
rect 8295 3690 8415 3810
rect 8470 3690 8590 3810
rect 8635 3690 8755 3810
rect 8800 3690 8920 3810
rect 8965 3690 9085 3810
rect 9140 3690 9260 3810
rect 9305 3690 9425 3810
rect 9470 3690 9590 3810
rect 9635 3690 9755 3810
rect 9810 3690 9930 3810
rect 9975 3690 10095 3810
rect 10140 3690 10260 3810
rect 10305 3690 10425 3810
rect 10480 3690 10600 3810
rect 10645 3690 10765 3810
rect 10810 3690 10930 3810
rect 10975 3690 11095 3810
rect 11150 3690 11270 3810
rect 11315 3690 11435 3810
rect 11480 3690 11600 3810
rect 11645 3690 11765 3810
rect 11820 3690 11940 3810
rect 11985 3690 12105 3810
rect 12150 3690 12270 3810
rect 12315 3690 12435 3810
rect 12490 3690 12610 3810
rect 7130 3515 7250 3635
rect 7295 3515 7415 3635
rect 7460 3515 7580 3635
rect 7625 3515 7745 3635
rect 7800 3515 7920 3635
rect 7965 3515 8085 3635
rect 8130 3515 8250 3635
rect 8295 3515 8415 3635
rect 8470 3515 8590 3635
rect 8635 3515 8755 3635
rect 8800 3515 8920 3635
rect 8965 3515 9085 3635
rect 9140 3515 9260 3635
rect 9305 3515 9425 3635
rect 9470 3515 9590 3635
rect 9635 3515 9755 3635
rect 9810 3515 9930 3635
rect 9975 3515 10095 3635
rect 10140 3515 10260 3635
rect 10305 3515 10425 3635
rect 10480 3515 10600 3635
rect 10645 3515 10765 3635
rect 10810 3515 10930 3635
rect 10975 3515 11095 3635
rect 11150 3515 11270 3635
rect 11315 3515 11435 3635
rect 11480 3515 11600 3635
rect 11645 3515 11765 3635
rect 11820 3515 11940 3635
rect 11985 3515 12105 3635
rect 12150 3515 12270 3635
rect 12315 3515 12435 3635
rect 12490 3515 12610 3635
rect 7130 3350 7250 3470
rect 7295 3350 7415 3470
rect 7460 3350 7580 3470
rect 7625 3350 7745 3470
rect 7800 3350 7920 3470
rect 7965 3350 8085 3470
rect 8130 3350 8250 3470
rect 8295 3350 8415 3470
rect 8470 3350 8590 3470
rect 8635 3350 8755 3470
rect 8800 3350 8920 3470
rect 8965 3350 9085 3470
rect 9140 3350 9260 3470
rect 9305 3350 9425 3470
rect 9470 3350 9590 3470
rect 9635 3350 9755 3470
rect 9810 3350 9930 3470
rect 9975 3350 10095 3470
rect 10140 3350 10260 3470
rect 10305 3350 10425 3470
rect 10480 3350 10600 3470
rect 10645 3350 10765 3470
rect 10810 3350 10930 3470
rect 10975 3350 11095 3470
rect 11150 3350 11270 3470
rect 11315 3350 11435 3470
rect 11480 3350 11600 3470
rect 11645 3350 11765 3470
rect 11820 3350 11940 3470
rect 11985 3350 12105 3470
rect 12150 3350 12270 3470
rect 12315 3350 12435 3470
rect 12490 3350 12610 3470
rect 7130 3185 7250 3305
rect 7295 3185 7415 3305
rect 7460 3185 7580 3305
rect 7625 3185 7745 3305
rect 7800 3185 7920 3305
rect 7965 3185 8085 3305
rect 8130 3185 8250 3305
rect 8295 3185 8415 3305
rect 8470 3185 8590 3305
rect 8635 3185 8755 3305
rect 8800 3185 8920 3305
rect 8965 3185 9085 3305
rect 9140 3185 9260 3305
rect 9305 3185 9425 3305
rect 9470 3185 9590 3305
rect 9635 3185 9755 3305
rect 9810 3185 9930 3305
rect 9975 3185 10095 3305
rect 10140 3185 10260 3305
rect 10305 3185 10425 3305
rect 10480 3185 10600 3305
rect 10645 3185 10765 3305
rect 10810 3185 10930 3305
rect 10975 3185 11095 3305
rect 11150 3185 11270 3305
rect 11315 3185 11435 3305
rect 11480 3185 11600 3305
rect 11645 3185 11765 3305
rect 11820 3185 11940 3305
rect 11985 3185 12105 3305
rect 12150 3185 12270 3305
rect 12315 3185 12435 3305
rect 12490 3185 12610 3305
rect 7130 3020 7250 3140
rect 7295 3020 7415 3140
rect 7460 3020 7580 3140
rect 7625 3020 7745 3140
rect 7800 3020 7920 3140
rect 7965 3020 8085 3140
rect 8130 3020 8250 3140
rect 8295 3020 8415 3140
rect 8470 3020 8590 3140
rect 8635 3020 8755 3140
rect 8800 3020 8920 3140
rect 8965 3020 9085 3140
rect 9140 3020 9260 3140
rect 9305 3020 9425 3140
rect 9470 3020 9590 3140
rect 9635 3020 9755 3140
rect 9810 3020 9930 3140
rect 9975 3020 10095 3140
rect 10140 3020 10260 3140
rect 10305 3020 10425 3140
rect 10480 3020 10600 3140
rect 10645 3020 10765 3140
rect 10810 3020 10930 3140
rect 10975 3020 11095 3140
rect 11150 3020 11270 3140
rect 11315 3020 11435 3140
rect 11480 3020 11600 3140
rect 11645 3020 11765 3140
rect 11820 3020 11940 3140
rect 11985 3020 12105 3140
rect 12150 3020 12270 3140
rect 12315 3020 12435 3140
rect 12490 3020 12610 3140
rect 7130 2845 7250 2965
rect 7295 2845 7415 2965
rect 7460 2845 7580 2965
rect 7625 2845 7745 2965
rect 7800 2845 7920 2965
rect 7965 2845 8085 2965
rect 8130 2845 8250 2965
rect 8295 2845 8415 2965
rect 8470 2845 8590 2965
rect 8635 2845 8755 2965
rect 8800 2845 8920 2965
rect 8965 2845 9085 2965
rect 9140 2845 9260 2965
rect 9305 2845 9425 2965
rect 9470 2845 9590 2965
rect 9635 2845 9755 2965
rect 9810 2845 9930 2965
rect 9975 2845 10095 2965
rect 10140 2845 10260 2965
rect 10305 2845 10425 2965
rect 10480 2845 10600 2965
rect 10645 2845 10765 2965
rect 10810 2845 10930 2965
rect 10975 2845 11095 2965
rect 11150 2845 11270 2965
rect 11315 2845 11435 2965
rect 11480 2845 11600 2965
rect 11645 2845 11765 2965
rect 11820 2845 11940 2965
rect 11985 2845 12105 2965
rect 12150 2845 12270 2965
rect 12315 2845 12435 2965
rect 12490 2845 12610 2965
rect 7130 2680 7250 2800
rect 7295 2680 7415 2800
rect 7460 2680 7580 2800
rect 7625 2680 7745 2800
rect 7800 2680 7920 2800
rect 7965 2680 8085 2800
rect 8130 2680 8250 2800
rect 8295 2680 8415 2800
rect 8470 2680 8590 2800
rect 8635 2680 8755 2800
rect 8800 2680 8920 2800
rect 8965 2680 9085 2800
rect 9140 2680 9260 2800
rect 9305 2680 9425 2800
rect 9470 2680 9590 2800
rect 9635 2680 9755 2800
rect 9810 2680 9930 2800
rect 9975 2680 10095 2800
rect 10140 2680 10260 2800
rect 10305 2680 10425 2800
rect 10480 2680 10600 2800
rect 10645 2680 10765 2800
rect 10810 2680 10930 2800
rect 10975 2680 11095 2800
rect 11150 2680 11270 2800
rect 11315 2680 11435 2800
rect 11480 2680 11600 2800
rect 11645 2680 11765 2800
rect 11820 2680 11940 2800
rect 11985 2680 12105 2800
rect 12150 2680 12270 2800
rect 12315 2680 12435 2800
rect 12490 2680 12610 2800
rect 7130 2515 7250 2635
rect 7295 2515 7415 2635
rect 7460 2515 7580 2635
rect 7625 2515 7745 2635
rect 7800 2515 7920 2635
rect 7965 2515 8085 2635
rect 8130 2515 8250 2635
rect 8295 2515 8415 2635
rect 8470 2515 8590 2635
rect 8635 2515 8755 2635
rect 8800 2515 8920 2635
rect 8965 2515 9085 2635
rect 9140 2515 9260 2635
rect 9305 2515 9425 2635
rect 9470 2515 9590 2635
rect 9635 2515 9755 2635
rect 9810 2515 9930 2635
rect 9975 2515 10095 2635
rect 10140 2515 10260 2635
rect 10305 2515 10425 2635
rect 10480 2515 10600 2635
rect 10645 2515 10765 2635
rect 10810 2515 10930 2635
rect 10975 2515 11095 2635
rect 11150 2515 11270 2635
rect 11315 2515 11435 2635
rect 11480 2515 11600 2635
rect 11645 2515 11765 2635
rect 11820 2515 11940 2635
rect 11985 2515 12105 2635
rect 12150 2515 12270 2635
rect 12315 2515 12435 2635
rect 12490 2515 12610 2635
rect 7130 2350 7250 2470
rect 7295 2350 7415 2470
rect 7460 2350 7580 2470
rect 7625 2350 7745 2470
rect 7800 2350 7920 2470
rect 7965 2350 8085 2470
rect 8130 2350 8250 2470
rect 8295 2350 8415 2470
rect 8470 2350 8590 2470
rect 8635 2350 8755 2470
rect 8800 2350 8920 2470
rect 8965 2350 9085 2470
rect 9140 2350 9260 2470
rect 9305 2350 9425 2470
rect 9470 2350 9590 2470
rect 9635 2350 9755 2470
rect 9810 2350 9930 2470
rect 9975 2350 10095 2470
rect 10140 2350 10260 2470
rect 10305 2350 10425 2470
rect 10480 2350 10600 2470
rect 10645 2350 10765 2470
rect 10810 2350 10930 2470
rect 10975 2350 11095 2470
rect 11150 2350 11270 2470
rect 11315 2350 11435 2470
rect 11480 2350 11600 2470
rect 11645 2350 11765 2470
rect 11820 2350 11940 2470
rect 11985 2350 12105 2470
rect 12150 2350 12270 2470
rect 12315 2350 12435 2470
rect 12490 2350 12610 2470
rect 7130 2175 7250 2295
rect 7295 2175 7415 2295
rect 7460 2175 7580 2295
rect 7625 2175 7745 2295
rect 7800 2175 7920 2295
rect 7965 2175 8085 2295
rect 8130 2175 8250 2295
rect 8295 2175 8415 2295
rect 8470 2175 8590 2295
rect 8635 2175 8755 2295
rect 8800 2175 8920 2295
rect 8965 2175 9085 2295
rect 9140 2175 9260 2295
rect 9305 2175 9425 2295
rect 9470 2175 9590 2295
rect 9635 2175 9755 2295
rect 9810 2175 9930 2295
rect 9975 2175 10095 2295
rect 10140 2175 10260 2295
rect 10305 2175 10425 2295
rect 10480 2175 10600 2295
rect 10645 2175 10765 2295
rect 10810 2175 10930 2295
rect 10975 2175 11095 2295
rect 11150 2175 11270 2295
rect 11315 2175 11435 2295
rect 11480 2175 11600 2295
rect 11645 2175 11765 2295
rect 11820 2175 11940 2295
rect 11985 2175 12105 2295
rect 12150 2175 12270 2295
rect 12315 2175 12435 2295
rect 12490 2175 12610 2295
rect 7130 2010 7250 2130
rect 7295 2010 7415 2130
rect 7460 2010 7580 2130
rect 7625 2010 7745 2130
rect 7800 2010 7920 2130
rect 7965 2010 8085 2130
rect 8130 2010 8250 2130
rect 8295 2010 8415 2130
rect 8470 2010 8590 2130
rect 8635 2010 8755 2130
rect 8800 2010 8920 2130
rect 8965 2010 9085 2130
rect 9140 2010 9260 2130
rect 9305 2010 9425 2130
rect 9470 2010 9590 2130
rect 9635 2010 9755 2130
rect 9810 2010 9930 2130
rect 9975 2010 10095 2130
rect 10140 2010 10260 2130
rect 10305 2010 10425 2130
rect 10480 2010 10600 2130
rect 10645 2010 10765 2130
rect 10810 2010 10930 2130
rect 10975 2010 11095 2130
rect 11150 2010 11270 2130
rect 11315 2010 11435 2130
rect 11480 2010 11600 2130
rect 11645 2010 11765 2130
rect 11820 2010 11940 2130
rect 11985 2010 12105 2130
rect 12150 2010 12270 2130
rect 12315 2010 12435 2130
rect 12490 2010 12610 2130
rect 7130 1845 7250 1965
rect 7295 1845 7415 1965
rect 7460 1845 7580 1965
rect 7625 1845 7745 1965
rect 7800 1845 7920 1965
rect 7965 1845 8085 1965
rect 8130 1845 8250 1965
rect 8295 1845 8415 1965
rect 8470 1845 8590 1965
rect 8635 1845 8755 1965
rect 8800 1845 8920 1965
rect 8965 1845 9085 1965
rect 9140 1845 9260 1965
rect 9305 1845 9425 1965
rect 9470 1845 9590 1965
rect 9635 1845 9755 1965
rect 9810 1845 9930 1965
rect 9975 1845 10095 1965
rect 10140 1845 10260 1965
rect 10305 1845 10425 1965
rect 10480 1845 10600 1965
rect 10645 1845 10765 1965
rect 10810 1845 10930 1965
rect 10975 1845 11095 1965
rect 11150 1845 11270 1965
rect 11315 1845 11435 1965
rect 11480 1845 11600 1965
rect 11645 1845 11765 1965
rect 11820 1845 11940 1965
rect 11985 1845 12105 1965
rect 12150 1845 12270 1965
rect 12315 1845 12435 1965
rect 12490 1845 12610 1965
rect 7130 1680 7250 1800
rect 7295 1680 7415 1800
rect 7460 1680 7580 1800
rect 7625 1680 7745 1800
rect 7800 1680 7920 1800
rect 7965 1680 8085 1800
rect 8130 1680 8250 1800
rect 8295 1680 8415 1800
rect 8470 1680 8590 1800
rect 8635 1680 8755 1800
rect 8800 1680 8920 1800
rect 8965 1680 9085 1800
rect 9140 1680 9260 1800
rect 9305 1680 9425 1800
rect 9470 1680 9590 1800
rect 9635 1680 9755 1800
rect 9810 1680 9930 1800
rect 9975 1680 10095 1800
rect 10140 1680 10260 1800
rect 10305 1680 10425 1800
rect 10480 1680 10600 1800
rect 10645 1680 10765 1800
rect 10810 1680 10930 1800
rect 10975 1680 11095 1800
rect 11150 1680 11270 1800
rect 11315 1680 11435 1800
rect 11480 1680 11600 1800
rect 11645 1680 11765 1800
rect 11820 1680 11940 1800
rect 11985 1680 12105 1800
rect 12150 1680 12270 1800
rect 12315 1680 12435 1800
rect 12490 1680 12610 1800
rect 12820 7040 12940 7160
rect 12985 7040 13105 7160
rect 13150 7040 13270 7160
rect 13315 7040 13435 7160
rect 13490 7040 13610 7160
rect 13655 7040 13775 7160
rect 13820 7040 13940 7160
rect 13985 7040 14105 7160
rect 14160 7040 14280 7160
rect 14325 7040 14445 7160
rect 14490 7040 14610 7160
rect 14655 7040 14775 7160
rect 14830 7040 14950 7160
rect 14995 7040 15115 7160
rect 15160 7040 15280 7160
rect 15325 7040 15445 7160
rect 15500 7040 15620 7160
rect 15665 7040 15785 7160
rect 15830 7040 15950 7160
rect 15995 7040 16115 7160
rect 16170 7040 16290 7160
rect 16335 7040 16455 7160
rect 16500 7040 16620 7160
rect 16665 7040 16785 7160
rect 16840 7040 16960 7160
rect 17005 7040 17125 7160
rect 17170 7040 17290 7160
rect 17335 7040 17455 7160
rect 17510 7040 17630 7160
rect 17675 7040 17795 7160
rect 17840 7040 17960 7160
rect 18005 7040 18125 7160
rect 18180 7040 18300 7160
rect 12820 6865 12940 6985
rect 12985 6865 13105 6985
rect 13150 6865 13270 6985
rect 13315 6865 13435 6985
rect 13490 6865 13610 6985
rect 13655 6865 13775 6985
rect 13820 6865 13940 6985
rect 13985 6865 14105 6985
rect 14160 6865 14280 6985
rect 14325 6865 14445 6985
rect 14490 6865 14610 6985
rect 14655 6865 14775 6985
rect 14830 6865 14950 6985
rect 14995 6865 15115 6985
rect 15160 6865 15280 6985
rect 15325 6865 15445 6985
rect 15500 6865 15620 6985
rect 15665 6865 15785 6985
rect 15830 6865 15950 6985
rect 15995 6865 16115 6985
rect 16170 6865 16290 6985
rect 16335 6865 16455 6985
rect 16500 6865 16620 6985
rect 16665 6865 16785 6985
rect 16840 6865 16960 6985
rect 17005 6865 17125 6985
rect 17170 6865 17290 6985
rect 17335 6865 17455 6985
rect 17510 6865 17630 6985
rect 17675 6865 17795 6985
rect 17840 6865 17960 6985
rect 18005 6865 18125 6985
rect 18180 6865 18300 6985
rect 12820 6700 12940 6820
rect 12985 6700 13105 6820
rect 13150 6700 13270 6820
rect 13315 6700 13435 6820
rect 13490 6700 13610 6820
rect 13655 6700 13775 6820
rect 13820 6700 13940 6820
rect 13985 6700 14105 6820
rect 14160 6700 14280 6820
rect 14325 6700 14445 6820
rect 14490 6700 14610 6820
rect 14655 6700 14775 6820
rect 14830 6700 14950 6820
rect 14995 6700 15115 6820
rect 15160 6700 15280 6820
rect 15325 6700 15445 6820
rect 15500 6700 15620 6820
rect 15665 6700 15785 6820
rect 15830 6700 15950 6820
rect 15995 6700 16115 6820
rect 16170 6700 16290 6820
rect 16335 6700 16455 6820
rect 16500 6700 16620 6820
rect 16665 6700 16785 6820
rect 16840 6700 16960 6820
rect 17005 6700 17125 6820
rect 17170 6700 17290 6820
rect 17335 6700 17455 6820
rect 17510 6700 17630 6820
rect 17675 6700 17795 6820
rect 17840 6700 17960 6820
rect 18005 6700 18125 6820
rect 18180 6700 18300 6820
rect 12820 6535 12940 6655
rect 12985 6535 13105 6655
rect 13150 6535 13270 6655
rect 13315 6535 13435 6655
rect 13490 6535 13610 6655
rect 13655 6535 13775 6655
rect 13820 6535 13940 6655
rect 13985 6535 14105 6655
rect 14160 6535 14280 6655
rect 14325 6535 14445 6655
rect 14490 6535 14610 6655
rect 14655 6535 14775 6655
rect 14830 6535 14950 6655
rect 14995 6535 15115 6655
rect 15160 6535 15280 6655
rect 15325 6535 15445 6655
rect 15500 6535 15620 6655
rect 15665 6535 15785 6655
rect 15830 6535 15950 6655
rect 15995 6535 16115 6655
rect 16170 6535 16290 6655
rect 16335 6535 16455 6655
rect 16500 6535 16620 6655
rect 16665 6535 16785 6655
rect 16840 6535 16960 6655
rect 17005 6535 17125 6655
rect 17170 6535 17290 6655
rect 17335 6535 17455 6655
rect 17510 6535 17630 6655
rect 17675 6535 17795 6655
rect 17840 6535 17960 6655
rect 18005 6535 18125 6655
rect 18180 6535 18300 6655
rect 12820 6370 12940 6490
rect 12985 6370 13105 6490
rect 13150 6370 13270 6490
rect 13315 6370 13435 6490
rect 13490 6370 13610 6490
rect 13655 6370 13775 6490
rect 13820 6370 13940 6490
rect 13985 6370 14105 6490
rect 14160 6370 14280 6490
rect 14325 6370 14445 6490
rect 14490 6370 14610 6490
rect 14655 6370 14775 6490
rect 14830 6370 14950 6490
rect 14995 6370 15115 6490
rect 15160 6370 15280 6490
rect 15325 6370 15445 6490
rect 15500 6370 15620 6490
rect 15665 6370 15785 6490
rect 15830 6370 15950 6490
rect 15995 6370 16115 6490
rect 16170 6370 16290 6490
rect 16335 6370 16455 6490
rect 16500 6370 16620 6490
rect 16665 6370 16785 6490
rect 16840 6370 16960 6490
rect 17005 6370 17125 6490
rect 17170 6370 17290 6490
rect 17335 6370 17455 6490
rect 17510 6370 17630 6490
rect 17675 6370 17795 6490
rect 17840 6370 17960 6490
rect 18005 6370 18125 6490
rect 18180 6370 18300 6490
rect 12820 6195 12940 6315
rect 12985 6195 13105 6315
rect 13150 6195 13270 6315
rect 13315 6195 13435 6315
rect 13490 6195 13610 6315
rect 13655 6195 13775 6315
rect 13820 6195 13940 6315
rect 13985 6195 14105 6315
rect 14160 6195 14280 6315
rect 14325 6195 14445 6315
rect 14490 6195 14610 6315
rect 14655 6195 14775 6315
rect 14830 6195 14950 6315
rect 14995 6195 15115 6315
rect 15160 6195 15280 6315
rect 15325 6195 15445 6315
rect 15500 6195 15620 6315
rect 15665 6195 15785 6315
rect 15830 6195 15950 6315
rect 15995 6195 16115 6315
rect 16170 6195 16290 6315
rect 16335 6195 16455 6315
rect 16500 6195 16620 6315
rect 16665 6195 16785 6315
rect 16840 6195 16960 6315
rect 17005 6195 17125 6315
rect 17170 6195 17290 6315
rect 17335 6195 17455 6315
rect 17510 6195 17630 6315
rect 17675 6195 17795 6315
rect 17840 6195 17960 6315
rect 18005 6195 18125 6315
rect 18180 6195 18300 6315
rect 12820 6030 12940 6150
rect 12985 6030 13105 6150
rect 13150 6030 13270 6150
rect 13315 6030 13435 6150
rect 13490 6030 13610 6150
rect 13655 6030 13775 6150
rect 13820 6030 13940 6150
rect 13985 6030 14105 6150
rect 14160 6030 14280 6150
rect 14325 6030 14445 6150
rect 14490 6030 14610 6150
rect 14655 6030 14775 6150
rect 14830 6030 14950 6150
rect 14995 6030 15115 6150
rect 15160 6030 15280 6150
rect 15325 6030 15445 6150
rect 15500 6030 15620 6150
rect 15665 6030 15785 6150
rect 15830 6030 15950 6150
rect 15995 6030 16115 6150
rect 16170 6030 16290 6150
rect 16335 6030 16455 6150
rect 16500 6030 16620 6150
rect 16665 6030 16785 6150
rect 16840 6030 16960 6150
rect 17005 6030 17125 6150
rect 17170 6030 17290 6150
rect 17335 6030 17455 6150
rect 17510 6030 17630 6150
rect 17675 6030 17795 6150
rect 17840 6030 17960 6150
rect 18005 6030 18125 6150
rect 18180 6030 18300 6150
rect 12820 5865 12940 5985
rect 12985 5865 13105 5985
rect 13150 5865 13270 5985
rect 13315 5865 13435 5985
rect 13490 5865 13610 5985
rect 13655 5865 13775 5985
rect 13820 5865 13940 5985
rect 13985 5865 14105 5985
rect 14160 5865 14280 5985
rect 14325 5865 14445 5985
rect 14490 5865 14610 5985
rect 14655 5865 14775 5985
rect 14830 5865 14950 5985
rect 14995 5865 15115 5985
rect 15160 5865 15280 5985
rect 15325 5865 15445 5985
rect 15500 5865 15620 5985
rect 15665 5865 15785 5985
rect 15830 5865 15950 5985
rect 15995 5865 16115 5985
rect 16170 5865 16290 5985
rect 16335 5865 16455 5985
rect 16500 5865 16620 5985
rect 16665 5865 16785 5985
rect 16840 5865 16960 5985
rect 17005 5865 17125 5985
rect 17170 5865 17290 5985
rect 17335 5865 17455 5985
rect 17510 5865 17630 5985
rect 17675 5865 17795 5985
rect 17840 5865 17960 5985
rect 18005 5865 18125 5985
rect 18180 5865 18300 5985
rect 12820 5700 12940 5820
rect 12985 5700 13105 5820
rect 13150 5700 13270 5820
rect 13315 5700 13435 5820
rect 13490 5700 13610 5820
rect 13655 5700 13775 5820
rect 13820 5700 13940 5820
rect 13985 5700 14105 5820
rect 14160 5700 14280 5820
rect 14325 5700 14445 5820
rect 14490 5700 14610 5820
rect 14655 5700 14775 5820
rect 14830 5700 14950 5820
rect 14995 5700 15115 5820
rect 15160 5700 15280 5820
rect 15325 5700 15445 5820
rect 15500 5700 15620 5820
rect 15665 5700 15785 5820
rect 15830 5700 15950 5820
rect 15995 5700 16115 5820
rect 16170 5700 16290 5820
rect 16335 5700 16455 5820
rect 16500 5700 16620 5820
rect 16665 5700 16785 5820
rect 16840 5700 16960 5820
rect 17005 5700 17125 5820
rect 17170 5700 17290 5820
rect 17335 5700 17455 5820
rect 17510 5700 17630 5820
rect 17675 5700 17795 5820
rect 17840 5700 17960 5820
rect 18005 5700 18125 5820
rect 18180 5700 18300 5820
rect 12820 5525 12940 5645
rect 12985 5525 13105 5645
rect 13150 5525 13270 5645
rect 13315 5525 13435 5645
rect 13490 5525 13610 5645
rect 13655 5525 13775 5645
rect 13820 5525 13940 5645
rect 13985 5525 14105 5645
rect 14160 5525 14280 5645
rect 14325 5525 14445 5645
rect 14490 5525 14610 5645
rect 14655 5525 14775 5645
rect 14830 5525 14950 5645
rect 14995 5525 15115 5645
rect 15160 5525 15280 5645
rect 15325 5525 15445 5645
rect 15500 5525 15620 5645
rect 15665 5525 15785 5645
rect 15830 5525 15950 5645
rect 15995 5525 16115 5645
rect 16170 5525 16290 5645
rect 16335 5525 16455 5645
rect 16500 5525 16620 5645
rect 16665 5525 16785 5645
rect 16840 5525 16960 5645
rect 17005 5525 17125 5645
rect 17170 5525 17290 5645
rect 17335 5525 17455 5645
rect 17510 5525 17630 5645
rect 17675 5525 17795 5645
rect 17840 5525 17960 5645
rect 18005 5525 18125 5645
rect 18180 5525 18300 5645
rect 12820 5360 12940 5480
rect 12985 5360 13105 5480
rect 13150 5360 13270 5480
rect 13315 5360 13435 5480
rect 13490 5360 13610 5480
rect 13655 5360 13775 5480
rect 13820 5360 13940 5480
rect 13985 5360 14105 5480
rect 14160 5360 14280 5480
rect 14325 5360 14445 5480
rect 14490 5360 14610 5480
rect 14655 5360 14775 5480
rect 14830 5360 14950 5480
rect 14995 5360 15115 5480
rect 15160 5360 15280 5480
rect 15325 5360 15445 5480
rect 15500 5360 15620 5480
rect 15665 5360 15785 5480
rect 15830 5360 15950 5480
rect 15995 5360 16115 5480
rect 16170 5360 16290 5480
rect 16335 5360 16455 5480
rect 16500 5360 16620 5480
rect 16665 5360 16785 5480
rect 16840 5360 16960 5480
rect 17005 5360 17125 5480
rect 17170 5360 17290 5480
rect 17335 5360 17455 5480
rect 17510 5360 17630 5480
rect 17675 5360 17795 5480
rect 17840 5360 17960 5480
rect 18005 5360 18125 5480
rect 18180 5360 18300 5480
rect 12820 5195 12940 5315
rect 12985 5195 13105 5315
rect 13150 5195 13270 5315
rect 13315 5195 13435 5315
rect 13490 5195 13610 5315
rect 13655 5195 13775 5315
rect 13820 5195 13940 5315
rect 13985 5195 14105 5315
rect 14160 5195 14280 5315
rect 14325 5195 14445 5315
rect 14490 5195 14610 5315
rect 14655 5195 14775 5315
rect 14830 5195 14950 5315
rect 14995 5195 15115 5315
rect 15160 5195 15280 5315
rect 15325 5195 15445 5315
rect 15500 5195 15620 5315
rect 15665 5195 15785 5315
rect 15830 5195 15950 5315
rect 15995 5195 16115 5315
rect 16170 5195 16290 5315
rect 16335 5195 16455 5315
rect 16500 5195 16620 5315
rect 16665 5195 16785 5315
rect 16840 5195 16960 5315
rect 17005 5195 17125 5315
rect 17170 5195 17290 5315
rect 17335 5195 17455 5315
rect 17510 5195 17630 5315
rect 17675 5195 17795 5315
rect 17840 5195 17960 5315
rect 18005 5195 18125 5315
rect 18180 5195 18300 5315
rect 12820 5030 12940 5150
rect 12985 5030 13105 5150
rect 13150 5030 13270 5150
rect 13315 5030 13435 5150
rect 13490 5030 13610 5150
rect 13655 5030 13775 5150
rect 13820 5030 13940 5150
rect 13985 5030 14105 5150
rect 14160 5030 14280 5150
rect 14325 5030 14445 5150
rect 14490 5030 14610 5150
rect 14655 5030 14775 5150
rect 14830 5030 14950 5150
rect 14995 5030 15115 5150
rect 15160 5030 15280 5150
rect 15325 5030 15445 5150
rect 15500 5030 15620 5150
rect 15665 5030 15785 5150
rect 15830 5030 15950 5150
rect 15995 5030 16115 5150
rect 16170 5030 16290 5150
rect 16335 5030 16455 5150
rect 16500 5030 16620 5150
rect 16665 5030 16785 5150
rect 16840 5030 16960 5150
rect 17005 5030 17125 5150
rect 17170 5030 17290 5150
rect 17335 5030 17455 5150
rect 17510 5030 17630 5150
rect 17675 5030 17795 5150
rect 17840 5030 17960 5150
rect 18005 5030 18125 5150
rect 18180 5030 18300 5150
rect 12820 4855 12940 4975
rect 12985 4855 13105 4975
rect 13150 4855 13270 4975
rect 13315 4855 13435 4975
rect 13490 4855 13610 4975
rect 13655 4855 13775 4975
rect 13820 4855 13940 4975
rect 13985 4855 14105 4975
rect 14160 4855 14280 4975
rect 14325 4855 14445 4975
rect 14490 4855 14610 4975
rect 14655 4855 14775 4975
rect 14830 4855 14950 4975
rect 14995 4855 15115 4975
rect 15160 4855 15280 4975
rect 15325 4855 15445 4975
rect 15500 4855 15620 4975
rect 15665 4855 15785 4975
rect 15830 4855 15950 4975
rect 15995 4855 16115 4975
rect 16170 4855 16290 4975
rect 16335 4855 16455 4975
rect 16500 4855 16620 4975
rect 16665 4855 16785 4975
rect 16840 4855 16960 4975
rect 17005 4855 17125 4975
rect 17170 4855 17290 4975
rect 17335 4855 17455 4975
rect 17510 4855 17630 4975
rect 17675 4855 17795 4975
rect 17840 4855 17960 4975
rect 18005 4855 18125 4975
rect 18180 4855 18300 4975
rect 12820 4690 12940 4810
rect 12985 4690 13105 4810
rect 13150 4690 13270 4810
rect 13315 4690 13435 4810
rect 13490 4690 13610 4810
rect 13655 4690 13775 4810
rect 13820 4690 13940 4810
rect 13985 4690 14105 4810
rect 14160 4690 14280 4810
rect 14325 4690 14445 4810
rect 14490 4690 14610 4810
rect 14655 4690 14775 4810
rect 14830 4690 14950 4810
rect 14995 4690 15115 4810
rect 15160 4690 15280 4810
rect 15325 4690 15445 4810
rect 15500 4690 15620 4810
rect 15665 4690 15785 4810
rect 15830 4690 15950 4810
rect 15995 4690 16115 4810
rect 16170 4690 16290 4810
rect 16335 4690 16455 4810
rect 16500 4690 16620 4810
rect 16665 4690 16785 4810
rect 16840 4690 16960 4810
rect 17005 4690 17125 4810
rect 17170 4690 17290 4810
rect 17335 4690 17455 4810
rect 17510 4690 17630 4810
rect 17675 4690 17795 4810
rect 17840 4690 17960 4810
rect 18005 4690 18125 4810
rect 18180 4690 18300 4810
rect 12820 4525 12940 4645
rect 12985 4525 13105 4645
rect 13150 4525 13270 4645
rect 13315 4525 13435 4645
rect 13490 4525 13610 4645
rect 13655 4525 13775 4645
rect 13820 4525 13940 4645
rect 13985 4525 14105 4645
rect 14160 4525 14280 4645
rect 14325 4525 14445 4645
rect 14490 4525 14610 4645
rect 14655 4525 14775 4645
rect 14830 4525 14950 4645
rect 14995 4525 15115 4645
rect 15160 4525 15280 4645
rect 15325 4525 15445 4645
rect 15500 4525 15620 4645
rect 15665 4525 15785 4645
rect 15830 4525 15950 4645
rect 15995 4525 16115 4645
rect 16170 4525 16290 4645
rect 16335 4525 16455 4645
rect 16500 4525 16620 4645
rect 16665 4525 16785 4645
rect 16840 4525 16960 4645
rect 17005 4525 17125 4645
rect 17170 4525 17290 4645
rect 17335 4525 17455 4645
rect 17510 4525 17630 4645
rect 17675 4525 17795 4645
rect 17840 4525 17960 4645
rect 18005 4525 18125 4645
rect 18180 4525 18300 4645
rect 12820 4360 12940 4480
rect 12985 4360 13105 4480
rect 13150 4360 13270 4480
rect 13315 4360 13435 4480
rect 13490 4360 13610 4480
rect 13655 4360 13775 4480
rect 13820 4360 13940 4480
rect 13985 4360 14105 4480
rect 14160 4360 14280 4480
rect 14325 4360 14445 4480
rect 14490 4360 14610 4480
rect 14655 4360 14775 4480
rect 14830 4360 14950 4480
rect 14995 4360 15115 4480
rect 15160 4360 15280 4480
rect 15325 4360 15445 4480
rect 15500 4360 15620 4480
rect 15665 4360 15785 4480
rect 15830 4360 15950 4480
rect 15995 4360 16115 4480
rect 16170 4360 16290 4480
rect 16335 4360 16455 4480
rect 16500 4360 16620 4480
rect 16665 4360 16785 4480
rect 16840 4360 16960 4480
rect 17005 4360 17125 4480
rect 17170 4360 17290 4480
rect 17335 4360 17455 4480
rect 17510 4360 17630 4480
rect 17675 4360 17795 4480
rect 17840 4360 17960 4480
rect 18005 4360 18125 4480
rect 18180 4360 18300 4480
rect 12820 4185 12940 4305
rect 12985 4185 13105 4305
rect 13150 4185 13270 4305
rect 13315 4185 13435 4305
rect 13490 4185 13610 4305
rect 13655 4185 13775 4305
rect 13820 4185 13940 4305
rect 13985 4185 14105 4305
rect 14160 4185 14280 4305
rect 14325 4185 14445 4305
rect 14490 4185 14610 4305
rect 14655 4185 14775 4305
rect 14830 4185 14950 4305
rect 14995 4185 15115 4305
rect 15160 4185 15280 4305
rect 15325 4185 15445 4305
rect 15500 4185 15620 4305
rect 15665 4185 15785 4305
rect 15830 4185 15950 4305
rect 15995 4185 16115 4305
rect 16170 4185 16290 4305
rect 16335 4185 16455 4305
rect 16500 4185 16620 4305
rect 16665 4185 16785 4305
rect 16840 4185 16960 4305
rect 17005 4185 17125 4305
rect 17170 4185 17290 4305
rect 17335 4185 17455 4305
rect 17510 4185 17630 4305
rect 17675 4185 17795 4305
rect 17840 4185 17960 4305
rect 18005 4185 18125 4305
rect 18180 4185 18300 4305
rect 12820 4020 12940 4140
rect 12985 4020 13105 4140
rect 13150 4020 13270 4140
rect 13315 4020 13435 4140
rect 13490 4020 13610 4140
rect 13655 4020 13775 4140
rect 13820 4020 13940 4140
rect 13985 4020 14105 4140
rect 14160 4020 14280 4140
rect 14325 4020 14445 4140
rect 14490 4020 14610 4140
rect 14655 4020 14775 4140
rect 14830 4020 14950 4140
rect 14995 4020 15115 4140
rect 15160 4020 15280 4140
rect 15325 4020 15445 4140
rect 15500 4020 15620 4140
rect 15665 4020 15785 4140
rect 15830 4020 15950 4140
rect 15995 4020 16115 4140
rect 16170 4020 16290 4140
rect 16335 4020 16455 4140
rect 16500 4020 16620 4140
rect 16665 4020 16785 4140
rect 16840 4020 16960 4140
rect 17005 4020 17125 4140
rect 17170 4020 17290 4140
rect 17335 4020 17455 4140
rect 17510 4020 17630 4140
rect 17675 4020 17795 4140
rect 17840 4020 17960 4140
rect 18005 4020 18125 4140
rect 18180 4020 18300 4140
rect 12820 3855 12940 3975
rect 12985 3855 13105 3975
rect 13150 3855 13270 3975
rect 13315 3855 13435 3975
rect 13490 3855 13610 3975
rect 13655 3855 13775 3975
rect 13820 3855 13940 3975
rect 13985 3855 14105 3975
rect 14160 3855 14280 3975
rect 14325 3855 14445 3975
rect 14490 3855 14610 3975
rect 14655 3855 14775 3975
rect 14830 3855 14950 3975
rect 14995 3855 15115 3975
rect 15160 3855 15280 3975
rect 15325 3855 15445 3975
rect 15500 3855 15620 3975
rect 15665 3855 15785 3975
rect 15830 3855 15950 3975
rect 15995 3855 16115 3975
rect 16170 3855 16290 3975
rect 16335 3855 16455 3975
rect 16500 3855 16620 3975
rect 16665 3855 16785 3975
rect 16840 3855 16960 3975
rect 17005 3855 17125 3975
rect 17170 3855 17290 3975
rect 17335 3855 17455 3975
rect 17510 3855 17630 3975
rect 17675 3855 17795 3975
rect 17840 3855 17960 3975
rect 18005 3855 18125 3975
rect 18180 3855 18300 3975
rect 12820 3690 12940 3810
rect 12985 3690 13105 3810
rect 13150 3690 13270 3810
rect 13315 3690 13435 3810
rect 13490 3690 13610 3810
rect 13655 3690 13775 3810
rect 13820 3690 13940 3810
rect 13985 3690 14105 3810
rect 14160 3690 14280 3810
rect 14325 3690 14445 3810
rect 14490 3690 14610 3810
rect 14655 3690 14775 3810
rect 14830 3690 14950 3810
rect 14995 3690 15115 3810
rect 15160 3690 15280 3810
rect 15325 3690 15445 3810
rect 15500 3690 15620 3810
rect 15665 3690 15785 3810
rect 15830 3690 15950 3810
rect 15995 3690 16115 3810
rect 16170 3690 16290 3810
rect 16335 3690 16455 3810
rect 16500 3690 16620 3810
rect 16665 3690 16785 3810
rect 16840 3690 16960 3810
rect 17005 3690 17125 3810
rect 17170 3690 17290 3810
rect 17335 3690 17455 3810
rect 17510 3690 17630 3810
rect 17675 3690 17795 3810
rect 17840 3690 17960 3810
rect 18005 3690 18125 3810
rect 18180 3690 18300 3810
rect 12820 3515 12940 3635
rect 12985 3515 13105 3635
rect 13150 3515 13270 3635
rect 13315 3515 13435 3635
rect 13490 3515 13610 3635
rect 13655 3515 13775 3635
rect 13820 3515 13940 3635
rect 13985 3515 14105 3635
rect 14160 3515 14280 3635
rect 14325 3515 14445 3635
rect 14490 3515 14610 3635
rect 14655 3515 14775 3635
rect 14830 3515 14950 3635
rect 14995 3515 15115 3635
rect 15160 3515 15280 3635
rect 15325 3515 15445 3635
rect 15500 3515 15620 3635
rect 15665 3515 15785 3635
rect 15830 3515 15950 3635
rect 15995 3515 16115 3635
rect 16170 3515 16290 3635
rect 16335 3515 16455 3635
rect 16500 3515 16620 3635
rect 16665 3515 16785 3635
rect 16840 3515 16960 3635
rect 17005 3515 17125 3635
rect 17170 3515 17290 3635
rect 17335 3515 17455 3635
rect 17510 3515 17630 3635
rect 17675 3515 17795 3635
rect 17840 3515 17960 3635
rect 18005 3515 18125 3635
rect 18180 3515 18300 3635
rect 12820 3350 12940 3470
rect 12985 3350 13105 3470
rect 13150 3350 13270 3470
rect 13315 3350 13435 3470
rect 13490 3350 13610 3470
rect 13655 3350 13775 3470
rect 13820 3350 13940 3470
rect 13985 3350 14105 3470
rect 14160 3350 14280 3470
rect 14325 3350 14445 3470
rect 14490 3350 14610 3470
rect 14655 3350 14775 3470
rect 14830 3350 14950 3470
rect 14995 3350 15115 3470
rect 15160 3350 15280 3470
rect 15325 3350 15445 3470
rect 15500 3350 15620 3470
rect 15665 3350 15785 3470
rect 15830 3350 15950 3470
rect 15995 3350 16115 3470
rect 16170 3350 16290 3470
rect 16335 3350 16455 3470
rect 16500 3350 16620 3470
rect 16665 3350 16785 3470
rect 16840 3350 16960 3470
rect 17005 3350 17125 3470
rect 17170 3350 17290 3470
rect 17335 3350 17455 3470
rect 17510 3350 17630 3470
rect 17675 3350 17795 3470
rect 17840 3350 17960 3470
rect 18005 3350 18125 3470
rect 18180 3350 18300 3470
rect 12820 3185 12940 3305
rect 12985 3185 13105 3305
rect 13150 3185 13270 3305
rect 13315 3185 13435 3305
rect 13490 3185 13610 3305
rect 13655 3185 13775 3305
rect 13820 3185 13940 3305
rect 13985 3185 14105 3305
rect 14160 3185 14280 3305
rect 14325 3185 14445 3305
rect 14490 3185 14610 3305
rect 14655 3185 14775 3305
rect 14830 3185 14950 3305
rect 14995 3185 15115 3305
rect 15160 3185 15280 3305
rect 15325 3185 15445 3305
rect 15500 3185 15620 3305
rect 15665 3185 15785 3305
rect 15830 3185 15950 3305
rect 15995 3185 16115 3305
rect 16170 3185 16290 3305
rect 16335 3185 16455 3305
rect 16500 3185 16620 3305
rect 16665 3185 16785 3305
rect 16840 3185 16960 3305
rect 17005 3185 17125 3305
rect 17170 3185 17290 3305
rect 17335 3185 17455 3305
rect 17510 3185 17630 3305
rect 17675 3185 17795 3305
rect 17840 3185 17960 3305
rect 18005 3185 18125 3305
rect 18180 3185 18300 3305
rect 12820 3020 12940 3140
rect 12985 3020 13105 3140
rect 13150 3020 13270 3140
rect 13315 3020 13435 3140
rect 13490 3020 13610 3140
rect 13655 3020 13775 3140
rect 13820 3020 13940 3140
rect 13985 3020 14105 3140
rect 14160 3020 14280 3140
rect 14325 3020 14445 3140
rect 14490 3020 14610 3140
rect 14655 3020 14775 3140
rect 14830 3020 14950 3140
rect 14995 3020 15115 3140
rect 15160 3020 15280 3140
rect 15325 3020 15445 3140
rect 15500 3020 15620 3140
rect 15665 3020 15785 3140
rect 15830 3020 15950 3140
rect 15995 3020 16115 3140
rect 16170 3020 16290 3140
rect 16335 3020 16455 3140
rect 16500 3020 16620 3140
rect 16665 3020 16785 3140
rect 16840 3020 16960 3140
rect 17005 3020 17125 3140
rect 17170 3020 17290 3140
rect 17335 3020 17455 3140
rect 17510 3020 17630 3140
rect 17675 3020 17795 3140
rect 17840 3020 17960 3140
rect 18005 3020 18125 3140
rect 18180 3020 18300 3140
rect 12820 2845 12940 2965
rect 12985 2845 13105 2965
rect 13150 2845 13270 2965
rect 13315 2845 13435 2965
rect 13490 2845 13610 2965
rect 13655 2845 13775 2965
rect 13820 2845 13940 2965
rect 13985 2845 14105 2965
rect 14160 2845 14280 2965
rect 14325 2845 14445 2965
rect 14490 2845 14610 2965
rect 14655 2845 14775 2965
rect 14830 2845 14950 2965
rect 14995 2845 15115 2965
rect 15160 2845 15280 2965
rect 15325 2845 15445 2965
rect 15500 2845 15620 2965
rect 15665 2845 15785 2965
rect 15830 2845 15950 2965
rect 15995 2845 16115 2965
rect 16170 2845 16290 2965
rect 16335 2845 16455 2965
rect 16500 2845 16620 2965
rect 16665 2845 16785 2965
rect 16840 2845 16960 2965
rect 17005 2845 17125 2965
rect 17170 2845 17290 2965
rect 17335 2845 17455 2965
rect 17510 2845 17630 2965
rect 17675 2845 17795 2965
rect 17840 2845 17960 2965
rect 18005 2845 18125 2965
rect 18180 2845 18300 2965
rect 12820 2680 12940 2800
rect 12985 2680 13105 2800
rect 13150 2680 13270 2800
rect 13315 2680 13435 2800
rect 13490 2680 13610 2800
rect 13655 2680 13775 2800
rect 13820 2680 13940 2800
rect 13985 2680 14105 2800
rect 14160 2680 14280 2800
rect 14325 2680 14445 2800
rect 14490 2680 14610 2800
rect 14655 2680 14775 2800
rect 14830 2680 14950 2800
rect 14995 2680 15115 2800
rect 15160 2680 15280 2800
rect 15325 2680 15445 2800
rect 15500 2680 15620 2800
rect 15665 2680 15785 2800
rect 15830 2680 15950 2800
rect 15995 2680 16115 2800
rect 16170 2680 16290 2800
rect 16335 2680 16455 2800
rect 16500 2680 16620 2800
rect 16665 2680 16785 2800
rect 16840 2680 16960 2800
rect 17005 2680 17125 2800
rect 17170 2680 17290 2800
rect 17335 2680 17455 2800
rect 17510 2680 17630 2800
rect 17675 2680 17795 2800
rect 17840 2680 17960 2800
rect 18005 2680 18125 2800
rect 18180 2680 18300 2800
rect 12820 2515 12940 2635
rect 12985 2515 13105 2635
rect 13150 2515 13270 2635
rect 13315 2515 13435 2635
rect 13490 2515 13610 2635
rect 13655 2515 13775 2635
rect 13820 2515 13940 2635
rect 13985 2515 14105 2635
rect 14160 2515 14280 2635
rect 14325 2515 14445 2635
rect 14490 2515 14610 2635
rect 14655 2515 14775 2635
rect 14830 2515 14950 2635
rect 14995 2515 15115 2635
rect 15160 2515 15280 2635
rect 15325 2515 15445 2635
rect 15500 2515 15620 2635
rect 15665 2515 15785 2635
rect 15830 2515 15950 2635
rect 15995 2515 16115 2635
rect 16170 2515 16290 2635
rect 16335 2515 16455 2635
rect 16500 2515 16620 2635
rect 16665 2515 16785 2635
rect 16840 2515 16960 2635
rect 17005 2515 17125 2635
rect 17170 2515 17290 2635
rect 17335 2515 17455 2635
rect 17510 2515 17630 2635
rect 17675 2515 17795 2635
rect 17840 2515 17960 2635
rect 18005 2515 18125 2635
rect 18180 2515 18300 2635
rect 12820 2350 12940 2470
rect 12985 2350 13105 2470
rect 13150 2350 13270 2470
rect 13315 2350 13435 2470
rect 13490 2350 13610 2470
rect 13655 2350 13775 2470
rect 13820 2350 13940 2470
rect 13985 2350 14105 2470
rect 14160 2350 14280 2470
rect 14325 2350 14445 2470
rect 14490 2350 14610 2470
rect 14655 2350 14775 2470
rect 14830 2350 14950 2470
rect 14995 2350 15115 2470
rect 15160 2350 15280 2470
rect 15325 2350 15445 2470
rect 15500 2350 15620 2470
rect 15665 2350 15785 2470
rect 15830 2350 15950 2470
rect 15995 2350 16115 2470
rect 16170 2350 16290 2470
rect 16335 2350 16455 2470
rect 16500 2350 16620 2470
rect 16665 2350 16785 2470
rect 16840 2350 16960 2470
rect 17005 2350 17125 2470
rect 17170 2350 17290 2470
rect 17335 2350 17455 2470
rect 17510 2350 17630 2470
rect 17675 2350 17795 2470
rect 17840 2350 17960 2470
rect 18005 2350 18125 2470
rect 18180 2350 18300 2470
rect 12820 2175 12940 2295
rect 12985 2175 13105 2295
rect 13150 2175 13270 2295
rect 13315 2175 13435 2295
rect 13490 2175 13610 2295
rect 13655 2175 13775 2295
rect 13820 2175 13940 2295
rect 13985 2175 14105 2295
rect 14160 2175 14280 2295
rect 14325 2175 14445 2295
rect 14490 2175 14610 2295
rect 14655 2175 14775 2295
rect 14830 2175 14950 2295
rect 14995 2175 15115 2295
rect 15160 2175 15280 2295
rect 15325 2175 15445 2295
rect 15500 2175 15620 2295
rect 15665 2175 15785 2295
rect 15830 2175 15950 2295
rect 15995 2175 16115 2295
rect 16170 2175 16290 2295
rect 16335 2175 16455 2295
rect 16500 2175 16620 2295
rect 16665 2175 16785 2295
rect 16840 2175 16960 2295
rect 17005 2175 17125 2295
rect 17170 2175 17290 2295
rect 17335 2175 17455 2295
rect 17510 2175 17630 2295
rect 17675 2175 17795 2295
rect 17840 2175 17960 2295
rect 18005 2175 18125 2295
rect 18180 2175 18300 2295
rect 12820 2010 12940 2130
rect 12985 2010 13105 2130
rect 13150 2010 13270 2130
rect 13315 2010 13435 2130
rect 13490 2010 13610 2130
rect 13655 2010 13775 2130
rect 13820 2010 13940 2130
rect 13985 2010 14105 2130
rect 14160 2010 14280 2130
rect 14325 2010 14445 2130
rect 14490 2010 14610 2130
rect 14655 2010 14775 2130
rect 14830 2010 14950 2130
rect 14995 2010 15115 2130
rect 15160 2010 15280 2130
rect 15325 2010 15445 2130
rect 15500 2010 15620 2130
rect 15665 2010 15785 2130
rect 15830 2010 15950 2130
rect 15995 2010 16115 2130
rect 16170 2010 16290 2130
rect 16335 2010 16455 2130
rect 16500 2010 16620 2130
rect 16665 2010 16785 2130
rect 16840 2010 16960 2130
rect 17005 2010 17125 2130
rect 17170 2010 17290 2130
rect 17335 2010 17455 2130
rect 17510 2010 17630 2130
rect 17675 2010 17795 2130
rect 17840 2010 17960 2130
rect 18005 2010 18125 2130
rect 18180 2010 18300 2130
rect 12820 1845 12940 1965
rect 12985 1845 13105 1965
rect 13150 1845 13270 1965
rect 13315 1845 13435 1965
rect 13490 1845 13610 1965
rect 13655 1845 13775 1965
rect 13820 1845 13940 1965
rect 13985 1845 14105 1965
rect 14160 1845 14280 1965
rect 14325 1845 14445 1965
rect 14490 1845 14610 1965
rect 14655 1845 14775 1965
rect 14830 1845 14950 1965
rect 14995 1845 15115 1965
rect 15160 1845 15280 1965
rect 15325 1845 15445 1965
rect 15500 1845 15620 1965
rect 15665 1845 15785 1965
rect 15830 1845 15950 1965
rect 15995 1845 16115 1965
rect 16170 1845 16290 1965
rect 16335 1845 16455 1965
rect 16500 1845 16620 1965
rect 16665 1845 16785 1965
rect 16840 1845 16960 1965
rect 17005 1845 17125 1965
rect 17170 1845 17290 1965
rect 17335 1845 17455 1965
rect 17510 1845 17630 1965
rect 17675 1845 17795 1965
rect 17840 1845 17960 1965
rect 18005 1845 18125 1965
rect 18180 1845 18300 1965
rect 12820 1680 12940 1800
rect 12985 1680 13105 1800
rect 13150 1680 13270 1800
rect 13315 1680 13435 1800
rect 13490 1680 13610 1800
rect 13655 1680 13775 1800
rect 13820 1680 13940 1800
rect 13985 1680 14105 1800
rect 14160 1680 14280 1800
rect 14325 1680 14445 1800
rect 14490 1680 14610 1800
rect 14655 1680 14775 1800
rect 14830 1680 14950 1800
rect 14995 1680 15115 1800
rect 15160 1680 15280 1800
rect 15325 1680 15445 1800
rect 15500 1680 15620 1800
rect 15665 1680 15785 1800
rect 15830 1680 15950 1800
rect 15995 1680 16115 1800
rect 16170 1680 16290 1800
rect 16335 1680 16455 1800
rect 16500 1680 16620 1800
rect 16665 1680 16785 1800
rect 16840 1680 16960 1800
rect 17005 1680 17125 1800
rect 17170 1680 17290 1800
rect 17335 1680 17455 1800
rect 17510 1680 17630 1800
rect 17675 1680 17795 1800
rect 17840 1680 17960 1800
rect 18005 1680 18125 1800
rect 18180 1680 18300 1800
rect 18510 7040 18630 7160
rect 18675 7040 18795 7160
rect 18840 7040 18960 7160
rect 19005 7040 19125 7160
rect 19180 7040 19300 7160
rect 19345 7040 19465 7160
rect 19510 7040 19630 7160
rect 19675 7040 19795 7160
rect 19850 7040 19970 7160
rect 20015 7040 20135 7160
rect 20180 7040 20300 7160
rect 20345 7040 20465 7160
rect 20520 7040 20640 7160
rect 20685 7040 20805 7160
rect 20850 7040 20970 7160
rect 21015 7040 21135 7160
rect 21190 7040 21310 7160
rect 21355 7040 21475 7160
rect 21520 7040 21640 7160
rect 21685 7040 21805 7160
rect 21860 7040 21980 7160
rect 22025 7040 22145 7160
rect 22190 7040 22310 7160
rect 22355 7040 22475 7160
rect 22530 7040 22650 7160
rect 22695 7040 22815 7160
rect 22860 7040 22980 7160
rect 23025 7040 23145 7160
rect 23200 7040 23320 7160
rect 23365 7040 23485 7160
rect 23530 7040 23650 7160
rect 23695 7040 23815 7160
rect 23870 7040 23990 7160
rect 18510 6865 18630 6985
rect 18675 6865 18795 6985
rect 18840 6865 18960 6985
rect 19005 6865 19125 6985
rect 19180 6865 19300 6985
rect 19345 6865 19465 6985
rect 19510 6865 19630 6985
rect 19675 6865 19795 6985
rect 19850 6865 19970 6985
rect 20015 6865 20135 6985
rect 20180 6865 20300 6985
rect 20345 6865 20465 6985
rect 20520 6865 20640 6985
rect 20685 6865 20805 6985
rect 20850 6865 20970 6985
rect 21015 6865 21135 6985
rect 21190 6865 21310 6985
rect 21355 6865 21475 6985
rect 21520 6865 21640 6985
rect 21685 6865 21805 6985
rect 21860 6865 21980 6985
rect 22025 6865 22145 6985
rect 22190 6865 22310 6985
rect 22355 6865 22475 6985
rect 22530 6865 22650 6985
rect 22695 6865 22815 6985
rect 22860 6865 22980 6985
rect 23025 6865 23145 6985
rect 23200 6865 23320 6985
rect 23365 6865 23485 6985
rect 23530 6865 23650 6985
rect 23695 6865 23815 6985
rect 23870 6865 23990 6985
rect 18510 6700 18630 6820
rect 18675 6700 18795 6820
rect 18840 6700 18960 6820
rect 19005 6700 19125 6820
rect 19180 6700 19300 6820
rect 19345 6700 19465 6820
rect 19510 6700 19630 6820
rect 19675 6700 19795 6820
rect 19850 6700 19970 6820
rect 20015 6700 20135 6820
rect 20180 6700 20300 6820
rect 20345 6700 20465 6820
rect 20520 6700 20640 6820
rect 20685 6700 20805 6820
rect 20850 6700 20970 6820
rect 21015 6700 21135 6820
rect 21190 6700 21310 6820
rect 21355 6700 21475 6820
rect 21520 6700 21640 6820
rect 21685 6700 21805 6820
rect 21860 6700 21980 6820
rect 22025 6700 22145 6820
rect 22190 6700 22310 6820
rect 22355 6700 22475 6820
rect 22530 6700 22650 6820
rect 22695 6700 22815 6820
rect 22860 6700 22980 6820
rect 23025 6700 23145 6820
rect 23200 6700 23320 6820
rect 23365 6700 23485 6820
rect 23530 6700 23650 6820
rect 23695 6700 23815 6820
rect 23870 6700 23990 6820
rect 18510 6535 18630 6655
rect 18675 6535 18795 6655
rect 18840 6535 18960 6655
rect 19005 6535 19125 6655
rect 19180 6535 19300 6655
rect 19345 6535 19465 6655
rect 19510 6535 19630 6655
rect 19675 6535 19795 6655
rect 19850 6535 19970 6655
rect 20015 6535 20135 6655
rect 20180 6535 20300 6655
rect 20345 6535 20465 6655
rect 20520 6535 20640 6655
rect 20685 6535 20805 6655
rect 20850 6535 20970 6655
rect 21015 6535 21135 6655
rect 21190 6535 21310 6655
rect 21355 6535 21475 6655
rect 21520 6535 21640 6655
rect 21685 6535 21805 6655
rect 21860 6535 21980 6655
rect 22025 6535 22145 6655
rect 22190 6535 22310 6655
rect 22355 6535 22475 6655
rect 22530 6535 22650 6655
rect 22695 6535 22815 6655
rect 22860 6535 22980 6655
rect 23025 6535 23145 6655
rect 23200 6535 23320 6655
rect 23365 6535 23485 6655
rect 23530 6535 23650 6655
rect 23695 6535 23815 6655
rect 23870 6535 23990 6655
rect 18510 6370 18630 6490
rect 18675 6370 18795 6490
rect 18840 6370 18960 6490
rect 19005 6370 19125 6490
rect 19180 6370 19300 6490
rect 19345 6370 19465 6490
rect 19510 6370 19630 6490
rect 19675 6370 19795 6490
rect 19850 6370 19970 6490
rect 20015 6370 20135 6490
rect 20180 6370 20300 6490
rect 20345 6370 20465 6490
rect 20520 6370 20640 6490
rect 20685 6370 20805 6490
rect 20850 6370 20970 6490
rect 21015 6370 21135 6490
rect 21190 6370 21310 6490
rect 21355 6370 21475 6490
rect 21520 6370 21640 6490
rect 21685 6370 21805 6490
rect 21860 6370 21980 6490
rect 22025 6370 22145 6490
rect 22190 6370 22310 6490
rect 22355 6370 22475 6490
rect 22530 6370 22650 6490
rect 22695 6370 22815 6490
rect 22860 6370 22980 6490
rect 23025 6370 23145 6490
rect 23200 6370 23320 6490
rect 23365 6370 23485 6490
rect 23530 6370 23650 6490
rect 23695 6370 23815 6490
rect 23870 6370 23990 6490
rect 18510 6195 18630 6315
rect 18675 6195 18795 6315
rect 18840 6195 18960 6315
rect 19005 6195 19125 6315
rect 19180 6195 19300 6315
rect 19345 6195 19465 6315
rect 19510 6195 19630 6315
rect 19675 6195 19795 6315
rect 19850 6195 19970 6315
rect 20015 6195 20135 6315
rect 20180 6195 20300 6315
rect 20345 6195 20465 6315
rect 20520 6195 20640 6315
rect 20685 6195 20805 6315
rect 20850 6195 20970 6315
rect 21015 6195 21135 6315
rect 21190 6195 21310 6315
rect 21355 6195 21475 6315
rect 21520 6195 21640 6315
rect 21685 6195 21805 6315
rect 21860 6195 21980 6315
rect 22025 6195 22145 6315
rect 22190 6195 22310 6315
rect 22355 6195 22475 6315
rect 22530 6195 22650 6315
rect 22695 6195 22815 6315
rect 22860 6195 22980 6315
rect 23025 6195 23145 6315
rect 23200 6195 23320 6315
rect 23365 6195 23485 6315
rect 23530 6195 23650 6315
rect 23695 6195 23815 6315
rect 23870 6195 23990 6315
rect 18510 6030 18630 6150
rect 18675 6030 18795 6150
rect 18840 6030 18960 6150
rect 19005 6030 19125 6150
rect 19180 6030 19300 6150
rect 19345 6030 19465 6150
rect 19510 6030 19630 6150
rect 19675 6030 19795 6150
rect 19850 6030 19970 6150
rect 20015 6030 20135 6150
rect 20180 6030 20300 6150
rect 20345 6030 20465 6150
rect 20520 6030 20640 6150
rect 20685 6030 20805 6150
rect 20850 6030 20970 6150
rect 21015 6030 21135 6150
rect 21190 6030 21310 6150
rect 21355 6030 21475 6150
rect 21520 6030 21640 6150
rect 21685 6030 21805 6150
rect 21860 6030 21980 6150
rect 22025 6030 22145 6150
rect 22190 6030 22310 6150
rect 22355 6030 22475 6150
rect 22530 6030 22650 6150
rect 22695 6030 22815 6150
rect 22860 6030 22980 6150
rect 23025 6030 23145 6150
rect 23200 6030 23320 6150
rect 23365 6030 23485 6150
rect 23530 6030 23650 6150
rect 23695 6030 23815 6150
rect 23870 6030 23990 6150
rect 18510 5865 18630 5985
rect 18675 5865 18795 5985
rect 18840 5865 18960 5985
rect 19005 5865 19125 5985
rect 19180 5865 19300 5985
rect 19345 5865 19465 5985
rect 19510 5865 19630 5985
rect 19675 5865 19795 5985
rect 19850 5865 19970 5985
rect 20015 5865 20135 5985
rect 20180 5865 20300 5985
rect 20345 5865 20465 5985
rect 20520 5865 20640 5985
rect 20685 5865 20805 5985
rect 20850 5865 20970 5985
rect 21015 5865 21135 5985
rect 21190 5865 21310 5985
rect 21355 5865 21475 5985
rect 21520 5865 21640 5985
rect 21685 5865 21805 5985
rect 21860 5865 21980 5985
rect 22025 5865 22145 5985
rect 22190 5865 22310 5985
rect 22355 5865 22475 5985
rect 22530 5865 22650 5985
rect 22695 5865 22815 5985
rect 22860 5865 22980 5985
rect 23025 5865 23145 5985
rect 23200 5865 23320 5985
rect 23365 5865 23485 5985
rect 23530 5865 23650 5985
rect 23695 5865 23815 5985
rect 23870 5865 23990 5985
rect 18510 5700 18630 5820
rect 18675 5700 18795 5820
rect 18840 5700 18960 5820
rect 19005 5700 19125 5820
rect 19180 5700 19300 5820
rect 19345 5700 19465 5820
rect 19510 5700 19630 5820
rect 19675 5700 19795 5820
rect 19850 5700 19970 5820
rect 20015 5700 20135 5820
rect 20180 5700 20300 5820
rect 20345 5700 20465 5820
rect 20520 5700 20640 5820
rect 20685 5700 20805 5820
rect 20850 5700 20970 5820
rect 21015 5700 21135 5820
rect 21190 5700 21310 5820
rect 21355 5700 21475 5820
rect 21520 5700 21640 5820
rect 21685 5700 21805 5820
rect 21860 5700 21980 5820
rect 22025 5700 22145 5820
rect 22190 5700 22310 5820
rect 22355 5700 22475 5820
rect 22530 5700 22650 5820
rect 22695 5700 22815 5820
rect 22860 5700 22980 5820
rect 23025 5700 23145 5820
rect 23200 5700 23320 5820
rect 23365 5700 23485 5820
rect 23530 5700 23650 5820
rect 23695 5700 23815 5820
rect 23870 5700 23990 5820
rect 18510 5525 18630 5645
rect 18675 5525 18795 5645
rect 18840 5525 18960 5645
rect 19005 5525 19125 5645
rect 19180 5525 19300 5645
rect 19345 5525 19465 5645
rect 19510 5525 19630 5645
rect 19675 5525 19795 5645
rect 19850 5525 19970 5645
rect 20015 5525 20135 5645
rect 20180 5525 20300 5645
rect 20345 5525 20465 5645
rect 20520 5525 20640 5645
rect 20685 5525 20805 5645
rect 20850 5525 20970 5645
rect 21015 5525 21135 5645
rect 21190 5525 21310 5645
rect 21355 5525 21475 5645
rect 21520 5525 21640 5645
rect 21685 5525 21805 5645
rect 21860 5525 21980 5645
rect 22025 5525 22145 5645
rect 22190 5525 22310 5645
rect 22355 5525 22475 5645
rect 22530 5525 22650 5645
rect 22695 5525 22815 5645
rect 22860 5525 22980 5645
rect 23025 5525 23145 5645
rect 23200 5525 23320 5645
rect 23365 5525 23485 5645
rect 23530 5525 23650 5645
rect 23695 5525 23815 5645
rect 23870 5525 23990 5645
rect 18510 5360 18630 5480
rect 18675 5360 18795 5480
rect 18840 5360 18960 5480
rect 19005 5360 19125 5480
rect 19180 5360 19300 5480
rect 19345 5360 19465 5480
rect 19510 5360 19630 5480
rect 19675 5360 19795 5480
rect 19850 5360 19970 5480
rect 20015 5360 20135 5480
rect 20180 5360 20300 5480
rect 20345 5360 20465 5480
rect 20520 5360 20640 5480
rect 20685 5360 20805 5480
rect 20850 5360 20970 5480
rect 21015 5360 21135 5480
rect 21190 5360 21310 5480
rect 21355 5360 21475 5480
rect 21520 5360 21640 5480
rect 21685 5360 21805 5480
rect 21860 5360 21980 5480
rect 22025 5360 22145 5480
rect 22190 5360 22310 5480
rect 22355 5360 22475 5480
rect 22530 5360 22650 5480
rect 22695 5360 22815 5480
rect 22860 5360 22980 5480
rect 23025 5360 23145 5480
rect 23200 5360 23320 5480
rect 23365 5360 23485 5480
rect 23530 5360 23650 5480
rect 23695 5360 23815 5480
rect 23870 5360 23990 5480
rect 18510 5195 18630 5315
rect 18675 5195 18795 5315
rect 18840 5195 18960 5315
rect 19005 5195 19125 5315
rect 19180 5195 19300 5315
rect 19345 5195 19465 5315
rect 19510 5195 19630 5315
rect 19675 5195 19795 5315
rect 19850 5195 19970 5315
rect 20015 5195 20135 5315
rect 20180 5195 20300 5315
rect 20345 5195 20465 5315
rect 20520 5195 20640 5315
rect 20685 5195 20805 5315
rect 20850 5195 20970 5315
rect 21015 5195 21135 5315
rect 21190 5195 21310 5315
rect 21355 5195 21475 5315
rect 21520 5195 21640 5315
rect 21685 5195 21805 5315
rect 21860 5195 21980 5315
rect 22025 5195 22145 5315
rect 22190 5195 22310 5315
rect 22355 5195 22475 5315
rect 22530 5195 22650 5315
rect 22695 5195 22815 5315
rect 22860 5195 22980 5315
rect 23025 5195 23145 5315
rect 23200 5195 23320 5315
rect 23365 5195 23485 5315
rect 23530 5195 23650 5315
rect 23695 5195 23815 5315
rect 23870 5195 23990 5315
rect 18510 5030 18630 5150
rect 18675 5030 18795 5150
rect 18840 5030 18960 5150
rect 19005 5030 19125 5150
rect 19180 5030 19300 5150
rect 19345 5030 19465 5150
rect 19510 5030 19630 5150
rect 19675 5030 19795 5150
rect 19850 5030 19970 5150
rect 20015 5030 20135 5150
rect 20180 5030 20300 5150
rect 20345 5030 20465 5150
rect 20520 5030 20640 5150
rect 20685 5030 20805 5150
rect 20850 5030 20970 5150
rect 21015 5030 21135 5150
rect 21190 5030 21310 5150
rect 21355 5030 21475 5150
rect 21520 5030 21640 5150
rect 21685 5030 21805 5150
rect 21860 5030 21980 5150
rect 22025 5030 22145 5150
rect 22190 5030 22310 5150
rect 22355 5030 22475 5150
rect 22530 5030 22650 5150
rect 22695 5030 22815 5150
rect 22860 5030 22980 5150
rect 23025 5030 23145 5150
rect 23200 5030 23320 5150
rect 23365 5030 23485 5150
rect 23530 5030 23650 5150
rect 23695 5030 23815 5150
rect 23870 5030 23990 5150
rect 18510 4855 18630 4975
rect 18675 4855 18795 4975
rect 18840 4855 18960 4975
rect 19005 4855 19125 4975
rect 19180 4855 19300 4975
rect 19345 4855 19465 4975
rect 19510 4855 19630 4975
rect 19675 4855 19795 4975
rect 19850 4855 19970 4975
rect 20015 4855 20135 4975
rect 20180 4855 20300 4975
rect 20345 4855 20465 4975
rect 20520 4855 20640 4975
rect 20685 4855 20805 4975
rect 20850 4855 20970 4975
rect 21015 4855 21135 4975
rect 21190 4855 21310 4975
rect 21355 4855 21475 4975
rect 21520 4855 21640 4975
rect 21685 4855 21805 4975
rect 21860 4855 21980 4975
rect 22025 4855 22145 4975
rect 22190 4855 22310 4975
rect 22355 4855 22475 4975
rect 22530 4855 22650 4975
rect 22695 4855 22815 4975
rect 22860 4855 22980 4975
rect 23025 4855 23145 4975
rect 23200 4855 23320 4975
rect 23365 4855 23485 4975
rect 23530 4855 23650 4975
rect 23695 4855 23815 4975
rect 23870 4855 23990 4975
rect 18510 4690 18630 4810
rect 18675 4690 18795 4810
rect 18840 4690 18960 4810
rect 19005 4690 19125 4810
rect 19180 4690 19300 4810
rect 19345 4690 19465 4810
rect 19510 4690 19630 4810
rect 19675 4690 19795 4810
rect 19850 4690 19970 4810
rect 20015 4690 20135 4810
rect 20180 4690 20300 4810
rect 20345 4690 20465 4810
rect 20520 4690 20640 4810
rect 20685 4690 20805 4810
rect 20850 4690 20970 4810
rect 21015 4690 21135 4810
rect 21190 4690 21310 4810
rect 21355 4690 21475 4810
rect 21520 4690 21640 4810
rect 21685 4690 21805 4810
rect 21860 4690 21980 4810
rect 22025 4690 22145 4810
rect 22190 4690 22310 4810
rect 22355 4690 22475 4810
rect 22530 4690 22650 4810
rect 22695 4690 22815 4810
rect 22860 4690 22980 4810
rect 23025 4690 23145 4810
rect 23200 4690 23320 4810
rect 23365 4690 23485 4810
rect 23530 4690 23650 4810
rect 23695 4690 23815 4810
rect 23870 4690 23990 4810
rect 18510 4525 18630 4645
rect 18675 4525 18795 4645
rect 18840 4525 18960 4645
rect 19005 4525 19125 4645
rect 19180 4525 19300 4645
rect 19345 4525 19465 4645
rect 19510 4525 19630 4645
rect 19675 4525 19795 4645
rect 19850 4525 19970 4645
rect 20015 4525 20135 4645
rect 20180 4525 20300 4645
rect 20345 4525 20465 4645
rect 20520 4525 20640 4645
rect 20685 4525 20805 4645
rect 20850 4525 20970 4645
rect 21015 4525 21135 4645
rect 21190 4525 21310 4645
rect 21355 4525 21475 4645
rect 21520 4525 21640 4645
rect 21685 4525 21805 4645
rect 21860 4525 21980 4645
rect 22025 4525 22145 4645
rect 22190 4525 22310 4645
rect 22355 4525 22475 4645
rect 22530 4525 22650 4645
rect 22695 4525 22815 4645
rect 22860 4525 22980 4645
rect 23025 4525 23145 4645
rect 23200 4525 23320 4645
rect 23365 4525 23485 4645
rect 23530 4525 23650 4645
rect 23695 4525 23815 4645
rect 23870 4525 23990 4645
rect 18510 4360 18630 4480
rect 18675 4360 18795 4480
rect 18840 4360 18960 4480
rect 19005 4360 19125 4480
rect 19180 4360 19300 4480
rect 19345 4360 19465 4480
rect 19510 4360 19630 4480
rect 19675 4360 19795 4480
rect 19850 4360 19970 4480
rect 20015 4360 20135 4480
rect 20180 4360 20300 4480
rect 20345 4360 20465 4480
rect 20520 4360 20640 4480
rect 20685 4360 20805 4480
rect 20850 4360 20970 4480
rect 21015 4360 21135 4480
rect 21190 4360 21310 4480
rect 21355 4360 21475 4480
rect 21520 4360 21640 4480
rect 21685 4360 21805 4480
rect 21860 4360 21980 4480
rect 22025 4360 22145 4480
rect 22190 4360 22310 4480
rect 22355 4360 22475 4480
rect 22530 4360 22650 4480
rect 22695 4360 22815 4480
rect 22860 4360 22980 4480
rect 23025 4360 23145 4480
rect 23200 4360 23320 4480
rect 23365 4360 23485 4480
rect 23530 4360 23650 4480
rect 23695 4360 23815 4480
rect 23870 4360 23990 4480
rect 18510 4185 18630 4305
rect 18675 4185 18795 4305
rect 18840 4185 18960 4305
rect 19005 4185 19125 4305
rect 19180 4185 19300 4305
rect 19345 4185 19465 4305
rect 19510 4185 19630 4305
rect 19675 4185 19795 4305
rect 19850 4185 19970 4305
rect 20015 4185 20135 4305
rect 20180 4185 20300 4305
rect 20345 4185 20465 4305
rect 20520 4185 20640 4305
rect 20685 4185 20805 4305
rect 20850 4185 20970 4305
rect 21015 4185 21135 4305
rect 21190 4185 21310 4305
rect 21355 4185 21475 4305
rect 21520 4185 21640 4305
rect 21685 4185 21805 4305
rect 21860 4185 21980 4305
rect 22025 4185 22145 4305
rect 22190 4185 22310 4305
rect 22355 4185 22475 4305
rect 22530 4185 22650 4305
rect 22695 4185 22815 4305
rect 22860 4185 22980 4305
rect 23025 4185 23145 4305
rect 23200 4185 23320 4305
rect 23365 4185 23485 4305
rect 23530 4185 23650 4305
rect 23695 4185 23815 4305
rect 23870 4185 23990 4305
rect 18510 4020 18630 4140
rect 18675 4020 18795 4140
rect 18840 4020 18960 4140
rect 19005 4020 19125 4140
rect 19180 4020 19300 4140
rect 19345 4020 19465 4140
rect 19510 4020 19630 4140
rect 19675 4020 19795 4140
rect 19850 4020 19970 4140
rect 20015 4020 20135 4140
rect 20180 4020 20300 4140
rect 20345 4020 20465 4140
rect 20520 4020 20640 4140
rect 20685 4020 20805 4140
rect 20850 4020 20970 4140
rect 21015 4020 21135 4140
rect 21190 4020 21310 4140
rect 21355 4020 21475 4140
rect 21520 4020 21640 4140
rect 21685 4020 21805 4140
rect 21860 4020 21980 4140
rect 22025 4020 22145 4140
rect 22190 4020 22310 4140
rect 22355 4020 22475 4140
rect 22530 4020 22650 4140
rect 22695 4020 22815 4140
rect 22860 4020 22980 4140
rect 23025 4020 23145 4140
rect 23200 4020 23320 4140
rect 23365 4020 23485 4140
rect 23530 4020 23650 4140
rect 23695 4020 23815 4140
rect 23870 4020 23990 4140
rect 18510 3855 18630 3975
rect 18675 3855 18795 3975
rect 18840 3855 18960 3975
rect 19005 3855 19125 3975
rect 19180 3855 19300 3975
rect 19345 3855 19465 3975
rect 19510 3855 19630 3975
rect 19675 3855 19795 3975
rect 19850 3855 19970 3975
rect 20015 3855 20135 3975
rect 20180 3855 20300 3975
rect 20345 3855 20465 3975
rect 20520 3855 20640 3975
rect 20685 3855 20805 3975
rect 20850 3855 20970 3975
rect 21015 3855 21135 3975
rect 21190 3855 21310 3975
rect 21355 3855 21475 3975
rect 21520 3855 21640 3975
rect 21685 3855 21805 3975
rect 21860 3855 21980 3975
rect 22025 3855 22145 3975
rect 22190 3855 22310 3975
rect 22355 3855 22475 3975
rect 22530 3855 22650 3975
rect 22695 3855 22815 3975
rect 22860 3855 22980 3975
rect 23025 3855 23145 3975
rect 23200 3855 23320 3975
rect 23365 3855 23485 3975
rect 23530 3855 23650 3975
rect 23695 3855 23815 3975
rect 23870 3855 23990 3975
rect 18510 3690 18630 3810
rect 18675 3690 18795 3810
rect 18840 3690 18960 3810
rect 19005 3690 19125 3810
rect 19180 3690 19300 3810
rect 19345 3690 19465 3810
rect 19510 3690 19630 3810
rect 19675 3690 19795 3810
rect 19850 3690 19970 3810
rect 20015 3690 20135 3810
rect 20180 3690 20300 3810
rect 20345 3690 20465 3810
rect 20520 3690 20640 3810
rect 20685 3690 20805 3810
rect 20850 3690 20970 3810
rect 21015 3690 21135 3810
rect 21190 3690 21310 3810
rect 21355 3690 21475 3810
rect 21520 3690 21640 3810
rect 21685 3690 21805 3810
rect 21860 3690 21980 3810
rect 22025 3690 22145 3810
rect 22190 3690 22310 3810
rect 22355 3690 22475 3810
rect 22530 3690 22650 3810
rect 22695 3690 22815 3810
rect 22860 3690 22980 3810
rect 23025 3690 23145 3810
rect 23200 3690 23320 3810
rect 23365 3690 23485 3810
rect 23530 3690 23650 3810
rect 23695 3690 23815 3810
rect 23870 3690 23990 3810
rect 18510 3515 18630 3635
rect 18675 3515 18795 3635
rect 18840 3515 18960 3635
rect 19005 3515 19125 3635
rect 19180 3515 19300 3635
rect 19345 3515 19465 3635
rect 19510 3515 19630 3635
rect 19675 3515 19795 3635
rect 19850 3515 19970 3635
rect 20015 3515 20135 3635
rect 20180 3515 20300 3635
rect 20345 3515 20465 3635
rect 20520 3515 20640 3635
rect 20685 3515 20805 3635
rect 20850 3515 20970 3635
rect 21015 3515 21135 3635
rect 21190 3515 21310 3635
rect 21355 3515 21475 3635
rect 21520 3515 21640 3635
rect 21685 3515 21805 3635
rect 21860 3515 21980 3635
rect 22025 3515 22145 3635
rect 22190 3515 22310 3635
rect 22355 3515 22475 3635
rect 22530 3515 22650 3635
rect 22695 3515 22815 3635
rect 22860 3515 22980 3635
rect 23025 3515 23145 3635
rect 23200 3515 23320 3635
rect 23365 3515 23485 3635
rect 23530 3515 23650 3635
rect 23695 3515 23815 3635
rect 23870 3515 23990 3635
rect 18510 3350 18630 3470
rect 18675 3350 18795 3470
rect 18840 3350 18960 3470
rect 19005 3350 19125 3470
rect 19180 3350 19300 3470
rect 19345 3350 19465 3470
rect 19510 3350 19630 3470
rect 19675 3350 19795 3470
rect 19850 3350 19970 3470
rect 20015 3350 20135 3470
rect 20180 3350 20300 3470
rect 20345 3350 20465 3470
rect 20520 3350 20640 3470
rect 20685 3350 20805 3470
rect 20850 3350 20970 3470
rect 21015 3350 21135 3470
rect 21190 3350 21310 3470
rect 21355 3350 21475 3470
rect 21520 3350 21640 3470
rect 21685 3350 21805 3470
rect 21860 3350 21980 3470
rect 22025 3350 22145 3470
rect 22190 3350 22310 3470
rect 22355 3350 22475 3470
rect 22530 3350 22650 3470
rect 22695 3350 22815 3470
rect 22860 3350 22980 3470
rect 23025 3350 23145 3470
rect 23200 3350 23320 3470
rect 23365 3350 23485 3470
rect 23530 3350 23650 3470
rect 23695 3350 23815 3470
rect 23870 3350 23990 3470
rect 18510 3185 18630 3305
rect 18675 3185 18795 3305
rect 18840 3185 18960 3305
rect 19005 3185 19125 3305
rect 19180 3185 19300 3305
rect 19345 3185 19465 3305
rect 19510 3185 19630 3305
rect 19675 3185 19795 3305
rect 19850 3185 19970 3305
rect 20015 3185 20135 3305
rect 20180 3185 20300 3305
rect 20345 3185 20465 3305
rect 20520 3185 20640 3305
rect 20685 3185 20805 3305
rect 20850 3185 20970 3305
rect 21015 3185 21135 3305
rect 21190 3185 21310 3305
rect 21355 3185 21475 3305
rect 21520 3185 21640 3305
rect 21685 3185 21805 3305
rect 21860 3185 21980 3305
rect 22025 3185 22145 3305
rect 22190 3185 22310 3305
rect 22355 3185 22475 3305
rect 22530 3185 22650 3305
rect 22695 3185 22815 3305
rect 22860 3185 22980 3305
rect 23025 3185 23145 3305
rect 23200 3185 23320 3305
rect 23365 3185 23485 3305
rect 23530 3185 23650 3305
rect 23695 3185 23815 3305
rect 23870 3185 23990 3305
rect 18510 3020 18630 3140
rect 18675 3020 18795 3140
rect 18840 3020 18960 3140
rect 19005 3020 19125 3140
rect 19180 3020 19300 3140
rect 19345 3020 19465 3140
rect 19510 3020 19630 3140
rect 19675 3020 19795 3140
rect 19850 3020 19970 3140
rect 20015 3020 20135 3140
rect 20180 3020 20300 3140
rect 20345 3020 20465 3140
rect 20520 3020 20640 3140
rect 20685 3020 20805 3140
rect 20850 3020 20970 3140
rect 21015 3020 21135 3140
rect 21190 3020 21310 3140
rect 21355 3020 21475 3140
rect 21520 3020 21640 3140
rect 21685 3020 21805 3140
rect 21860 3020 21980 3140
rect 22025 3020 22145 3140
rect 22190 3020 22310 3140
rect 22355 3020 22475 3140
rect 22530 3020 22650 3140
rect 22695 3020 22815 3140
rect 22860 3020 22980 3140
rect 23025 3020 23145 3140
rect 23200 3020 23320 3140
rect 23365 3020 23485 3140
rect 23530 3020 23650 3140
rect 23695 3020 23815 3140
rect 23870 3020 23990 3140
rect 18510 2845 18630 2965
rect 18675 2845 18795 2965
rect 18840 2845 18960 2965
rect 19005 2845 19125 2965
rect 19180 2845 19300 2965
rect 19345 2845 19465 2965
rect 19510 2845 19630 2965
rect 19675 2845 19795 2965
rect 19850 2845 19970 2965
rect 20015 2845 20135 2965
rect 20180 2845 20300 2965
rect 20345 2845 20465 2965
rect 20520 2845 20640 2965
rect 20685 2845 20805 2965
rect 20850 2845 20970 2965
rect 21015 2845 21135 2965
rect 21190 2845 21310 2965
rect 21355 2845 21475 2965
rect 21520 2845 21640 2965
rect 21685 2845 21805 2965
rect 21860 2845 21980 2965
rect 22025 2845 22145 2965
rect 22190 2845 22310 2965
rect 22355 2845 22475 2965
rect 22530 2845 22650 2965
rect 22695 2845 22815 2965
rect 22860 2845 22980 2965
rect 23025 2845 23145 2965
rect 23200 2845 23320 2965
rect 23365 2845 23485 2965
rect 23530 2845 23650 2965
rect 23695 2845 23815 2965
rect 23870 2845 23990 2965
rect 18510 2680 18630 2800
rect 18675 2680 18795 2800
rect 18840 2680 18960 2800
rect 19005 2680 19125 2800
rect 19180 2680 19300 2800
rect 19345 2680 19465 2800
rect 19510 2680 19630 2800
rect 19675 2680 19795 2800
rect 19850 2680 19970 2800
rect 20015 2680 20135 2800
rect 20180 2680 20300 2800
rect 20345 2680 20465 2800
rect 20520 2680 20640 2800
rect 20685 2680 20805 2800
rect 20850 2680 20970 2800
rect 21015 2680 21135 2800
rect 21190 2680 21310 2800
rect 21355 2680 21475 2800
rect 21520 2680 21640 2800
rect 21685 2680 21805 2800
rect 21860 2680 21980 2800
rect 22025 2680 22145 2800
rect 22190 2680 22310 2800
rect 22355 2680 22475 2800
rect 22530 2680 22650 2800
rect 22695 2680 22815 2800
rect 22860 2680 22980 2800
rect 23025 2680 23145 2800
rect 23200 2680 23320 2800
rect 23365 2680 23485 2800
rect 23530 2680 23650 2800
rect 23695 2680 23815 2800
rect 23870 2680 23990 2800
rect 18510 2515 18630 2635
rect 18675 2515 18795 2635
rect 18840 2515 18960 2635
rect 19005 2515 19125 2635
rect 19180 2515 19300 2635
rect 19345 2515 19465 2635
rect 19510 2515 19630 2635
rect 19675 2515 19795 2635
rect 19850 2515 19970 2635
rect 20015 2515 20135 2635
rect 20180 2515 20300 2635
rect 20345 2515 20465 2635
rect 20520 2515 20640 2635
rect 20685 2515 20805 2635
rect 20850 2515 20970 2635
rect 21015 2515 21135 2635
rect 21190 2515 21310 2635
rect 21355 2515 21475 2635
rect 21520 2515 21640 2635
rect 21685 2515 21805 2635
rect 21860 2515 21980 2635
rect 22025 2515 22145 2635
rect 22190 2515 22310 2635
rect 22355 2515 22475 2635
rect 22530 2515 22650 2635
rect 22695 2515 22815 2635
rect 22860 2515 22980 2635
rect 23025 2515 23145 2635
rect 23200 2515 23320 2635
rect 23365 2515 23485 2635
rect 23530 2515 23650 2635
rect 23695 2515 23815 2635
rect 23870 2515 23990 2635
rect 18510 2350 18630 2470
rect 18675 2350 18795 2470
rect 18840 2350 18960 2470
rect 19005 2350 19125 2470
rect 19180 2350 19300 2470
rect 19345 2350 19465 2470
rect 19510 2350 19630 2470
rect 19675 2350 19795 2470
rect 19850 2350 19970 2470
rect 20015 2350 20135 2470
rect 20180 2350 20300 2470
rect 20345 2350 20465 2470
rect 20520 2350 20640 2470
rect 20685 2350 20805 2470
rect 20850 2350 20970 2470
rect 21015 2350 21135 2470
rect 21190 2350 21310 2470
rect 21355 2350 21475 2470
rect 21520 2350 21640 2470
rect 21685 2350 21805 2470
rect 21860 2350 21980 2470
rect 22025 2350 22145 2470
rect 22190 2350 22310 2470
rect 22355 2350 22475 2470
rect 22530 2350 22650 2470
rect 22695 2350 22815 2470
rect 22860 2350 22980 2470
rect 23025 2350 23145 2470
rect 23200 2350 23320 2470
rect 23365 2350 23485 2470
rect 23530 2350 23650 2470
rect 23695 2350 23815 2470
rect 23870 2350 23990 2470
rect 18510 2175 18630 2295
rect 18675 2175 18795 2295
rect 18840 2175 18960 2295
rect 19005 2175 19125 2295
rect 19180 2175 19300 2295
rect 19345 2175 19465 2295
rect 19510 2175 19630 2295
rect 19675 2175 19795 2295
rect 19850 2175 19970 2295
rect 20015 2175 20135 2295
rect 20180 2175 20300 2295
rect 20345 2175 20465 2295
rect 20520 2175 20640 2295
rect 20685 2175 20805 2295
rect 20850 2175 20970 2295
rect 21015 2175 21135 2295
rect 21190 2175 21310 2295
rect 21355 2175 21475 2295
rect 21520 2175 21640 2295
rect 21685 2175 21805 2295
rect 21860 2175 21980 2295
rect 22025 2175 22145 2295
rect 22190 2175 22310 2295
rect 22355 2175 22475 2295
rect 22530 2175 22650 2295
rect 22695 2175 22815 2295
rect 22860 2175 22980 2295
rect 23025 2175 23145 2295
rect 23200 2175 23320 2295
rect 23365 2175 23485 2295
rect 23530 2175 23650 2295
rect 23695 2175 23815 2295
rect 23870 2175 23990 2295
rect 18510 2010 18630 2130
rect 18675 2010 18795 2130
rect 18840 2010 18960 2130
rect 19005 2010 19125 2130
rect 19180 2010 19300 2130
rect 19345 2010 19465 2130
rect 19510 2010 19630 2130
rect 19675 2010 19795 2130
rect 19850 2010 19970 2130
rect 20015 2010 20135 2130
rect 20180 2010 20300 2130
rect 20345 2010 20465 2130
rect 20520 2010 20640 2130
rect 20685 2010 20805 2130
rect 20850 2010 20970 2130
rect 21015 2010 21135 2130
rect 21190 2010 21310 2130
rect 21355 2010 21475 2130
rect 21520 2010 21640 2130
rect 21685 2010 21805 2130
rect 21860 2010 21980 2130
rect 22025 2010 22145 2130
rect 22190 2010 22310 2130
rect 22355 2010 22475 2130
rect 22530 2010 22650 2130
rect 22695 2010 22815 2130
rect 22860 2010 22980 2130
rect 23025 2010 23145 2130
rect 23200 2010 23320 2130
rect 23365 2010 23485 2130
rect 23530 2010 23650 2130
rect 23695 2010 23815 2130
rect 23870 2010 23990 2130
rect 18510 1845 18630 1965
rect 18675 1845 18795 1965
rect 18840 1845 18960 1965
rect 19005 1845 19125 1965
rect 19180 1845 19300 1965
rect 19345 1845 19465 1965
rect 19510 1845 19630 1965
rect 19675 1845 19795 1965
rect 19850 1845 19970 1965
rect 20015 1845 20135 1965
rect 20180 1845 20300 1965
rect 20345 1845 20465 1965
rect 20520 1845 20640 1965
rect 20685 1845 20805 1965
rect 20850 1845 20970 1965
rect 21015 1845 21135 1965
rect 21190 1845 21310 1965
rect 21355 1845 21475 1965
rect 21520 1845 21640 1965
rect 21685 1845 21805 1965
rect 21860 1845 21980 1965
rect 22025 1845 22145 1965
rect 22190 1845 22310 1965
rect 22355 1845 22475 1965
rect 22530 1845 22650 1965
rect 22695 1845 22815 1965
rect 22860 1845 22980 1965
rect 23025 1845 23145 1965
rect 23200 1845 23320 1965
rect 23365 1845 23485 1965
rect 23530 1845 23650 1965
rect 23695 1845 23815 1965
rect 23870 1845 23990 1965
rect 18510 1680 18630 1800
rect 18675 1680 18795 1800
rect 18840 1680 18960 1800
rect 19005 1680 19125 1800
rect 19180 1680 19300 1800
rect 19345 1680 19465 1800
rect 19510 1680 19630 1800
rect 19675 1680 19795 1800
rect 19850 1680 19970 1800
rect 20015 1680 20135 1800
rect 20180 1680 20300 1800
rect 20345 1680 20465 1800
rect 20520 1680 20640 1800
rect 20685 1680 20805 1800
rect 20850 1680 20970 1800
rect 21015 1680 21135 1800
rect 21190 1680 21310 1800
rect 21355 1680 21475 1800
rect 21520 1680 21640 1800
rect 21685 1680 21805 1800
rect 21860 1680 21980 1800
rect 22025 1680 22145 1800
rect 22190 1680 22310 1800
rect 22355 1680 22475 1800
rect 22530 1680 22650 1800
rect 22695 1680 22815 1800
rect 22860 1680 22980 1800
rect 23025 1680 23145 1800
rect 23200 1680 23320 1800
rect 23365 1680 23485 1800
rect 23530 1680 23650 1800
rect 23695 1680 23815 1800
rect 23870 1680 23990 1800
rect 24200 7040 24320 7160
rect 24365 7040 24485 7160
rect 24530 7040 24650 7160
rect 24695 7040 24815 7160
rect 24870 7040 24990 7160
rect 25035 7040 25155 7160
rect 25200 7040 25320 7160
rect 25365 7040 25485 7160
rect 25540 7040 25660 7160
rect 25705 7040 25825 7160
rect 25870 7040 25990 7160
rect 26035 7040 26155 7160
rect 26210 7040 26330 7160
rect 26375 7040 26495 7160
rect 26540 7040 26660 7160
rect 26705 7040 26825 7160
rect 26880 7040 27000 7160
rect 27045 7040 27165 7160
rect 27210 7040 27330 7160
rect 27375 7040 27495 7160
rect 27550 7040 27670 7160
rect 27715 7040 27835 7160
rect 27880 7040 28000 7160
rect 28045 7040 28165 7160
rect 28220 7040 28340 7160
rect 28385 7040 28505 7160
rect 28550 7040 28670 7160
rect 28715 7040 28835 7160
rect 28890 7040 29010 7160
rect 29055 7040 29175 7160
rect 29220 7040 29340 7160
rect 29385 7040 29505 7160
rect 29560 7040 29680 7160
rect 24200 6865 24320 6985
rect 24365 6865 24485 6985
rect 24530 6865 24650 6985
rect 24695 6865 24815 6985
rect 24870 6865 24990 6985
rect 25035 6865 25155 6985
rect 25200 6865 25320 6985
rect 25365 6865 25485 6985
rect 25540 6865 25660 6985
rect 25705 6865 25825 6985
rect 25870 6865 25990 6985
rect 26035 6865 26155 6985
rect 26210 6865 26330 6985
rect 26375 6865 26495 6985
rect 26540 6865 26660 6985
rect 26705 6865 26825 6985
rect 26880 6865 27000 6985
rect 27045 6865 27165 6985
rect 27210 6865 27330 6985
rect 27375 6865 27495 6985
rect 27550 6865 27670 6985
rect 27715 6865 27835 6985
rect 27880 6865 28000 6985
rect 28045 6865 28165 6985
rect 28220 6865 28340 6985
rect 28385 6865 28505 6985
rect 28550 6865 28670 6985
rect 28715 6865 28835 6985
rect 28890 6865 29010 6985
rect 29055 6865 29175 6985
rect 29220 6865 29340 6985
rect 29385 6865 29505 6985
rect 29560 6865 29680 6985
rect 24200 6700 24320 6820
rect 24365 6700 24485 6820
rect 24530 6700 24650 6820
rect 24695 6700 24815 6820
rect 24870 6700 24990 6820
rect 25035 6700 25155 6820
rect 25200 6700 25320 6820
rect 25365 6700 25485 6820
rect 25540 6700 25660 6820
rect 25705 6700 25825 6820
rect 25870 6700 25990 6820
rect 26035 6700 26155 6820
rect 26210 6700 26330 6820
rect 26375 6700 26495 6820
rect 26540 6700 26660 6820
rect 26705 6700 26825 6820
rect 26880 6700 27000 6820
rect 27045 6700 27165 6820
rect 27210 6700 27330 6820
rect 27375 6700 27495 6820
rect 27550 6700 27670 6820
rect 27715 6700 27835 6820
rect 27880 6700 28000 6820
rect 28045 6700 28165 6820
rect 28220 6700 28340 6820
rect 28385 6700 28505 6820
rect 28550 6700 28670 6820
rect 28715 6700 28835 6820
rect 28890 6700 29010 6820
rect 29055 6700 29175 6820
rect 29220 6700 29340 6820
rect 29385 6700 29505 6820
rect 29560 6700 29680 6820
rect 24200 6535 24320 6655
rect 24365 6535 24485 6655
rect 24530 6535 24650 6655
rect 24695 6535 24815 6655
rect 24870 6535 24990 6655
rect 25035 6535 25155 6655
rect 25200 6535 25320 6655
rect 25365 6535 25485 6655
rect 25540 6535 25660 6655
rect 25705 6535 25825 6655
rect 25870 6535 25990 6655
rect 26035 6535 26155 6655
rect 26210 6535 26330 6655
rect 26375 6535 26495 6655
rect 26540 6535 26660 6655
rect 26705 6535 26825 6655
rect 26880 6535 27000 6655
rect 27045 6535 27165 6655
rect 27210 6535 27330 6655
rect 27375 6535 27495 6655
rect 27550 6535 27670 6655
rect 27715 6535 27835 6655
rect 27880 6535 28000 6655
rect 28045 6535 28165 6655
rect 28220 6535 28340 6655
rect 28385 6535 28505 6655
rect 28550 6535 28670 6655
rect 28715 6535 28835 6655
rect 28890 6535 29010 6655
rect 29055 6535 29175 6655
rect 29220 6535 29340 6655
rect 29385 6535 29505 6655
rect 29560 6535 29680 6655
rect 24200 6370 24320 6490
rect 24365 6370 24485 6490
rect 24530 6370 24650 6490
rect 24695 6370 24815 6490
rect 24870 6370 24990 6490
rect 25035 6370 25155 6490
rect 25200 6370 25320 6490
rect 25365 6370 25485 6490
rect 25540 6370 25660 6490
rect 25705 6370 25825 6490
rect 25870 6370 25990 6490
rect 26035 6370 26155 6490
rect 26210 6370 26330 6490
rect 26375 6370 26495 6490
rect 26540 6370 26660 6490
rect 26705 6370 26825 6490
rect 26880 6370 27000 6490
rect 27045 6370 27165 6490
rect 27210 6370 27330 6490
rect 27375 6370 27495 6490
rect 27550 6370 27670 6490
rect 27715 6370 27835 6490
rect 27880 6370 28000 6490
rect 28045 6370 28165 6490
rect 28220 6370 28340 6490
rect 28385 6370 28505 6490
rect 28550 6370 28670 6490
rect 28715 6370 28835 6490
rect 28890 6370 29010 6490
rect 29055 6370 29175 6490
rect 29220 6370 29340 6490
rect 29385 6370 29505 6490
rect 29560 6370 29680 6490
rect 24200 6195 24320 6315
rect 24365 6195 24485 6315
rect 24530 6195 24650 6315
rect 24695 6195 24815 6315
rect 24870 6195 24990 6315
rect 25035 6195 25155 6315
rect 25200 6195 25320 6315
rect 25365 6195 25485 6315
rect 25540 6195 25660 6315
rect 25705 6195 25825 6315
rect 25870 6195 25990 6315
rect 26035 6195 26155 6315
rect 26210 6195 26330 6315
rect 26375 6195 26495 6315
rect 26540 6195 26660 6315
rect 26705 6195 26825 6315
rect 26880 6195 27000 6315
rect 27045 6195 27165 6315
rect 27210 6195 27330 6315
rect 27375 6195 27495 6315
rect 27550 6195 27670 6315
rect 27715 6195 27835 6315
rect 27880 6195 28000 6315
rect 28045 6195 28165 6315
rect 28220 6195 28340 6315
rect 28385 6195 28505 6315
rect 28550 6195 28670 6315
rect 28715 6195 28835 6315
rect 28890 6195 29010 6315
rect 29055 6195 29175 6315
rect 29220 6195 29340 6315
rect 29385 6195 29505 6315
rect 29560 6195 29680 6315
rect 24200 6030 24320 6150
rect 24365 6030 24485 6150
rect 24530 6030 24650 6150
rect 24695 6030 24815 6150
rect 24870 6030 24990 6150
rect 25035 6030 25155 6150
rect 25200 6030 25320 6150
rect 25365 6030 25485 6150
rect 25540 6030 25660 6150
rect 25705 6030 25825 6150
rect 25870 6030 25990 6150
rect 26035 6030 26155 6150
rect 26210 6030 26330 6150
rect 26375 6030 26495 6150
rect 26540 6030 26660 6150
rect 26705 6030 26825 6150
rect 26880 6030 27000 6150
rect 27045 6030 27165 6150
rect 27210 6030 27330 6150
rect 27375 6030 27495 6150
rect 27550 6030 27670 6150
rect 27715 6030 27835 6150
rect 27880 6030 28000 6150
rect 28045 6030 28165 6150
rect 28220 6030 28340 6150
rect 28385 6030 28505 6150
rect 28550 6030 28670 6150
rect 28715 6030 28835 6150
rect 28890 6030 29010 6150
rect 29055 6030 29175 6150
rect 29220 6030 29340 6150
rect 29385 6030 29505 6150
rect 29560 6030 29680 6150
rect 24200 5865 24320 5985
rect 24365 5865 24485 5985
rect 24530 5865 24650 5985
rect 24695 5865 24815 5985
rect 24870 5865 24990 5985
rect 25035 5865 25155 5985
rect 25200 5865 25320 5985
rect 25365 5865 25485 5985
rect 25540 5865 25660 5985
rect 25705 5865 25825 5985
rect 25870 5865 25990 5985
rect 26035 5865 26155 5985
rect 26210 5865 26330 5985
rect 26375 5865 26495 5985
rect 26540 5865 26660 5985
rect 26705 5865 26825 5985
rect 26880 5865 27000 5985
rect 27045 5865 27165 5985
rect 27210 5865 27330 5985
rect 27375 5865 27495 5985
rect 27550 5865 27670 5985
rect 27715 5865 27835 5985
rect 27880 5865 28000 5985
rect 28045 5865 28165 5985
rect 28220 5865 28340 5985
rect 28385 5865 28505 5985
rect 28550 5865 28670 5985
rect 28715 5865 28835 5985
rect 28890 5865 29010 5985
rect 29055 5865 29175 5985
rect 29220 5865 29340 5985
rect 29385 5865 29505 5985
rect 29560 5865 29680 5985
rect 24200 5700 24320 5820
rect 24365 5700 24485 5820
rect 24530 5700 24650 5820
rect 24695 5700 24815 5820
rect 24870 5700 24990 5820
rect 25035 5700 25155 5820
rect 25200 5700 25320 5820
rect 25365 5700 25485 5820
rect 25540 5700 25660 5820
rect 25705 5700 25825 5820
rect 25870 5700 25990 5820
rect 26035 5700 26155 5820
rect 26210 5700 26330 5820
rect 26375 5700 26495 5820
rect 26540 5700 26660 5820
rect 26705 5700 26825 5820
rect 26880 5700 27000 5820
rect 27045 5700 27165 5820
rect 27210 5700 27330 5820
rect 27375 5700 27495 5820
rect 27550 5700 27670 5820
rect 27715 5700 27835 5820
rect 27880 5700 28000 5820
rect 28045 5700 28165 5820
rect 28220 5700 28340 5820
rect 28385 5700 28505 5820
rect 28550 5700 28670 5820
rect 28715 5700 28835 5820
rect 28890 5700 29010 5820
rect 29055 5700 29175 5820
rect 29220 5700 29340 5820
rect 29385 5700 29505 5820
rect 29560 5700 29680 5820
rect 24200 5525 24320 5645
rect 24365 5525 24485 5645
rect 24530 5525 24650 5645
rect 24695 5525 24815 5645
rect 24870 5525 24990 5645
rect 25035 5525 25155 5645
rect 25200 5525 25320 5645
rect 25365 5525 25485 5645
rect 25540 5525 25660 5645
rect 25705 5525 25825 5645
rect 25870 5525 25990 5645
rect 26035 5525 26155 5645
rect 26210 5525 26330 5645
rect 26375 5525 26495 5645
rect 26540 5525 26660 5645
rect 26705 5525 26825 5645
rect 26880 5525 27000 5645
rect 27045 5525 27165 5645
rect 27210 5525 27330 5645
rect 27375 5525 27495 5645
rect 27550 5525 27670 5645
rect 27715 5525 27835 5645
rect 27880 5525 28000 5645
rect 28045 5525 28165 5645
rect 28220 5525 28340 5645
rect 28385 5525 28505 5645
rect 28550 5525 28670 5645
rect 28715 5525 28835 5645
rect 28890 5525 29010 5645
rect 29055 5525 29175 5645
rect 29220 5525 29340 5645
rect 29385 5525 29505 5645
rect 29560 5525 29680 5645
rect 24200 5360 24320 5480
rect 24365 5360 24485 5480
rect 24530 5360 24650 5480
rect 24695 5360 24815 5480
rect 24870 5360 24990 5480
rect 25035 5360 25155 5480
rect 25200 5360 25320 5480
rect 25365 5360 25485 5480
rect 25540 5360 25660 5480
rect 25705 5360 25825 5480
rect 25870 5360 25990 5480
rect 26035 5360 26155 5480
rect 26210 5360 26330 5480
rect 26375 5360 26495 5480
rect 26540 5360 26660 5480
rect 26705 5360 26825 5480
rect 26880 5360 27000 5480
rect 27045 5360 27165 5480
rect 27210 5360 27330 5480
rect 27375 5360 27495 5480
rect 27550 5360 27670 5480
rect 27715 5360 27835 5480
rect 27880 5360 28000 5480
rect 28045 5360 28165 5480
rect 28220 5360 28340 5480
rect 28385 5360 28505 5480
rect 28550 5360 28670 5480
rect 28715 5360 28835 5480
rect 28890 5360 29010 5480
rect 29055 5360 29175 5480
rect 29220 5360 29340 5480
rect 29385 5360 29505 5480
rect 29560 5360 29680 5480
rect 24200 5195 24320 5315
rect 24365 5195 24485 5315
rect 24530 5195 24650 5315
rect 24695 5195 24815 5315
rect 24870 5195 24990 5315
rect 25035 5195 25155 5315
rect 25200 5195 25320 5315
rect 25365 5195 25485 5315
rect 25540 5195 25660 5315
rect 25705 5195 25825 5315
rect 25870 5195 25990 5315
rect 26035 5195 26155 5315
rect 26210 5195 26330 5315
rect 26375 5195 26495 5315
rect 26540 5195 26660 5315
rect 26705 5195 26825 5315
rect 26880 5195 27000 5315
rect 27045 5195 27165 5315
rect 27210 5195 27330 5315
rect 27375 5195 27495 5315
rect 27550 5195 27670 5315
rect 27715 5195 27835 5315
rect 27880 5195 28000 5315
rect 28045 5195 28165 5315
rect 28220 5195 28340 5315
rect 28385 5195 28505 5315
rect 28550 5195 28670 5315
rect 28715 5195 28835 5315
rect 28890 5195 29010 5315
rect 29055 5195 29175 5315
rect 29220 5195 29340 5315
rect 29385 5195 29505 5315
rect 29560 5195 29680 5315
rect 24200 5030 24320 5150
rect 24365 5030 24485 5150
rect 24530 5030 24650 5150
rect 24695 5030 24815 5150
rect 24870 5030 24990 5150
rect 25035 5030 25155 5150
rect 25200 5030 25320 5150
rect 25365 5030 25485 5150
rect 25540 5030 25660 5150
rect 25705 5030 25825 5150
rect 25870 5030 25990 5150
rect 26035 5030 26155 5150
rect 26210 5030 26330 5150
rect 26375 5030 26495 5150
rect 26540 5030 26660 5150
rect 26705 5030 26825 5150
rect 26880 5030 27000 5150
rect 27045 5030 27165 5150
rect 27210 5030 27330 5150
rect 27375 5030 27495 5150
rect 27550 5030 27670 5150
rect 27715 5030 27835 5150
rect 27880 5030 28000 5150
rect 28045 5030 28165 5150
rect 28220 5030 28340 5150
rect 28385 5030 28505 5150
rect 28550 5030 28670 5150
rect 28715 5030 28835 5150
rect 28890 5030 29010 5150
rect 29055 5030 29175 5150
rect 29220 5030 29340 5150
rect 29385 5030 29505 5150
rect 29560 5030 29680 5150
rect 24200 4855 24320 4975
rect 24365 4855 24485 4975
rect 24530 4855 24650 4975
rect 24695 4855 24815 4975
rect 24870 4855 24990 4975
rect 25035 4855 25155 4975
rect 25200 4855 25320 4975
rect 25365 4855 25485 4975
rect 25540 4855 25660 4975
rect 25705 4855 25825 4975
rect 25870 4855 25990 4975
rect 26035 4855 26155 4975
rect 26210 4855 26330 4975
rect 26375 4855 26495 4975
rect 26540 4855 26660 4975
rect 26705 4855 26825 4975
rect 26880 4855 27000 4975
rect 27045 4855 27165 4975
rect 27210 4855 27330 4975
rect 27375 4855 27495 4975
rect 27550 4855 27670 4975
rect 27715 4855 27835 4975
rect 27880 4855 28000 4975
rect 28045 4855 28165 4975
rect 28220 4855 28340 4975
rect 28385 4855 28505 4975
rect 28550 4855 28670 4975
rect 28715 4855 28835 4975
rect 28890 4855 29010 4975
rect 29055 4855 29175 4975
rect 29220 4855 29340 4975
rect 29385 4855 29505 4975
rect 29560 4855 29680 4975
rect 24200 4690 24320 4810
rect 24365 4690 24485 4810
rect 24530 4690 24650 4810
rect 24695 4690 24815 4810
rect 24870 4690 24990 4810
rect 25035 4690 25155 4810
rect 25200 4690 25320 4810
rect 25365 4690 25485 4810
rect 25540 4690 25660 4810
rect 25705 4690 25825 4810
rect 25870 4690 25990 4810
rect 26035 4690 26155 4810
rect 26210 4690 26330 4810
rect 26375 4690 26495 4810
rect 26540 4690 26660 4810
rect 26705 4690 26825 4810
rect 26880 4690 27000 4810
rect 27045 4690 27165 4810
rect 27210 4690 27330 4810
rect 27375 4690 27495 4810
rect 27550 4690 27670 4810
rect 27715 4690 27835 4810
rect 27880 4690 28000 4810
rect 28045 4690 28165 4810
rect 28220 4690 28340 4810
rect 28385 4690 28505 4810
rect 28550 4690 28670 4810
rect 28715 4690 28835 4810
rect 28890 4690 29010 4810
rect 29055 4690 29175 4810
rect 29220 4690 29340 4810
rect 29385 4690 29505 4810
rect 29560 4690 29680 4810
rect 24200 4525 24320 4645
rect 24365 4525 24485 4645
rect 24530 4525 24650 4645
rect 24695 4525 24815 4645
rect 24870 4525 24990 4645
rect 25035 4525 25155 4645
rect 25200 4525 25320 4645
rect 25365 4525 25485 4645
rect 25540 4525 25660 4645
rect 25705 4525 25825 4645
rect 25870 4525 25990 4645
rect 26035 4525 26155 4645
rect 26210 4525 26330 4645
rect 26375 4525 26495 4645
rect 26540 4525 26660 4645
rect 26705 4525 26825 4645
rect 26880 4525 27000 4645
rect 27045 4525 27165 4645
rect 27210 4525 27330 4645
rect 27375 4525 27495 4645
rect 27550 4525 27670 4645
rect 27715 4525 27835 4645
rect 27880 4525 28000 4645
rect 28045 4525 28165 4645
rect 28220 4525 28340 4645
rect 28385 4525 28505 4645
rect 28550 4525 28670 4645
rect 28715 4525 28835 4645
rect 28890 4525 29010 4645
rect 29055 4525 29175 4645
rect 29220 4525 29340 4645
rect 29385 4525 29505 4645
rect 29560 4525 29680 4645
rect 24200 4360 24320 4480
rect 24365 4360 24485 4480
rect 24530 4360 24650 4480
rect 24695 4360 24815 4480
rect 24870 4360 24990 4480
rect 25035 4360 25155 4480
rect 25200 4360 25320 4480
rect 25365 4360 25485 4480
rect 25540 4360 25660 4480
rect 25705 4360 25825 4480
rect 25870 4360 25990 4480
rect 26035 4360 26155 4480
rect 26210 4360 26330 4480
rect 26375 4360 26495 4480
rect 26540 4360 26660 4480
rect 26705 4360 26825 4480
rect 26880 4360 27000 4480
rect 27045 4360 27165 4480
rect 27210 4360 27330 4480
rect 27375 4360 27495 4480
rect 27550 4360 27670 4480
rect 27715 4360 27835 4480
rect 27880 4360 28000 4480
rect 28045 4360 28165 4480
rect 28220 4360 28340 4480
rect 28385 4360 28505 4480
rect 28550 4360 28670 4480
rect 28715 4360 28835 4480
rect 28890 4360 29010 4480
rect 29055 4360 29175 4480
rect 29220 4360 29340 4480
rect 29385 4360 29505 4480
rect 29560 4360 29680 4480
rect 24200 4185 24320 4305
rect 24365 4185 24485 4305
rect 24530 4185 24650 4305
rect 24695 4185 24815 4305
rect 24870 4185 24990 4305
rect 25035 4185 25155 4305
rect 25200 4185 25320 4305
rect 25365 4185 25485 4305
rect 25540 4185 25660 4305
rect 25705 4185 25825 4305
rect 25870 4185 25990 4305
rect 26035 4185 26155 4305
rect 26210 4185 26330 4305
rect 26375 4185 26495 4305
rect 26540 4185 26660 4305
rect 26705 4185 26825 4305
rect 26880 4185 27000 4305
rect 27045 4185 27165 4305
rect 27210 4185 27330 4305
rect 27375 4185 27495 4305
rect 27550 4185 27670 4305
rect 27715 4185 27835 4305
rect 27880 4185 28000 4305
rect 28045 4185 28165 4305
rect 28220 4185 28340 4305
rect 28385 4185 28505 4305
rect 28550 4185 28670 4305
rect 28715 4185 28835 4305
rect 28890 4185 29010 4305
rect 29055 4185 29175 4305
rect 29220 4185 29340 4305
rect 29385 4185 29505 4305
rect 29560 4185 29680 4305
rect 24200 4020 24320 4140
rect 24365 4020 24485 4140
rect 24530 4020 24650 4140
rect 24695 4020 24815 4140
rect 24870 4020 24990 4140
rect 25035 4020 25155 4140
rect 25200 4020 25320 4140
rect 25365 4020 25485 4140
rect 25540 4020 25660 4140
rect 25705 4020 25825 4140
rect 25870 4020 25990 4140
rect 26035 4020 26155 4140
rect 26210 4020 26330 4140
rect 26375 4020 26495 4140
rect 26540 4020 26660 4140
rect 26705 4020 26825 4140
rect 26880 4020 27000 4140
rect 27045 4020 27165 4140
rect 27210 4020 27330 4140
rect 27375 4020 27495 4140
rect 27550 4020 27670 4140
rect 27715 4020 27835 4140
rect 27880 4020 28000 4140
rect 28045 4020 28165 4140
rect 28220 4020 28340 4140
rect 28385 4020 28505 4140
rect 28550 4020 28670 4140
rect 28715 4020 28835 4140
rect 28890 4020 29010 4140
rect 29055 4020 29175 4140
rect 29220 4020 29340 4140
rect 29385 4020 29505 4140
rect 29560 4020 29680 4140
rect 24200 3855 24320 3975
rect 24365 3855 24485 3975
rect 24530 3855 24650 3975
rect 24695 3855 24815 3975
rect 24870 3855 24990 3975
rect 25035 3855 25155 3975
rect 25200 3855 25320 3975
rect 25365 3855 25485 3975
rect 25540 3855 25660 3975
rect 25705 3855 25825 3975
rect 25870 3855 25990 3975
rect 26035 3855 26155 3975
rect 26210 3855 26330 3975
rect 26375 3855 26495 3975
rect 26540 3855 26660 3975
rect 26705 3855 26825 3975
rect 26880 3855 27000 3975
rect 27045 3855 27165 3975
rect 27210 3855 27330 3975
rect 27375 3855 27495 3975
rect 27550 3855 27670 3975
rect 27715 3855 27835 3975
rect 27880 3855 28000 3975
rect 28045 3855 28165 3975
rect 28220 3855 28340 3975
rect 28385 3855 28505 3975
rect 28550 3855 28670 3975
rect 28715 3855 28835 3975
rect 28890 3855 29010 3975
rect 29055 3855 29175 3975
rect 29220 3855 29340 3975
rect 29385 3855 29505 3975
rect 29560 3855 29680 3975
rect 24200 3690 24320 3810
rect 24365 3690 24485 3810
rect 24530 3690 24650 3810
rect 24695 3690 24815 3810
rect 24870 3690 24990 3810
rect 25035 3690 25155 3810
rect 25200 3690 25320 3810
rect 25365 3690 25485 3810
rect 25540 3690 25660 3810
rect 25705 3690 25825 3810
rect 25870 3690 25990 3810
rect 26035 3690 26155 3810
rect 26210 3690 26330 3810
rect 26375 3690 26495 3810
rect 26540 3690 26660 3810
rect 26705 3690 26825 3810
rect 26880 3690 27000 3810
rect 27045 3690 27165 3810
rect 27210 3690 27330 3810
rect 27375 3690 27495 3810
rect 27550 3690 27670 3810
rect 27715 3690 27835 3810
rect 27880 3690 28000 3810
rect 28045 3690 28165 3810
rect 28220 3690 28340 3810
rect 28385 3690 28505 3810
rect 28550 3690 28670 3810
rect 28715 3690 28835 3810
rect 28890 3690 29010 3810
rect 29055 3690 29175 3810
rect 29220 3690 29340 3810
rect 29385 3690 29505 3810
rect 29560 3690 29680 3810
rect 24200 3515 24320 3635
rect 24365 3515 24485 3635
rect 24530 3515 24650 3635
rect 24695 3515 24815 3635
rect 24870 3515 24990 3635
rect 25035 3515 25155 3635
rect 25200 3515 25320 3635
rect 25365 3515 25485 3635
rect 25540 3515 25660 3635
rect 25705 3515 25825 3635
rect 25870 3515 25990 3635
rect 26035 3515 26155 3635
rect 26210 3515 26330 3635
rect 26375 3515 26495 3635
rect 26540 3515 26660 3635
rect 26705 3515 26825 3635
rect 26880 3515 27000 3635
rect 27045 3515 27165 3635
rect 27210 3515 27330 3635
rect 27375 3515 27495 3635
rect 27550 3515 27670 3635
rect 27715 3515 27835 3635
rect 27880 3515 28000 3635
rect 28045 3515 28165 3635
rect 28220 3515 28340 3635
rect 28385 3515 28505 3635
rect 28550 3515 28670 3635
rect 28715 3515 28835 3635
rect 28890 3515 29010 3635
rect 29055 3515 29175 3635
rect 29220 3515 29340 3635
rect 29385 3515 29505 3635
rect 29560 3515 29680 3635
rect 24200 3350 24320 3470
rect 24365 3350 24485 3470
rect 24530 3350 24650 3470
rect 24695 3350 24815 3470
rect 24870 3350 24990 3470
rect 25035 3350 25155 3470
rect 25200 3350 25320 3470
rect 25365 3350 25485 3470
rect 25540 3350 25660 3470
rect 25705 3350 25825 3470
rect 25870 3350 25990 3470
rect 26035 3350 26155 3470
rect 26210 3350 26330 3470
rect 26375 3350 26495 3470
rect 26540 3350 26660 3470
rect 26705 3350 26825 3470
rect 26880 3350 27000 3470
rect 27045 3350 27165 3470
rect 27210 3350 27330 3470
rect 27375 3350 27495 3470
rect 27550 3350 27670 3470
rect 27715 3350 27835 3470
rect 27880 3350 28000 3470
rect 28045 3350 28165 3470
rect 28220 3350 28340 3470
rect 28385 3350 28505 3470
rect 28550 3350 28670 3470
rect 28715 3350 28835 3470
rect 28890 3350 29010 3470
rect 29055 3350 29175 3470
rect 29220 3350 29340 3470
rect 29385 3350 29505 3470
rect 29560 3350 29680 3470
rect 24200 3185 24320 3305
rect 24365 3185 24485 3305
rect 24530 3185 24650 3305
rect 24695 3185 24815 3305
rect 24870 3185 24990 3305
rect 25035 3185 25155 3305
rect 25200 3185 25320 3305
rect 25365 3185 25485 3305
rect 25540 3185 25660 3305
rect 25705 3185 25825 3305
rect 25870 3185 25990 3305
rect 26035 3185 26155 3305
rect 26210 3185 26330 3305
rect 26375 3185 26495 3305
rect 26540 3185 26660 3305
rect 26705 3185 26825 3305
rect 26880 3185 27000 3305
rect 27045 3185 27165 3305
rect 27210 3185 27330 3305
rect 27375 3185 27495 3305
rect 27550 3185 27670 3305
rect 27715 3185 27835 3305
rect 27880 3185 28000 3305
rect 28045 3185 28165 3305
rect 28220 3185 28340 3305
rect 28385 3185 28505 3305
rect 28550 3185 28670 3305
rect 28715 3185 28835 3305
rect 28890 3185 29010 3305
rect 29055 3185 29175 3305
rect 29220 3185 29340 3305
rect 29385 3185 29505 3305
rect 29560 3185 29680 3305
rect 24200 3020 24320 3140
rect 24365 3020 24485 3140
rect 24530 3020 24650 3140
rect 24695 3020 24815 3140
rect 24870 3020 24990 3140
rect 25035 3020 25155 3140
rect 25200 3020 25320 3140
rect 25365 3020 25485 3140
rect 25540 3020 25660 3140
rect 25705 3020 25825 3140
rect 25870 3020 25990 3140
rect 26035 3020 26155 3140
rect 26210 3020 26330 3140
rect 26375 3020 26495 3140
rect 26540 3020 26660 3140
rect 26705 3020 26825 3140
rect 26880 3020 27000 3140
rect 27045 3020 27165 3140
rect 27210 3020 27330 3140
rect 27375 3020 27495 3140
rect 27550 3020 27670 3140
rect 27715 3020 27835 3140
rect 27880 3020 28000 3140
rect 28045 3020 28165 3140
rect 28220 3020 28340 3140
rect 28385 3020 28505 3140
rect 28550 3020 28670 3140
rect 28715 3020 28835 3140
rect 28890 3020 29010 3140
rect 29055 3020 29175 3140
rect 29220 3020 29340 3140
rect 29385 3020 29505 3140
rect 29560 3020 29680 3140
rect 24200 2845 24320 2965
rect 24365 2845 24485 2965
rect 24530 2845 24650 2965
rect 24695 2845 24815 2965
rect 24870 2845 24990 2965
rect 25035 2845 25155 2965
rect 25200 2845 25320 2965
rect 25365 2845 25485 2965
rect 25540 2845 25660 2965
rect 25705 2845 25825 2965
rect 25870 2845 25990 2965
rect 26035 2845 26155 2965
rect 26210 2845 26330 2965
rect 26375 2845 26495 2965
rect 26540 2845 26660 2965
rect 26705 2845 26825 2965
rect 26880 2845 27000 2965
rect 27045 2845 27165 2965
rect 27210 2845 27330 2965
rect 27375 2845 27495 2965
rect 27550 2845 27670 2965
rect 27715 2845 27835 2965
rect 27880 2845 28000 2965
rect 28045 2845 28165 2965
rect 28220 2845 28340 2965
rect 28385 2845 28505 2965
rect 28550 2845 28670 2965
rect 28715 2845 28835 2965
rect 28890 2845 29010 2965
rect 29055 2845 29175 2965
rect 29220 2845 29340 2965
rect 29385 2845 29505 2965
rect 29560 2845 29680 2965
rect 24200 2680 24320 2800
rect 24365 2680 24485 2800
rect 24530 2680 24650 2800
rect 24695 2680 24815 2800
rect 24870 2680 24990 2800
rect 25035 2680 25155 2800
rect 25200 2680 25320 2800
rect 25365 2680 25485 2800
rect 25540 2680 25660 2800
rect 25705 2680 25825 2800
rect 25870 2680 25990 2800
rect 26035 2680 26155 2800
rect 26210 2680 26330 2800
rect 26375 2680 26495 2800
rect 26540 2680 26660 2800
rect 26705 2680 26825 2800
rect 26880 2680 27000 2800
rect 27045 2680 27165 2800
rect 27210 2680 27330 2800
rect 27375 2680 27495 2800
rect 27550 2680 27670 2800
rect 27715 2680 27835 2800
rect 27880 2680 28000 2800
rect 28045 2680 28165 2800
rect 28220 2680 28340 2800
rect 28385 2680 28505 2800
rect 28550 2680 28670 2800
rect 28715 2680 28835 2800
rect 28890 2680 29010 2800
rect 29055 2680 29175 2800
rect 29220 2680 29340 2800
rect 29385 2680 29505 2800
rect 29560 2680 29680 2800
rect 24200 2515 24320 2635
rect 24365 2515 24485 2635
rect 24530 2515 24650 2635
rect 24695 2515 24815 2635
rect 24870 2515 24990 2635
rect 25035 2515 25155 2635
rect 25200 2515 25320 2635
rect 25365 2515 25485 2635
rect 25540 2515 25660 2635
rect 25705 2515 25825 2635
rect 25870 2515 25990 2635
rect 26035 2515 26155 2635
rect 26210 2515 26330 2635
rect 26375 2515 26495 2635
rect 26540 2515 26660 2635
rect 26705 2515 26825 2635
rect 26880 2515 27000 2635
rect 27045 2515 27165 2635
rect 27210 2515 27330 2635
rect 27375 2515 27495 2635
rect 27550 2515 27670 2635
rect 27715 2515 27835 2635
rect 27880 2515 28000 2635
rect 28045 2515 28165 2635
rect 28220 2515 28340 2635
rect 28385 2515 28505 2635
rect 28550 2515 28670 2635
rect 28715 2515 28835 2635
rect 28890 2515 29010 2635
rect 29055 2515 29175 2635
rect 29220 2515 29340 2635
rect 29385 2515 29505 2635
rect 29560 2515 29680 2635
rect 24200 2350 24320 2470
rect 24365 2350 24485 2470
rect 24530 2350 24650 2470
rect 24695 2350 24815 2470
rect 24870 2350 24990 2470
rect 25035 2350 25155 2470
rect 25200 2350 25320 2470
rect 25365 2350 25485 2470
rect 25540 2350 25660 2470
rect 25705 2350 25825 2470
rect 25870 2350 25990 2470
rect 26035 2350 26155 2470
rect 26210 2350 26330 2470
rect 26375 2350 26495 2470
rect 26540 2350 26660 2470
rect 26705 2350 26825 2470
rect 26880 2350 27000 2470
rect 27045 2350 27165 2470
rect 27210 2350 27330 2470
rect 27375 2350 27495 2470
rect 27550 2350 27670 2470
rect 27715 2350 27835 2470
rect 27880 2350 28000 2470
rect 28045 2350 28165 2470
rect 28220 2350 28340 2470
rect 28385 2350 28505 2470
rect 28550 2350 28670 2470
rect 28715 2350 28835 2470
rect 28890 2350 29010 2470
rect 29055 2350 29175 2470
rect 29220 2350 29340 2470
rect 29385 2350 29505 2470
rect 29560 2350 29680 2470
rect 24200 2175 24320 2295
rect 24365 2175 24485 2295
rect 24530 2175 24650 2295
rect 24695 2175 24815 2295
rect 24870 2175 24990 2295
rect 25035 2175 25155 2295
rect 25200 2175 25320 2295
rect 25365 2175 25485 2295
rect 25540 2175 25660 2295
rect 25705 2175 25825 2295
rect 25870 2175 25990 2295
rect 26035 2175 26155 2295
rect 26210 2175 26330 2295
rect 26375 2175 26495 2295
rect 26540 2175 26660 2295
rect 26705 2175 26825 2295
rect 26880 2175 27000 2295
rect 27045 2175 27165 2295
rect 27210 2175 27330 2295
rect 27375 2175 27495 2295
rect 27550 2175 27670 2295
rect 27715 2175 27835 2295
rect 27880 2175 28000 2295
rect 28045 2175 28165 2295
rect 28220 2175 28340 2295
rect 28385 2175 28505 2295
rect 28550 2175 28670 2295
rect 28715 2175 28835 2295
rect 28890 2175 29010 2295
rect 29055 2175 29175 2295
rect 29220 2175 29340 2295
rect 29385 2175 29505 2295
rect 29560 2175 29680 2295
rect 24200 2010 24320 2130
rect 24365 2010 24485 2130
rect 24530 2010 24650 2130
rect 24695 2010 24815 2130
rect 24870 2010 24990 2130
rect 25035 2010 25155 2130
rect 25200 2010 25320 2130
rect 25365 2010 25485 2130
rect 25540 2010 25660 2130
rect 25705 2010 25825 2130
rect 25870 2010 25990 2130
rect 26035 2010 26155 2130
rect 26210 2010 26330 2130
rect 26375 2010 26495 2130
rect 26540 2010 26660 2130
rect 26705 2010 26825 2130
rect 26880 2010 27000 2130
rect 27045 2010 27165 2130
rect 27210 2010 27330 2130
rect 27375 2010 27495 2130
rect 27550 2010 27670 2130
rect 27715 2010 27835 2130
rect 27880 2010 28000 2130
rect 28045 2010 28165 2130
rect 28220 2010 28340 2130
rect 28385 2010 28505 2130
rect 28550 2010 28670 2130
rect 28715 2010 28835 2130
rect 28890 2010 29010 2130
rect 29055 2010 29175 2130
rect 29220 2010 29340 2130
rect 29385 2010 29505 2130
rect 29560 2010 29680 2130
rect 24200 1845 24320 1965
rect 24365 1845 24485 1965
rect 24530 1845 24650 1965
rect 24695 1845 24815 1965
rect 24870 1845 24990 1965
rect 25035 1845 25155 1965
rect 25200 1845 25320 1965
rect 25365 1845 25485 1965
rect 25540 1845 25660 1965
rect 25705 1845 25825 1965
rect 25870 1845 25990 1965
rect 26035 1845 26155 1965
rect 26210 1845 26330 1965
rect 26375 1845 26495 1965
rect 26540 1845 26660 1965
rect 26705 1845 26825 1965
rect 26880 1845 27000 1965
rect 27045 1845 27165 1965
rect 27210 1845 27330 1965
rect 27375 1845 27495 1965
rect 27550 1845 27670 1965
rect 27715 1845 27835 1965
rect 27880 1845 28000 1965
rect 28045 1845 28165 1965
rect 28220 1845 28340 1965
rect 28385 1845 28505 1965
rect 28550 1845 28670 1965
rect 28715 1845 28835 1965
rect 28890 1845 29010 1965
rect 29055 1845 29175 1965
rect 29220 1845 29340 1965
rect 29385 1845 29505 1965
rect 29560 1845 29680 1965
rect 24200 1680 24320 1800
rect 24365 1680 24485 1800
rect 24530 1680 24650 1800
rect 24695 1680 24815 1800
rect 24870 1680 24990 1800
rect 25035 1680 25155 1800
rect 25200 1680 25320 1800
rect 25365 1680 25485 1800
rect 25540 1680 25660 1800
rect 25705 1680 25825 1800
rect 25870 1680 25990 1800
rect 26035 1680 26155 1800
rect 26210 1680 26330 1800
rect 26375 1680 26495 1800
rect 26540 1680 26660 1800
rect 26705 1680 26825 1800
rect 26880 1680 27000 1800
rect 27045 1680 27165 1800
rect 27210 1680 27330 1800
rect 27375 1680 27495 1800
rect 27550 1680 27670 1800
rect 27715 1680 27835 1800
rect 27880 1680 28000 1800
rect 28045 1680 28165 1800
rect 28220 1680 28340 1800
rect 28385 1680 28505 1800
rect 28550 1680 28670 1800
rect 28715 1680 28835 1800
rect 28890 1680 29010 1800
rect 29055 1680 29175 1800
rect 29220 1680 29340 1800
rect 29385 1680 29505 1800
rect 29560 1680 29680 1800
rect 7130 1260 7250 1380
rect 7305 1260 7425 1380
rect 7470 1260 7590 1380
rect 7635 1260 7755 1380
rect 7800 1260 7920 1380
rect 7975 1260 8095 1380
rect 8140 1260 8260 1380
rect 8305 1260 8425 1380
rect 8470 1260 8590 1380
rect 8645 1260 8765 1380
rect 8810 1260 8930 1380
rect 8975 1260 9095 1380
rect 9140 1260 9260 1380
rect 9315 1260 9435 1380
rect 9480 1260 9600 1380
rect 9645 1260 9765 1380
rect 9810 1260 9930 1380
rect 9985 1260 10105 1380
rect 10150 1260 10270 1380
rect 10315 1260 10435 1380
rect 10480 1260 10600 1380
rect 10655 1260 10775 1380
rect 10820 1260 10940 1380
rect 10985 1260 11105 1380
rect 11150 1260 11270 1380
rect 11325 1260 11445 1380
rect 11490 1260 11610 1380
rect 11655 1260 11775 1380
rect 11820 1260 11940 1380
rect 11995 1260 12115 1380
rect 12160 1260 12280 1380
rect 12325 1260 12445 1380
rect 12490 1260 12610 1380
rect 7130 1095 7250 1215
rect 7305 1095 7425 1215
rect 7470 1095 7590 1215
rect 7635 1095 7755 1215
rect 7800 1095 7920 1215
rect 7975 1095 8095 1215
rect 8140 1095 8260 1215
rect 8305 1095 8425 1215
rect 8470 1095 8590 1215
rect 8645 1095 8765 1215
rect 8810 1095 8930 1215
rect 8975 1095 9095 1215
rect 9140 1095 9260 1215
rect 9315 1095 9435 1215
rect 9480 1095 9600 1215
rect 9645 1095 9765 1215
rect 9810 1095 9930 1215
rect 9985 1095 10105 1215
rect 10150 1095 10270 1215
rect 10315 1095 10435 1215
rect 10480 1095 10600 1215
rect 10655 1095 10775 1215
rect 10820 1095 10940 1215
rect 10985 1095 11105 1215
rect 11150 1095 11270 1215
rect 11325 1095 11445 1215
rect 11490 1095 11610 1215
rect 11655 1095 11775 1215
rect 11820 1095 11940 1215
rect 11995 1095 12115 1215
rect 12160 1095 12280 1215
rect 12325 1095 12445 1215
rect 12490 1095 12610 1215
rect 7130 930 7250 1050
rect 7305 930 7425 1050
rect 7470 930 7590 1050
rect 7635 930 7755 1050
rect 7800 930 7920 1050
rect 7975 930 8095 1050
rect 8140 930 8260 1050
rect 8305 930 8425 1050
rect 8470 930 8590 1050
rect 8645 930 8765 1050
rect 8810 930 8930 1050
rect 8975 930 9095 1050
rect 9140 930 9260 1050
rect 9315 930 9435 1050
rect 9480 930 9600 1050
rect 9645 930 9765 1050
rect 9810 930 9930 1050
rect 9985 930 10105 1050
rect 10150 930 10270 1050
rect 10315 930 10435 1050
rect 10480 930 10600 1050
rect 10655 930 10775 1050
rect 10820 930 10940 1050
rect 10985 930 11105 1050
rect 11150 930 11270 1050
rect 11325 930 11445 1050
rect 11490 930 11610 1050
rect 11655 930 11775 1050
rect 11820 930 11940 1050
rect 11995 930 12115 1050
rect 12160 930 12280 1050
rect 12325 930 12445 1050
rect 12490 930 12610 1050
rect 7130 765 7250 885
rect 7305 765 7425 885
rect 7470 765 7590 885
rect 7635 765 7755 885
rect 7800 765 7920 885
rect 7975 765 8095 885
rect 8140 765 8260 885
rect 8305 765 8425 885
rect 8470 765 8590 885
rect 8645 765 8765 885
rect 8810 765 8930 885
rect 8975 765 9095 885
rect 9140 765 9260 885
rect 9315 765 9435 885
rect 9480 765 9600 885
rect 9645 765 9765 885
rect 9810 765 9930 885
rect 9985 765 10105 885
rect 10150 765 10270 885
rect 10315 765 10435 885
rect 10480 765 10600 885
rect 10655 765 10775 885
rect 10820 765 10940 885
rect 10985 765 11105 885
rect 11150 765 11270 885
rect 11325 765 11445 885
rect 11490 765 11610 885
rect 11655 765 11775 885
rect 11820 765 11940 885
rect 11995 765 12115 885
rect 12160 765 12280 885
rect 12325 765 12445 885
rect 12490 765 12610 885
rect 7130 590 7250 710
rect 7305 590 7425 710
rect 7470 590 7590 710
rect 7635 590 7755 710
rect 7800 590 7920 710
rect 7975 590 8095 710
rect 8140 590 8260 710
rect 8305 590 8425 710
rect 8470 590 8590 710
rect 8645 590 8765 710
rect 8810 590 8930 710
rect 8975 590 9095 710
rect 9140 590 9260 710
rect 9315 590 9435 710
rect 9480 590 9600 710
rect 9645 590 9765 710
rect 9810 590 9930 710
rect 9985 590 10105 710
rect 10150 590 10270 710
rect 10315 590 10435 710
rect 10480 590 10600 710
rect 10655 590 10775 710
rect 10820 590 10940 710
rect 10985 590 11105 710
rect 11150 590 11270 710
rect 11325 590 11445 710
rect 11490 590 11610 710
rect 11655 590 11775 710
rect 11820 590 11940 710
rect 11995 590 12115 710
rect 12160 590 12280 710
rect 12325 590 12445 710
rect 12490 590 12610 710
rect 7130 425 7250 545
rect 7305 425 7425 545
rect 7470 425 7590 545
rect 7635 425 7755 545
rect 7800 425 7920 545
rect 7975 425 8095 545
rect 8140 425 8260 545
rect 8305 425 8425 545
rect 8470 425 8590 545
rect 8645 425 8765 545
rect 8810 425 8930 545
rect 8975 425 9095 545
rect 9140 425 9260 545
rect 9315 425 9435 545
rect 9480 425 9600 545
rect 9645 425 9765 545
rect 9810 425 9930 545
rect 9985 425 10105 545
rect 10150 425 10270 545
rect 10315 425 10435 545
rect 10480 425 10600 545
rect 10655 425 10775 545
rect 10820 425 10940 545
rect 10985 425 11105 545
rect 11150 425 11270 545
rect 11325 425 11445 545
rect 11490 425 11610 545
rect 11655 425 11775 545
rect 11820 425 11940 545
rect 11995 425 12115 545
rect 12160 425 12280 545
rect 12325 425 12445 545
rect 12490 425 12610 545
rect 7130 260 7250 380
rect 7305 260 7425 380
rect 7470 260 7590 380
rect 7635 260 7755 380
rect 7800 260 7920 380
rect 7975 260 8095 380
rect 8140 260 8260 380
rect 8305 260 8425 380
rect 8470 260 8590 380
rect 8645 260 8765 380
rect 8810 260 8930 380
rect 8975 260 9095 380
rect 9140 260 9260 380
rect 9315 260 9435 380
rect 9480 260 9600 380
rect 9645 260 9765 380
rect 9810 260 9930 380
rect 9985 260 10105 380
rect 10150 260 10270 380
rect 10315 260 10435 380
rect 10480 260 10600 380
rect 10655 260 10775 380
rect 10820 260 10940 380
rect 10985 260 11105 380
rect 11150 260 11270 380
rect 11325 260 11445 380
rect 11490 260 11610 380
rect 11655 260 11775 380
rect 11820 260 11940 380
rect 11995 260 12115 380
rect 12160 260 12280 380
rect 12325 260 12445 380
rect 12490 260 12610 380
rect 7130 95 7250 215
rect 7305 95 7425 215
rect 7470 95 7590 215
rect 7635 95 7755 215
rect 7800 95 7920 215
rect 7975 95 8095 215
rect 8140 95 8260 215
rect 8305 95 8425 215
rect 8470 95 8590 215
rect 8645 95 8765 215
rect 8810 95 8930 215
rect 8975 95 9095 215
rect 9140 95 9260 215
rect 9315 95 9435 215
rect 9480 95 9600 215
rect 9645 95 9765 215
rect 9810 95 9930 215
rect 9985 95 10105 215
rect 10150 95 10270 215
rect 10315 95 10435 215
rect 10480 95 10600 215
rect 10655 95 10775 215
rect 10820 95 10940 215
rect 10985 95 11105 215
rect 11150 95 11270 215
rect 11325 95 11445 215
rect 11490 95 11610 215
rect 11655 95 11775 215
rect 11820 95 11940 215
rect 11995 95 12115 215
rect 12160 95 12280 215
rect 12325 95 12445 215
rect 12490 95 12610 215
rect 7130 -80 7250 40
rect 7305 -80 7425 40
rect 7470 -80 7590 40
rect 7635 -80 7755 40
rect 7800 -80 7920 40
rect 7975 -80 8095 40
rect 8140 -80 8260 40
rect 8305 -80 8425 40
rect 8470 -80 8590 40
rect 8645 -80 8765 40
rect 8810 -80 8930 40
rect 8975 -80 9095 40
rect 9140 -80 9260 40
rect 9315 -80 9435 40
rect 9480 -80 9600 40
rect 9645 -80 9765 40
rect 9810 -80 9930 40
rect 9985 -80 10105 40
rect 10150 -80 10270 40
rect 10315 -80 10435 40
rect 10480 -80 10600 40
rect 10655 -80 10775 40
rect 10820 -80 10940 40
rect 10985 -80 11105 40
rect 11150 -80 11270 40
rect 11325 -80 11445 40
rect 11490 -80 11610 40
rect 11655 -80 11775 40
rect 11820 -80 11940 40
rect 11995 -80 12115 40
rect 12160 -80 12280 40
rect 12325 -80 12445 40
rect 12490 -80 12610 40
rect 7130 -245 7250 -125
rect 7305 -245 7425 -125
rect 7470 -245 7590 -125
rect 7635 -245 7755 -125
rect 7800 -245 7920 -125
rect 7975 -245 8095 -125
rect 8140 -245 8260 -125
rect 8305 -245 8425 -125
rect 8470 -245 8590 -125
rect 8645 -245 8765 -125
rect 8810 -245 8930 -125
rect 8975 -245 9095 -125
rect 9140 -245 9260 -125
rect 9315 -245 9435 -125
rect 9480 -245 9600 -125
rect 9645 -245 9765 -125
rect 9810 -245 9930 -125
rect 9985 -245 10105 -125
rect 10150 -245 10270 -125
rect 10315 -245 10435 -125
rect 10480 -245 10600 -125
rect 10655 -245 10775 -125
rect 10820 -245 10940 -125
rect 10985 -245 11105 -125
rect 11150 -245 11270 -125
rect 11325 -245 11445 -125
rect 11490 -245 11610 -125
rect 11655 -245 11775 -125
rect 11820 -245 11940 -125
rect 11995 -245 12115 -125
rect 12160 -245 12280 -125
rect 12325 -245 12445 -125
rect 12490 -245 12610 -125
rect 7130 -410 7250 -290
rect 7305 -410 7425 -290
rect 7470 -410 7590 -290
rect 7635 -410 7755 -290
rect 7800 -410 7920 -290
rect 7975 -410 8095 -290
rect 8140 -410 8260 -290
rect 8305 -410 8425 -290
rect 8470 -410 8590 -290
rect 8645 -410 8765 -290
rect 8810 -410 8930 -290
rect 8975 -410 9095 -290
rect 9140 -410 9260 -290
rect 9315 -410 9435 -290
rect 9480 -410 9600 -290
rect 9645 -410 9765 -290
rect 9810 -410 9930 -290
rect 9985 -410 10105 -290
rect 10150 -410 10270 -290
rect 10315 -410 10435 -290
rect 10480 -410 10600 -290
rect 10655 -410 10775 -290
rect 10820 -410 10940 -290
rect 10985 -410 11105 -290
rect 11150 -410 11270 -290
rect 11325 -410 11445 -290
rect 11490 -410 11610 -290
rect 11655 -410 11775 -290
rect 11820 -410 11940 -290
rect 11995 -410 12115 -290
rect 12160 -410 12280 -290
rect 12325 -410 12445 -290
rect 12490 -410 12610 -290
rect 7130 -575 7250 -455
rect 7305 -575 7425 -455
rect 7470 -575 7590 -455
rect 7635 -575 7755 -455
rect 7800 -575 7920 -455
rect 7975 -575 8095 -455
rect 8140 -575 8260 -455
rect 8305 -575 8425 -455
rect 8470 -575 8590 -455
rect 8645 -575 8765 -455
rect 8810 -575 8930 -455
rect 8975 -575 9095 -455
rect 9140 -575 9260 -455
rect 9315 -575 9435 -455
rect 9480 -575 9600 -455
rect 9645 -575 9765 -455
rect 9810 -575 9930 -455
rect 9985 -575 10105 -455
rect 10150 -575 10270 -455
rect 10315 -575 10435 -455
rect 10480 -575 10600 -455
rect 10655 -575 10775 -455
rect 10820 -575 10940 -455
rect 10985 -575 11105 -455
rect 11150 -575 11270 -455
rect 11325 -575 11445 -455
rect 11490 -575 11610 -455
rect 11655 -575 11775 -455
rect 11820 -575 11940 -455
rect 11995 -575 12115 -455
rect 12160 -575 12280 -455
rect 12325 -575 12445 -455
rect 12490 -575 12610 -455
rect 7130 -750 7250 -630
rect 7305 -750 7425 -630
rect 7470 -750 7590 -630
rect 7635 -750 7755 -630
rect 7800 -750 7920 -630
rect 7975 -750 8095 -630
rect 8140 -750 8260 -630
rect 8305 -750 8425 -630
rect 8470 -750 8590 -630
rect 8645 -750 8765 -630
rect 8810 -750 8930 -630
rect 8975 -750 9095 -630
rect 9140 -750 9260 -630
rect 9315 -750 9435 -630
rect 9480 -750 9600 -630
rect 9645 -750 9765 -630
rect 9810 -750 9930 -630
rect 9985 -750 10105 -630
rect 10150 -750 10270 -630
rect 10315 -750 10435 -630
rect 10480 -750 10600 -630
rect 10655 -750 10775 -630
rect 10820 -750 10940 -630
rect 10985 -750 11105 -630
rect 11150 -750 11270 -630
rect 11325 -750 11445 -630
rect 11490 -750 11610 -630
rect 11655 -750 11775 -630
rect 11820 -750 11940 -630
rect 11995 -750 12115 -630
rect 12160 -750 12280 -630
rect 12325 -750 12445 -630
rect 12490 -750 12610 -630
rect 7130 -915 7250 -795
rect 7305 -915 7425 -795
rect 7470 -915 7590 -795
rect 7635 -915 7755 -795
rect 7800 -915 7920 -795
rect 7975 -915 8095 -795
rect 8140 -915 8260 -795
rect 8305 -915 8425 -795
rect 8470 -915 8590 -795
rect 8645 -915 8765 -795
rect 8810 -915 8930 -795
rect 8975 -915 9095 -795
rect 9140 -915 9260 -795
rect 9315 -915 9435 -795
rect 9480 -915 9600 -795
rect 9645 -915 9765 -795
rect 9810 -915 9930 -795
rect 9985 -915 10105 -795
rect 10150 -915 10270 -795
rect 10315 -915 10435 -795
rect 10480 -915 10600 -795
rect 10655 -915 10775 -795
rect 10820 -915 10940 -795
rect 10985 -915 11105 -795
rect 11150 -915 11270 -795
rect 11325 -915 11445 -795
rect 11490 -915 11610 -795
rect 11655 -915 11775 -795
rect 11820 -915 11940 -795
rect 11995 -915 12115 -795
rect 12160 -915 12280 -795
rect 12325 -915 12445 -795
rect 12490 -915 12610 -795
rect 7130 -1080 7250 -960
rect 7305 -1080 7425 -960
rect 7470 -1080 7590 -960
rect 7635 -1080 7755 -960
rect 7800 -1080 7920 -960
rect 7975 -1080 8095 -960
rect 8140 -1080 8260 -960
rect 8305 -1080 8425 -960
rect 8470 -1080 8590 -960
rect 8645 -1080 8765 -960
rect 8810 -1080 8930 -960
rect 8975 -1080 9095 -960
rect 9140 -1080 9260 -960
rect 9315 -1080 9435 -960
rect 9480 -1080 9600 -960
rect 9645 -1080 9765 -960
rect 9810 -1080 9930 -960
rect 9985 -1080 10105 -960
rect 10150 -1080 10270 -960
rect 10315 -1080 10435 -960
rect 10480 -1080 10600 -960
rect 10655 -1080 10775 -960
rect 10820 -1080 10940 -960
rect 10985 -1080 11105 -960
rect 11150 -1080 11270 -960
rect 11325 -1080 11445 -960
rect 11490 -1080 11610 -960
rect 11655 -1080 11775 -960
rect 11820 -1080 11940 -960
rect 11995 -1080 12115 -960
rect 12160 -1080 12280 -960
rect 12325 -1080 12445 -960
rect 12490 -1080 12610 -960
rect 7130 -1245 7250 -1125
rect 7305 -1245 7425 -1125
rect 7470 -1245 7590 -1125
rect 7635 -1245 7755 -1125
rect 7800 -1245 7920 -1125
rect 7975 -1245 8095 -1125
rect 8140 -1245 8260 -1125
rect 8305 -1245 8425 -1125
rect 8470 -1245 8590 -1125
rect 8645 -1245 8765 -1125
rect 8810 -1245 8930 -1125
rect 8975 -1245 9095 -1125
rect 9140 -1245 9260 -1125
rect 9315 -1245 9435 -1125
rect 9480 -1245 9600 -1125
rect 9645 -1245 9765 -1125
rect 9810 -1245 9930 -1125
rect 9985 -1245 10105 -1125
rect 10150 -1245 10270 -1125
rect 10315 -1245 10435 -1125
rect 10480 -1245 10600 -1125
rect 10655 -1245 10775 -1125
rect 10820 -1245 10940 -1125
rect 10985 -1245 11105 -1125
rect 11150 -1245 11270 -1125
rect 11325 -1245 11445 -1125
rect 11490 -1245 11610 -1125
rect 11655 -1245 11775 -1125
rect 11820 -1245 11940 -1125
rect 11995 -1245 12115 -1125
rect 12160 -1245 12280 -1125
rect 12325 -1245 12445 -1125
rect 12490 -1245 12610 -1125
rect 7130 -1420 7250 -1300
rect 7305 -1420 7425 -1300
rect 7470 -1420 7590 -1300
rect 7635 -1420 7755 -1300
rect 7800 -1420 7920 -1300
rect 7975 -1420 8095 -1300
rect 8140 -1420 8260 -1300
rect 8305 -1420 8425 -1300
rect 8470 -1420 8590 -1300
rect 8645 -1420 8765 -1300
rect 8810 -1420 8930 -1300
rect 8975 -1420 9095 -1300
rect 9140 -1420 9260 -1300
rect 9315 -1420 9435 -1300
rect 9480 -1420 9600 -1300
rect 9645 -1420 9765 -1300
rect 9810 -1420 9930 -1300
rect 9985 -1420 10105 -1300
rect 10150 -1420 10270 -1300
rect 10315 -1420 10435 -1300
rect 10480 -1420 10600 -1300
rect 10655 -1420 10775 -1300
rect 10820 -1420 10940 -1300
rect 10985 -1420 11105 -1300
rect 11150 -1420 11270 -1300
rect 11325 -1420 11445 -1300
rect 11490 -1420 11610 -1300
rect 11655 -1420 11775 -1300
rect 11820 -1420 11940 -1300
rect 11995 -1420 12115 -1300
rect 12160 -1420 12280 -1300
rect 12325 -1420 12445 -1300
rect 12490 -1420 12610 -1300
rect 7130 -1585 7250 -1465
rect 7305 -1585 7425 -1465
rect 7470 -1585 7590 -1465
rect 7635 -1585 7755 -1465
rect 7800 -1585 7920 -1465
rect 7975 -1585 8095 -1465
rect 8140 -1585 8260 -1465
rect 8305 -1585 8425 -1465
rect 8470 -1585 8590 -1465
rect 8645 -1585 8765 -1465
rect 8810 -1585 8930 -1465
rect 8975 -1585 9095 -1465
rect 9140 -1585 9260 -1465
rect 9315 -1585 9435 -1465
rect 9480 -1585 9600 -1465
rect 9645 -1585 9765 -1465
rect 9810 -1585 9930 -1465
rect 9985 -1585 10105 -1465
rect 10150 -1585 10270 -1465
rect 10315 -1585 10435 -1465
rect 10480 -1585 10600 -1465
rect 10655 -1585 10775 -1465
rect 10820 -1585 10940 -1465
rect 10985 -1585 11105 -1465
rect 11150 -1585 11270 -1465
rect 11325 -1585 11445 -1465
rect 11490 -1585 11610 -1465
rect 11655 -1585 11775 -1465
rect 11820 -1585 11940 -1465
rect 11995 -1585 12115 -1465
rect 12160 -1585 12280 -1465
rect 12325 -1585 12445 -1465
rect 12490 -1585 12610 -1465
rect 7130 -1750 7250 -1630
rect 7305 -1750 7425 -1630
rect 7470 -1750 7590 -1630
rect 7635 -1750 7755 -1630
rect 7800 -1750 7920 -1630
rect 7975 -1750 8095 -1630
rect 8140 -1750 8260 -1630
rect 8305 -1750 8425 -1630
rect 8470 -1750 8590 -1630
rect 8645 -1750 8765 -1630
rect 8810 -1750 8930 -1630
rect 8975 -1750 9095 -1630
rect 9140 -1750 9260 -1630
rect 9315 -1750 9435 -1630
rect 9480 -1750 9600 -1630
rect 9645 -1750 9765 -1630
rect 9810 -1750 9930 -1630
rect 9985 -1750 10105 -1630
rect 10150 -1750 10270 -1630
rect 10315 -1750 10435 -1630
rect 10480 -1750 10600 -1630
rect 10655 -1750 10775 -1630
rect 10820 -1750 10940 -1630
rect 10985 -1750 11105 -1630
rect 11150 -1750 11270 -1630
rect 11325 -1750 11445 -1630
rect 11490 -1750 11610 -1630
rect 11655 -1750 11775 -1630
rect 11820 -1750 11940 -1630
rect 11995 -1750 12115 -1630
rect 12160 -1750 12280 -1630
rect 12325 -1750 12445 -1630
rect 12490 -1750 12610 -1630
rect 7130 -1915 7250 -1795
rect 7305 -1915 7425 -1795
rect 7470 -1915 7590 -1795
rect 7635 -1915 7755 -1795
rect 7800 -1915 7920 -1795
rect 7975 -1915 8095 -1795
rect 8140 -1915 8260 -1795
rect 8305 -1915 8425 -1795
rect 8470 -1915 8590 -1795
rect 8645 -1915 8765 -1795
rect 8810 -1915 8930 -1795
rect 8975 -1915 9095 -1795
rect 9140 -1915 9260 -1795
rect 9315 -1915 9435 -1795
rect 9480 -1915 9600 -1795
rect 9645 -1915 9765 -1795
rect 9810 -1915 9930 -1795
rect 9985 -1915 10105 -1795
rect 10150 -1915 10270 -1795
rect 10315 -1915 10435 -1795
rect 10480 -1915 10600 -1795
rect 10655 -1915 10775 -1795
rect 10820 -1915 10940 -1795
rect 10985 -1915 11105 -1795
rect 11150 -1915 11270 -1795
rect 11325 -1915 11445 -1795
rect 11490 -1915 11610 -1795
rect 11655 -1915 11775 -1795
rect 11820 -1915 11940 -1795
rect 11995 -1915 12115 -1795
rect 12160 -1915 12280 -1795
rect 12325 -1915 12445 -1795
rect 12490 -1915 12610 -1795
rect 7130 -2090 7250 -1970
rect 7305 -2090 7425 -1970
rect 7470 -2090 7590 -1970
rect 7635 -2090 7755 -1970
rect 7800 -2090 7920 -1970
rect 7975 -2090 8095 -1970
rect 8140 -2090 8260 -1970
rect 8305 -2090 8425 -1970
rect 8470 -2090 8590 -1970
rect 8645 -2090 8765 -1970
rect 8810 -2090 8930 -1970
rect 8975 -2090 9095 -1970
rect 9140 -2090 9260 -1970
rect 9315 -2090 9435 -1970
rect 9480 -2090 9600 -1970
rect 9645 -2090 9765 -1970
rect 9810 -2090 9930 -1970
rect 9985 -2090 10105 -1970
rect 10150 -2090 10270 -1970
rect 10315 -2090 10435 -1970
rect 10480 -2090 10600 -1970
rect 10655 -2090 10775 -1970
rect 10820 -2090 10940 -1970
rect 10985 -2090 11105 -1970
rect 11150 -2090 11270 -1970
rect 11325 -2090 11445 -1970
rect 11490 -2090 11610 -1970
rect 11655 -2090 11775 -1970
rect 11820 -2090 11940 -1970
rect 11995 -2090 12115 -1970
rect 12160 -2090 12280 -1970
rect 12325 -2090 12445 -1970
rect 12490 -2090 12610 -1970
rect 7130 -2255 7250 -2135
rect 7305 -2255 7425 -2135
rect 7470 -2255 7590 -2135
rect 7635 -2255 7755 -2135
rect 7800 -2255 7920 -2135
rect 7975 -2255 8095 -2135
rect 8140 -2255 8260 -2135
rect 8305 -2255 8425 -2135
rect 8470 -2255 8590 -2135
rect 8645 -2255 8765 -2135
rect 8810 -2255 8930 -2135
rect 8975 -2255 9095 -2135
rect 9140 -2255 9260 -2135
rect 9315 -2255 9435 -2135
rect 9480 -2255 9600 -2135
rect 9645 -2255 9765 -2135
rect 9810 -2255 9930 -2135
rect 9985 -2255 10105 -2135
rect 10150 -2255 10270 -2135
rect 10315 -2255 10435 -2135
rect 10480 -2255 10600 -2135
rect 10655 -2255 10775 -2135
rect 10820 -2255 10940 -2135
rect 10985 -2255 11105 -2135
rect 11150 -2255 11270 -2135
rect 11325 -2255 11445 -2135
rect 11490 -2255 11610 -2135
rect 11655 -2255 11775 -2135
rect 11820 -2255 11940 -2135
rect 11995 -2255 12115 -2135
rect 12160 -2255 12280 -2135
rect 12325 -2255 12445 -2135
rect 12490 -2255 12610 -2135
rect 7130 -2420 7250 -2300
rect 7305 -2420 7425 -2300
rect 7470 -2420 7590 -2300
rect 7635 -2420 7755 -2300
rect 7800 -2420 7920 -2300
rect 7975 -2420 8095 -2300
rect 8140 -2420 8260 -2300
rect 8305 -2420 8425 -2300
rect 8470 -2420 8590 -2300
rect 8645 -2420 8765 -2300
rect 8810 -2420 8930 -2300
rect 8975 -2420 9095 -2300
rect 9140 -2420 9260 -2300
rect 9315 -2420 9435 -2300
rect 9480 -2420 9600 -2300
rect 9645 -2420 9765 -2300
rect 9810 -2420 9930 -2300
rect 9985 -2420 10105 -2300
rect 10150 -2420 10270 -2300
rect 10315 -2420 10435 -2300
rect 10480 -2420 10600 -2300
rect 10655 -2420 10775 -2300
rect 10820 -2420 10940 -2300
rect 10985 -2420 11105 -2300
rect 11150 -2420 11270 -2300
rect 11325 -2420 11445 -2300
rect 11490 -2420 11610 -2300
rect 11655 -2420 11775 -2300
rect 11820 -2420 11940 -2300
rect 11995 -2420 12115 -2300
rect 12160 -2420 12280 -2300
rect 12325 -2420 12445 -2300
rect 12490 -2420 12610 -2300
rect 7130 -2585 7250 -2465
rect 7305 -2585 7425 -2465
rect 7470 -2585 7590 -2465
rect 7635 -2585 7755 -2465
rect 7800 -2585 7920 -2465
rect 7975 -2585 8095 -2465
rect 8140 -2585 8260 -2465
rect 8305 -2585 8425 -2465
rect 8470 -2585 8590 -2465
rect 8645 -2585 8765 -2465
rect 8810 -2585 8930 -2465
rect 8975 -2585 9095 -2465
rect 9140 -2585 9260 -2465
rect 9315 -2585 9435 -2465
rect 9480 -2585 9600 -2465
rect 9645 -2585 9765 -2465
rect 9810 -2585 9930 -2465
rect 9985 -2585 10105 -2465
rect 10150 -2585 10270 -2465
rect 10315 -2585 10435 -2465
rect 10480 -2585 10600 -2465
rect 10655 -2585 10775 -2465
rect 10820 -2585 10940 -2465
rect 10985 -2585 11105 -2465
rect 11150 -2585 11270 -2465
rect 11325 -2585 11445 -2465
rect 11490 -2585 11610 -2465
rect 11655 -2585 11775 -2465
rect 11820 -2585 11940 -2465
rect 11995 -2585 12115 -2465
rect 12160 -2585 12280 -2465
rect 12325 -2585 12445 -2465
rect 12490 -2585 12610 -2465
rect 7130 -2760 7250 -2640
rect 7305 -2760 7425 -2640
rect 7470 -2760 7590 -2640
rect 7635 -2760 7755 -2640
rect 7800 -2760 7920 -2640
rect 7975 -2760 8095 -2640
rect 8140 -2760 8260 -2640
rect 8305 -2760 8425 -2640
rect 8470 -2760 8590 -2640
rect 8645 -2760 8765 -2640
rect 8810 -2760 8930 -2640
rect 8975 -2760 9095 -2640
rect 9140 -2760 9260 -2640
rect 9315 -2760 9435 -2640
rect 9480 -2760 9600 -2640
rect 9645 -2760 9765 -2640
rect 9810 -2760 9930 -2640
rect 9985 -2760 10105 -2640
rect 10150 -2760 10270 -2640
rect 10315 -2760 10435 -2640
rect 10480 -2760 10600 -2640
rect 10655 -2760 10775 -2640
rect 10820 -2760 10940 -2640
rect 10985 -2760 11105 -2640
rect 11150 -2760 11270 -2640
rect 11325 -2760 11445 -2640
rect 11490 -2760 11610 -2640
rect 11655 -2760 11775 -2640
rect 11820 -2760 11940 -2640
rect 11995 -2760 12115 -2640
rect 12160 -2760 12280 -2640
rect 12325 -2760 12445 -2640
rect 12490 -2760 12610 -2640
rect 7130 -2925 7250 -2805
rect 7305 -2925 7425 -2805
rect 7470 -2925 7590 -2805
rect 7635 -2925 7755 -2805
rect 7800 -2925 7920 -2805
rect 7975 -2925 8095 -2805
rect 8140 -2925 8260 -2805
rect 8305 -2925 8425 -2805
rect 8470 -2925 8590 -2805
rect 8645 -2925 8765 -2805
rect 8810 -2925 8930 -2805
rect 8975 -2925 9095 -2805
rect 9140 -2925 9260 -2805
rect 9315 -2925 9435 -2805
rect 9480 -2925 9600 -2805
rect 9645 -2925 9765 -2805
rect 9810 -2925 9930 -2805
rect 9985 -2925 10105 -2805
rect 10150 -2925 10270 -2805
rect 10315 -2925 10435 -2805
rect 10480 -2925 10600 -2805
rect 10655 -2925 10775 -2805
rect 10820 -2925 10940 -2805
rect 10985 -2925 11105 -2805
rect 11150 -2925 11270 -2805
rect 11325 -2925 11445 -2805
rect 11490 -2925 11610 -2805
rect 11655 -2925 11775 -2805
rect 11820 -2925 11940 -2805
rect 11995 -2925 12115 -2805
rect 12160 -2925 12280 -2805
rect 12325 -2925 12445 -2805
rect 12490 -2925 12610 -2805
rect 7130 -3090 7250 -2970
rect 7305 -3090 7425 -2970
rect 7470 -3090 7590 -2970
rect 7635 -3090 7755 -2970
rect 7800 -3090 7920 -2970
rect 7975 -3090 8095 -2970
rect 8140 -3090 8260 -2970
rect 8305 -3090 8425 -2970
rect 8470 -3090 8590 -2970
rect 8645 -3090 8765 -2970
rect 8810 -3090 8930 -2970
rect 8975 -3090 9095 -2970
rect 9140 -3090 9260 -2970
rect 9315 -3090 9435 -2970
rect 9480 -3090 9600 -2970
rect 9645 -3090 9765 -2970
rect 9810 -3090 9930 -2970
rect 9985 -3090 10105 -2970
rect 10150 -3090 10270 -2970
rect 10315 -3090 10435 -2970
rect 10480 -3090 10600 -2970
rect 10655 -3090 10775 -2970
rect 10820 -3090 10940 -2970
rect 10985 -3090 11105 -2970
rect 11150 -3090 11270 -2970
rect 11325 -3090 11445 -2970
rect 11490 -3090 11610 -2970
rect 11655 -3090 11775 -2970
rect 11820 -3090 11940 -2970
rect 11995 -3090 12115 -2970
rect 12160 -3090 12280 -2970
rect 12325 -3090 12445 -2970
rect 12490 -3090 12610 -2970
rect 7130 -3255 7250 -3135
rect 7305 -3255 7425 -3135
rect 7470 -3255 7590 -3135
rect 7635 -3255 7755 -3135
rect 7800 -3255 7920 -3135
rect 7975 -3255 8095 -3135
rect 8140 -3255 8260 -3135
rect 8305 -3255 8425 -3135
rect 8470 -3255 8590 -3135
rect 8645 -3255 8765 -3135
rect 8810 -3255 8930 -3135
rect 8975 -3255 9095 -3135
rect 9140 -3255 9260 -3135
rect 9315 -3255 9435 -3135
rect 9480 -3255 9600 -3135
rect 9645 -3255 9765 -3135
rect 9810 -3255 9930 -3135
rect 9985 -3255 10105 -3135
rect 10150 -3255 10270 -3135
rect 10315 -3255 10435 -3135
rect 10480 -3255 10600 -3135
rect 10655 -3255 10775 -3135
rect 10820 -3255 10940 -3135
rect 10985 -3255 11105 -3135
rect 11150 -3255 11270 -3135
rect 11325 -3255 11445 -3135
rect 11490 -3255 11610 -3135
rect 11655 -3255 11775 -3135
rect 11820 -3255 11940 -3135
rect 11995 -3255 12115 -3135
rect 12160 -3255 12280 -3135
rect 12325 -3255 12445 -3135
rect 12490 -3255 12610 -3135
rect 7130 -3430 7250 -3310
rect 7305 -3430 7425 -3310
rect 7470 -3430 7590 -3310
rect 7635 -3430 7755 -3310
rect 7800 -3430 7920 -3310
rect 7975 -3430 8095 -3310
rect 8140 -3430 8260 -3310
rect 8305 -3430 8425 -3310
rect 8470 -3430 8590 -3310
rect 8645 -3430 8765 -3310
rect 8810 -3430 8930 -3310
rect 8975 -3430 9095 -3310
rect 9140 -3430 9260 -3310
rect 9315 -3430 9435 -3310
rect 9480 -3430 9600 -3310
rect 9645 -3430 9765 -3310
rect 9810 -3430 9930 -3310
rect 9985 -3430 10105 -3310
rect 10150 -3430 10270 -3310
rect 10315 -3430 10435 -3310
rect 10480 -3430 10600 -3310
rect 10655 -3430 10775 -3310
rect 10820 -3430 10940 -3310
rect 10985 -3430 11105 -3310
rect 11150 -3430 11270 -3310
rect 11325 -3430 11445 -3310
rect 11490 -3430 11610 -3310
rect 11655 -3430 11775 -3310
rect 11820 -3430 11940 -3310
rect 11995 -3430 12115 -3310
rect 12160 -3430 12280 -3310
rect 12325 -3430 12445 -3310
rect 12490 -3430 12610 -3310
rect 7130 -3595 7250 -3475
rect 7305 -3595 7425 -3475
rect 7470 -3595 7590 -3475
rect 7635 -3595 7755 -3475
rect 7800 -3595 7920 -3475
rect 7975 -3595 8095 -3475
rect 8140 -3595 8260 -3475
rect 8305 -3595 8425 -3475
rect 8470 -3595 8590 -3475
rect 8645 -3595 8765 -3475
rect 8810 -3595 8930 -3475
rect 8975 -3595 9095 -3475
rect 9140 -3595 9260 -3475
rect 9315 -3595 9435 -3475
rect 9480 -3595 9600 -3475
rect 9645 -3595 9765 -3475
rect 9810 -3595 9930 -3475
rect 9985 -3595 10105 -3475
rect 10150 -3595 10270 -3475
rect 10315 -3595 10435 -3475
rect 10480 -3595 10600 -3475
rect 10655 -3595 10775 -3475
rect 10820 -3595 10940 -3475
rect 10985 -3595 11105 -3475
rect 11150 -3595 11270 -3475
rect 11325 -3595 11445 -3475
rect 11490 -3595 11610 -3475
rect 11655 -3595 11775 -3475
rect 11820 -3595 11940 -3475
rect 11995 -3595 12115 -3475
rect 12160 -3595 12280 -3475
rect 12325 -3595 12445 -3475
rect 12490 -3595 12610 -3475
rect 7130 -3760 7250 -3640
rect 7305 -3760 7425 -3640
rect 7470 -3760 7590 -3640
rect 7635 -3760 7755 -3640
rect 7800 -3760 7920 -3640
rect 7975 -3760 8095 -3640
rect 8140 -3760 8260 -3640
rect 8305 -3760 8425 -3640
rect 8470 -3760 8590 -3640
rect 8645 -3760 8765 -3640
rect 8810 -3760 8930 -3640
rect 8975 -3760 9095 -3640
rect 9140 -3760 9260 -3640
rect 9315 -3760 9435 -3640
rect 9480 -3760 9600 -3640
rect 9645 -3760 9765 -3640
rect 9810 -3760 9930 -3640
rect 9985 -3760 10105 -3640
rect 10150 -3760 10270 -3640
rect 10315 -3760 10435 -3640
rect 10480 -3760 10600 -3640
rect 10655 -3760 10775 -3640
rect 10820 -3760 10940 -3640
rect 10985 -3760 11105 -3640
rect 11150 -3760 11270 -3640
rect 11325 -3760 11445 -3640
rect 11490 -3760 11610 -3640
rect 11655 -3760 11775 -3640
rect 11820 -3760 11940 -3640
rect 11995 -3760 12115 -3640
rect 12160 -3760 12280 -3640
rect 12325 -3760 12445 -3640
rect 12490 -3760 12610 -3640
rect 7130 -3925 7250 -3805
rect 7305 -3925 7425 -3805
rect 7470 -3925 7590 -3805
rect 7635 -3925 7755 -3805
rect 7800 -3925 7920 -3805
rect 7975 -3925 8095 -3805
rect 8140 -3925 8260 -3805
rect 8305 -3925 8425 -3805
rect 8470 -3925 8590 -3805
rect 8645 -3925 8765 -3805
rect 8810 -3925 8930 -3805
rect 8975 -3925 9095 -3805
rect 9140 -3925 9260 -3805
rect 9315 -3925 9435 -3805
rect 9480 -3925 9600 -3805
rect 9645 -3925 9765 -3805
rect 9810 -3925 9930 -3805
rect 9985 -3925 10105 -3805
rect 10150 -3925 10270 -3805
rect 10315 -3925 10435 -3805
rect 10480 -3925 10600 -3805
rect 10655 -3925 10775 -3805
rect 10820 -3925 10940 -3805
rect 10985 -3925 11105 -3805
rect 11150 -3925 11270 -3805
rect 11325 -3925 11445 -3805
rect 11490 -3925 11610 -3805
rect 11655 -3925 11775 -3805
rect 11820 -3925 11940 -3805
rect 11995 -3925 12115 -3805
rect 12160 -3925 12280 -3805
rect 12325 -3925 12445 -3805
rect 12490 -3925 12610 -3805
rect 7130 -4100 7250 -3980
rect 7305 -4100 7425 -3980
rect 7470 -4100 7590 -3980
rect 7635 -4100 7755 -3980
rect 7800 -4100 7920 -3980
rect 7975 -4100 8095 -3980
rect 8140 -4100 8260 -3980
rect 8305 -4100 8425 -3980
rect 8470 -4100 8590 -3980
rect 8645 -4100 8765 -3980
rect 8810 -4100 8930 -3980
rect 8975 -4100 9095 -3980
rect 9140 -4100 9260 -3980
rect 9315 -4100 9435 -3980
rect 9480 -4100 9600 -3980
rect 9645 -4100 9765 -3980
rect 9810 -4100 9930 -3980
rect 9985 -4100 10105 -3980
rect 10150 -4100 10270 -3980
rect 10315 -4100 10435 -3980
rect 10480 -4100 10600 -3980
rect 10655 -4100 10775 -3980
rect 10820 -4100 10940 -3980
rect 10985 -4100 11105 -3980
rect 11150 -4100 11270 -3980
rect 11325 -4100 11445 -3980
rect 11490 -4100 11610 -3980
rect 11655 -4100 11775 -3980
rect 11820 -4100 11940 -3980
rect 11995 -4100 12115 -3980
rect 12160 -4100 12280 -3980
rect 12325 -4100 12445 -3980
rect 12490 -4100 12610 -3980
rect 12820 1260 12940 1380
rect 12995 1260 13115 1380
rect 13160 1260 13280 1380
rect 13325 1260 13445 1380
rect 13490 1260 13610 1380
rect 13665 1260 13785 1380
rect 13830 1260 13950 1380
rect 13995 1260 14115 1380
rect 14160 1260 14280 1380
rect 14335 1260 14455 1380
rect 14500 1260 14620 1380
rect 14665 1260 14785 1380
rect 14830 1260 14950 1380
rect 15005 1260 15125 1380
rect 15170 1260 15290 1380
rect 15335 1260 15455 1380
rect 15500 1260 15620 1380
rect 15675 1260 15795 1380
rect 15840 1260 15960 1380
rect 16005 1260 16125 1380
rect 16170 1260 16290 1380
rect 16345 1260 16465 1380
rect 16510 1260 16630 1380
rect 16675 1260 16795 1380
rect 16840 1260 16960 1380
rect 17015 1260 17135 1380
rect 17180 1260 17300 1380
rect 17345 1260 17465 1380
rect 17510 1260 17630 1380
rect 17685 1260 17805 1380
rect 17850 1260 17970 1380
rect 18015 1260 18135 1380
rect 18180 1260 18300 1380
rect 12820 1095 12940 1215
rect 12995 1095 13115 1215
rect 13160 1095 13280 1215
rect 13325 1095 13445 1215
rect 13490 1095 13610 1215
rect 13665 1095 13785 1215
rect 13830 1095 13950 1215
rect 13995 1095 14115 1215
rect 14160 1095 14280 1215
rect 14335 1095 14455 1215
rect 14500 1095 14620 1215
rect 14665 1095 14785 1215
rect 14830 1095 14950 1215
rect 15005 1095 15125 1215
rect 15170 1095 15290 1215
rect 15335 1095 15455 1215
rect 15500 1095 15620 1215
rect 15675 1095 15795 1215
rect 15840 1095 15960 1215
rect 16005 1095 16125 1215
rect 16170 1095 16290 1215
rect 16345 1095 16465 1215
rect 16510 1095 16630 1215
rect 16675 1095 16795 1215
rect 16840 1095 16960 1215
rect 17015 1095 17135 1215
rect 17180 1095 17300 1215
rect 17345 1095 17465 1215
rect 17510 1095 17630 1215
rect 17685 1095 17805 1215
rect 17850 1095 17970 1215
rect 18015 1095 18135 1215
rect 18180 1095 18300 1215
rect 12820 930 12940 1050
rect 12995 930 13115 1050
rect 13160 930 13280 1050
rect 13325 930 13445 1050
rect 13490 930 13610 1050
rect 13665 930 13785 1050
rect 13830 930 13950 1050
rect 13995 930 14115 1050
rect 14160 930 14280 1050
rect 14335 930 14455 1050
rect 14500 930 14620 1050
rect 14665 930 14785 1050
rect 14830 930 14950 1050
rect 15005 930 15125 1050
rect 15170 930 15290 1050
rect 15335 930 15455 1050
rect 15500 930 15620 1050
rect 15675 930 15795 1050
rect 15840 930 15960 1050
rect 16005 930 16125 1050
rect 16170 930 16290 1050
rect 16345 930 16465 1050
rect 16510 930 16630 1050
rect 16675 930 16795 1050
rect 16840 930 16960 1050
rect 17015 930 17135 1050
rect 17180 930 17300 1050
rect 17345 930 17465 1050
rect 17510 930 17630 1050
rect 17685 930 17805 1050
rect 17850 930 17970 1050
rect 18015 930 18135 1050
rect 18180 930 18300 1050
rect 12820 765 12940 885
rect 12995 765 13115 885
rect 13160 765 13280 885
rect 13325 765 13445 885
rect 13490 765 13610 885
rect 13665 765 13785 885
rect 13830 765 13950 885
rect 13995 765 14115 885
rect 14160 765 14280 885
rect 14335 765 14455 885
rect 14500 765 14620 885
rect 14665 765 14785 885
rect 14830 765 14950 885
rect 15005 765 15125 885
rect 15170 765 15290 885
rect 15335 765 15455 885
rect 15500 765 15620 885
rect 15675 765 15795 885
rect 15840 765 15960 885
rect 16005 765 16125 885
rect 16170 765 16290 885
rect 16345 765 16465 885
rect 16510 765 16630 885
rect 16675 765 16795 885
rect 16840 765 16960 885
rect 17015 765 17135 885
rect 17180 765 17300 885
rect 17345 765 17465 885
rect 17510 765 17630 885
rect 17685 765 17805 885
rect 17850 765 17970 885
rect 18015 765 18135 885
rect 18180 765 18300 885
rect 12820 590 12940 710
rect 12995 590 13115 710
rect 13160 590 13280 710
rect 13325 590 13445 710
rect 13490 590 13610 710
rect 13665 590 13785 710
rect 13830 590 13950 710
rect 13995 590 14115 710
rect 14160 590 14280 710
rect 14335 590 14455 710
rect 14500 590 14620 710
rect 14665 590 14785 710
rect 14830 590 14950 710
rect 15005 590 15125 710
rect 15170 590 15290 710
rect 15335 590 15455 710
rect 15500 590 15620 710
rect 15675 590 15795 710
rect 15840 590 15960 710
rect 16005 590 16125 710
rect 16170 590 16290 710
rect 16345 590 16465 710
rect 16510 590 16630 710
rect 16675 590 16795 710
rect 16840 590 16960 710
rect 17015 590 17135 710
rect 17180 590 17300 710
rect 17345 590 17465 710
rect 17510 590 17630 710
rect 17685 590 17805 710
rect 17850 590 17970 710
rect 18015 590 18135 710
rect 18180 590 18300 710
rect 12820 425 12940 545
rect 12995 425 13115 545
rect 13160 425 13280 545
rect 13325 425 13445 545
rect 13490 425 13610 545
rect 13665 425 13785 545
rect 13830 425 13950 545
rect 13995 425 14115 545
rect 14160 425 14280 545
rect 14335 425 14455 545
rect 14500 425 14620 545
rect 14665 425 14785 545
rect 14830 425 14950 545
rect 15005 425 15125 545
rect 15170 425 15290 545
rect 15335 425 15455 545
rect 15500 425 15620 545
rect 15675 425 15795 545
rect 15840 425 15960 545
rect 16005 425 16125 545
rect 16170 425 16290 545
rect 16345 425 16465 545
rect 16510 425 16630 545
rect 16675 425 16795 545
rect 16840 425 16960 545
rect 17015 425 17135 545
rect 17180 425 17300 545
rect 17345 425 17465 545
rect 17510 425 17630 545
rect 17685 425 17805 545
rect 17850 425 17970 545
rect 18015 425 18135 545
rect 18180 425 18300 545
rect 12820 260 12940 380
rect 12995 260 13115 380
rect 13160 260 13280 380
rect 13325 260 13445 380
rect 13490 260 13610 380
rect 13665 260 13785 380
rect 13830 260 13950 380
rect 13995 260 14115 380
rect 14160 260 14280 380
rect 14335 260 14455 380
rect 14500 260 14620 380
rect 14665 260 14785 380
rect 14830 260 14950 380
rect 15005 260 15125 380
rect 15170 260 15290 380
rect 15335 260 15455 380
rect 15500 260 15620 380
rect 15675 260 15795 380
rect 15840 260 15960 380
rect 16005 260 16125 380
rect 16170 260 16290 380
rect 16345 260 16465 380
rect 16510 260 16630 380
rect 16675 260 16795 380
rect 16840 260 16960 380
rect 17015 260 17135 380
rect 17180 260 17300 380
rect 17345 260 17465 380
rect 17510 260 17630 380
rect 17685 260 17805 380
rect 17850 260 17970 380
rect 18015 260 18135 380
rect 18180 260 18300 380
rect 12820 95 12940 215
rect 12995 95 13115 215
rect 13160 95 13280 215
rect 13325 95 13445 215
rect 13490 95 13610 215
rect 13665 95 13785 215
rect 13830 95 13950 215
rect 13995 95 14115 215
rect 14160 95 14280 215
rect 14335 95 14455 215
rect 14500 95 14620 215
rect 14665 95 14785 215
rect 14830 95 14950 215
rect 15005 95 15125 215
rect 15170 95 15290 215
rect 15335 95 15455 215
rect 15500 95 15620 215
rect 15675 95 15795 215
rect 15840 95 15960 215
rect 16005 95 16125 215
rect 16170 95 16290 215
rect 16345 95 16465 215
rect 16510 95 16630 215
rect 16675 95 16795 215
rect 16840 95 16960 215
rect 17015 95 17135 215
rect 17180 95 17300 215
rect 17345 95 17465 215
rect 17510 95 17630 215
rect 17685 95 17805 215
rect 17850 95 17970 215
rect 18015 95 18135 215
rect 18180 95 18300 215
rect 12820 -80 12940 40
rect 12995 -80 13115 40
rect 13160 -80 13280 40
rect 13325 -80 13445 40
rect 13490 -80 13610 40
rect 13665 -80 13785 40
rect 13830 -80 13950 40
rect 13995 -80 14115 40
rect 14160 -80 14280 40
rect 14335 -80 14455 40
rect 14500 -80 14620 40
rect 14665 -80 14785 40
rect 14830 -80 14950 40
rect 15005 -80 15125 40
rect 15170 -80 15290 40
rect 15335 -80 15455 40
rect 15500 -80 15620 40
rect 15675 -80 15795 40
rect 15840 -80 15960 40
rect 16005 -80 16125 40
rect 16170 -80 16290 40
rect 16345 -80 16465 40
rect 16510 -80 16630 40
rect 16675 -80 16795 40
rect 16840 -80 16960 40
rect 17015 -80 17135 40
rect 17180 -80 17300 40
rect 17345 -80 17465 40
rect 17510 -80 17630 40
rect 17685 -80 17805 40
rect 17850 -80 17970 40
rect 18015 -80 18135 40
rect 18180 -80 18300 40
rect 12820 -245 12940 -125
rect 12995 -245 13115 -125
rect 13160 -245 13280 -125
rect 13325 -245 13445 -125
rect 13490 -245 13610 -125
rect 13665 -245 13785 -125
rect 13830 -245 13950 -125
rect 13995 -245 14115 -125
rect 14160 -245 14280 -125
rect 14335 -245 14455 -125
rect 14500 -245 14620 -125
rect 14665 -245 14785 -125
rect 14830 -245 14950 -125
rect 15005 -245 15125 -125
rect 15170 -245 15290 -125
rect 15335 -245 15455 -125
rect 15500 -245 15620 -125
rect 15675 -245 15795 -125
rect 15840 -245 15960 -125
rect 16005 -245 16125 -125
rect 16170 -245 16290 -125
rect 16345 -245 16465 -125
rect 16510 -245 16630 -125
rect 16675 -245 16795 -125
rect 16840 -245 16960 -125
rect 17015 -245 17135 -125
rect 17180 -245 17300 -125
rect 17345 -245 17465 -125
rect 17510 -245 17630 -125
rect 17685 -245 17805 -125
rect 17850 -245 17970 -125
rect 18015 -245 18135 -125
rect 18180 -245 18300 -125
rect 12820 -410 12940 -290
rect 12995 -410 13115 -290
rect 13160 -410 13280 -290
rect 13325 -410 13445 -290
rect 13490 -410 13610 -290
rect 13665 -410 13785 -290
rect 13830 -410 13950 -290
rect 13995 -410 14115 -290
rect 14160 -410 14280 -290
rect 14335 -410 14455 -290
rect 14500 -410 14620 -290
rect 14665 -410 14785 -290
rect 14830 -410 14950 -290
rect 15005 -410 15125 -290
rect 15170 -410 15290 -290
rect 15335 -410 15455 -290
rect 15500 -410 15620 -290
rect 15675 -410 15795 -290
rect 15840 -410 15960 -290
rect 16005 -410 16125 -290
rect 16170 -410 16290 -290
rect 16345 -410 16465 -290
rect 16510 -410 16630 -290
rect 16675 -410 16795 -290
rect 16840 -410 16960 -290
rect 17015 -410 17135 -290
rect 17180 -410 17300 -290
rect 17345 -410 17465 -290
rect 17510 -410 17630 -290
rect 17685 -410 17805 -290
rect 17850 -410 17970 -290
rect 18015 -410 18135 -290
rect 18180 -410 18300 -290
rect 12820 -575 12940 -455
rect 12995 -575 13115 -455
rect 13160 -575 13280 -455
rect 13325 -575 13445 -455
rect 13490 -575 13610 -455
rect 13665 -575 13785 -455
rect 13830 -575 13950 -455
rect 13995 -575 14115 -455
rect 14160 -575 14280 -455
rect 14335 -575 14455 -455
rect 14500 -575 14620 -455
rect 14665 -575 14785 -455
rect 14830 -575 14950 -455
rect 15005 -575 15125 -455
rect 15170 -575 15290 -455
rect 15335 -575 15455 -455
rect 15500 -575 15620 -455
rect 15675 -575 15795 -455
rect 15840 -575 15960 -455
rect 16005 -575 16125 -455
rect 16170 -575 16290 -455
rect 16345 -575 16465 -455
rect 16510 -575 16630 -455
rect 16675 -575 16795 -455
rect 16840 -575 16960 -455
rect 17015 -575 17135 -455
rect 17180 -575 17300 -455
rect 17345 -575 17465 -455
rect 17510 -575 17630 -455
rect 17685 -575 17805 -455
rect 17850 -575 17970 -455
rect 18015 -575 18135 -455
rect 18180 -575 18300 -455
rect 12820 -750 12940 -630
rect 12995 -750 13115 -630
rect 13160 -750 13280 -630
rect 13325 -750 13445 -630
rect 13490 -750 13610 -630
rect 13665 -750 13785 -630
rect 13830 -750 13950 -630
rect 13995 -750 14115 -630
rect 14160 -750 14280 -630
rect 14335 -750 14455 -630
rect 14500 -750 14620 -630
rect 14665 -750 14785 -630
rect 14830 -750 14950 -630
rect 15005 -750 15125 -630
rect 15170 -750 15290 -630
rect 15335 -750 15455 -630
rect 15500 -750 15620 -630
rect 15675 -750 15795 -630
rect 15840 -750 15960 -630
rect 16005 -750 16125 -630
rect 16170 -750 16290 -630
rect 16345 -750 16465 -630
rect 16510 -750 16630 -630
rect 16675 -750 16795 -630
rect 16840 -750 16960 -630
rect 17015 -750 17135 -630
rect 17180 -750 17300 -630
rect 17345 -750 17465 -630
rect 17510 -750 17630 -630
rect 17685 -750 17805 -630
rect 17850 -750 17970 -630
rect 18015 -750 18135 -630
rect 18180 -750 18300 -630
rect 12820 -915 12940 -795
rect 12995 -915 13115 -795
rect 13160 -915 13280 -795
rect 13325 -915 13445 -795
rect 13490 -915 13610 -795
rect 13665 -915 13785 -795
rect 13830 -915 13950 -795
rect 13995 -915 14115 -795
rect 14160 -915 14280 -795
rect 14335 -915 14455 -795
rect 14500 -915 14620 -795
rect 14665 -915 14785 -795
rect 14830 -915 14950 -795
rect 15005 -915 15125 -795
rect 15170 -915 15290 -795
rect 15335 -915 15455 -795
rect 15500 -915 15620 -795
rect 15675 -915 15795 -795
rect 15840 -915 15960 -795
rect 16005 -915 16125 -795
rect 16170 -915 16290 -795
rect 16345 -915 16465 -795
rect 16510 -915 16630 -795
rect 16675 -915 16795 -795
rect 16840 -915 16960 -795
rect 17015 -915 17135 -795
rect 17180 -915 17300 -795
rect 17345 -915 17465 -795
rect 17510 -915 17630 -795
rect 17685 -915 17805 -795
rect 17850 -915 17970 -795
rect 18015 -915 18135 -795
rect 18180 -915 18300 -795
rect 12820 -1080 12940 -960
rect 12995 -1080 13115 -960
rect 13160 -1080 13280 -960
rect 13325 -1080 13445 -960
rect 13490 -1080 13610 -960
rect 13665 -1080 13785 -960
rect 13830 -1080 13950 -960
rect 13995 -1080 14115 -960
rect 14160 -1080 14280 -960
rect 14335 -1080 14455 -960
rect 14500 -1080 14620 -960
rect 14665 -1080 14785 -960
rect 14830 -1080 14950 -960
rect 15005 -1080 15125 -960
rect 15170 -1080 15290 -960
rect 15335 -1080 15455 -960
rect 15500 -1080 15620 -960
rect 15675 -1080 15795 -960
rect 15840 -1080 15960 -960
rect 16005 -1080 16125 -960
rect 16170 -1080 16290 -960
rect 16345 -1080 16465 -960
rect 16510 -1080 16630 -960
rect 16675 -1080 16795 -960
rect 16840 -1080 16960 -960
rect 17015 -1080 17135 -960
rect 17180 -1080 17300 -960
rect 17345 -1080 17465 -960
rect 17510 -1080 17630 -960
rect 17685 -1080 17805 -960
rect 17850 -1080 17970 -960
rect 18015 -1080 18135 -960
rect 18180 -1080 18300 -960
rect 12820 -1245 12940 -1125
rect 12995 -1245 13115 -1125
rect 13160 -1245 13280 -1125
rect 13325 -1245 13445 -1125
rect 13490 -1245 13610 -1125
rect 13665 -1245 13785 -1125
rect 13830 -1245 13950 -1125
rect 13995 -1245 14115 -1125
rect 14160 -1245 14280 -1125
rect 14335 -1245 14455 -1125
rect 14500 -1245 14620 -1125
rect 14665 -1245 14785 -1125
rect 14830 -1245 14950 -1125
rect 15005 -1245 15125 -1125
rect 15170 -1245 15290 -1125
rect 15335 -1245 15455 -1125
rect 15500 -1245 15620 -1125
rect 15675 -1245 15795 -1125
rect 15840 -1245 15960 -1125
rect 16005 -1245 16125 -1125
rect 16170 -1245 16290 -1125
rect 16345 -1245 16465 -1125
rect 16510 -1245 16630 -1125
rect 16675 -1245 16795 -1125
rect 16840 -1245 16960 -1125
rect 17015 -1245 17135 -1125
rect 17180 -1245 17300 -1125
rect 17345 -1245 17465 -1125
rect 17510 -1245 17630 -1125
rect 17685 -1245 17805 -1125
rect 17850 -1245 17970 -1125
rect 18015 -1245 18135 -1125
rect 18180 -1245 18300 -1125
rect 12820 -1420 12940 -1300
rect 12995 -1420 13115 -1300
rect 13160 -1420 13280 -1300
rect 13325 -1420 13445 -1300
rect 13490 -1420 13610 -1300
rect 13665 -1420 13785 -1300
rect 13830 -1420 13950 -1300
rect 13995 -1420 14115 -1300
rect 14160 -1420 14280 -1300
rect 14335 -1420 14455 -1300
rect 14500 -1420 14620 -1300
rect 14665 -1420 14785 -1300
rect 14830 -1420 14950 -1300
rect 15005 -1420 15125 -1300
rect 15170 -1420 15290 -1300
rect 15335 -1420 15455 -1300
rect 15500 -1420 15620 -1300
rect 15675 -1420 15795 -1300
rect 15840 -1420 15960 -1300
rect 16005 -1420 16125 -1300
rect 16170 -1420 16290 -1300
rect 16345 -1420 16465 -1300
rect 16510 -1420 16630 -1300
rect 16675 -1420 16795 -1300
rect 16840 -1420 16960 -1300
rect 17015 -1420 17135 -1300
rect 17180 -1420 17300 -1300
rect 17345 -1420 17465 -1300
rect 17510 -1420 17630 -1300
rect 17685 -1420 17805 -1300
rect 17850 -1420 17970 -1300
rect 18015 -1420 18135 -1300
rect 18180 -1420 18300 -1300
rect 12820 -1585 12940 -1465
rect 12995 -1585 13115 -1465
rect 13160 -1585 13280 -1465
rect 13325 -1585 13445 -1465
rect 13490 -1585 13610 -1465
rect 13665 -1585 13785 -1465
rect 13830 -1585 13950 -1465
rect 13995 -1585 14115 -1465
rect 14160 -1585 14280 -1465
rect 14335 -1585 14455 -1465
rect 14500 -1585 14620 -1465
rect 14665 -1585 14785 -1465
rect 14830 -1585 14950 -1465
rect 15005 -1585 15125 -1465
rect 15170 -1585 15290 -1465
rect 15335 -1585 15455 -1465
rect 15500 -1585 15620 -1465
rect 15675 -1585 15795 -1465
rect 15840 -1585 15960 -1465
rect 16005 -1585 16125 -1465
rect 16170 -1585 16290 -1465
rect 16345 -1585 16465 -1465
rect 16510 -1585 16630 -1465
rect 16675 -1585 16795 -1465
rect 16840 -1585 16960 -1465
rect 17015 -1585 17135 -1465
rect 17180 -1585 17300 -1465
rect 17345 -1585 17465 -1465
rect 17510 -1585 17630 -1465
rect 17685 -1585 17805 -1465
rect 17850 -1585 17970 -1465
rect 18015 -1585 18135 -1465
rect 18180 -1585 18300 -1465
rect 12820 -1750 12940 -1630
rect 12995 -1750 13115 -1630
rect 13160 -1750 13280 -1630
rect 13325 -1750 13445 -1630
rect 13490 -1750 13610 -1630
rect 13665 -1750 13785 -1630
rect 13830 -1750 13950 -1630
rect 13995 -1750 14115 -1630
rect 14160 -1750 14280 -1630
rect 14335 -1750 14455 -1630
rect 14500 -1750 14620 -1630
rect 14665 -1750 14785 -1630
rect 14830 -1750 14950 -1630
rect 15005 -1750 15125 -1630
rect 15170 -1750 15290 -1630
rect 15335 -1750 15455 -1630
rect 15500 -1750 15620 -1630
rect 15675 -1750 15795 -1630
rect 15840 -1750 15960 -1630
rect 16005 -1750 16125 -1630
rect 16170 -1750 16290 -1630
rect 16345 -1750 16465 -1630
rect 16510 -1750 16630 -1630
rect 16675 -1750 16795 -1630
rect 16840 -1750 16960 -1630
rect 17015 -1750 17135 -1630
rect 17180 -1750 17300 -1630
rect 17345 -1750 17465 -1630
rect 17510 -1750 17630 -1630
rect 17685 -1750 17805 -1630
rect 17850 -1750 17970 -1630
rect 18015 -1750 18135 -1630
rect 18180 -1750 18300 -1630
rect 12820 -1915 12940 -1795
rect 12995 -1915 13115 -1795
rect 13160 -1915 13280 -1795
rect 13325 -1915 13445 -1795
rect 13490 -1915 13610 -1795
rect 13665 -1915 13785 -1795
rect 13830 -1915 13950 -1795
rect 13995 -1915 14115 -1795
rect 14160 -1915 14280 -1795
rect 14335 -1915 14455 -1795
rect 14500 -1915 14620 -1795
rect 14665 -1915 14785 -1795
rect 14830 -1915 14950 -1795
rect 15005 -1915 15125 -1795
rect 15170 -1915 15290 -1795
rect 15335 -1915 15455 -1795
rect 15500 -1915 15620 -1795
rect 15675 -1915 15795 -1795
rect 15840 -1915 15960 -1795
rect 16005 -1915 16125 -1795
rect 16170 -1915 16290 -1795
rect 16345 -1915 16465 -1795
rect 16510 -1915 16630 -1795
rect 16675 -1915 16795 -1795
rect 16840 -1915 16960 -1795
rect 17015 -1915 17135 -1795
rect 17180 -1915 17300 -1795
rect 17345 -1915 17465 -1795
rect 17510 -1915 17630 -1795
rect 17685 -1915 17805 -1795
rect 17850 -1915 17970 -1795
rect 18015 -1915 18135 -1795
rect 18180 -1915 18300 -1795
rect 12820 -2090 12940 -1970
rect 12995 -2090 13115 -1970
rect 13160 -2090 13280 -1970
rect 13325 -2090 13445 -1970
rect 13490 -2090 13610 -1970
rect 13665 -2090 13785 -1970
rect 13830 -2090 13950 -1970
rect 13995 -2090 14115 -1970
rect 14160 -2090 14280 -1970
rect 14335 -2090 14455 -1970
rect 14500 -2090 14620 -1970
rect 14665 -2090 14785 -1970
rect 14830 -2090 14950 -1970
rect 15005 -2090 15125 -1970
rect 15170 -2090 15290 -1970
rect 15335 -2090 15455 -1970
rect 15500 -2090 15620 -1970
rect 15675 -2090 15795 -1970
rect 15840 -2090 15960 -1970
rect 16005 -2090 16125 -1970
rect 16170 -2090 16290 -1970
rect 16345 -2090 16465 -1970
rect 16510 -2090 16630 -1970
rect 16675 -2090 16795 -1970
rect 16840 -2090 16960 -1970
rect 17015 -2090 17135 -1970
rect 17180 -2090 17300 -1970
rect 17345 -2090 17465 -1970
rect 17510 -2090 17630 -1970
rect 17685 -2090 17805 -1970
rect 17850 -2090 17970 -1970
rect 18015 -2090 18135 -1970
rect 18180 -2090 18300 -1970
rect 12820 -2255 12940 -2135
rect 12995 -2255 13115 -2135
rect 13160 -2255 13280 -2135
rect 13325 -2255 13445 -2135
rect 13490 -2255 13610 -2135
rect 13665 -2255 13785 -2135
rect 13830 -2255 13950 -2135
rect 13995 -2255 14115 -2135
rect 14160 -2255 14280 -2135
rect 14335 -2255 14455 -2135
rect 14500 -2255 14620 -2135
rect 14665 -2255 14785 -2135
rect 14830 -2255 14950 -2135
rect 15005 -2255 15125 -2135
rect 15170 -2255 15290 -2135
rect 15335 -2255 15455 -2135
rect 15500 -2255 15620 -2135
rect 15675 -2255 15795 -2135
rect 15840 -2255 15960 -2135
rect 16005 -2255 16125 -2135
rect 16170 -2255 16290 -2135
rect 16345 -2255 16465 -2135
rect 16510 -2255 16630 -2135
rect 16675 -2255 16795 -2135
rect 16840 -2255 16960 -2135
rect 17015 -2255 17135 -2135
rect 17180 -2255 17300 -2135
rect 17345 -2255 17465 -2135
rect 17510 -2255 17630 -2135
rect 17685 -2255 17805 -2135
rect 17850 -2255 17970 -2135
rect 18015 -2255 18135 -2135
rect 18180 -2255 18300 -2135
rect 12820 -2420 12940 -2300
rect 12995 -2420 13115 -2300
rect 13160 -2420 13280 -2300
rect 13325 -2420 13445 -2300
rect 13490 -2420 13610 -2300
rect 13665 -2420 13785 -2300
rect 13830 -2420 13950 -2300
rect 13995 -2420 14115 -2300
rect 14160 -2420 14280 -2300
rect 14335 -2420 14455 -2300
rect 14500 -2420 14620 -2300
rect 14665 -2420 14785 -2300
rect 14830 -2420 14950 -2300
rect 15005 -2420 15125 -2300
rect 15170 -2420 15290 -2300
rect 15335 -2420 15455 -2300
rect 15500 -2420 15620 -2300
rect 15675 -2420 15795 -2300
rect 15840 -2420 15960 -2300
rect 16005 -2420 16125 -2300
rect 16170 -2420 16290 -2300
rect 16345 -2420 16465 -2300
rect 16510 -2420 16630 -2300
rect 16675 -2420 16795 -2300
rect 16840 -2420 16960 -2300
rect 17015 -2420 17135 -2300
rect 17180 -2420 17300 -2300
rect 17345 -2420 17465 -2300
rect 17510 -2420 17630 -2300
rect 17685 -2420 17805 -2300
rect 17850 -2420 17970 -2300
rect 18015 -2420 18135 -2300
rect 18180 -2420 18300 -2300
rect 12820 -2585 12940 -2465
rect 12995 -2585 13115 -2465
rect 13160 -2585 13280 -2465
rect 13325 -2585 13445 -2465
rect 13490 -2585 13610 -2465
rect 13665 -2585 13785 -2465
rect 13830 -2585 13950 -2465
rect 13995 -2585 14115 -2465
rect 14160 -2585 14280 -2465
rect 14335 -2585 14455 -2465
rect 14500 -2585 14620 -2465
rect 14665 -2585 14785 -2465
rect 14830 -2585 14950 -2465
rect 15005 -2585 15125 -2465
rect 15170 -2585 15290 -2465
rect 15335 -2585 15455 -2465
rect 15500 -2585 15620 -2465
rect 15675 -2585 15795 -2465
rect 15840 -2585 15960 -2465
rect 16005 -2585 16125 -2465
rect 16170 -2585 16290 -2465
rect 16345 -2585 16465 -2465
rect 16510 -2585 16630 -2465
rect 16675 -2585 16795 -2465
rect 16840 -2585 16960 -2465
rect 17015 -2585 17135 -2465
rect 17180 -2585 17300 -2465
rect 17345 -2585 17465 -2465
rect 17510 -2585 17630 -2465
rect 17685 -2585 17805 -2465
rect 17850 -2585 17970 -2465
rect 18015 -2585 18135 -2465
rect 18180 -2585 18300 -2465
rect 12820 -2760 12940 -2640
rect 12995 -2760 13115 -2640
rect 13160 -2760 13280 -2640
rect 13325 -2760 13445 -2640
rect 13490 -2760 13610 -2640
rect 13665 -2760 13785 -2640
rect 13830 -2760 13950 -2640
rect 13995 -2760 14115 -2640
rect 14160 -2760 14280 -2640
rect 14335 -2760 14455 -2640
rect 14500 -2760 14620 -2640
rect 14665 -2760 14785 -2640
rect 14830 -2760 14950 -2640
rect 15005 -2760 15125 -2640
rect 15170 -2760 15290 -2640
rect 15335 -2760 15455 -2640
rect 15500 -2760 15620 -2640
rect 15675 -2760 15795 -2640
rect 15840 -2760 15960 -2640
rect 16005 -2760 16125 -2640
rect 16170 -2760 16290 -2640
rect 16345 -2760 16465 -2640
rect 16510 -2760 16630 -2640
rect 16675 -2760 16795 -2640
rect 16840 -2760 16960 -2640
rect 17015 -2760 17135 -2640
rect 17180 -2760 17300 -2640
rect 17345 -2760 17465 -2640
rect 17510 -2760 17630 -2640
rect 17685 -2760 17805 -2640
rect 17850 -2760 17970 -2640
rect 18015 -2760 18135 -2640
rect 18180 -2760 18300 -2640
rect 12820 -2925 12940 -2805
rect 12995 -2925 13115 -2805
rect 13160 -2925 13280 -2805
rect 13325 -2925 13445 -2805
rect 13490 -2925 13610 -2805
rect 13665 -2925 13785 -2805
rect 13830 -2925 13950 -2805
rect 13995 -2925 14115 -2805
rect 14160 -2925 14280 -2805
rect 14335 -2925 14455 -2805
rect 14500 -2925 14620 -2805
rect 14665 -2925 14785 -2805
rect 14830 -2925 14950 -2805
rect 15005 -2925 15125 -2805
rect 15170 -2925 15290 -2805
rect 15335 -2925 15455 -2805
rect 15500 -2925 15620 -2805
rect 15675 -2925 15795 -2805
rect 15840 -2925 15960 -2805
rect 16005 -2925 16125 -2805
rect 16170 -2925 16290 -2805
rect 16345 -2925 16465 -2805
rect 16510 -2925 16630 -2805
rect 16675 -2925 16795 -2805
rect 16840 -2925 16960 -2805
rect 17015 -2925 17135 -2805
rect 17180 -2925 17300 -2805
rect 17345 -2925 17465 -2805
rect 17510 -2925 17630 -2805
rect 17685 -2925 17805 -2805
rect 17850 -2925 17970 -2805
rect 18015 -2925 18135 -2805
rect 18180 -2925 18300 -2805
rect 12820 -3090 12940 -2970
rect 12995 -3090 13115 -2970
rect 13160 -3090 13280 -2970
rect 13325 -3090 13445 -2970
rect 13490 -3090 13610 -2970
rect 13665 -3090 13785 -2970
rect 13830 -3090 13950 -2970
rect 13995 -3090 14115 -2970
rect 14160 -3090 14280 -2970
rect 14335 -3090 14455 -2970
rect 14500 -3090 14620 -2970
rect 14665 -3090 14785 -2970
rect 14830 -3090 14950 -2970
rect 15005 -3090 15125 -2970
rect 15170 -3090 15290 -2970
rect 15335 -3090 15455 -2970
rect 15500 -3090 15620 -2970
rect 15675 -3090 15795 -2970
rect 15840 -3090 15960 -2970
rect 16005 -3090 16125 -2970
rect 16170 -3090 16290 -2970
rect 16345 -3090 16465 -2970
rect 16510 -3090 16630 -2970
rect 16675 -3090 16795 -2970
rect 16840 -3090 16960 -2970
rect 17015 -3090 17135 -2970
rect 17180 -3090 17300 -2970
rect 17345 -3090 17465 -2970
rect 17510 -3090 17630 -2970
rect 17685 -3090 17805 -2970
rect 17850 -3090 17970 -2970
rect 18015 -3090 18135 -2970
rect 18180 -3090 18300 -2970
rect 12820 -3255 12940 -3135
rect 12995 -3255 13115 -3135
rect 13160 -3255 13280 -3135
rect 13325 -3255 13445 -3135
rect 13490 -3255 13610 -3135
rect 13665 -3255 13785 -3135
rect 13830 -3255 13950 -3135
rect 13995 -3255 14115 -3135
rect 14160 -3255 14280 -3135
rect 14335 -3255 14455 -3135
rect 14500 -3255 14620 -3135
rect 14665 -3255 14785 -3135
rect 14830 -3255 14950 -3135
rect 15005 -3255 15125 -3135
rect 15170 -3255 15290 -3135
rect 15335 -3255 15455 -3135
rect 15500 -3255 15620 -3135
rect 15675 -3255 15795 -3135
rect 15840 -3255 15960 -3135
rect 16005 -3255 16125 -3135
rect 16170 -3255 16290 -3135
rect 16345 -3255 16465 -3135
rect 16510 -3255 16630 -3135
rect 16675 -3255 16795 -3135
rect 16840 -3255 16960 -3135
rect 17015 -3255 17135 -3135
rect 17180 -3255 17300 -3135
rect 17345 -3255 17465 -3135
rect 17510 -3255 17630 -3135
rect 17685 -3255 17805 -3135
rect 17850 -3255 17970 -3135
rect 18015 -3255 18135 -3135
rect 18180 -3255 18300 -3135
rect 12820 -3430 12940 -3310
rect 12995 -3430 13115 -3310
rect 13160 -3430 13280 -3310
rect 13325 -3430 13445 -3310
rect 13490 -3430 13610 -3310
rect 13665 -3430 13785 -3310
rect 13830 -3430 13950 -3310
rect 13995 -3430 14115 -3310
rect 14160 -3430 14280 -3310
rect 14335 -3430 14455 -3310
rect 14500 -3430 14620 -3310
rect 14665 -3430 14785 -3310
rect 14830 -3430 14950 -3310
rect 15005 -3430 15125 -3310
rect 15170 -3430 15290 -3310
rect 15335 -3430 15455 -3310
rect 15500 -3430 15620 -3310
rect 15675 -3430 15795 -3310
rect 15840 -3430 15960 -3310
rect 16005 -3430 16125 -3310
rect 16170 -3430 16290 -3310
rect 16345 -3430 16465 -3310
rect 16510 -3430 16630 -3310
rect 16675 -3430 16795 -3310
rect 16840 -3430 16960 -3310
rect 17015 -3430 17135 -3310
rect 17180 -3430 17300 -3310
rect 17345 -3430 17465 -3310
rect 17510 -3430 17630 -3310
rect 17685 -3430 17805 -3310
rect 17850 -3430 17970 -3310
rect 18015 -3430 18135 -3310
rect 18180 -3430 18300 -3310
rect 12820 -3595 12940 -3475
rect 12995 -3595 13115 -3475
rect 13160 -3595 13280 -3475
rect 13325 -3595 13445 -3475
rect 13490 -3595 13610 -3475
rect 13665 -3595 13785 -3475
rect 13830 -3595 13950 -3475
rect 13995 -3595 14115 -3475
rect 14160 -3595 14280 -3475
rect 14335 -3595 14455 -3475
rect 14500 -3595 14620 -3475
rect 14665 -3595 14785 -3475
rect 14830 -3595 14950 -3475
rect 15005 -3595 15125 -3475
rect 15170 -3595 15290 -3475
rect 15335 -3595 15455 -3475
rect 15500 -3595 15620 -3475
rect 15675 -3595 15795 -3475
rect 15840 -3595 15960 -3475
rect 16005 -3595 16125 -3475
rect 16170 -3595 16290 -3475
rect 16345 -3595 16465 -3475
rect 16510 -3595 16630 -3475
rect 16675 -3595 16795 -3475
rect 16840 -3595 16960 -3475
rect 17015 -3595 17135 -3475
rect 17180 -3595 17300 -3475
rect 17345 -3595 17465 -3475
rect 17510 -3595 17630 -3475
rect 17685 -3595 17805 -3475
rect 17850 -3595 17970 -3475
rect 18015 -3595 18135 -3475
rect 18180 -3595 18300 -3475
rect 12820 -3760 12940 -3640
rect 12995 -3760 13115 -3640
rect 13160 -3760 13280 -3640
rect 13325 -3760 13445 -3640
rect 13490 -3760 13610 -3640
rect 13665 -3760 13785 -3640
rect 13830 -3760 13950 -3640
rect 13995 -3760 14115 -3640
rect 14160 -3760 14280 -3640
rect 14335 -3760 14455 -3640
rect 14500 -3760 14620 -3640
rect 14665 -3760 14785 -3640
rect 14830 -3760 14950 -3640
rect 15005 -3760 15125 -3640
rect 15170 -3760 15290 -3640
rect 15335 -3760 15455 -3640
rect 15500 -3760 15620 -3640
rect 15675 -3760 15795 -3640
rect 15840 -3760 15960 -3640
rect 16005 -3760 16125 -3640
rect 16170 -3760 16290 -3640
rect 16345 -3760 16465 -3640
rect 16510 -3760 16630 -3640
rect 16675 -3760 16795 -3640
rect 16840 -3760 16960 -3640
rect 17015 -3760 17135 -3640
rect 17180 -3760 17300 -3640
rect 17345 -3760 17465 -3640
rect 17510 -3760 17630 -3640
rect 17685 -3760 17805 -3640
rect 17850 -3760 17970 -3640
rect 18015 -3760 18135 -3640
rect 18180 -3760 18300 -3640
rect 12820 -3925 12940 -3805
rect 12995 -3925 13115 -3805
rect 13160 -3925 13280 -3805
rect 13325 -3925 13445 -3805
rect 13490 -3925 13610 -3805
rect 13665 -3925 13785 -3805
rect 13830 -3925 13950 -3805
rect 13995 -3925 14115 -3805
rect 14160 -3925 14280 -3805
rect 14335 -3925 14455 -3805
rect 14500 -3925 14620 -3805
rect 14665 -3925 14785 -3805
rect 14830 -3925 14950 -3805
rect 15005 -3925 15125 -3805
rect 15170 -3925 15290 -3805
rect 15335 -3925 15455 -3805
rect 15500 -3925 15620 -3805
rect 15675 -3925 15795 -3805
rect 15840 -3925 15960 -3805
rect 16005 -3925 16125 -3805
rect 16170 -3925 16290 -3805
rect 16345 -3925 16465 -3805
rect 16510 -3925 16630 -3805
rect 16675 -3925 16795 -3805
rect 16840 -3925 16960 -3805
rect 17015 -3925 17135 -3805
rect 17180 -3925 17300 -3805
rect 17345 -3925 17465 -3805
rect 17510 -3925 17630 -3805
rect 17685 -3925 17805 -3805
rect 17850 -3925 17970 -3805
rect 18015 -3925 18135 -3805
rect 18180 -3925 18300 -3805
rect 12820 -4100 12940 -3980
rect 12995 -4100 13115 -3980
rect 13160 -4100 13280 -3980
rect 13325 -4100 13445 -3980
rect 13490 -4100 13610 -3980
rect 13665 -4100 13785 -3980
rect 13830 -4100 13950 -3980
rect 13995 -4100 14115 -3980
rect 14160 -4100 14280 -3980
rect 14335 -4100 14455 -3980
rect 14500 -4100 14620 -3980
rect 14665 -4100 14785 -3980
rect 14830 -4100 14950 -3980
rect 15005 -4100 15125 -3980
rect 15170 -4100 15290 -3980
rect 15335 -4100 15455 -3980
rect 15500 -4100 15620 -3980
rect 15675 -4100 15795 -3980
rect 15840 -4100 15960 -3980
rect 16005 -4100 16125 -3980
rect 16170 -4100 16290 -3980
rect 16345 -4100 16465 -3980
rect 16510 -4100 16630 -3980
rect 16675 -4100 16795 -3980
rect 16840 -4100 16960 -3980
rect 17015 -4100 17135 -3980
rect 17180 -4100 17300 -3980
rect 17345 -4100 17465 -3980
rect 17510 -4100 17630 -3980
rect 17685 -4100 17805 -3980
rect 17850 -4100 17970 -3980
rect 18015 -4100 18135 -3980
rect 18180 -4100 18300 -3980
rect 18510 1260 18630 1380
rect 18685 1260 18805 1380
rect 18850 1260 18970 1380
rect 19015 1260 19135 1380
rect 19180 1260 19300 1380
rect 19355 1260 19475 1380
rect 19520 1260 19640 1380
rect 19685 1260 19805 1380
rect 19850 1260 19970 1380
rect 20025 1260 20145 1380
rect 20190 1260 20310 1380
rect 20355 1260 20475 1380
rect 20520 1260 20640 1380
rect 20695 1260 20815 1380
rect 20860 1260 20980 1380
rect 21025 1260 21145 1380
rect 21190 1260 21310 1380
rect 21365 1260 21485 1380
rect 21530 1260 21650 1380
rect 21695 1260 21815 1380
rect 21860 1260 21980 1380
rect 22035 1260 22155 1380
rect 22200 1260 22320 1380
rect 22365 1260 22485 1380
rect 22530 1260 22650 1380
rect 22705 1260 22825 1380
rect 22870 1260 22990 1380
rect 23035 1260 23155 1380
rect 23200 1260 23320 1380
rect 23375 1260 23495 1380
rect 23540 1260 23660 1380
rect 23705 1260 23825 1380
rect 23870 1260 23990 1380
rect 18510 1095 18630 1215
rect 18685 1095 18805 1215
rect 18850 1095 18970 1215
rect 19015 1095 19135 1215
rect 19180 1095 19300 1215
rect 19355 1095 19475 1215
rect 19520 1095 19640 1215
rect 19685 1095 19805 1215
rect 19850 1095 19970 1215
rect 20025 1095 20145 1215
rect 20190 1095 20310 1215
rect 20355 1095 20475 1215
rect 20520 1095 20640 1215
rect 20695 1095 20815 1215
rect 20860 1095 20980 1215
rect 21025 1095 21145 1215
rect 21190 1095 21310 1215
rect 21365 1095 21485 1215
rect 21530 1095 21650 1215
rect 21695 1095 21815 1215
rect 21860 1095 21980 1215
rect 22035 1095 22155 1215
rect 22200 1095 22320 1215
rect 22365 1095 22485 1215
rect 22530 1095 22650 1215
rect 22705 1095 22825 1215
rect 22870 1095 22990 1215
rect 23035 1095 23155 1215
rect 23200 1095 23320 1215
rect 23375 1095 23495 1215
rect 23540 1095 23660 1215
rect 23705 1095 23825 1215
rect 23870 1095 23990 1215
rect 18510 930 18630 1050
rect 18685 930 18805 1050
rect 18850 930 18970 1050
rect 19015 930 19135 1050
rect 19180 930 19300 1050
rect 19355 930 19475 1050
rect 19520 930 19640 1050
rect 19685 930 19805 1050
rect 19850 930 19970 1050
rect 20025 930 20145 1050
rect 20190 930 20310 1050
rect 20355 930 20475 1050
rect 20520 930 20640 1050
rect 20695 930 20815 1050
rect 20860 930 20980 1050
rect 21025 930 21145 1050
rect 21190 930 21310 1050
rect 21365 930 21485 1050
rect 21530 930 21650 1050
rect 21695 930 21815 1050
rect 21860 930 21980 1050
rect 22035 930 22155 1050
rect 22200 930 22320 1050
rect 22365 930 22485 1050
rect 22530 930 22650 1050
rect 22705 930 22825 1050
rect 22870 930 22990 1050
rect 23035 930 23155 1050
rect 23200 930 23320 1050
rect 23375 930 23495 1050
rect 23540 930 23660 1050
rect 23705 930 23825 1050
rect 23870 930 23990 1050
rect 18510 765 18630 885
rect 18685 765 18805 885
rect 18850 765 18970 885
rect 19015 765 19135 885
rect 19180 765 19300 885
rect 19355 765 19475 885
rect 19520 765 19640 885
rect 19685 765 19805 885
rect 19850 765 19970 885
rect 20025 765 20145 885
rect 20190 765 20310 885
rect 20355 765 20475 885
rect 20520 765 20640 885
rect 20695 765 20815 885
rect 20860 765 20980 885
rect 21025 765 21145 885
rect 21190 765 21310 885
rect 21365 765 21485 885
rect 21530 765 21650 885
rect 21695 765 21815 885
rect 21860 765 21980 885
rect 22035 765 22155 885
rect 22200 765 22320 885
rect 22365 765 22485 885
rect 22530 765 22650 885
rect 22705 765 22825 885
rect 22870 765 22990 885
rect 23035 765 23155 885
rect 23200 765 23320 885
rect 23375 765 23495 885
rect 23540 765 23660 885
rect 23705 765 23825 885
rect 23870 765 23990 885
rect 18510 590 18630 710
rect 18685 590 18805 710
rect 18850 590 18970 710
rect 19015 590 19135 710
rect 19180 590 19300 710
rect 19355 590 19475 710
rect 19520 590 19640 710
rect 19685 590 19805 710
rect 19850 590 19970 710
rect 20025 590 20145 710
rect 20190 590 20310 710
rect 20355 590 20475 710
rect 20520 590 20640 710
rect 20695 590 20815 710
rect 20860 590 20980 710
rect 21025 590 21145 710
rect 21190 590 21310 710
rect 21365 590 21485 710
rect 21530 590 21650 710
rect 21695 590 21815 710
rect 21860 590 21980 710
rect 22035 590 22155 710
rect 22200 590 22320 710
rect 22365 590 22485 710
rect 22530 590 22650 710
rect 22705 590 22825 710
rect 22870 590 22990 710
rect 23035 590 23155 710
rect 23200 590 23320 710
rect 23375 590 23495 710
rect 23540 590 23660 710
rect 23705 590 23825 710
rect 23870 590 23990 710
rect 18510 425 18630 545
rect 18685 425 18805 545
rect 18850 425 18970 545
rect 19015 425 19135 545
rect 19180 425 19300 545
rect 19355 425 19475 545
rect 19520 425 19640 545
rect 19685 425 19805 545
rect 19850 425 19970 545
rect 20025 425 20145 545
rect 20190 425 20310 545
rect 20355 425 20475 545
rect 20520 425 20640 545
rect 20695 425 20815 545
rect 20860 425 20980 545
rect 21025 425 21145 545
rect 21190 425 21310 545
rect 21365 425 21485 545
rect 21530 425 21650 545
rect 21695 425 21815 545
rect 21860 425 21980 545
rect 22035 425 22155 545
rect 22200 425 22320 545
rect 22365 425 22485 545
rect 22530 425 22650 545
rect 22705 425 22825 545
rect 22870 425 22990 545
rect 23035 425 23155 545
rect 23200 425 23320 545
rect 23375 425 23495 545
rect 23540 425 23660 545
rect 23705 425 23825 545
rect 23870 425 23990 545
rect 18510 260 18630 380
rect 18685 260 18805 380
rect 18850 260 18970 380
rect 19015 260 19135 380
rect 19180 260 19300 380
rect 19355 260 19475 380
rect 19520 260 19640 380
rect 19685 260 19805 380
rect 19850 260 19970 380
rect 20025 260 20145 380
rect 20190 260 20310 380
rect 20355 260 20475 380
rect 20520 260 20640 380
rect 20695 260 20815 380
rect 20860 260 20980 380
rect 21025 260 21145 380
rect 21190 260 21310 380
rect 21365 260 21485 380
rect 21530 260 21650 380
rect 21695 260 21815 380
rect 21860 260 21980 380
rect 22035 260 22155 380
rect 22200 260 22320 380
rect 22365 260 22485 380
rect 22530 260 22650 380
rect 22705 260 22825 380
rect 22870 260 22990 380
rect 23035 260 23155 380
rect 23200 260 23320 380
rect 23375 260 23495 380
rect 23540 260 23660 380
rect 23705 260 23825 380
rect 23870 260 23990 380
rect 18510 95 18630 215
rect 18685 95 18805 215
rect 18850 95 18970 215
rect 19015 95 19135 215
rect 19180 95 19300 215
rect 19355 95 19475 215
rect 19520 95 19640 215
rect 19685 95 19805 215
rect 19850 95 19970 215
rect 20025 95 20145 215
rect 20190 95 20310 215
rect 20355 95 20475 215
rect 20520 95 20640 215
rect 20695 95 20815 215
rect 20860 95 20980 215
rect 21025 95 21145 215
rect 21190 95 21310 215
rect 21365 95 21485 215
rect 21530 95 21650 215
rect 21695 95 21815 215
rect 21860 95 21980 215
rect 22035 95 22155 215
rect 22200 95 22320 215
rect 22365 95 22485 215
rect 22530 95 22650 215
rect 22705 95 22825 215
rect 22870 95 22990 215
rect 23035 95 23155 215
rect 23200 95 23320 215
rect 23375 95 23495 215
rect 23540 95 23660 215
rect 23705 95 23825 215
rect 23870 95 23990 215
rect 18510 -80 18630 40
rect 18685 -80 18805 40
rect 18850 -80 18970 40
rect 19015 -80 19135 40
rect 19180 -80 19300 40
rect 19355 -80 19475 40
rect 19520 -80 19640 40
rect 19685 -80 19805 40
rect 19850 -80 19970 40
rect 20025 -80 20145 40
rect 20190 -80 20310 40
rect 20355 -80 20475 40
rect 20520 -80 20640 40
rect 20695 -80 20815 40
rect 20860 -80 20980 40
rect 21025 -80 21145 40
rect 21190 -80 21310 40
rect 21365 -80 21485 40
rect 21530 -80 21650 40
rect 21695 -80 21815 40
rect 21860 -80 21980 40
rect 22035 -80 22155 40
rect 22200 -80 22320 40
rect 22365 -80 22485 40
rect 22530 -80 22650 40
rect 22705 -80 22825 40
rect 22870 -80 22990 40
rect 23035 -80 23155 40
rect 23200 -80 23320 40
rect 23375 -80 23495 40
rect 23540 -80 23660 40
rect 23705 -80 23825 40
rect 23870 -80 23990 40
rect 18510 -245 18630 -125
rect 18685 -245 18805 -125
rect 18850 -245 18970 -125
rect 19015 -245 19135 -125
rect 19180 -245 19300 -125
rect 19355 -245 19475 -125
rect 19520 -245 19640 -125
rect 19685 -245 19805 -125
rect 19850 -245 19970 -125
rect 20025 -245 20145 -125
rect 20190 -245 20310 -125
rect 20355 -245 20475 -125
rect 20520 -245 20640 -125
rect 20695 -245 20815 -125
rect 20860 -245 20980 -125
rect 21025 -245 21145 -125
rect 21190 -245 21310 -125
rect 21365 -245 21485 -125
rect 21530 -245 21650 -125
rect 21695 -245 21815 -125
rect 21860 -245 21980 -125
rect 22035 -245 22155 -125
rect 22200 -245 22320 -125
rect 22365 -245 22485 -125
rect 22530 -245 22650 -125
rect 22705 -245 22825 -125
rect 22870 -245 22990 -125
rect 23035 -245 23155 -125
rect 23200 -245 23320 -125
rect 23375 -245 23495 -125
rect 23540 -245 23660 -125
rect 23705 -245 23825 -125
rect 23870 -245 23990 -125
rect 18510 -410 18630 -290
rect 18685 -410 18805 -290
rect 18850 -410 18970 -290
rect 19015 -410 19135 -290
rect 19180 -410 19300 -290
rect 19355 -410 19475 -290
rect 19520 -410 19640 -290
rect 19685 -410 19805 -290
rect 19850 -410 19970 -290
rect 20025 -410 20145 -290
rect 20190 -410 20310 -290
rect 20355 -410 20475 -290
rect 20520 -410 20640 -290
rect 20695 -410 20815 -290
rect 20860 -410 20980 -290
rect 21025 -410 21145 -290
rect 21190 -410 21310 -290
rect 21365 -410 21485 -290
rect 21530 -410 21650 -290
rect 21695 -410 21815 -290
rect 21860 -410 21980 -290
rect 22035 -410 22155 -290
rect 22200 -410 22320 -290
rect 22365 -410 22485 -290
rect 22530 -410 22650 -290
rect 22705 -410 22825 -290
rect 22870 -410 22990 -290
rect 23035 -410 23155 -290
rect 23200 -410 23320 -290
rect 23375 -410 23495 -290
rect 23540 -410 23660 -290
rect 23705 -410 23825 -290
rect 23870 -410 23990 -290
rect 18510 -575 18630 -455
rect 18685 -575 18805 -455
rect 18850 -575 18970 -455
rect 19015 -575 19135 -455
rect 19180 -575 19300 -455
rect 19355 -575 19475 -455
rect 19520 -575 19640 -455
rect 19685 -575 19805 -455
rect 19850 -575 19970 -455
rect 20025 -575 20145 -455
rect 20190 -575 20310 -455
rect 20355 -575 20475 -455
rect 20520 -575 20640 -455
rect 20695 -575 20815 -455
rect 20860 -575 20980 -455
rect 21025 -575 21145 -455
rect 21190 -575 21310 -455
rect 21365 -575 21485 -455
rect 21530 -575 21650 -455
rect 21695 -575 21815 -455
rect 21860 -575 21980 -455
rect 22035 -575 22155 -455
rect 22200 -575 22320 -455
rect 22365 -575 22485 -455
rect 22530 -575 22650 -455
rect 22705 -575 22825 -455
rect 22870 -575 22990 -455
rect 23035 -575 23155 -455
rect 23200 -575 23320 -455
rect 23375 -575 23495 -455
rect 23540 -575 23660 -455
rect 23705 -575 23825 -455
rect 23870 -575 23990 -455
rect 18510 -750 18630 -630
rect 18685 -750 18805 -630
rect 18850 -750 18970 -630
rect 19015 -750 19135 -630
rect 19180 -750 19300 -630
rect 19355 -750 19475 -630
rect 19520 -750 19640 -630
rect 19685 -750 19805 -630
rect 19850 -750 19970 -630
rect 20025 -750 20145 -630
rect 20190 -750 20310 -630
rect 20355 -750 20475 -630
rect 20520 -750 20640 -630
rect 20695 -750 20815 -630
rect 20860 -750 20980 -630
rect 21025 -750 21145 -630
rect 21190 -750 21310 -630
rect 21365 -750 21485 -630
rect 21530 -750 21650 -630
rect 21695 -750 21815 -630
rect 21860 -750 21980 -630
rect 22035 -750 22155 -630
rect 22200 -750 22320 -630
rect 22365 -750 22485 -630
rect 22530 -750 22650 -630
rect 22705 -750 22825 -630
rect 22870 -750 22990 -630
rect 23035 -750 23155 -630
rect 23200 -750 23320 -630
rect 23375 -750 23495 -630
rect 23540 -750 23660 -630
rect 23705 -750 23825 -630
rect 23870 -750 23990 -630
rect 18510 -915 18630 -795
rect 18685 -915 18805 -795
rect 18850 -915 18970 -795
rect 19015 -915 19135 -795
rect 19180 -915 19300 -795
rect 19355 -915 19475 -795
rect 19520 -915 19640 -795
rect 19685 -915 19805 -795
rect 19850 -915 19970 -795
rect 20025 -915 20145 -795
rect 20190 -915 20310 -795
rect 20355 -915 20475 -795
rect 20520 -915 20640 -795
rect 20695 -915 20815 -795
rect 20860 -915 20980 -795
rect 21025 -915 21145 -795
rect 21190 -915 21310 -795
rect 21365 -915 21485 -795
rect 21530 -915 21650 -795
rect 21695 -915 21815 -795
rect 21860 -915 21980 -795
rect 22035 -915 22155 -795
rect 22200 -915 22320 -795
rect 22365 -915 22485 -795
rect 22530 -915 22650 -795
rect 22705 -915 22825 -795
rect 22870 -915 22990 -795
rect 23035 -915 23155 -795
rect 23200 -915 23320 -795
rect 23375 -915 23495 -795
rect 23540 -915 23660 -795
rect 23705 -915 23825 -795
rect 23870 -915 23990 -795
rect 18510 -1080 18630 -960
rect 18685 -1080 18805 -960
rect 18850 -1080 18970 -960
rect 19015 -1080 19135 -960
rect 19180 -1080 19300 -960
rect 19355 -1080 19475 -960
rect 19520 -1080 19640 -960
rect 19685 -1080 19805 -960
rect 19850 -1080 19970 -960
rect 20025 -1080 20145 -960
rect 20190 -1080 20310 -960
rect 20355 -1080 20475 -960
rect 20520 -1080 20640 -960
rect 20695 -1080 20815 -960
rect 20860 -1080 20980 -960
rect 21025 -1080 21145 -960
rect 21190 -1080 21310 -960
rect 21365 -1080 21485 -960
rect 21530 -1080 21650 -960
rect 21695 -1080 21815 -960
rect 21860 -1080 21980 -960
rect 22035 -1080 22155 -960
rect 22200 -1080 22320 -960
rect 22365 -1080 22485 -960
rect 22530 -1080 22650 -960
rect 22705 -1080 22825 -960
rect 22870 -1080 22990 -960
rect 23035 -1080 23155 -960
rect 23200 -1080 23320 -960
rect 23375 -1080 23495 -960
rect 23540 -1080 23660 -960
rect 23705 -1080 23825 -960
rect 23870 -1080 23990 -960
rect 18510 -1245 18630 -1125
rect 18685 -1245 18805 -1125
rect 18850 -1245 18970 -1125
rect 19015 -1245 19135 -1125
rect 19180 -1245 19300 -1125
rect 19355 -1245 19475 -1125
rect 19520 -1245 19640 -1125
rect 19685 -1245 19805 -1125
rect 19850 -1245 19970 -1125
rect 20025 -1245 20145 -1125
rect 20190 -1245 20310 -1125
rect 20355 -1245 20475 -1125
rect 20520 -1245 20640 -1125
rect 20695 -1245 20815 -1125
rect 20860 -1245 20980 -1125
rect 21025 -1245 21145 -1125
rect 21190 -1245 21310 -1125
rect 21365 -1245 21485 -1125
rect 21530 -1245 21650 -1125
rect 21695 -1245 21815 -1125
rect 21860 -1245 21980 -1125
rect 22035 -1245 22155 -1125
rect 22200 -1245 22320 -1125
rect 22365 -1245 22485 -1125
rect 22530 -1245 22650 -1125
rect 22705 -1245 22825 -1125
rect 22870 -1245 22990 -1125
rect 23035 -1245 23155 -1125
rect 23200 -1245 23320 -1125
rect 23375 -1245 23495 -1125
rect 23540 -1245 23660 -1125
rect 23705 -1245 23825 -1125
rect 23870 -1245 23990 -1125
rect 18510 -1420 18630 -1300
rect 18685 -1420 18805 -1300
rect 18850 -1420 18970 -1300
rect 19015 -1420 19135 -1300
rect 19180 -1420 19300 -1300
rect 19355 -1420 19475 -1300
rect 19520 -1420 19640 -1300
rect 19685 -1420 19805 -1300
rect 19850 -1420 19970 -1300
rect 20025 -1420 20145 -1300
rect 20190 -1420 20310 -1300
rect 20355 -1420 20475 -1300
rect 20520 -1420 20640 -1300
rect 20695 -1420 20815 -1300
rect 20860 -1420 20980 -1300
rect 21025 -1420 21145 -1300
rect 21190 -1420 21310 -1300
rect 21365 -1420 21485 -1300
rect 21530 -1420 21650 -1300
rect 21695 -1420 21815 -1300
rect 21860 -1420 21980 -1300
rect 22035 -1420 22155 -1300
rect 22200 -1420 22320 -1300
rect 22365 -1420 22485 -1300
rect 22530 -1420 22650 -1300
rect 22705 -1420 22825 -1300
rect 22870 -1420 22990 -1300
rect 23035 -1420 23155 -1300
rect 23200 -1420 23320 -1300
rect 23375 -1420 23495 -1300
rect 23540 -1420 23660 -1300
rect 23705 -1420 23825 -1300
rect 23870 -1420 23990 -1300
rect 18510 -1585 18630 -1465
rect 18685 -1585 18805 -1465
rect 18850 -1585 18970 -1465
rect 19015 -1585 19135 -1465
rect 19180 -1585 19300 -1465
rect 19355 -1585 19475 -1465
rect 19520 -1585 19640 -1465
rect 19685 -1585 19805 -1465
rect 19850 -1585 19970 -1465
rect 20025 -1585 20145 -1465
rect 20190 -1585 20310 -1465
rect 20355 -1585 20475 -1465
rect 20520 -1585 20640 -1465
rect 20695 -1585 20815 -1465
rect 20860 -1585 20980 -1465
rect 21025 -1585 21145 -1465
rect 21190 -1585 21310 -1465
rect 21365 -1585 21485 -1465
rect 21530 -1585 21650 -1465
rect 21695 -1585 21815 -1465
rect 21860 -1585 21980 -1465
rect 22035 -1585 22155 -1465
rect 22200 -1585 22320 -1465
rect 22365 -1585 22485 -1465
rect 22530 -1585 22650 -1465
rect 22705 -1585 22825 -1465
rect 22870 -1585 22990 -1465
rect 23035 -1585 23155 -1465
rect 23200 -1585 23320 -1465
rect 23375 -1585 23495 -1465
rect 23540 -1585 23660 -1465
rect 23705 -1585 23825 -1465
rect 23870 -1585 23990 -1465
rect 18510 -1750 18630 -1630
rect 18685 -1750 18805 -1630
rect 18850 -1750 18970 -1630
rect 19015 -1750 19135 -1630
rect 19180 -1750 19300 -1630
rect 19355 -1750 19475 -1630
rect 19520 -1750 19640 -1630
rect 19685 -1750 19805 -1630
rect 19850 -1750 19970 -1630
rect 20025 -1750 20145 -1630
rect 20190 -1750 20310 -1630
rect 20355 -1750 20475 -1630
rect 20520 -1750 20640 -1630
rect 20695 -1750 20815 -1630
rect 20860 -1750 20980 -1630
rect 21025 -1750 21145 -1630
rect 21190 -1750 21310 -1630
rect 21365 -1750 21485 -1630
rect 21530 -1750 21650 -1630
rect 21695 -1750 21815 -1630
rect 21860 -1750 21980 -1630
rect 22035 -1750 22155 -1630
rect 22200 -1750 22320 -1630
rect 22365 -1750 22485 -1630
rect 22530 -1750 22650 -1630
rect 22705 -1750 22825 -1630
rect 22870 -1750 22990 -1630
rect 23035 -1750 23155 -1630
rect 23200 -1750 23320 -1630
rect 23375 -1750 23495 -1630
rect 23540 -1750 23660 -1630
rect 23705 -1750 23825 -1630
rect 23870 -1750 23990 -1630
rect 18510 -1915 18630 -1795
rect 18685 -1915 18805 -1795
rect 18850 -1915 18970 -1795
rect 19015 -1915 19135 -1795
rect 19180 -1915 19300 -1795
rect 19355 -1915 19475 -1795
rect 19520 -1915 19640 -1795
rect 19685 -1915 19805 -1795
rect 19850 -1915 19970 -1795
rect 20025 -1915 20145 -1795
rect 20190 -1915 20310 -1795
rect 20355 -1915 20475 -1795
rect 20520 -1915 20640 -1795
rect 20695 -1915 20815 -1795
rect 20860 -1915 20980 -1795
rect 21025 -1915 21145 -1795
rect 21190 -1915 21310 -1795
rect 21365 -1915 21485 -1795
rect 21530 -1915 21650 -1795
rect 21695 -1915 21815 -1795
rect 21860 -1915 21980 -1795
rect 22035 -1915 22155 -1795
rect 22200 -1915 22320 -1795
rect 22365 -1915 22485 -1795
rect 22530 -1915 22650 -1795
rect 22705 -1915 22825 -1795
rect 22870 -1915 22990 -1795
rect 23035 -1915 23155 -1795
rect 23200 -1915 23320 -1795
rect 23375 -1915 23495 -1795
rect 23540 -1915 23660 -1795
rect 23705 -1915 23825 -1795
rect 23870 -1915 23990 -1795
rect 18510 -2090 18630 -1970
rect 18685 -2090 18805 -1970
rect 18850 -2090 18970 -1970
rect 19015 -2090 19135 -1970
rect 19180 -2090 19300 -1970
rect 19355 -2090 19475 -1970
rect 19520 -2090 19640 -1970
rect 19685 -2090 19805 -1970
rect 19850 -2090 19970 -1970
rect 20025 -2090 20145 -1970
rect 20190 -2090 20310 -1970
rect 20355 -2090 20475 -1970
rect 20520 -2090 20640 -1970
rect 20695 -2090 20815 -1970
rect 20860 -2090 20980 -1970
rect 21025 -2090 21145 -1970
rect 21190 -2090 21310 -1970
rect 21365 -2090 21485 -1970
rect 21530 -2090 21650 -1970
rect 21695 -2090 21815 -1970
rect 21860 -2090 21980 -1970
rect 22035 -2090 22155 -1970
rect 22200 -2090 22320 -1970
rect 22365 -2090 22485 -1970
rect 22530 -2090 22650 -1970
rect 22705 -2090 22825 -1970
rect 22870 -2090 22990 -1970
rect 23035 -2090 23155 -1970
rect 23200 -2090 23320 -1970
rect 23375 -2090 23495 -1970
rect 23540 -2090 23660 -1970
rect 23705 -2090 23825 -1970
rect 23870 -2090 23990 -1970
rect 18510 -2255 18630 -2135
rect 18685 -2255 18805 -2135
rect 18850 -2255 18970 -2135
rect 19015 -2255 19135 -2135
rect 19180 -2255 19300 -2135
rect 19355 -2255 19475 -2135
rect 19520 -2255 19640 -2135
rect 19685 -2255 19805 -2135
rect 19850 -2255 19970 -2135
rect 20025 -2255 20145 -2135
rect 20190 -2255 20310 -2135
rect 20355 -2255 20475 -2135
rect 20520 -2255 20640 -2135
rect 20695 -2255 20815 -2135
rect 20860 -2255 20980 -2135
rect 21025 -2255 21145 -2135
rect 21190 -2255 21310 -2135
rect 21365 -2255 21485 -2135
rect 21530 -2255 21650 -2135
rect 21695 -2255 21815 -2135
rect 21860 -2255 21980 -2135
rect 22035 -2255 22155 -2135
rect 22200 -2255 22320 -2135
rect 22365 -2255 22485 -2135
rect 22530 -2255 22650 -2135
rect 22705 -2255 22825 -2135
rect 22870 -2255 22990 -2135
rect 23035 -2255 23155 -2135
rect 23200 -2255 23320 -2135
rect 23375 -2255 23495 -2135
rect 23540 -2255 23660 -2135
rect 23705 -2255 23825 -2135
rect 23870 -2255 23990 -2135
rect 18510 -2420 18630 -2300
rect 18685 -2420 18805 -2300
rect 18850 -2420 18970 -2300
rect 19015 -2420 19135 -2300
rect 19180 -2420 19300 -2300
rect 19355 -2420 19475 -2300
rect 19520 -2420 19640 -2300
rect 19685 -2420 19805 -2300
rect 19850 -2420 19970 -2300
rect 20025 -2420 20145 -2300
rect 20190 -2420 20310 -2300
rect 20355 -2420 20475 -2300
rect 20520 -2420 20640 -2300
rect 20695 -2420 20815 -2300
rect 20860 -2420 20980 -2300
rect 21025 -2420 21145 -2300
rect 21190 -2420 21310 -2300
rect 21365 -2420 21485 -2300
rect 21530 -2420 21650 -2300
rect 21695 -2420 21815 -2300
rect 21860 -2420 21980 -2300
rect 22035 -2420 22155 -2300
rect 22200 -2420 22320 -2300
rect 22365 -2420 22485 -2300
rect 22530 -2420 22650 -2300
rect 22705 -2420 22825 -2300
rect 22870 -2420 22990 -2300
rect 23035 -2420 23155 -2300
rect 23200 -2420 23320 -2300
rect 23375 -2420 23495 -2300
rect 23540 -2420 23660 -2300
rect 23705 -2420 23825 -2300
rect 23870 -2420 23990 -2300
rect 18510 -2585 18630 -2465
rect 18685 -2585 18805 -2465
rect 18850 -2585 18970 -2465
rect 19015 -2585 19135 -2465
rect 19180 -2585 19300 -2465
rect 19355 -2585 19475 -2465
rect 19520 -2585 19640 -2465
rect 19685 -2585 19805 -2465
rect 19850 -2585 19970 -2465
rect 20025 -2585 20145 -2465
rect 20190 -2585 20310 -2465
rect 20355 -2585 20475 -2465
rect 20520 -2585 20640 -2465
rect 20695 -2585 20815 -2465
rect 20860 -2585 20980 -2465
rect 21025 -2585 21145 -2465
rect 21190 -2585 21310 -2465
rect 21365 -2585 21485 -2465
rect 21530 -2585 21650 -2465
rect 21695 -2585 21815 -2465
rect 21860 -2585 21980 -2465
rect 22035 -2585 22155 -2465
rect 22200 -2585 22320 -2465
rect 22365 -2585 22485 -2465
rect 22530 -2585 22650 -2465
rect 22705 -2585 22825 -2465
rect 22870 -2585 22990 -2465
rect 23035 -2585 23155 -2465
rect 23200 -2585 23320 -2465
rect 23375 -2585 23495 -2465
rect 23540 -2585 23660 -2465
rect 23705 -2585 23825 -2465
rect 23870 -2585 23990 -2465
rect 18510 -2760 18630 -2640
rect 18685 -2760 18805 -2640
rect 18850 -2760 18970 -2640
rect 19015 -2760 19135 -2640
rect 19180 -2760 19300 -2640
rect 19355 -2760 19475 -2640
rect 19520 -2760 19640 -2640
rect 19685 -2760 19805 -2640
rect 19850 -2760 19970 -2640
rect 20025 -2760 20145 -2640
rect 20190 -2760 20310 -2640
rect 20355 -2760 20475 -2640
rect 20520 -2760 20640 -2640
rect 20695 -2760 20815 -2640
rect 20860 -2760 20980 -2640
rect 21025 -2760 21145 -2640
rect 21190 -2760 21310 -2640
rect 21365 -2760 21485 -2640
rect 21530 -2760 21650 -2640
rect 21695 -2760 21815 -2640
rect 21860 -2760 21980 -2640
rect 22035 -2760 22155 -2640
rect 22200 -2760 22320 -2640
rect 22365 -2760 22485 -2640
rect 22530 -2760 22650 -2640
rect 22705 -2760 22825 -2640
rect 22870 -2760 22990 -2640
rect 23035 -2760 23155 -2640
rect 23200 -2760 23320 -2640
rect 23375 -2760 23495 -2640
rect 23540 -2760 23660 -2640
rect 23705 -2760 23825 -2640
rect 23870 -2760 23990 -2640
rect 18510 -2925 18630 -2805
rect 18685 -2925 18805 -2805
rect 18850 -2925 18970 -2805
rect 19015 -2925 19135 -2805
rect 19180 -2925 19300 -2805
rect 19355 -2925 19475 -2805
rect 19520 -2925 19640 -2805
rect 19685 -2925 19805 -2805
rect 19850 -2925 19970 -2805
rect 20025 -2925 20145 -2805
rect 20190 -2925 20310 -2805
rect 20355 -2925 20475 -2805
rect 20520 -2925 20640 -2805
rect 20695 -2925 20815 -2805
rect 20860 -2925 20980 -2805
rect 21025 -2925 21145 -2805
rect 21190 -2925 21310 -2805
rect 21365 -2925 21485 -2805
rect 21530 -2925 21650 -2805
rect 21695 -2925 21815 -2805
rect 21860 -2925 21980 -2805
rect 22035 -2925 22155 -2805
rect 22200 -2925 22320 -2805
rect 22365 -2925 22485 -2805
rect 22530 -2925 22650 -2805
rect 22705 -2925 22825 -2805
rect 22870 -2925 22990 -2805
rect 23035 -2925 23155 -2805
rect 23200 -2925 23320 -2805
rect 23375 -2925 23495 -2805
rect 23540 -2925 23660 -2805
rect 23705 -2925 23825 -2805
rect 23870 -2925 23990 -2805
rect 18510 -3090 18630 -2970
rect 18685 -3090 18805 -2970
rect 18850 -3090 18970 -2970
rect 19015 -3090 19135 -2970
rect 19180 -3090 19300 -2970
rect 19355 -3090 19475 -2970
rect 19520 -3090 19640 -2970
rect 19685 -3090 19805 -2970
rect 19850 -3090 19970 -2970
rect 20025 -3090 20145 -2970
rect 20190 -3090 20310 -2970
rect 20355 -3090 20475 -2970
rect 20520 -3090 20640 -2970
rect 20695 -3090 20815 -2970
rect 20860 -3090 20980 -2970
rect 21025 -3090 21145 -2970
rect 21190 -3090 21310 -2970
rect 21365 -3090 21485 -2970
rect 21530 -3090 21650 -2970
rect 21695 -3090 21815 -2970
rect 21860 -3090 21980 -2970
rect 22035 -3090 22155 -2970
rect 22200 -3090 22320 -2970
rect 22365 -3090 22485 -2970
rect 22530 -3090 22650 -2970
rect 22705 -3090 22825 -2970
rect 22870 -3090 22990 -2970
rect 23035 -3090 23155 -2970
rect 23200 -3090 23320 -2970
rect 23375 -3090 23495 -2970
rect 23540 -3090 23660 -2970
rect 23705 -3090 23825 -2970
rect 23870 -3090 23990 -2970
rect 18510 -3255 18630 -3135
rect 18685 -3255 18805 -3135
rect 18850 -3255 18970 -3135
rect 19015 -3255 19135 -3135
rect 19180 -3255 19300 -3135
rect 19355 -3255 19475 -3135
rect 19520 -3255 19640 -3135
rect 19685 -3255 19805 -3135
rect 19850 -3255 19970 -3135
rect 20025 -3255 20145 -3135
rect 20190 -3255 20310 -3135
rect 20355 -3255 20475 -3135
rect 20520 -3255 20640 -3135
rect 20695 -3255 20815 -3135
rect 20860 -3255 20980 -3135
rect 21025 -3255 21145 -3135
rect 21190 -3255 21310 -3135
rect 21365 -3255 21485 -3135
rect 21530 -3255 21650 -3135
rect 21695 -3255 21815 -3135
rect 21860 -3255 21980 -3135
rect 22035 -3255 22155 -3135
rect 22200 -3255 22320 -3135
rect 22365 -3255 22485 -3135
rect 22530 -3255 22650 -3135
rect 22705 -3255 22825 -3135
rect 22870 -3255 22990 -3135
rect 23035 -3255 23155 -3135
rect 23200 -3255 23320 -3135
rect 23375 -3255 23495 -3135
rect 23540 -3255 23660 -3135
rect 23705 -3255 23825 -3135
rect 23870 -3255 23990 -3135
rect 18510 -3430 18630 -3310
rect 18685 -3430 18805 -3310
rect 18850 -3430 18970 -3310
rect 19015 -3430 19135 -3310
rect 19180 -3430 19300 -3310
rect 19355 -3430 19475 -3310
rect 19520 -3430 19640 -3310
rect 19685 -3430 19805 -3310
rect 19850 -3430 19970 -3310
rect 20025 -3430 20145 -3310
rect 20190 -3430 20310 -3310
rect 20355 -3430 20475 -3310
rect 20520 -3430 20640 -3310
rect 20695 -3430 20815 -3310
rect 20860 -3430 20980 -3310
rect 21025 -3430 21145 -3310
rect 21190 -3430 21310 -3310
rect 21365 -3430 21485 -3310
rect 21530 -3430 21650 -3310
rect 21695 -3430 21815 -3310
rect 21860 -3430 21980 -3310
rect 22035 -3430 22155 -3310
rect 22200 -3430 22320 -3310
rect 22365 -3430 22485 -3310
rect 22530 -3430 22650 -3310
rect 22705 -3430 22825 -3310
rect 22870 -3430 22990 -3310
rect 23035 -3430 23155 -3310
rect 23200 -3430 23320 -3310
rect 23375 -3430 23495 -3310
rect 23540 -3430 23660 -3310
rect 23705 -3430 23825 -3310
rect 23870 -3430 23990 -3310
rect 18510 -3595 18630 -3475
rect 18685 -3595 18805 -3475
rect 18850 -3595 18970 -3475
rect 19015 -3595 19135 -3475
rect 19180 -3595 19300 -3475
rect 19355 -3595 19475 -3475
rect 19520 -3595 19640 -3475
rect 19685 -3595 19805 -3475
rect 19850 -3595 19970 -3475
rect 20025 -3595 20145 -3475
rect 20190 -3595 20310 -3475
rect 20355 -3595 20475 -3475
rect 20520 -3595 20640 -3475
rect 20695 -3595 20815 -3475
rect 20860 -3595 20980 -3475
rect 21025 -3595 21145 -3475
rect 21190 -3595 21310 -3475
rect 21365 -3595 21485 -3475
rect 21530 -3595 21650 -3475
rect 21695 -3595 21815 -3475
rect 21860 -3595 21980 -3475
rect 22035 -3595 22155 -3475
rect 22200 -3595 22320 -3475
rect 22365 -3595 22485 -3475
rect 22530 -3595 22650 -3475
rect 22705 -3595 22825 -3475
rect 22870 -3595 22990 -3475
rect 23035 -3595 23155 -3475
rect 23200 -3595 23320 -3475
rect 23375 -3595 23495 -3475
rect 23540 -3595 23660 -3475
rect 23705 -3595 23825 -3475
rect 23870 -3595 23990 -3475
rect 18510 -3760 18630 -3640
rect 18685 -3760 18805 -3640
rect 18850 -3760 18970 -3640
rect 19015 -3760 19135 -3640
rect 19180 -3760 19300 -3640
rect 19355 -3760 19475 -3640
rect 19520 -3760 19640 -3640
rect 19685 -3760 19805 -3640
rect 19850 -3760 19970 -3640
rect 20025 -3760 20145 -3640
rect 20190 -3760 20310 -3640
rect 20355 -3760 20475 -3640
rect 20520 -3760 20640 -3640
rect 20695 -3760 20815 -3640
rect 20860 -3760 20980 -3640
rect 21025 -3760 21145 -3640
rect 21190 -3760 21310 -3640
rect 21365 -3760 21485 -3640
rect 21530 -3760 21650 -3640
rect 21695 -3760 21815 -3640
rect 21860 -3760 21980 -3640
rect 22035 -3760 22155 -3640
rect 22200 -3760 22320 -3640
rect 22365 -3760 22485 -3640
rect 22530 -3760 22650 -3640
rect 22705 -3760 22825 -3640
rect 22870 -3760 22990 -3640
rect 23035 -3760 23155 -3640
rect 23200 -3760 23320 -3640
rect 23375 -3760 23495 -3640
rect 23540 -3760 23660 -3640
rect 23705 -3760 23825 -3640
rect 23870 -3760 23990 -3640
rect 18510 -3925 18630 -3805
rect 18685 -3925 18805 -3805
rect 18850 -3925 18970 -3805
rect 19015 -3925 19135 -3805
rect 19180 -3925 19300 -3805
rect 19355 -3925 19475 -3805
rect 19520 -3925 19640 -3805
rect 19685 -3925 19805 -3805
rect 19850 -3925 19970 -3805
rect 20025 -3925 20145 -3805
rect 20190 -3925 20310 -3805
rect 20355 -3925 20475 -3805
rect 20520 -3925 20640 -3805
rect 20695 -3925 20815 -3805
rect 20860 -3925 20980 -3805
rect 21025 -3925 21145 -3805
rect 21190 -3925 21310 -3805
rect 21365 -3925 21485 -3805
rect 21530 -3925 21650 -3805
rect 21695 -3925 21815 -3805
rect 21860 -3925 21980 -3805
rect 22035 -3925 22155 -3805
rect 22200 -3925 22320 -3805
rect 22365 -3925 22485 -3805
rect 22530 -3925 22650 -3805
rect 22705 -3925 22825 -3805
rect 22870 -3925 22990 -3805
rect 23035 -3925 23155 -3805
rect 23200 -3925 23320 -3805
rect 23375 -3925 23495 -3805
rect 23540 -3925 23660 -3805
rect 23705 -3925 23825 -3805
rect 23870 -3925 23990 -3805
rect 18510 -4100 18630 -3980
rect 18685 -4100 18805 -3980
rect 18850 -4100 18970 -3980
rect 19015 -4100 19135 -3980
rect 19180 -4100 19300 -3980
rect 19355 -4100 19475 -3980
rect 19520 -4100 19640 -3980
rect 19685 -4100 19805 -3980
rect 19850 -4100 19970 -3980
rect 20025 -4100 20145 -3980
rect 20190 -4100 20310 -3980
rect 20355 -4100 20475 -3980
rect 20520 -4100 20640 -3980
rect 20695 -4100 20815 -3980
rect 20860 -4100 20980 -3980
rect 21025 -4100 21145 -3980
rect 21190 -4100 21310 -3980
rect 21365 -4100 21485 -3980
rect 21530 -4100 21650 -3980
rect 21695 -4100 21815 -3980
rect 21860 -4100 21980 -3980
rect 22035 -4100 22155 -3980
rect 22200 -4100 22320 -3980
rect 22365 -4100 22485 -3980
rect 22530 -4100 22650 -3980
rect 22705 -4100 22825 -3980
rect 22870 -4100 22990 -3980
rect 23035 -4100 23155 -3980
rect 23200 -4100 23320 -3980
rect 23375 -4100 23495 -3980
rect 23540 -4100 23660 -3980
rect 23705 -4100 23825 -3980
rect 23870 -4100 23990 -3980
rect 24200 1260 24320 1380
rect 24375 1260 24495 1380
rect 24540 1260 24660 1380
rect 24705 1260 24825 1380
rect 24870 1260 24990 1380
rect 25045 1260 25165 1380
rect 25210 1260 25330 1380
rect 25375 1260 25495 1380
rect 25540 1260 25660 1380
rect 25715 1260 25835 1380
rect 25880 1260 26000 1380
rect 26045 1260 26165 1380
rect 26210 1260 26330 1380
rect 26385 1260 26505 1380
rect 26550 1260 26670 1380
rect 26715 1260 26835 1380
rect 26880 1260 27000 1380
rect 27055 1260 27175 1380
rect 27220 1260 27340 1380
rect 27385 1260 27505 1380
rect 27550 1260 27670 1380
rect 27725 1260 27845 1380
rect 27890 1260 28010 1380
rect 28055 1260 28175 1380
rect 28220 1260 28340 1380
rect 28395 1260 28515 1380
rect 28560 1260 28680 1380
rect 28725 1260 28845 1380
rect 28890 1260 29010 1380
rect 29065 1260 29185 1380
rect 29230 1260 29350 1380
rect 29395 1260 29515 1380
rect 29560 1260 29680 1380
rect 24200 1095 24320 1215
rect 24375 1095 24495 1215
rect 24540 1095 24660 1215
rect 24705 1095 24825 1215
rect 24870 1095 24990 1215
rect 25045 1095 25165 1215
rect 25210 1095 25330 1215
rect 25375 1095 25495 1215
rect 25540 1095 25660 1215
rect 25715 1095 25835 1215
rect 25880 1095 26000 1215
rect 26045 1095 26165 1215
rect 26210 1095 26330 1215
rect 26385 1095 26505 1215
rect 26550 1095 26670 1215
rect 26715 1095 26835 1215
rect 26880 1095 27000 1215
rect 27055 1095 27175 1215
rect 27220 1095 27340 1215
rect 27385 1095 27505 1215
rect 27550 1095 27670 1215
rect 27725 1095 27845 1215
rect 27890 1095 28010 1215
rect 28055 1095 28175 1215
rect 28220 1095 28340 1215
rect 28395 1095 28515 1215
rect 28560 1095 28680 1215
rect 28725 1095 28845 1215
rect 28890 1095 29010 1215
rect 29065 1095 29185 1215
rect 29230 1095 29350 1215
rect 29395 1095 29515 1215
rect 29560 1095 29680 1215
rect 24200 930 24320 1050
rect 24375 930 24495 1050
rect 24540 930 24660 1050
rect 24705 930 24825 1050
rect 24870 930 24990 1050
rect 25045 930 25165 1050
rect 25210 930 25330 1050
rect 25375 930 25495 1050
rect 25540 930 25660 1050
rect 25715 930 25835 1050
rect 25880 930 26000 1050
rect 26045 930 26165 1050
rect 26210 930 26330 1050
rect 26385 930 26505 1050
rect 26550 930 26670 1050
rect 26715 930 26835 1050
rect 26880 930 27000 1050
rect 27055 930 27175 1050
rect 27220 930 27340 1050
rect 27385 930 27505 1050
rect 27550 930 27670 1050
rect 27725 930 27845 1050
rect 27890 930 28010 1050
rect 28055 930 28175 1050
rect 28220 930 28340 1050
rect 28395 930 28515 1050
rect 28560 930 28680 1050
rect 28725 930 28845 1050
rect 28890 930 29010 1050
rect 29065 930 29185 1050
rect 29230 930 29350 1050
rect 29395 930 29515 1050
rect 29560 930 29680 1050
rect 24200 765 24320 885
rect 24375 765 24495 885
rect 24540 765 24660 885
rect 24705 765 24825 885
rect 24870 765 24990 885
rect 25045 765 25165 885
rect 25210 765 25330 885
rect 25375 765 25495 885
rect 25540 765 25660 885
rect 25715 765 25835 885
rect 25880 765 26000 885
rect 26045 765 26165 885
rect 26210 765 26330 885
rect 26385 765 26505 885
rect 26550 765 26670 885
rect 26715 765 26835 885
rect 26880 765 27000 885
rect 27055 765 27175 885
rect 27220 765 27340 885
rect 27385 765 27505 885
rect 27550 765 27670 885
rect 27725 765 27845 885
rect 27890 765 28010 885
rect 28055 765 28175 885
rect 28220 765 28340 885
rect 28395 765 28515 885
rect 28560 765 28680 885
rect 28725 765 28845 885
rect 28890 765 29010 885
rect 29065 765 29185 885
rect 29230 765 29350 885
rect 29395 765 29515 885
rect 29560 765 29680 885
rect 24200 590 24320 710
rect 24375 590 24495 710
rect 24540 590 24660 710
rect 24705 590 24825 710
rect 24870 590 24990 710
rect 25045 590 25165 710
rect 25210 590 25330 710
rect 25375 590 25495 710
rect 25540 590 25660 710
rect 25715 590 25835 710
rect 25880 590 26000 710
rect 26045 590 26165 710
rect 26210 590 26330 710
rect 26385 590 26505 710
rect 26550 590 26670 710
rect 26715 590 26835 710
rect 26880 590 27000 710
rect 27055 590 27175 710
rect 27220 590 27340 710
rect 27385 590 27505 710
rect 27550 590 27670 710
rect 27725 590 27845 710
rect 27890 590 28010 710
rect 28055 590 28175 710
rect 28220 590 28340 710
rect 28395 590 28515 710
rect 28560 590 28680 710
rect 28725 590 28845 710
rect 28890 590 29010 710
rect 29065 590 29185 710
rect 29230 590 29350 710
rect 29395 590 29515 710
rect 29560 590 29680 710
rect 24200 425 24320 545
rect 24375 425 24495 545
rect 24540 425 24660 545
rect 24705 425 24825 545
rect 24870 425 24990 545
rect 25045 425 25165 545
rect 25210 425 25330 545
rect 25375 425 25495 545
rect 25540 425 25660 545
rect 25715 425 25835 545
rect 25880 425 26000 545
rect 26045 425 26165 545
rect 26210 425 26330 545
rect 26385 425 26505 545
rect 26550 425 26670 545
rect 26715 425 26835 545
rect 26880 425 27000 545
rect 27055 425 27175 545
rect 27220 425 27340 545
rect 27385 425 27505 545
rect 27550 425 27670 545
rect 27725 425 27845 545
rect 27890 425 28010 545
rect 28055 425 28175 545
rect 28220 425 28340 545
rect 28395 425 28515 545
rect 28560 425 28680 545
rect 28725 425 28845 545
rect 28890 425 29010 545
rect 29065 425 29185 545
rect 29230 425 29350 545
rect 29395 425 29515 545
rect 29560 425 29680 545
rect 24200 260 24320 380
rect 24375 260 24495 380
rect 24540 260 24660 380
rect 24705 260 24825 380
rect 24870 260 24990 380
rect 25045 260 25165 380
rect 25210 260 25330 380
rect 25375 260 25495 380
rect 25540 260 25660 380
rect 25715 260 25835 380
rect 25880 260 26000 380
rect 26045 260 26165 380
rect 26210 260 26330 380
rect 26385 260 26505 380
rect 26550 260 26670 380
rect 26715 260 26835 380
rect 26880 260 27000 380
rect 27055 260 27175 380
rect 27220 260 27340 380
rect 27385 260 27505 380
rect 27550 260 27670 380
rect 27725 260 27845 380
rect 27890 260 28010 380
rect 28055 260 28175 380
rect 28220 260 28340 380
rect 28395 260 28515 380
rect 28560 260 28680 380
rect 28725 260 28845 380
rect 28890 260 29010 380
rect 29065 260 29185 380
rect 29230 260 29350 380
rect 29395 260 29515 380
rect 29560 260 29680 380
rect 24200 95 24320 215
rect 24375 95 24495 215
rect 24540 95 24660 215
rect 24705 95 24825 215
rect 24870 95 24990 215
rect 25045 95 25165 215
rect 25210 95 25330 215
rect 25375 95 25495 215
rect 25540 95 25660 215
rect 25715 95 25835 215
rect 25880 95 26000 215
rect 26045 95 26165 215
rect 26210 95 26330 215
rect 26385 95 26505 215
rect 26550 95 26670 215
rect 26715 95 26835 215
rect 26880 95 27000 215
rect 27055 95 27175 215
rect 27220 95 27340 215
rect 27385 95 27505 215
rect 27550 95 27670 215
rect 27725 95 27845 215
rect 27890 95 28010 215
rect 28055 95 28175 215
rect 28220 95 28340 215
rect 28395 95 28515 215
rect 28560 95 28680 215
rect 28725 95 28845 215
rect 28890 95 29010 215
rect 29065 95 29185 215
rect 29230 95 29350 215
rect 29395 95 29515 215
rect 29560 95 29680 215
rect 24200 -80 24320 40
rect 24375 -80 24495 40
rect 24540 -80 24660 40
rect 24705 -80 24825 40
rect 24870 -80 24990 40
rect 25045 -80 25165 40
rect 25210 -80 25330 40
rect 25375 -80 25495 40
rect 25540 -80 25660 40
rect 25715 -80 25835 40
rect 25880 -80 26000 40
rect 26045 -80 26165 40
rect 26210 -80 26330 40
rect 26385 -80 26505 40
rect 26550 -80 26670 40
rect 26715 -80 26835 40
rect 26880 -80 27000 40
rect 27055 -80 27175 40
rect 27220 -80 27340 40
rect 27385 -80 27505 40
rect 27550 -80 27670 40
rect 27725 -80 27845 40
rect 27890 -80 28010 40
rect 28055 -80 28175 40
rect 28220 -80 28340 40
rect 28395 -80 28515 40
rect 28560 -80 28680 40
rect 28725 -80 28845 40
rect 28890 -80 29010 40
rect 29065 -80 29185 40
rect 29230 -80 29350 40
rect 29395 -80 29515 40
rect 29560 -80 29680 40
rect 24200 -245 24320 -125
rect 24375 -245 24495 -125
rect 24540 -245 24660 -125
rect 24705 -245 24825 -125
rect 24870 -245 24990 -125
rect 25045 -245 25165 -125
rect 25210 -245 25330 -125
rect 25375 -245 25495 -125
rect 25540 -245 25660 -125
rect 25715 -245 25835 -125
rect 25880 -245 26000 -125
rect 26045 -245 26165 -125
rect 26210 -245 26330 -125
rect 26385 -245 26505 -125
rect 26550 -245 26670 -125
rect 26715 -245 26835 -125
rect 26880 -245 27000 -125
rect 27055 -245 27175 -125
rect 27220 -245 27340 -125
rect 27385 -245 27505 -125
rect 27550 -245 27670 -125
rect 27725 -245 27845 -125
rect 27890 -245 28010 -125
rect 28055 -245 28175 -125
rect 28220 -245 28340 -125
rect 28395 -245 28515 -125
rect 28560 -245 28680 -125
rect 28725 -245 28845 -125
rect 28890 -245 29010 -125
rect 29065 -245 29185 -125
rect 29230 -245 29350 -125
rect 29395 -245 29515 -125
rect 29560 -245 29680 -125
rect 24200 -410 24320 -290
rect 24375 -410 24495 -290
rect 24540 -410 24660 -290
rect 24705 -410 24825 -290
rect 24870 -410 24990 -290
rect 25045 -410 25165 -290
rect 25210 -410 25330 -290
rect 25375 -410 25495 -290
rect 25540 -410 25660 -290
rect 25715 -410 25835 -290
rect 25880 -410 26000 -290
rect 26045 -410 26165 -290
rect 26210 -410 26330 -290
rect 26385 -410 26505 -290
rect 26550 -410 26670 -290
rect 26715 -410 26835 -290
rect 26880 -410 27000 -290
rect 27055 -410 27175 -290
rect 27220 -410 27340 -290
rect 27385 -410 27505 -290
rect 27550 -410 27670 -290
rect 27725 -410 27845 -290
rect 27890 -410 28010 -290
rect 28055 -410 28175 -290
rect 28220 -410 28340 -290
rect 28395 -410 28515 -290
rect 28560 -410 28680 -290
rect 28725 -410 28845 -290
rect 28890 -410 29010 -290
rect 29065 -410 29185 -290
rect 29230 -410 29350 -290
rect 29395 -410 29515 -290
rect 29560 -410 29680 -290
rect 24200 -575 24320 -455
rect 24375 -575 24495 -455
rect 24540 -575 24660 -455
rect 24705 -575 24825 -455
rect 24870 -575 24990 -455
rect 25045 -575 25165 -455
rect 25210 -575 25330 -455
rect 25375 -575 25495 -455
rect 25540 -575 25660 -455
rect 25715 -575 25835 -455
rect 25880 -575 26000 -455
rect 26045 -575 26165 -455
rect 26210 -575 26330 -455
rect 26385 -575 26505 -455
rect 26550 -575 26670 -455
rect 26715 -575 26835 -455
rect 26880 -575 27000 -455
rect 27055 -575 27175 -455
rect 27220 -575 27340 -455
rect 27385 -575 27505 -455
rect 27550 -575 27670 -455
rect 27725 -575 27845 -455
rect 27890 -575 28010 -455
rect 28055 -575 28175 -455
rect 28220 -575 28340 -455
rect 28395 -575 28515 -455
rect 28560 -575 28680 -455
rect 28725 -575 28845 -455
rect 28890 -575 29010 -455
rect 29065 -575 29185 -455
rect 29230 -575 29350 -455
rect 29395 -575 29515 -455
rect 29560 -575 29680 -455
rect 24200 -750 24320 -630
rect 24375 -750 24495 -630
rect 24540 -750 24660 -630
rect 24705 -750 24825 -630
rect 24870 -750 24990 -630
rect 25045 -750 25165 -630
rect 25210 -750 25330 -630
rect 25375 -750 25495 -630
rect 25540 -750 25660 -630
rect 25715 -750 25835 -630
rect 25880 -750 26000 -630
rect 26045 -750 26165 -630
rect 26210 -750 26330 -630
rect 26385 -750 26505 -630
rect 26550 -750 26670 -630
rect 26715 -750 26835 -630
rect 26880 -750 27000 -630
rect 27055 -750 27175 -630
rect 27220 -750 27340 -630
rect 27385 -750 27505 -630
rect 27550 -750 27670 -630
rect 27725 -750 27845 -630
rect 27890 -750 28010 -630
rect 28055 -750 28175 -630
rect 28220 -750 28340 -630
rect 28395 -750 28515 -630
rect 28560 -750 28680 -630
rect 28725 -750 28845 -630
rect 28890 -750 29010 -630
rect 29065 -750 29185 -630
rect 29230 -750 29350 -630
rect 29395 -750 29515 -630
rect 29560 -750 29680 -630
rect 24200 -915 24320 -795
rect 24375 -915 24495 -795
rect 24540 -915 24660 -795
rect 24705 -915 24825 -795
rect 24870 -915 24990 -795
rect 25045 -915 25165 -795
rect 25210 -915 25330 -795
rect 25375 -915 25495 -795
rect 25540 -915 25660 -795
rect 25715 -915 25835 -795
rect 25880 -915 26000 -795
rect 26045 -915 26165 -795
rect 26210 -915 26330 -795
rect 26385 -915 26505 -795
rect 26550 -915 26670 -795
rect 26715 -915 26835 -795
rect 26880 -915 27000 -795
rect 27055 -915 27175 -795
rect 27220 -915 27340 -795
rect 27385 -915 27505 -795
rect 27550 -915 27670 -795
rect 27725 -915 27845 -795
rect 27890 -915 28010 -795
rect 28055 -915 28175 -795
rect 28220 -915 28340 -795
rect 28395 -915 28515 -795
rect 28560 -915 28680 -795
rect 28725 -915 28845 -795
rect 28890 -915 29010 -795
rect 29065 -915 29185 -795
rect 29230 -915 29350 -795
rect 29395 -915 29515 -795
rect 29560 -915 29680 -795
rect 24200 -1080 24320 -960
rect 24375 -1080 24495 -960
rect 24540 -1080 24660 -960
rect 24705 -1080 24825 -960
rect 24870 -1080 24990 -960
rect 25045 -1080 25165 -960
rect 25210 -1080 25330 -960
rect 25375 -1080 25495 -960
rect 25540 -1080 25660 -960
rect 25715 -1080 25835 -960
rect 25880 -1080 26000 -960
rect 26045 -1080 26165 -960
rect 26210 -1080 26330 -960
rect 26385 -1080 26505 -960
rect 26550 -1080 26670 -960
rect 26715 -1080 26835 -960
rect 26880 -1080 27000 -960
rect 27055 -1080 27175 -960
rect 27220 -1080 27340 -960
rect 27385 -1080 27505 -960
rect 27550 -1080 27670 -960
rect 27725 -1080 27845 -960
rect 27890 -1080 28010 -960
rect 28055 -1080 28175 -960
rect 28220 -1080 28340 -960
rect 28395 -1080 28515 -960
rect 28560 -1080 28680 -960
rect 28725 -1080 28845 -960
rect 28890 -1080 29010 -960
rect 29065 -1080 29185 -960
rect 29230 -1080 29350 -960
rect 29395 -1080 29515 -960
rect 29560 -1080 29680 -960
rect 24200 -1245 24320 -1125
rect 24375 -1245 24495 -1125
rect 24540 -1245 24660 -1125
rect 24705 -1245 24825 -1125
rect 24870 -1245 24990 -1125
rect 25045 -1245 25165 -1125
rect 25210 -1245 25330 -1125
rect 25375 -1245 25495 -1125
rect 25540 -1245 25660 -1125
rect 25715 -1245 25835 -1125
rect 25880 -1245 26000 -1125
rect 26045 -1245 26165 -1125
rect 26210 -1245 26330 -1125
rect 26385 -1245 26505 -1125
rect 26550 -1245 26670 -1125
rect 26715 -1245 26835 -1125
rect 26880 -1245 27000 -1125
rect 27055 -1245 27175 -1125
rect 27220 -1245 27340 -1125
rect 27385 -1245 27505 -1125
rect 27550 -1245 27670 -1125
rect 27725 -1245 27845 -1125
rect 27890 -1245 28010 -1125
rect 28055 -1245 28175 -1125
rect 28220 -1245 28340 -1125
rect 28395 -1245 28515 -1125
rect 28560 -1245 28680 -1125
rect 28725 -1245 28845 -1125
rect 28890 -1245 29010 -1125
rect 29065 -1245 29185 -1125
rect 29230 -1245 29350 -1125
rect 29395 -1245 29515 -1125
rect 29560 -1245 29680 -1125
rect 24200 -1420 24320 -1300
rect 24375 -1420 24495 -1300
rect 24540 -1420 24660 -1300
rect 24705 -1420 24825 -1300
rect 24870 -1420 24990 -1300
rect 25045 -1420 25165 -1300
rect 25210 -1420 25330 -1300
rect 25375 -1420 25495 -1300
rect 25540 -1420 25660 -1300
rect 25715 -1420 25835 -1300
rect 25880 -1420 26000 -1300
rect 26045 -1420 26165 -1300
rect 26210 -1420 26330 -1300
rect 26385 -1420 26505 -1300
rect 26550 -1420 26670 -1300
rect 26715 -1420 26835 -1300
rect 26880 -1420 27000 -1300
rect 27055 -1420 27175 -1300
rect 27220 -1420 27340 -1300
rect 27385 -1420 27505 -1300
rect 27550 -1420 27670 -1300
rect 27725 -1420 27845 -1300
rect 27890 -1420 28010 -1300
rect 28055 -1420 28175 -1300
rect 28220 -1420 28340 -1300
rect 28395 -1420 28515 -1300
rect 28560 -1420 28680 -1300
rect 28725 -1420 28845 -1300
rect 28890 -1420 29010 -1300
rect 29065 -1420 29185 -1300
rect 29230 -1420 29350 -1300
rect 29395 -1420 29515 -1300
rect 29560 -1420 29680 -1300
rect 24200 -1585 24320 -1465
rect 24375 -1585 24495 -1465
rect 24540 -1585 24660 -1465
rect 24705 -1585 24825 -1465
rect 24870 -1585 24990 -1465
rect 25045 -1585 25165 -1465
rect 25210 -1585 25330 -1465
rect 25375 -1585 25495 -1465
rect 25540 -1585 25660 -1465
rect 25715 -1585 25835 -1465
rect 25880 -1585 26000 -1465
rect 26045 -1585 26165 -1465
rect 26210 -1585 26330 -1465
rect 26385 -1585 26505 -1465
rect 26550 -1585 26670 -1465
rect 26715 -1585 26835 -1465
rect 26880 -1585 27000 -1465
rect 27055 -1585 27175 -1465
rect 27220 -1585 27340 -1465
rect 27385 -1585 27505 -1465
rect 27550 -1585 27670 -1465
rect 27725 -1585 27845 -1465
rect 27890 -1585 28010 -1465
rect 28055 -1585 28175 -1465
rect 28220 -1585 28340 -1465
rect 28395 -1585 28515 -1465
rect 28560 -1585 28680 -1465
rect 28725 -1585 28845 -1465
rect 28890 -1585 29010 -1465
rect 29065 -1585 29185 -1465
rect 29230 -1585 29350 -1465
rect 29395 -1585 29515 -1465
rect 29560 -1585 29680 -1465
rect 24200 -1750 24320 -1630
rect 24375 -1750 24495 -1630
rect 24540 -1750 24660 -1630
rect 24705 -1750 24825 -1630
rect 24870 -1750 24990 -1630
rect 25045 -1750 25165 -1630
rect 25210 -1750 25330 -1630
rect 25375 -1750 25495 -1630
rect 25540 -1750 25660 -1630
rect 25715 -1750 25835 -1630
rect 25880 -1750 26000 -1630
rect 26045 -1750 26165 -1630
rect 26210 -1750 26330 -1630
rect 26385 -1750 26505 -1630
rect 26550 -1750 26670 -1630
rect 26715 -1750 26835 -1630
rect 26880 -1750 27000 -1630
rect 27055 -1750 27175 -1630
rect 27220 -1750 27340 -1630
rect 27385 -1750 27505 -1630
rect 27550 -1750 27670 -1630
rect 27725 -1750 27845 -1630
rect 27890 -1750 28010 -1630
rect 28055 -1750 28175 -1630
rect 28220 -1750 28340 -1630
rect 28395 -1750 28515 -1630
rect 28560 -1750 28680 -1630
rect 28725 -1750 28845 -1630
rect 28890 -1750 29010 -1630
rect 29065 -1750 29185 -1630
rect 29230 -1750 29350 -1630
rect 29395 -1750 29515 -1630
rect 29560 -1750 29680 -1630
rect 24200 -1915 24320 -1795
rect 24375 -1915 24495 -1795
rect 24540 -1915 24660 -1795
rect 24705 -1915 24825 -1795
rect 24870 -1915 24990 -1795
rect 25045 -1915 25165 -1795
rect 25210 -1915 25330 -1795
rect 25375 -1915 25495 -1795
rect 25540 -1915 25660 -1795
rect 25715 -1915 25835 -1795
rect 25880 -1915 26000 -1795
rect 26045 -1915 26165 -1795
rect 26210 -1915 26330 -1795
rect 26385 -1915 26505 -1795
rect 26550 -1915 26670 -1795
rect 26715 -1915 26835 -1795
rect 26880 -1915 27000 -1795
rect 27055 -1915 27175 -1795
rect 27220 -1915 27340 -1795
rect 27385 -1915 27505 -1795
rect 27550 -1915 27670 -1795
rect 27725 -1915 27845 -1795
rect 27890 -1915 28010 -1795
rect 28055 -1915 28175 -1795
rect 28220 -1915 28340 -1795
rect 28395 -1915 28515 -1795
rect 28560 -1915 28680 -1795
rect 28725 -1915 28845 -1795
rect 28890 -1915 29010 -1795
rect 29065 -1915 29185 -1795
rect 29230 -1915 29350 -1795
rect 29395 -1915 29515 -1795
rect 29560 -1915 29680 -1795
rect 24200 -2090 24320 -1970
rect 24375 -2090 24495 -1970
rect 24540 -2090 24660 -1970
rect 24705 -2090 24825 -1970
rect 24870 -2090 24990 -1970
rect 25045 -2090 25165 -1970
rect 25210 -2090 25330 -1970
rect 25375 -2090 25495 -1970
rect 25540 -2090 25660 -1970
rect 25715 -2090 25835 -1970
rect 25880 -2090 26000 -1970
rect 26045 -2090 26165 -1970
rect 26210 -2090 26330 -1970
rect 26385 -2090 26505 -1970
rect 26550 -2090 26670 -1970
rect 26715 -2090 26835 -1970
rect 26880 -2090 27000 -1970
rect 27055 -2090 27175 -1970
rect 27220 -2090 27340 -1970
rect 27385 -2090 27505 -1970
rect 27550 -2090 27670 -1970
rect 27725 -2090 27845 -1970
rect 27890 -2090 28010 -1970
rect 28055 -2090 28175 -1970
rect 28220 -2090 28340 -1970
rect 28395 -2090 28515 -1970
rect 28560 -2090 28680 -1970
rect 28725 -2090 28845 -1970
rect 28890 -2090 29010 -1970
rect 29065 -2090 29185 -1970
rect 29230 -2090 29350 -1970
rect 29395 -2090 29515 -1970
rect 29560 -2090 29680 -1970
rect 24200 -2255 24320 -2135
rect 24375 -2255 24495 -2135
rect 24540 -2255 24660 -2135
rect 24705 -2255 24825 -2135
rect 24870 -2255 24990 -2135
rect 25045 -2255 25165 -2135
rect 25210 -2255 25330 -2135
rect 25375 -2255 25495 -2135
rect 25540 -2255 25660 -2135
rect 25715 -2255 25835 -2135
rect 25880 -2255 26000 -2135
rect 26045 -2255 26165 -2135
rect 26210 -2255 26330 -2135
rect 26385 -2255 26505 -2135
rect 26550 -2255 26670 -2135
rect 26715 -2255 26835 -2135
rect 26880 -2255 27000 -2135
rect 27055 -2255 27175 -2135
rect 27220 -2255 27340 -2135
rect 27385 -2255 27505 -2135
rect 27550 -2255 27670 -2135
rect 27725 -2255 27845 -2135
rect 27890 -2255 28010 -2135
rect 28055 -2255 28175 -2135
rect 28220 -2255 28340 -2135
rect 28395 -2255 28515 -2135
rect 28560 -2255 28680 -2135
rect 28725 -2255 28845 -2135
rect 28890 -2255 29010 -2135
rect 29065 -2255 29185 -2135
rect 29230 -2255 29350 -2135
rect 29395 -2255 29515 -2135
rect 29560 -2255 29680 -2135
rect 24200 -2420 24320 -2300
rect 24375 -2420 24495 -2300
rect 24540 -2420 24660 -2300
rect 24705 -2420 24825 -2300
rect 24870 -2420 24990 -2300
rect 25045 -2420 25165 -2300
rect 25210 -2420 25330 -2300
rect 25375 -2420 25495 -2300
rect 25540 -2420 25660 -2300
rect 25715 -2420 25835 -2300
rect 25880 -2420 26000 -2300
rect 26045 -2420 26165 -2300
rect 26210 -2420 26330 -2300
rect 26385 -2420 26505 -2300
rect 26550 -2420 26670 -2300
rect 26715 -2420 26835 -2300
rect 26880 -2420 27000 -2300
rect 27055 -2420 27175 -2300
rect 27220 -2420 27340 -2300
rect 27385 -2420 27505 -2300
rect 27550 -2420 27670 -2300
rect 27725 -2420 27845 -2300
rect 27890 -2420 28010 -2300
rect 28055 -2420 28175 -2300
rect 28220 -2420 28340 -2300
rect 28395 -2420 28515 -2300
rect 28560 -2420 28680 -2300
rect 28725 -2420 28845 -2300
rect 28890 -2420 29010 -2300
rect 29065 -2420 29185 -2300
rect 29230 -2420 29350 -2300
rect 29395 -2420 29515 -2300
rect 29560 -2420 29680 -2300
rect 24200 -2585 24320 -2465
rect 24375 -2585 24495 -2465
rect 24540 -2585 24660 -2465
rect 24705 -2585 24825 -2465
rect 24870 -2585 24990 -2465
rect 25045 -2585 25165 -2465
rect 25210 -2585 25330 -2465
rect 25375 -2585 25495 -2465
rect 25540 -2585 25660 -2465
rect 25715 -2585 25835 -2465
rect 25880 -2585 26000 -2465
rect 26045 -2585 26165 -2465
rect 26210 -2585 26330 -2465
rect 26385 -2585 26505 -2465
rect 26550 -2585 26670 -2465
rect 26715 -2585 26835 -2465
rect 26880 -2585 27000 -2465
rect 27055 -2585 27175 -2465
rect 27220 -2585 27340 -2465
rect 27385 -2585 27505 -2465
rect 27550 -2585 27670 -2465
rect 27725 -2585 27845 -2465
rect 27890 -2585 28010 -2465
rect 28055 -2585 28175 -2465
rect 28220 -2585 28340 -2465
rect 28395 -2585 28515 -2465
rect 28560 -2585 28680 -2465
rect 28725 -2585 28845 -2465
rect 28890 -2585 29010 -2465
rect 29065 -2585 29185 -2465
rect 29230 -2585 29350 -2465
rect 29395 -2585 29515 -2465
rect 29560 -2585 29680 -2465
rect 24200 -2760 24320 -2640
rect 24375 -2760 24495 -2640
rect 24540 -2760 24660 -2640
rect 24705 -2760 24825 -2640
rect 24870 -2760 24990 -2640
rect 25045 -2760 25165 -2640
rect 25210 -2760 25330 -2640
rect 25375 -2760 25495 -2640
rect 25540 -2760 25660 -2640
rect 25715 -2760 25835 -2640
rect 25880 -2760 26000 -2640
rect 26045 -2760 26165 -2640
rect 26210 -2760 26330 -2640
rect 26385 -2760 26505 -2640
rect 26550 -2760 26670 -2640
rect 26715 -2760 26835 -2640
rect 26880 -2760 27000 -2640
rect 27055 -2760 27175 -2640
rect 27220 -2760 27340 -2640
rect 27385 -2760 27505 -2640
rect 27550 -2760 27670 -2640
rect 27725 -2760 27845 -2640
rect 27890 -2760 28010 -2640
rect 28055 -2760 28175 -2640
rect 28220 -2760 28340 -2640
rect 28395 -2760 28515 -2640
rect 28560 -2760 28680 -2640
rect 28725 -2760 28845 -2640
rect 28890 -2760 29010 -2640
rect 29065 -2760 29185 -2640
rect 29230 -2760 29350 -2640
rect 29395 -2760 29515 -2640
rect 29560 -2760 29680 -2640
rect 24200 -2925 24320 -2805
rect 24375 -2925 24495 -2805
rect 24540 -2925 24660 -2805
rect 24705 -2925 24825 -2805
rect 24870 -2925 24990 -2805
rect 25045 -2925 25165 -2805
rect 25210 -2925 25330 -2805
rect 25375 -2925 25495 -2805
rect 25540 -2925 25660 -2805
rect 25715 -2925 25835 -2805
rect 25880 -2925 26000 -2805
rect 26045 -2925 26165 -2805
rect 26210 -2925 26330 -2805
rect 26385 -2925 26505 -2805
rect 26550 -2925 26670 -2805
rect 26715 -2925 26835 -2805
rect 26880 -2925 27000 -2805
rect 27055 -2925 27175 -2805
rect 27220 -2925 27340 -2805
rect 27385 -2925 27505 -2805
rect 27550 -2925 27670 -2805
rect 27725 -2925 27845 -2805
rect 27890 -2925 28010 -2805
rect 28055 -2925 28175 -2805
rect 28220 -2925 28340 -2805
rect 28395 -2925 28515 -2805
rect 28560 -2925 28680 -2805
rect 28725 -2925 28845 -2805
rect 28890 -2925 29010 -2805
rect 29065 -2925 29185 -2805
rect 29230 -2925 29350 -2805
rect 29395 -2925 29515 -2805
rect 29560 -2925 29680 -2805
rect 24200 -3090 24320 -2970
rect 24375 -3090 24495 -2970
rect 24540 -3090 24660 -2970
rect 24705 -3090 24825 -2970
rect 24870 -3090 24990 -2970
rect 25045 -3090 25165 -2970
rect 25210 -3090 25330 -2970
rect 25375 -3090 25495 -2970
rect 25540 -3090 25660 -2970
rect 25715 -3090 25835 -2970
rect 25880 -3090 26000 -2970
rect 26045 -3090 26165 -2970
rect 26210 -3090 26330 -2970
rect 26385 -3090 26505 -2970
rect 26550 -3090 26670 -2970
rect 26715 -3090 26835 -2970
rect 26880 -3090 27000 -2970
rect 27055 -3090 27175 -2970
rect 27220 -3090 27340 -2970
rect 27385 -3090 27505 -2970
rect 27550 -3090 27670 -2970
rect 27725 -3090 27845 -2970
rect 27890 -3090 28010 -2970
rect 28055 -3090 28175 -2970
rect 28220 -3090 28340 -2970
rect 28395 -3090 28515 -2970
rect 28560 -3090 28680 -2970
rect 28725 -3090 28845 -2970
rect 28890 -3090 29010 -2970
rect 29065 -3090 29185 -2970
rect 29230 -3090 29350 -2970
rect 29395 -3090 29515 -2970
rect 29560 -3090 29680 -2970
rect 24200 -3255 24320 -3135
rect 24375 -3255 24495 -3135
rect 24540 -3255 24660 -3135
rect 24705 -3255 24825 -3135
rect 24870 -3255 24990 -3135
rect 25045 -3255 25165 -3135
rect 25210 -3255 25330 -3135
rect 25375 -3255 25495 -3135
rect 25540 -3255 25660 -3135
rect 25715 -3255 25835 -3135
rect 25880 -3255 26000 -3135
rect 26045 -3255 26165 -3135
rect 26210 -3255 26330 -3135
rect 26385 -3255 26505 -3135
rect 26550 -3255 26670 -3135
rect 26715 -3255 26835 -3135
rect 26880 -3255 27000 -3135
rect 27055 -3255 27175 -3135
rect 27220 -3255 27340 -3135
rect 27385 -3255 27505 -3135
rect 27550 -3255 27670 -3135
rect 27725 -3255 27845 -3135
rect 27890 -3255 28010 -3135
rect 28055 -3255 28175 -3135
rect 28220 -3255 28340 -3135
rect 28395 -3255 28515 -3135
rect 28560 -3255 28680 -3135
rect 28725 -3255 28845 -3135
rect 28890 -3255 29010 -3135
rect 29065 -3255 29185 -3135
rect 29230 -3255 29350 -3135
rect 29395 -3255 29515 -3135
rect 29560 -3255 29680 -3135
rect 24200 -3430 24320 -3310
rect 24375 -3430 24495 -3310
rect 24540 -3430 24660 -3310
rect 24705 -3430 24825 -3310
rect 24870 -3430 24990 -3310
rect 25045 -3430 25165 -3310
rect 25210 -3430 25330 -3310
rect 25375 -3430 25495 -3310
rect 25540 -3430 25660 -3310
rect 25715 -3430 25835 -3310
rect 25880 -3430 26000 -3310
rect 26045 -3430 26165 -3310
rect 26210 -3430 26330 -3310
rect 26385 -3430 26505 -3310
rect 26550 -3430 26670 -3310
rect 26715 -3430 26835 -3310
rect 26880 -3430 27000 -3310
rect 27055 -3430 27175 -3310
rect 27220 -3430 27340 -3310
rect 27385 -3430 27505 -3310
rect 27550 -3430 27670 -3310
rect 27725 -3430 27845 -3310
rect 27890 -3430 28010 -3310
rect 28055 -3430 28175 -3310
rect 28220 -3430 28340 -3310
rect 28395 -3430 28515 -3310
rect 28560 -3430 28680 -3310
rect 28725 -3430 28845 -3310
rect 28890 -3430 29010 -3310
rect 29065 -3430 29185 -3310
rect 29230 -3430 29350 -3310
rect 29395 -3430 29515 -3310
rect 29560 -3430 29680 -3310
rect 24200 -3595 24320 -3475
rect 24375 -3595 24495 -3475
rect 24540 -3595 24660 -3475
rect 24705 -3595 24825 -3475
rect 24870 -3595 24990 -3475
rect 25045 -3595 25165 -3475
rect 25210 -3595 25330 -3475
rect 25375 -3595 25495 -3475
rect 25540 -3595 25660 -3475
rect 25715 -3595 25835 -3475
rect 25880 -3595 26000 -3475
rect 26045 -3595 26165 -3475
rect 26210 -3595 26330 -3475
rect 26385 -3595 26505 -3475
rect 26550 -3595 26670 -3475
rect 26715 -3595 26835 -3475
rect 26880 -3595 27000 -3475
rect 27055 -3595 27175 -3475
rect 27220 -3595 27340 -3475
rect 27385 -3595 27505 -3475
rect 27550 -3595 27670 -3475
rect 27725 -3595 27845 -3475
rect 27890 -3595 28010 -3475
rect 28055 -3595 28175 -3475
rect 28220 -3595 28340 -3475
rect 28395 -3595 28515 -3475
rect 28560 -3595 28680 -3475
rect 28725 -3595 28845 -3475
rect 28890 -3595 29010 -3475
rect 29065 -3595 29185 -3475
rect 29230 -3595 29350 -3475
rect 29395 -3595 29515 -3475
rect 29560 -3595 29680 -3475
rect 24200 -3760 24320 -3640
rect 24375 -3760 24495 -3640
rect 24540 -3760 24660 -3640
rect 24705 -3760 24825 -3640
rect 24870 -3760 24990 -3640
rect 25045 -3760 25165 -3640
rect 25210 -3760 25330 -3640
rect 25375 -3760 25495 -3640
rect 25540 -3760 25660 -3640
rect 25715 -3760 25835 -3640
rect 25880 -3760 26000 -3640
rect 26045 -3760 26165 -3640
rect 26210 -3760 26330 -3640
rect 26385 -3760 26505 -3640
rect 26550 -3760 26670 -3640
rect 26715 -3760 26835 -3640
rect 26880 -3760 27000 -3640
rect 27055 -3760 27175 -3640
rect 27220 -3760 27340 -3640
rect 27385 -3760 27505 -3640
rect 27550 -3760 27670 -3640
rect 27725 -3760 27845 -3640
rect 27890 -3760 28010 -3640
rect 28055 -3760 28175 -3640
rect 28220 -3760 28340 -3640
rect 28395 -3760 28515 -3640
rect 28560 -3760 28680 -3640
rect 28725 -3760 28845 -3640
rect 28890 -3760 29010 -3640
rect 29065 -3760 29185 -3640
rect 29230 -3760 29350 -3640
rect 29395 -3760 29515 -3640
rect 29560 -3760 29680 -3640
rect 24200 -3925 24320 -3805
rect 24375 -3925 24495 -3805
rect 24540 -3925 24660 -3805
rect 24705 -3925 24825 -3805
rect 24870 -3925 24990 -3805
rect 25045 -3925 25165 -3805
rect 25210 -3925 25330 -3805
rect 25375 -3925 25495 -3805
rect 25540 -3925 25660 -3805
rect 25715 -3925 25835 -3805
rect 25880 -3925 26000 -3805
rect 26045 -3925 26165 -3805
rect 26210 -3925 26330 -3805
rect 26385 -3925 26505 -3805
rect 26550 -3925 26670 -3805
rect 26715 -3925 26835 -3805
rect 26880 -3925 27000 -3805
rect 27055 -3925 27175 -3805
rect 27220 -3925 27340 -3805
rect 27385 -3925 27505 -3805
rect 27550 -3925 27670 -3805
rect 27725 -3925 27845 -3805
rect 27890 -3925 28010 -3805
rect 28055 -3925 28175 -3805
rect 28220 -3925 28340 -3805
rect 28395 -3925 28515 -3805
rect 28560 -3925 28680 -3805
rect 28725 -3925 28845 -3805
rect 28890 -3925 29010 -3805
rect 29065 -3925 29185 -3805
rect 29230 -3925 29350 -3805
rect 29395 -3925 29515 -3805
rect 29560 -3925 29680 -3805
rect 24200 -4100 24320 -3980
rect 24375 -4100 24495 -3980
rect 24540 -4100 24660 -3980
rect 24705 -4100 24825 -3980
rect 24870 -4100 24990 -3980
rect 25045 -4100 25165 -3980
rect 25210 -4100 25330 -3980
rect 25375 -4100 25495 -3980
rect 25540 -4100 25660 -3980
rect 25715 -4100 25835 -3980
rect 25880 -4100 26000 -3980
rect 26045 -4100 26165 -3980
rect 26210 -4100 26330 -3980
rect 26385 -4100 26505 -3980
rect 26550 -4100 26670 -3980
rect 26715 -4100 26835 -3980
rect 26880 -4100 27000 -3980
rect 27055 -4100 27175 -3980
rect 27220 -4100 27340 -3980
rect 27385 -4100 27505 -3980
rect 27550 -4100 27670 -3980
rect 27725 -4100 27845 -3980
rect 27890 -4100 28010 -3980
rect 28055 -4100 28175 -3980
rect 28220 -4100 28340 -3980
rect 28395 -4100 28515 -3980
rect 28560 -4100 28680 -3980
rect 28725 -4100 28845 -3980
rect 28890 -4100 29010 -3980
rect 29065 -4100 29185 -3980
rect 29230 -4100 29350 -3980
rect 29395 -4100 29515 -3980
rect 29560 -4100 29680 -3980
rect 7130 -4430 7250 -4310
rect 7295 -4430 7415 -4310
rect 7460 -4430 7580 -4310
rect 7625 -4430 7745 -4310
rect 7800 -4430 7920 -4310
rect 7965 -4430 8085 -4310
rect 8130 -4430 8250 -4310
rect 8295 -4430 8415 -4310
rect 8470 -4430 8590 -4310
rect 8635 -4430 8755 -4310
rect 8800 -4430 8920 -4310
rect 8965 -4430 9085 -4310
rect 9140 -4430 9260 -4310
rect 9305 -4430 9425 -4310
rect 9470 -4430 9590 -4310
rect 9635 -4430 9755 -4310
rect 9810 -4430 9930 -4310
rect 9975 -4430 10095 -4310
rect 10140 -4430 10260 -4310
rect 10305 -4430 10425 -4310
rect 10480 -4430 10600 -4310
rect 10645 -4430 10765 -4310
rect 10810 -4430 10930 -4310
rect 10975 -4430 11095 -4310
rect 11150 -4430 11270 -4310
rect 11315 -4430 11435 -4310
rect 11480 -4430 11600 -4310
rect 11645 -4430 11765 -4310
rect 11820 -4430 11940 -4310
rect 11985 -4430 12105 -4310
rect 12150 -4430 12270 -4310
rect 12315 -4430 12435 -4310
rect 12490 -4430 12610 -4310
rect 7130 -4605 7250 -4485
rect 7295 -4605 7415 -4485
rect 7460 -4605 7580 -4485
rect 7625 -4605 7745 -4485
rect 7800 -4605 7920 -4485
rect 7965 -4605 8085 -4485
rect 8130 -4605 8250 -4485
rect 8295 -4605 8415 -4485
rect 8470 -4605 8590 -4485
rect 8635 -4605 8755 -4485
rect 8800 -4605 8920 -4485
rect 8965 -4605 9085 -4485
rect 9140 -4605 9260 -4485
rect 9305 -4605 9425 -4485
rect 9470 -4605 9590 -4485
rect 9635 -4605 9755 -4485
rect 9810 -4605 9930 -4485
rect 9975 -4605 10095 -4485
rect 10140 -4605 10260 -4485
rect 10305 -4605 10425 -4485
rect 10480 -4605 10600 -4485
rect 10645 -4605 10765 -4485
rect 10810 -4605 10930 -4485
rect 10975 -4605 11095 -4485
rect 11150 -4605 11270 -4485
rect 11315 -4605 11435 -4485
rect 11480 -4605 11600 -4485
rect 11645 -4605 11765 -4485
rect 11820 -4605 11940 -4485
rect 11985 -4605 12105 -4485
rect 12150 -4605 12270 -4485
rect 12315 -4605 12435 -4485
rect 12490 -4605 12610 -4485
rect 7130 -4770 7250 -4650
rect 7295 -4770 7415 -4650
rect 7460 -4770 7580 -4650
rect 7625 -4770 7745 -4650
rect 7800 -4770 7920 -4650
rect 7965 -4770 8085 -4650
rect 8130 -4770 8250 -4650
rect 8295 -4770 8415 -4650
rect 8470 -4770 8590 -4650
rect 8635 -4770 8755 -4650
rect 8800 -4770 8920 -4650
rect 8965 -4770 9085 -4650
rect 9140 -4770 9260 -4650
rect 9305 -4770 9425 -4650
rect 9470 -4770 9590 -4650
rect 9635 -4770 9755 -4650
rect 9810 -4770 9930 -4650
rect 9975 -4770 10095 -4650
rect 10140 -4770 10260 -4650
rect 10305 -4770 10425 -4650
rect 10480 -4770 10600 -4650
rect 10645 -4770 10765 -4650
rect 10810 -4770 10930 -4650
rect 10975 -4770 11095 -4650
rect 11150 -4770 11270 -4650
rect 11315 -4770 11435 -4650
rect 11480 -4770 11600 -4650
rect 11645 -4770 11765 -4650
rect 11820 -4770 11940 -4650
rect 11985 -4770 12105 -4650
rect 12150 -4770 12270 -4650
rect 12315 -4770 12435 -4650
rect 12490 -4770 12610 -4650
rect 7130 -4935 7250 -4815
rect 7295 -4935 7415 -4815
rect 7460 -4935 7580 -4815
rect 7625 -4935 7745 -4815
rect 7800 -4935 7920 -4815
rect 7965 -4935 8085 -4815
rect 8130 -4935 8250 -4815
rect 8295 -4935 8415 -4815
rect 8470 -4935 8590 -4815
rect 8635 -4935 8755 -4815
rect 8800 -4935 8920 -4815
rect 8965 -4935 9085 -4815
rect 9140 -4935 9260 -4815
rect 9305 -4935 9425 -4815
rect 9470 -4935 9590 -4815
rect 9635 -4935 9755 -4815
rect 9810 -4935 9930 -4815
rect 9975 -4935 10095 -4815
rect 10140 -4935 10260 -4815
rect 10305 -4935 10425 -4815
rect 10480 -4935 10600 -4815
rect 10645 -4935 10765 -4815
rect 10810 -4935 10930 -4815
rect 10975 -4935 11095 -4815
rect 11150 -4935 11270 -4815
rect 11315 -4935 11435 -4815
rect 11480 -4935 11600 -4815
rect 11645 -4935 11765 -4815
rect 11820 -4935 11940 -4815
rect 11985 -4935 12105 -4815
rect 12150 -4935 12270 -4815
rect 12315 -4935 12435 -4815
rect 12490 -4935 12610 -4815
rect 7130 -5100 7250 -4980
rect 7295 -5100 7415 -4980
rect 7460 -5100 7580 -4980
rect 7625 -5100 7745 -4980
rect 7800 -5100 7920 -4980
rect 7965 -5100 8085 -4980
rect 8130 -5100 8250 -4980
rect 8295 -5100 8415 -4980
rect 8470 -5100 8590 -4980
rect 8635 -5100 8755 -4980
rect 8800 -5100 8920 -4980
rect 8965 -5100 9085 -4980
rect 9140 -5100 9260 -4980
rect 9305 -5100 9425 -4980
rect 9470 -5100 9590 -4980
rect 9635 -5100 9755 -4980
rect 9810 -5100 9930 -4980
rect 9975 -5100 10095 -4980
rect 10140 -5100 10260 -4980
rect 10305 -5100 10425 -4980
rect 10480 -5100 10600 -4980
rect 10645 -5100 10765 -4980
rect 10810 -5100 10930 -4980
rect 10975 -5100 11095 -4980
rect 11150 -5100 11270 -4980
rect 11315 -5100 11435 -4980
rect 11480 -5100 11600 -4980
rect 11645 -5100 11765 -4980
rect 11820 -5100 11940 -4980
rect 11985 -5100 12105 -4980
rect 12150 -5100 12270 -4980
rect 12315 -5100 12435 -4980
rect 12490 -5100 12610 -4980
rect 7130 -5275 7250 -5155
rect 7295 -5275 7415 -5155
rect 7460 -5275 7580 -5155
rect 7625 -5275 7745 -5155
rect 7800 -5275 7920 -5155
rect 7965 -5275 8085 -5155
rect 8130 -5275 8250 -5155
rect 8295 -5275 8415 -5155
rect 8470 -5275 8590 -5155
rect 8635 -5275 8755 -5155
rect 8800 -5275 8920 -5155
rect 8965 -5275 9085 -5155
rect 9140 -5275 9260 -5155
rect 9305 -5275 9425 -5155
rect 9470 -5275 9590 -5155
rect 9635 -5275 9755 -5155
rect 9810 -5275 9930 -5155
rect 9975 -5275 10095 -5155
rect 10140 -5275 10260 -5155
rect 10305 -5275 10425 -5155
rect 10480 -5275 10600 -5155
rect 10645 -5275 10765 -5155
rect 10810 -5275 10930 -5155
rect 10975 -5275 11095 -5155
rect 11150 -5275 11270 -5155
rect 11315 -5275 11435 -5155
rect 11480 -5275 11600 -5155
rect 11645 -5275 11765 -5155
rect 11820 -5275 11940 -5155
rect 11985 -5275 12105 -5155
rect 12150 -5275 12270 -5155
rect 12315 -5275 12435 -5155
rect 12490 -5275 12610 -5155
rect 7130 -5440 7250 -5320
rect 7295 -5440 7415 -5320
rect 7460 -5440 7580 -5320
rect 7625 -5440 7745 -5320
rect 7800 -5440 7920 -5320
rect 7965 -5440 8085 -5320
rect 8130 -5440 8250 -5320
rect 8295 -5440 8415 -5320
rect 8470 -5440 8590 -5320
rect 8635 -5440 8755 -5320
rect 8800 -5440 8920 -5320
rect 8965 -5440 9085 -5320
rect 9140 -5440 9260 -5320
rect 9305 -5440 9425 -5320
rect 9470 -5440 9590 -5320
rect 9635 -5440 9755 -5320
rect 9810 -5440 9930 -5320
rect 9975 -5440 10095 -5320
rect 10140 -5440 10260 -5320
rect 10305 -5440 10425 -5320
rect 10480 -5440 10600 -5320
rect 10645 -5440 10765 -5320
rect 10810 -5440 10930 -5320
rect 10975 -5440 11095 -5320
rect 11150 -5440 11270 -5320
rect 11315 -5440 11435 -5320
rect 11480 -5440 11600 -5320
rect 11645 -5440 11765 -5320
rect 11820 -5440 11940 -5320
rect 11985 -5440 12105 -5320
rect 12150 -5440 12270 -5320
rect 12315 -5440 12435 -5320
rect 12490 -5440 12610 -5320
rect 7130 -5605 7250 -5485
rect 7295 -5605 7415 -5485
rect 7460 -5605 7580 -5485
rect 7625 -5605 7745 -5485
rect 7800 -5605 7920 -5485
rect 7965 -5605 8085 -5485
rect 8130 -5605 8250 -5485
rect 8295 -5605 8415 -5485
rect 8470 -5605 8590 -5485
rect 8635 -5605 8755 -5485
rect 8800 -5605 8920 -5485
rect 8965 -5605 9085 -5485
rect 9140 -5605 9260 -5485
rect 9305 -5605 9425 -5485
rect 9470 -5605 9590 -5485
rect 9635 -5605 9755 -5485
rect 9810 -5605 9930 -5485
rect 9975 -5605 10095 -5485
rect 10140 -5605 10260 -5485
rect 10305 -5605 10425 -5485
rect 10480 -5605 10600 -5485
rect 10645 -5605 10765 -5485
rect 10810 -5605 10930 -5485
rect 10975 -5605 11095 -5485
rect 11150 -5605 11270 -5485
rect 11315 -5605 11435 -5485
rect 11480 -5605 11600 -5485
rect 11645 -5605 11765 -5485
rect 11820 -5605 11940 -5485
rect 11985 -5605 12105 -5485
rect 12150 -5605 12270 -5485
rect 12315 -5605 12435 -5485
rect 12490 -5605 12610 -5485
rect 7130 -5770 7250 -5650
rect 7295 -5770 7415 -5650
rect 7460 -5770 7580 -5650
rect 7625 -5770 7745 -5650
rect 7800 -5770 7920 -5650
rect 7965 -5770 8085 -5650
rect 8130 -5770 8250 -5650
rect 8295 -5770 8415 -5650
rect 8470 -5770 8590 -5650
rect 8635 -5770 8755 -5650
rect 8800 -5770 8920 -5650
rect 8965 -5770 9085 -5650
rect 9140 -5770 9260 -5650
rect 9305 -5770 9425 -5650
rect 9470 -5770 9590 -5650
rect 9635 -5770 9755 -5650
rect 9810 -5770 9930 -5650
rect 9975 -5770 10095 -5650
rect 10140 -5770 10260 -5650
rect 10305 -5770 10425 -5650
rect 10480 -5770 10600 -5650
rect 10645 -5770 10765 -5650
rect 10810 -5770 10930 -5650
rect 10975 -5770 11095 -5650
rect 11150 -5770 11270 -5650
rect 11315 -5770 11435 -5650
rect 11480 -5770 11600 -5650
rect 11645 -5770 11765 -5650
rect 11820 -5770 11940 -5650
rect 11985 -5770 12105 -5650
rect 12150 -5770 12270 -5650
rect 12315 -5770 12435 -5650
rect 12490 -5770 12610 -5650
rect 7130 -5945 7250 -5825
rect 7295 -5945 7415 -5825
rect 7460 -5945 7580 -5825
rect 7625 -5945 7745 -5825
rect 7800 -5945 7920 -5825
rect 7965 -5945 8085 -5825
rect 8130 -5945 8250 -5825
rect 8295 -5945 8415 -5825
rect 8470 -5945 8590 -5825
rect 8635 -5945 8755 -5825
rect 8800 -5945 8920 -5825
rect 8965 -5945 9085 -5825
rect 9140 -5945 9260 -5825
rect 9305 -5945 9425 -5825
rect 9470 -5945 9590 -5825
rect 9635 -5945 9755 -5825
rect 9810 -5945 9930 -5825
rect 9975 -5945 10095 -5825
rect 10140 -5945 10260 -5825
rect 10305 -5945 10425 -5825
rect 10480 -5945 10600 -5825
rect 10645 -5945 10765 -5825
rect 10810 -5945 10930 -5825
rect 10975 -5945 11095 -5825
rect 11150 -5945 11270 -5825
rect 11315 -5945 11435 -5825
rect 11480 -5945 11600 -5825
rect 11645 -5945 11765 -5825
rect 11820 -5945 11940 -5825
rect 11985 -5945 12105 -5825
rect 12150 -5945 12270 -5825
rect 12315 -5945 12435 -5825
rect 12490 -5945 12610 -5825
rect 7130 -6110 7250 -5990
rect 7295 -6110 7415 -5990
rect 7460 -6110 7580 -5990
rect 7625 -6110 7745 -5990
rect 7800 -6110 7920 -5990
rect 7965 -6110 8085 -5990
rect 8130 -6110 8250 -5990
rect 8295 -6110 8415 -5990
rect 8470 -6110 8590 -5990
rect 8635 -6110 8755 -5990
rect 8800 -6110 8920 -5990
rect 8965 -6110 9085 -5990
rect 9140 -6110 9260 -5990
rect 9305 -6110 9425 -5990
rect 9470 -6110 9590 -5990
rect 9635 -6110 9755 -5990
rect 9810 -6110 9930 -5990
rect 9975 -6110 10095 -5990
rect 10140 -6110 10260 -5990
rect 10305 -6110 10425 -5990
rect 10480 -6110 10600 -5990
rect 10645 -6110 10765 -5990
rect 10810 -6110 10930 -5990
rect 10975 -6110 11095 -5990
rect 11150 -6110 11270 -5990
rect 11315 -6110 11435 -5990
rect 11480 -6110 11600 -5990
rect 11645 -6110 11765 -5990
rect 11820 -6110 11940 -5990
rect 11985 -6110 12105 -5990
rect 12150 -6110 12270 -5990
rect 12315 -6110 12435 -5990
rect 12490 -6110 12610 -5990
rect 7130 -6275 7250 -6155
rect 7295 -6275 7415 -6155
rect 7460 -6275 7580 -6155
rect 7625 -6275 7745 -6155
rect 7800 -6275 7920 -6155
rect 7965 -6275 8085 -6155
rect 8130 -6275 8250 -6155
rect 8295 -6275 8415 -6155
rect 8470 -6275 8590 -6155
rect 8635 -6275 8755 -6155
rect 8800 -6275 8920 -6155
rect 8965 -6275 9085 -6155
rect 9140 -6275 9260 -6155
rect 9305 -6275 9425 -6155
rect 9470 -6275 9590 -6155
rect 9635 -6275 9755 -6155
rect 9810 -6275 9930 -6155
rect 9975 -6275 10095 -6155
rect 10140 -6275 10260 -6155
rect 10305 -6275 10425 -6155
rect 10480 -6275 10600 -6155
rect 10645 -6275 10765 -6155
rect 10810 -6275 10930 -6155
rect 10975 -6275 11095 -6155
rect 11150 -6275 11270 -6155
rect 11315 -6275 11435 -6155
rect 11480 -6275 11600 -6155
rect 11645 -6275 11765 -6155
rect 11820 -6275 11940 -6155
rect 11985 -6275 12105 -6155
rect 12150 -6275 12270 -6155
rect 12315 -6275 12435 -6155
rect 12490 -6275 12610 -6155
rect 7130 -6440 7250 -6320
rect 7295 -6440 7415 -6320
rect 7460 -6440 7580 -6320
rect 7625 -6440 7745 -6320
rect 7800 -6440 7920 -6320
rect 7965 -6440 8085 -6320
rect 8130 -6440 8250 -6320
rect 8295 -6440 8415 -6320
rect 8470 -6440 8590 -6320
rect 8635 -6440 8755 -6320
rect 8800 -6440 8920 -6320
rect 8965 -6440 9085 -6320
rect 9140 -6440 9260 -6320
rect 9305 -6440 9425 -6320
rect 9470 -6440 9590 -6320
rect 9635 -6440 9755 -6320
rect 9810 -6440 9930 -6320
rect 9975 -6440 10095 -6320
rect 10140 -6440 10260 -6320
rect 10305 -6440 10425 -6320
rect 10480 -6440 10600 -6320
rect 10645 -6440 10765 -6320
rect 10810 -6440 10930 -6320
rect 10975 -6440 11095 -6320
rect 11150 -6440 11270 -6320
rect 11315 -6440 11435 -6320
rect 11480 -6440 11600 -6320
rect 11645 -6440 11765 -6320
rect 11820 -6440 11940 -6320
rect 11985 -6440 12105 -6320
rect 12150 -6440 12270 -6320
rect 12315 -6440 12435 -6320
rect 12490 -6440 12610 -6320
rect 7130 -6615 7250 -6495
rect 7295 -6615 7415 -6495
rect 7460 -6615 7580 -6495
rect 7625 -6615 7745 -6495
rect 7800 -6615 7920 -6495
rect 7965 -6615 8085 -6495
rect 8130 -6615 8250 -6495
rect 8295 -6615 8415 -6495
rect 8470 -6615 8590 -6495
rect 8635 -6615 8755 -6495
rect 8800 -6615 8920 -6495
rect 8965 -6615 9085 -6495
rect 9140 -6615 9260 -6495
rect 9305 -6615 9425 -6495
rect 9470 -6615 9590 -6495
rect 9635 -6615 9755 -6495
rect 9810 -6615 9930 -6495
rect 9975 -6615 10095 -6495
rect 10140 -6615 10260 -6495
rect 10305 -6615 10425 -6495
rect 10480 -6615 10600 -6495
rect 10645 -6615 10765 -6495
rect 10810 -6615 10930 -6495
rect 10975 -6615 11095 -6495
rect 11150 -6615 11270 -6495
rect 11315 -6615 11435 -6495
rect 11480 -6615 11600 -6495
rect 11645 -6615 11765 -6495
rect 11820 -6615 11940 -6495
rect 11985 -6615 12105 -6495
rect 12150 -6615 12270 -6495
rect 12315 -6615 12435 -6495
rect 12490 -6615 12610 -6495
rect 7130 -6780 7250 -6660
rect 7295 -6780 7415 -6660
rect 7460 -6780 7580 -6660
rect 7625 -6780 7745 -6660
rect 7800 -6780 7920 -6660
rect 7965 -6780 8085 -6660
rect 8130 -6780 8250 -6660
rect 8295 -6780 8415 -6660
rect 8470 -6780 8590 -6660
rect 8635 -6780 8755 -6660
rect 8800 -6780 8920 -6660
rect 8965 -6780 9085 -6660
rect 9140 -6780 9260 -6660
rect 9305 -6780 9425 -6660
rect 9470 -6780 9590 -6660
rect 9635 -6780 9755 -6660
rect 9810 -6780 9930 -6660
rect 9975 -6780 10095 -6660
rect 10140 -6780 10260 -6660
rect 10305 -6780 10425 -6660
rect 10480 -6780 10600 -6660
rect 10645 -6780 10765 -6660
rect 10810 -6780 10930 -6660
rect 10975 -6780 11095 -6660
rect 11150 -6780 11270 -6660
rect 11315 -6780 11435 -6660
rect 11480 -6780 11600 -6660
rect 11645 -6780 11765 -6660
rect 11820 -6780 11940 -6660
rect 11985 -6780 12105 -6660
rect 12150 -6780 12270 -6660
rect 12315 -6780 12435 -6660
rect 12490 -6780 12610 -6660
rect 7130 -6945 7250 -6825
rect 7295 -6945 7415 -6825
rect 7460 -6945 7580 -6825
rect 7625 -6945 7745 -6825
rect 7800 -6945 7920 -6825
rect 7965 -6945 8085 -6825
rect 8130 -6945 8250 -6825
rect 8295 -6945 8415 -6825
rect 8470 -6945 8590 -6825
rect 8635 -6945 8755 -6825
rect 8800 -6945 8920 -6825
rect 8965 -6945 9085 -6825
rect 9140 -6945 9260 -6825
rect 9305 -6945 9425 -6825
rect 9470 -6945 9590 -6825
rect 9635 -6945 9755 -6825
rect 9810 -6945 9930 -6825
rect 9975 -6945 10095 -6825
rect 10140 -6945 10260 -6825
rect 10305 -6945 10425 -6825
rect 10480 -6945 10600 -6825
rect 10645 -6945 10765 -6825
rect 10810 -6945 10930 -6825
rect 10975 -6945 11095 -6825
rect 11150 -6945 11270 -6825
rect 11315 -6945 11435 -6825
rect 11480 -6945 11600 -6825
rect 11645 -6945 11765 -6825
rect 11820 -6945 11940 -6825
rect 11985 -6945 12105 -6825
rect 12150 -6945 12270 -6825
rect 12315 -6945 12435 -6825
rect 12490 -6945 12610 -6825
rect 7130 -7110 7250 -6990
rect 7295 -7110 7415 -6990
rect 7460 -7110 7580 -6990
rect 7625 -7110 7745 -6990
rect 7800 -7110 7920 -6990
rect 7965 -7110 8085 -6990
rect 8130 -7110 8250 -6990
rect 8295 -7110 8415 -6990
rect 8470 -7110 8590 -6990
rect 8635 -7110 8755 -6990
rect 8800 -7110 8920 -6990
rect 8965 -7110 9085 -6990
rect 9140 -7110 9260 -6990
rect 9305 -7110 9425 -6990
rect 9470 -7110 9590 -6990
rect 9635 -7110 9755 -6990
rect 9810 -7110 9930 -6990
rect 9975 -7110 10095 -6990
rect 10140 -7110 10260 -6990
rect 10305 -7110 10425 -6990
rect 10480 -7110 10600 -6990
rect 10645 -7110 10765 -6990
rect 10810 -7110 10930 -6990
rect 10975 -7110 11095 -6990
rect 11150 -7110 11270 -6990
rect 11315 -7110 11435 -6990
rect 11480 -7110 11600 -6990
rect 11645 -7110 11765 -6990
rect 11820 -7110 11940 -6990
rect 11985 -7110 12105 -6990
rect 12150 -7110 12270 -6990
rect 12315 -7110 12435 -6990
rect 12490 -7110 12610 -6990
rect 7130 -7285 7250 -7165
rect 7295 -7285 7415 -7165
rect 7460 -7285 7580 -7165
rect 7625 -7285 7745 -7165
rect 7800 -7285 7920 -7165
rect 7965 -7285 8085 -7165
rect 8130 -7285 8250 -7165
rect 8295 -7285 8415 -7165
rect 8470 -7285 8590 -7165
rect 8635 -7285 8755 -7165
rect 8800 -7285 8920 -7165
rect 8965 -7285 9085 -7165
rect 9140 -7285 9260 -7165
rect 9305 -7285 9425 -7165
rect 9470 -7285 9590 -7165
rect 9635 -7285 9755 -7165
rect 9810 -7285 9930 -7165
rect 9975 -7285 10095 -7165
rect 10140 -7285 10260 -7165
rect 10305 -7285 10425 -7165
rect 10480 -7285 10600 -7165
rect 10645 -7285 10765 -7165
rect 10810 -7285 10930 -7165
rect 10975 -7285 11095 -7165
rect 11150 -7285 11270 -7165
rect 11315 -7285 11435 -7165
rect 11480 -7285 11600 -7165
rect 11645 -7285 11765 -7165
rect 11820 -7285 11940 -7165
rect 11985 -7285 12105 -7165
rect 12150 -7285 12270 -7165
rect 12315 -7285 12435 -7165
rect 12490 -7285 12610 -7165
rect 7130 -7450 7250 -7330
rect 7295 -7450 7415 -7330
rect 7460 -7450 7580 -7330
rect 7625 -7450 7745 -7330
rect 7800 -7450 7920 -7330
rect 7965 -7450 8085 -7330
rect 8130 -7450 8250 -7330
rect 8295 -7450 8415 -7330
rect 8470 -7450 8590 -7330
rect 8635 -7450 8755 -7330
rect 8800 -7450 8920 -7330
rect 8965 -7450 9085 -7330
rect 9140 -7450 9260 -7330
rect 9305 -7450 9425 -7330
rect 9470 -7450 9590 -7330
rect 9635 -7450 9755 -7330
rect 9810 -7450 9930 -7330
rect 9975 -7450 10095 -7330
rect 10140 -7450 10260 -7330
rect 10305 -7450 10425 -7330
rect 10480 -7450 10600 -7330
rect 10645 -7450 10765 -7330
rect 10810 -7450 10930 -7330
rect 10975 -7450 11095 -7330
rect 11150 -7450 11270 -7330
rect 11315 -7450 11435 -7330
rect 11480 -7450 11600 -7330
rect 11645 -7450 11765 -7330
rect 11820 -7450 11940 -7330
rect 11985 -7450 12105 -7330
rect 12150 -7450 12270 -7330
rect 12315 -7450 12435 -7330
rect 12490 -7450 12610 -7330
rect 7130 -7615 7250 -7495
rect 7295 -7615 7415 -7495
rect 7460 -7615 7580 -7495
rect 7625 -7615 7745 -7495
rect 7800 -7615 7920 -7495
rect 7965 -7615 8085 -7495
rect 8130 -7615 8250 -7495
rect 8295 -7615 8415 -7495
rect 8470 -7615 8590 -7495
rect 8635 -7615 8755 -7495
rect 8800 -7615 8920 -7495
rect 8965 -7615 9085 -7495
rect 9140 -7615 9260 -7495
rect 9305 -7615 9425 -7495
rect 9470 -7615 9590 -7495
rect 9635 -7615 9755 -7495
rect 9810 -7615 9930 -7495
rect 9975 -7615 10095 -7495
rect 10140 -7615 10260 -7495
rect 10305 -7615 10425 -7495
rect 10480 -7615 10600 -7495
rect 10645 -7615 10765 -7495
rect 10810 -7615 10930 -7495
rect 10975 -7615 11095 -7495
rect 11150 -7615 11270 -7495
rect 11315 -7615 11435 -7495
rect 11480 -7615 11600 -7495
rect 11645 -7615 11765 -7495
rect 11820 -7615 11940 -7495
rect 11985 -7615 12105 -7495
rect 12150 -7615 12270 -7495
rect 12315 -7615 12435 -7495
rect 12490 -7615 12610 -7495
rect 7130 -7780 7250 -7660
rect 7295 -7780 7415 -7660
rect 7460 -7780 7580 -7660
rect 7625 -7780 7745 -7660
rect 7800 -7780 7920 -7660
rect 7965 -7780 8085 -7660
rect 8130 -7780 8250 -7660
rect 8295 -7780 8415 -7660
rect 8470 -7780 8590 -7660
rect 8635 -7780 8755 -7660
rect 8800 -7780 8920 -7660
rect 8965 -7780 9085 -7660
rect 9140 -7780 9260 -7660
rect 9305 -7780 9425 -7660
rect 9470 -7780 9590 -7660
rect 9635 -7780 9755 -7660
rect 9810 -7780 9930 -7660
rect 9975 -7780 10095 -7660
rect 10140 -7780 10260 -7660
rect 10305 -7780 10425 -7660
rect 10480 -7780 10600 -7660
rect 10645 -7780 10765 -7660
rect 10810 -7780 10930 -7660
rect 10975 -7780 11095 -7660
rect 11150 -7780 11270 -7660
rect 11315 -7780 11435 -7660
rect 11480 -7780 11600 -7660
rect 11645 -7780 11765 -7660
rect 11820 -7780 11940 -7660
rect 11985 -7780 12105 -7660
rect 12150 -7780 12270 -7660
rect 12315 -7780 12435 -7660
rect 12490 -7780 12610 -7660
rect 7130 -7955 7250 -7835
rect 7295 -7955 7415 -7835
rect 7460 -7955 7580 -7835
rect 7625 -7955 7745 -7835
rect 7800 -7955 7920 -7835
rect 7965 -7955 8085 -7835
rect 8130 -7955 8250 -7835
rect 8295 -7955 8415 -7835
rect 8470 -7955 8590 -7835
rect 8635 -7955 8755 -7835
rect 8800 -7955 8920 -7835
rect 8965 -7955 9085 -7835
rect 9140 -7955 9260 -7835
rect 9305 -7955 9425 -7835
rect 9470 -7955 9590 -7835
rect 9635 -7955 9755 -7835
rect 9810 -7955 9930 -7835
rect 9975 -7955 10095 -7835
rect 10140 -7955 10260 -7835
rect 10305 -7955 10425 -7835
rect 10480 -7955 10600 -7835
rect 10645 -7955 10765 -7835
rect 10810 -7955 10930 -7835
rect 10975 -7955 11095 -7835
rect 11150 -7955 11270 -7835
rect 11315 -7955 11435 -7835
rect 11480 -7955 11600 -7835
rect 11645 -7955 11765 -7835
rect 11820 -7955 11940 -7835
rect 11985 -7955 12105 -7835
rect 12150 -7955 12270 -7835
rect 12315 -7955 12435 -7835
rect 12490 -7955 12610 -7835
rect 7130 -8120 7250 -8000
rect 7295 -8120 7415 -8000
rect 7460 -8120 7580 -8000
rect 7625 -8120 7745 -8000
rect 7800 -8120 7920 -8000
rect 7965 -8120 8085 -8000
rect 8130 -8120 8250 -8000
rect 8295 -8120 8415 -8000
rect 8470 -8120 8590 -8000
rect 8635 -8120 8755 -8000
rect 8800 -8120 8920 -8000
rect 8965 -8120 9085 -8000
rect 9140 -8120 9260 -8000
rect 9305 -8120 9425 -8000
rect 9470 -8120 9590 -8000
rect 9635 -8120 9755 -8000
rect 9810 -8120 9930 -8000
rect 9975 -8120 10095 -8000
rect 10140 -8120 10260 -8000
rect 10305 -8120 10425 -8000
rect 10480 -8120 10600 -8000
rect 10645 -8120 10765 -8000
rect 10810 -8120 10930 -8000
rect 10975 -8120 11095 -8000
rect 11150 -8120 11270 -8000
rect 11315 -8120 11435 -8000
rect 11480 -8120 11600 -8000
rect 11645 -8120 11765 -8000
rect 11820 -8120 11940 -8000
rect 11985 -8120 12105 -8000
rect 12150 -8120 12270 -8000
rect 12315 -8120 12435 -8000
rect 12490 -8120 12610 -8000
rect 7130 -8285 7250 -8165
rect 7295 -8285 7415 -8165
rect 7460 -8285 7580 -8165
rect 7625 -8285 7745 -8165
rect 7800 -8285 7920 -8165
rect 7965 -8285 8085 -8165
rect 8130 -8285 8250 -8165
rect 8295 -8285 8415 -8165
rect 8470 -8285 8590 -8165
rect 8635 -8285 8755 -8165
rect 8800 -8285 8920 -8165
rect 8965 -8285 9085 -8165
rect 9140 -8285 9260 -8165
rect 9305 -8285 9425 -8165
rect 9470 -8285 9590 -8165
rect 9635 -8285 9755 -8165
rect 9810 -8285 9930 -8165
rect 9975 -8285 10095 -8165
rect 10140 -8285 10260 -8165
rect 10305 -8285 10425 -8165
rect 10480 -8285 10600 -8165
rect 10645 -8285 10765 -8165
rect 10810 -8285 10930 -8165
rect 10975 -8285 11095 -8165
rect 11150 -8285 11270 -8165
rect 11315 -8285 11435 -8165
rect 11480 -8285 11600 -8165
rect 11645 -8285 11765 -8165
rect 11820 -8285 11940 -8165
rect 11985 -8285 12105 -8165
rect 12150 -8285 12270 -8165
rect 12315 -8285 12435 -8165
rect 12490 -8285 12610 -8165
rect 7130 -8450 7250 -8330
rect 7295 -8450 7415 -8330
rect 7460 -8450 7580 -8330
rect 7625 -8450 7745 -8330
rect 7800 -8450 7920 -8330
rect 7965 -8450 8085 -8330
rect 8130 -8450 8250 -8330
rect 8295 -8450 8415 -8330
rect 8470 -8450 8590 -8330
rect 8635 -8450 8755 -8330
rect 8800 -8450 8920 -8330
rect 8965 -8450 9085 -8330
rect 9140 -8450 9260 -8330
rect 9305 -8450 9425 -8330
rect 9470 -8450 9590 -8330
rect 9635 -8450 9755 -8330
rect 9810 -8450 9930 -8330
rect 9975 -8450 10095 -8330
rect 10140 -8450 10260 -8330
rect 10305 -8450 10425 -8330
rect 10480 -8450 10600 -8330
rect 10645 -8450 10765 -8330
rect 10810 -8450 10930 -8330
rect 10975 -8450 11095 -8330
rect 11150 -8450 11270 -8330
rect 11315 -8450 11435 -8330
rect 11480 -8450 11600 -8330
rect 11645 -8450 11765 -8330
rect 11820 -8450 11940 -8330
rect 11985 -8450 12105 -8330
rect 12150 -8450 12270 -8330
rect 12315 -8450 12435 -8330
rect 12490 -8450 12610 -8330
rect 7130 -8625 7250 -8505
rect 7295 -8625 7415 -8505
rect 7460 -8625 7580 -8505
rect 7625 -8625 7745 -8505
rect 7800 -8625 7920 -8505
rect 7965 -8625 8085 -8505
rect 8130 -8625 8250 -8505
rect 8295 -8625 8415 -8505
rect 8470 -8625 8590 -8505
rect 8635 -8625 8755 -8505
rect 8800 -8625 8920 -8505
rect 8965 -8625 9085 -8505
rect 9140 -8625 9260 -8505
rect 9305 -8625 9425 -8505
rect 9470 -8625 9590 -8505
rect 9635 -8625 9755 -8505
rect 9810 -8625 9930 -8505
rect 9975 -8625 10095 -8505
rect 10140 -8625 10260 -8505
rect 10305 -8625 10425 -8505
rect 10480 -8625 10600 -8505
rect 10645 -8625 10765 -8505
rect 10810 -8625 10930 -8505
rect 10975 -8625 11095 -8505
rect 11150 -8625 11270 -8505
rect 11315 -8625 11435 -8505
rect 11480 -8625 11600 -8505
rect 11645 -8625 11765 -8505
rect 11820 -8625 11940 -8505
rect 11985 -8625 12105 -8505
rect 12150 -8625 12270 -8505
rect 12315 -8625 12435 -8505
rect 12490 -8625 12610 -8505
rect 7130 -8790 7250 -8670
rect 7295 -8790 7415 -8670
rect 7460 -8790 7580 -8670
rect 7625 -8790 7745 -8670
rect 7800 -8790 7920 -8670
rect 7965 -8790 8085 -8670
rect 8130 -8790 8250 -8670
rect 8295 -8790 8415 -8670
rect 8470 -8790 8590 -8670
rect 8635 -8790 8755 -8670
rect 8800 -8790 8920 -8670
rect 8965 -8790 9085 -8670
rect 9140 -8790 9260 -8670
rect 9305 -8790 9425 -8670
rect 9470 -8790 9590 -8670
rect 9635 -8790 9755 -8670
rect 9810 -8790 9930 -8670
rect 9975 -8790 10095 -8670
rect 10140 -8790 10260 -8670
rect 10305 -8790 10425 -8670
rect 10480 -8790 10600 -8670
rect 10645 -8790 10765 -8670
rect 10810 -8790 10930 -8670
rect 10975 -8790 11095 -8670
rect 11150 -8790 11270 -8670
rect 11315 -8790 11435 -8670
rect 11480 -8790 11600 -8670
rect 11645 -8790 11765 -8670
rect 11820 -8790 11940 -8670
rect 11985 -8790 12105 -8670
rect 12150 -8790 12270 -8670
rect 12315 -8790 12435 -8670
rect 12490 -8790 12610 -8670
rect 7130 -8955 7250 -8835
rect 7295 -8955 7415 -8835
rect 7460 -8955 7580 -8835
rect 7625 -8955 7745 -8835
rect 7800 -8955 7920 -8835
rect 7965 -8955 8085 -8835
rect 8130 -8955 8250 -8835
rect 8295 -8955 8415 -8835
rect 8470 -8955 8590 -8835
rect 8635 -8955 8755 -8835
rect 8800 -8955 8920 -8835
rect 8965 -8955 9085 -8835
rect 9140 -8955 9260 -8835
rect 9305 -8955 9425 -8835
rect 9470 -8955 9590 -8835
rect 9635 -8955 9755 -8835
rect 9810 -8955 9930 -8835
rect 9975 -8955 10095 -8835
rect 10140 -8955 10260 -8835
rect 10305 -8955 10425 -8835
rect 10480 -8955 10600 -8835
rect 10645 -8955 10765 -8835
rect 10810 -8955 10930 -8835
rect 10975 -8955 11095 -8835
rect 11150 -8955 11270 -8835
rect 11315 -8955 11435 -8835
rect 11480 -8955 11600 -8835
rect 11645 -8955 11765 -8835
rect 11820 -8955 11940 -8835
rect 11985 -8955 12105 -8835
rect 12150 -8955 12270 -8835
rect 12315 -8955 12435 -8835
rect 12490 -8955 12610 -8835
rect 7130 -9120 7250 -9000
rect 7295 -9120 7415 -9000
rect 7460 -9120 7580 -9000
rect 7625 -9120 7745 -9000
rect 7800 -9120 7920 -9000
rect 7965 -9120 8085 -9000
rect 8130 -9120 8250 -9000
rect 8295 -9120 8415 -9000
rect 8470 -9120 8590 -9000
rect 8635 -9120 8755 -9000
rect 8800 -9120 8920 -9000
rect 8965 -9120 9085 -9000
rect 9140 -9120 9260 -9000
rect 9305 -9120 9425 -9000
rect 9470 -9120 9590 -9000
rect 9635 -9120 9755 -9000
rect 9810 -9120 9930 -9000
rect 9975 -9120 10095 -9000
rect 10140 -9120 10260 -9000
rect 10305 -9120 10425 -9000
rect 10480 -9120 10600 -9000
rect 10645 -9120 10765 -9000
rect 10810 -9120 10930 -9000
rect 10975 -9120 11095 -9000
rect 11150 -9120 11270 -9000
rect 11315 -9120 11435 -9000
rect 11480 -9120 11600 -9000
rect 11645 -9120 11765 -9000
rect 11820 -9120 11940 -9000
rect 11985 -9120 12105 -9000
rect 12150 -9120 12270 -9000
rect 12315 -9120 12435 -9000
rect 12490 -9120 12610 -9000
rect 7130 -9295 7250 -9175
rect 7295 -9295 7415 -9175
rect 7460 -9295 7580 -9175
rect 7625 -9295 7745 -9175
rect 7800 -9295 7920 -9175
rect 7965 -9295 8085 -9175
rect 8130 -9295 8250 -9175
rect 8295 -9295 8415 -9175
rect 8470 -9295 8590 -9175
rect 8635 -9295 8755 -9175
rect 8800 -9295 8920 -9175
rect 8965 -9295 9085 -9175
rect 9140 -9295 9260 -9175
rect 9305 -9295 9425 -9175
rect 9470 -9295 9590 -9175
rect 9635 -9295 9755 -9175
rect 9810 -9295 9930 -9175
rect 9975 -9295 10095 -9175
rect 10140 -9295 10260 -9175
rect 10305 -9295 10425 -9175
rect 10480 -9295 10600 -9175
rect 10645 -9295 10765 -9175
rect 10810 -9295 10930 -9175
rect 10975 -9295 11095 -9175
rect 11150 -9295 11270 -9175
rect 11315 -9295 11435 -9175
rect 11480 -9295 11600 -9175
rect 11645 -9295 11765 -9175
rect 11820 -9295 11940 -9175
rect 11985 -9295 12105 -9175
rect 12150 -9295 12270 -9175
rect 12315 -9295 12435 -9175
rect 12490 -9295 12610 -9175
rect 7130 -9460 7250 -9340
rect 7295 -9460 7415 -9340
rect 7460 -9460 7580 -9340
rect 7625 -9460 7745 -9340
rect 7800 -9460 7920 -9340
rect 7965 -9460 8085 -9340
rect 8130 -9460 8250 -9340
rect 8295 -9460 8415 -9340
rect 8470 -9460 8590 -9340
rect 8635 -9460 8755 -9340
rect 8800 -9460 8920 -9340
rect 8965 -9460 9085 -9340
rect 9140 -9460 9260 -9340
rect 9305 -9460 9425 -9340
rect 9470 -9460 9590 -9340
rect 9635 -9460 9755 -9340
rect 9810 -9460 9930 -9340
rect 9975 -9460 10095 -9340
rect 10140 -9460 10260 -9340
rect 10305 -9460 10425 -9340
rect 10480 -9460 10600 -9340
rect 10645 -9460 10765 -9340
rect 10810 -9460 10930 -9340
rect 10975 -9460 11095 -9340
rect 11150 -9460 11270 -9340
rect 11315 -9460 11435 -9340
rect 11480 -9460 11600 -9340
rect 11645 -9460 11765 -9340
rect 11820 -9460 11940 -9340
rect 11985 -9460 12105 -9340
rect 12150 -9460 12270 -9340
rect 12315 -9460 12435 -9340
rect 12490 -9460 12610 -9340
rect 7130 -9625 7250 -9505
rect 7295 -9625 7415 -9505
rect 7460 -9625 7580 -9505
rect 7625 -9625 7745 -9505
rect 7800 -9625 7920 -9505
rect 7965 -9625 8085 -9505
rect 8130 -9625 8250 -9505
rect 8295 -9625 8415 -9505
rect 8470 -9625 8590 -9505
rect 8635 -9625 8755 -9505
rect 8800 -9625 8920 -9505
rect 8965 -9625 9085 -9505
rect 9140 -9625 9260 -9505
rect 9305 -9625 9425 -9505
rect 9470 -9625 9590 -9505
rect 9635 -9625 9755 -9505
rect 9810 -9625 9930 -9505
rect 9975 -9625 10095 -9505
rect 10140 -9625 10260 -9505
rect 10305 -9625 10425 -9505
rect 10480 -9625 10600 -9505
rect 10645 -9625 10765 -9505
rect 10810 -9625 10930 -9505
rect 10975 -9625 11095 -9505
rect 11150 -9625 11270 -9505
rect 11315 -9625 11435 -9505
rect 11480 -9625 11600 -9505
rect 11645 -9625 11765 -9505
rect 11820 -9625 11940 -9505
rect 11985 -9625 12105 -9505
rect 12150 -9625 12270 -9505
rect 12315 -9625 12435 -9505
rect 12490 -9625 12610 -9505
rect 7130 -9790 7250 -9670
rect 7295 -9790 7415 -9670
rect 7460 -9790 7580 -9670
rect 7625 -9790 7745 -9670
rect 7800 -9790 7920 -9670
rect 7965 -9790 8085 -9670
rect 8130 -9790 8250 -9670
rect 8295 -9790 8415 -9670
rect 8470 -9790 8590 -9670
rect 8635 -9790 8755 -9670
rect 8800 -9790 8920 -9670
rect 8965 -9790 9085 -9670
rect 9140 -9790 9260 -9670
rect 9305 -9790 9425 -9670
rect 9470 -9790 9590 -9670
rect 9635 -9790 9755 -9670
rect 9810 -9790 9930 -9670
rect 9975 -9790 10095 -9670
rect 10140 -9790 10260 -9670
rect 10305 -9790 10425 -9670
rect 10480 -9790 10600 -9670
rect 10645 -9790 10765 -9670
rect 10810 -9790 10930 -9670
rect 10975 -9790 11095 -9670
rect 11150 -9790 11270 -9670
rect 11315 -9790 11435 -9670
rect 11480 -9790 11600 -9670
rect 11645 -9790 11765 -9670
rect 11820 -9790 11940 -9670
rect 11985 -9790 12105 -9670
rect 12150 -9790 12270 -9670
rect 12315 -9790 12435 -9670
rect 12490 -9790 12610 -9670
rect 12820 -4430 12940 -4310
rect 12985 -4430 13105 -4310
rect 13150 -4430 13270 -4310
rect 13315 -4430 13435 -4310
rect 13490 -4430 13610 -4310
rect 13655 -4430 13775 -4310
rect 13820 -4430 13940 -4310
rect 13985 -4430 14105 -4310
rect 14160 -4430 14280 -4310
rect 14325 -4430 14445 -4310
rect 14490 -4430 14610 -4310
rect 14655 -4430 14775 -4310
rect 14830 -4430 14950 -4310
rect 14995 -4430 15115 -4310
rect 15160 -4430 15280 -4310
rect 15325 -4430 15445 -4310
rect 15500 -4430 15620 -4310
rect 15665 -4430 15785 -4310
rect 15830 -4430 15950 -4310
rect 15995 -4430 16115 -4310
rect 16170 -4430 16290 -4310
rect 16335 -4430 16455 -4310
rect 16500 -4430 16620 -4310
rect 16665 -4430 16785 -4310
rect 16840 -4430 16960 -4310
rect 17005 -4430 17125 -4310
rect 17170 -4430 17290 -4310
rect 17335 -4430 17455 -4310
rect 17510 -4430 17630 -4310
rect 17675 -4430 17795 -4310
rect 17840 -4430 17960 -4310
rect 18005 -4430 18125 -4310
rect 18180 -4430 18300 -4310
rect 12820 -4605 12940 -4485
rect 12985 -4605 13105 -4485
rect 13150 -4605 13270 -4485
rect 13315 -4605 13435 -4485
rect 13490 -4605 13610 -4485
rect 13655 -4605 13775 -4485
rect 13820 -4605 13940 -4485
rect 13985 -4605 14105 -4485
rect 14160 -4605 14280 -4485
rect 14325 -4605 14445 -4485
rect 14490 -4605 14610 -4485
rect 14655 -4605 14775 -4485
rect 14830 -4605 14950 -4485
rect 14995 -4605 15115 -4485
rect 15160 -4605 15280 -4485
rect 15325 -4605 15445 -4485
rect 15500 -4605 15620 -4485
rect 15665 -4605 15785 -4485
rect 15830 -4605 15950 -4485
rect 15995 -4605 16115 -4485
rect 16170 -4605 16290 -4485
rect 16335 -4605 16455 -4485
rect 16500 -4605 16620 -4485
rect 16665 -4605 16785 -4485
rect 16840 -4605 16960 -4485
rect 17005 -4605 17125 -4485
rect 17170 -4605 17290 -4485
rect 17335 -4605 17455 -4485
rect 17510 -4605 17630 -4485
rect 17675 -4605 17795 -4485
rect 17840 -4605 17960 -4485
rect 18005 -4605 18125 -4485
rect 18180 -4605 18300 -4485
rect 12820 -4770 12940 -4650
rect 12985 -4770 13105 -4650
rect 13150 -4770 13270 -4650
rect 13315 -4770 13435 -4650
rect 13490 -4770 13610 -4650
rect 13655 -4770 13775 -4650
rect 13820 -4770 13940 -4650
rect 13985 -4770 14105 -4650
rect 14160 -4770 14280 -4650
rect 14325 -4770 14445 -4650
rect 14490 -4770 14610 -4650
rect 14655 -4770 14775 -4650
rect 14830 -4770 14950 -4650
rect 14995 -4770 15115 -4650
rect 15160 -4770 15280 -4650
rect 15325 -4770 15445 -4650
rect 15500 -4770 15620 -4650
rect 15665 -4770 15785 -4650
rect 15830 -4770 15950 -4650
rect 15995 -4770 16115 -4650
rect 16170 -4770 16290 -4650
rect 16335 -4770 16455 -4650
rect 16500 -4770 16620 -4650
rect 16665 -4770 16785 -4650
rect 16840 -4770 16960 -4650
rect 17005 -4770 17125 -4650
rect 17170 -4770 17290 -4650
rect 17335 -4770 17455 -4650
rect 17510 -4770 17630 -4650
rect 17675 -4770 17795 -4650
rect 17840 -4770 17960 -4650
rect 18005 -4770 18125 -4650
rect 18180 -4770 18300 -4650
rect 12820 -4935 12940 -4815
rect 12985 -4935 13105 -4815
rect 13150 -4935 13270 -4815
rect 13315 -4935 13435 -4815
rect 13490 -4935 13610 -4815
rect 13655 -4935 13775 -4815
rect 13820 -4935 13940 -4815
rect 13985 -4935 14105 -4815
rect 14160 -4935 14280 -4815
rect 14325 -4935 14445 -4815
rect 14490 -4935 14610 -4815
rect 14655 -4935 14775 -4815
rect 14830 -4935 14950 -4815
rect 14995 -4935 15115 -4815
rect 15160 -4935 15280 -4815
rect 15325 -4935 15445 -4815
rect 15500 -4935 15620 -4815
rect 15665 -4935 15785 -4815
rect 15830 -4935 15950 -4815
rect 15995 -4935 16115 -4815
rect 16170 -4935 16290 -4815
rect 16335 -4935 16455 -4815
rect 16500 -4935 16620 -4815
rect 16665 -4935 16785 -4815
rect 16840 -4935 16960 -4815
rect 17005 -4935 17125 -4815
rect 17170 -4935 17290 -4815
rect 17335 -4935 17455 -4815
rect 17510 -4935 17630 -4815
rect 17675 -4935 17795 -4815
rect 17840 -4935 17960 -4815
rect 18005 -4935 18125 -4815
rect 18180 -4935 18300 -4815
rect 12820 -5100 12940 -4980
rect 12985 -5100 13105 -4980
rect 13150 -5100 13270 -4980
rect 13315 -5100 13435 -4980
rect 13490 -5100 13610 -4980
rect 13655 -5100 13775 -4980
rect 13820 -5100 13940 -4980
rect 13985 -5100 14105 -4980
rect 14160 -5100 14280 -4980
rect 14325 -5100 14445 -4980
rect 14490 -5100 14610 -4980
rect 14655 -5100 14775 -4980
rect 14830 -5100 14950 -4980
rect 14995 -5100 15115 -4980
rect 15160 -5100 15280 -4980
rect 15325 -5100 15445 -4980
rect 15500 -5100 15620 -4980
rect 15665 -5100 15785 -4980
rect 15830 -5100 15950 -4980
rect 15995 -5100 16115 -4980
rect 16170 -5100 16290 -4980
rect 16335 -5100 16455 -4980
rect 16500 -5100 16620 -4980
rect 16665 -5100 16785 -4980
rect 16840 -5100 16960 -4980
rect 17005 -5100 17125 -4980
rect 17170 -5100 17290 -4980
rect 17335 -5100 17455 -4980
rect 17510 -5100 17630 -4980
rect 17675 -5100 17795 -4980
rect 17840 -5100 17960 -4980
rect 18005 -5100 18125 -4980
rect 18180 -5100 18300 -4980
rect 12820 -5275 12940 -5155
rect 12985 -5275 13105 -5155
rect 13150 -5275 13270 -5155
rect 13315 -5275 13435 -5155
rect 13490 -5275 13610 -5155
rect 13655 -5275 13775 -5155
rect 13820 -5275 13940 -5155
rect 13985 -5275 14105 -5155
rect 14160 -5275 14280 -5155
rect 14325 -5275 14445 -5155
rect 14490 -5275 14610 -5155
rect 14655 -5275 14775 -5155
rect 14830 -5275 14950 -5155
rect 14995 -5275 15115 -5155
rect 15160 -5275 15280 -5155
rect 15325 -5275 15445 -5155
rect 15500 -5275 15620 -5155
rect 15665 -5275 15785 -5155
rect 15830 -5275 15950 -5155
rect 15995 -5275 16115 -5155
rect 16170 -5275 16290 -5155
rect 16335 -5275 16455 -5155
rect 16500 -5275 16620 -5155
rect 16665 -5275 16785 -5155
rect 16840 -5275 16960 -5155
rect 17005 -5275 17125 -5155
rect 17170 -5275 17290 -5155
rect 17335 -5275 17455 -5155
rect 17510 -5275 17630 -5155
rect 17675 -5275 17795 -5155
rect 17840 -5275 17960 -5155
rect 18005 -5275 18125 -5155
rect 18180 -5275 18300 -5155
rect 12820 -5440 12940 -5320
rect 12985 -5440 13105 -5320
rect 13150 -5440 13270 -5320
rect 13315 -5440 13435 -5320
rect 13490 -5440 13610 -5320
rect 13655 -5440 13775 -5320
rect 13820 -5440 13940 -5320
rect 13985 -5440 14105 -5320
rect 14160 -5440 14280 -5320
rect 14325 -5440 14445 -5320
rect 14490 -5440 14610 -5320
rect 14655 -5440 14775 -5320
rect 14830 -5440 14950 -5320
rect 14995 -5440 15115 -5320
rect 15160 -5440 15280 -5320
rect 15325 -5440 15445 -5320
rect 15500 -5440 15620 -5320
rect 15665 -5440 15785 -5320
rect 15830 -5440 15950 -5320
rect 15995 -5440 16115 -5320
rect 16170 -5440 16290 -5320
rect 16335 -5440 16455 -5320
rect 16500 -5440 16620 -5320
rect 16665 -5440 16785 -5320
rect 16840 -5440 16960 -5320
rect 17005 -5440 17125 -5320
rect 17170 -5440 17290 -5320
rect 17335 -5440 17455 -5320
rect 17510 -5440 17630 -5320
rect 17675 -5440 17795 -5320
rect 17840 -5440 17960 -5320
rect 18005 -5440 18125 -5320
rect 18180 -5440 18300 -5320
rect 12820 -5605 12940 -5485
rect 12985 -5605 13105 -5485
rect 13150 -5605 13270 -5485
rect 13315 -5605 13435 -5485
rect 13490 -5605 13610 -5485
rect 13655 -5605 13775 -5485
rect 13820 -5605 13940 -5485
rect 13985 -5605 14105 -5485
rect 14160 -5605 14280 -5485
rect 14325 -5605 14445 -5485
rect 14490 -5605 14610 -5485
rect 14655 -5605 14775 -5485
rect 14830 -5605 14950 -5485
rect 14995 -5605 15115 -5485
rect 15160 -5605 15280 -5485
rect 15325 -5605 15445 -5485
rect 15500 -5605 15620 -5485
rect 15665 -5605 15785 -5485
rect 15830 -5605 15950 -5485
rect 15995 -5605 16115 -5485
rect 16170 -5605 16290 -5485
rect 16335 -5605 16455 -5485
rect 16500 -5605 16620 -5485
rect 16665 -5605 16785 -5485
rect 16840 -5605 16960 -5485
rect 17005 -5605 17125 -5485
rect 17170 -5605 17290 -5485
rect 17335 -5605 17455 -5485
rect 17510 -5605 17630 -5485
rect 17675 -5605 17795 -5485
rect 17840 -5605 17960 -5485
rect 18005 -5605 18125 -5485
rect 18180 -5605 18300 -5485
rect 12820 -5770 12940 -5650
rect 12985 -5770 13105 -5650
rect 13150 -5770 13270 -5650
rect 13315 -5770 13435 -5650
rect 13490 -5770 13610 -5650
rect 13655 -5770 13775 -5650
rect 13820 -5770 13940 -5650
rect 13985 -5770 14105 -5650
rect 14160 -5770 14280 -5650
rect 14325 -5770 14445 -5650
rect 14490 -5770 14610 -5650
rect 14655 -5770 14775 -5650
rect 14830 -5770 14950 -5650
rect 14995 -5770 15115 -5650
rect 15160 -5770 15280 -5650
rect 15325 -5770 15445 -5650
rect 15500 -5770 15620 -5650
rect 15665 -5770 15785 -5650
rect 15830 -5770 15950 -5650
rect 15995 -5770 16115 -5650
rect 16170 -5770 16290 -5650
rect 16335 -5770 16455 -5650
rect 16500 -5770 16620 -5650
rect 16665 -5770 16785 -5650
rect 16840 -5770 16960 -5650
rect 17005 -5770 17125 -5650
rect 17170 -5770 17290 -5650
rect 17335 -5770 17455 -5650
rect 17510 -5770 17630 -5650
rect 17675 -5770 17795 -5650
rect 17840 -5770 17960 -5650
rect 18005 -5770 18125 -5650
rect 18180 -5770 18300 -5650
rect 12820 -5945 12940 -5825
rect 12985 -5945 13105 -5825
rect 13150 -5945 13270 -5825
rect 13315 -5945 13435 -5825
rect 13490 -5945 13610 -5825
rect 13655 -5945 13775 -5825
rect 13820 -5945 13940 -5825
rect 13985 -5945 14105 -5825
rect 14160 -5945 14280 -5825
rect 14325 -5945 14445 -5825
rect 14490 -5945 14610 -5825
rect 14655 -5945 14775 -5825
rect 14830 -5945 14950 -5825
rect 14995 -5945 15115 -5825
rect 15160 -5945 15280 -5825
rect 15325 -5945 15445 -5825
rect 15500 -5945 15620 -5825
rect 15665 -5945 15785 -5825
rect 15830 -5945 15950 -5825
rect 15995 -5945 16115 -5825
rect 16170 -5945 16290 -5825
rect 16335 -5945 16455 -5825
rect 16500 -5945 16620 -5825
rect 16665 -5945 16785 -5825
rect 16840 -5945 16960 -5825
rect 17005 -5945 17125 -5825
rect 17170 -5945 17290 -5825
rect 17335 -5945 17455 -5825
rect 17510 -5945 17630 -5825
rect 17675 -5945 17795 -5825
rect 17840 -5945 17960 -5825
rect 18005 -5945 18125 -5825
rect 18180 -5945 18300 -5825
rect 12820 -6110 12940 -5990
rect 12985 -6110 13105 -5990
rect 13150 -6110 13270 -5990
rect 13315 -6110 13435 -5990
rect 13490 -6110 13610 -5990
rect 13655 -6110 13775 -5990
rect 13820 -6110 13940 -5990
rect 13985 -6110 14105 -5990
rect 14160 -6110 14280 -5990
rect 14325 -6110 14445 -5990
rect 14490 -6110 14610 -5990
rect 14655 -6110 14775 -5990
rect 14830 -6110 14950 -5990
rect 14995 -6110 15115 -5990
rect 15160 -6110 15280 -5990
rect 15325 -6110 15445 -5990
rect 15500 -6110 15620 -5990
rect 15665 -6110 15785 -5990
rect 15830 -6110 15950 -5990
rect 15995 -6110 16115 -5990
rect 16170 -6110 16290 -5990
rect 16335 -6110 16455 -5990
rect 16500 -6110 16620 -5990
rect 16665 -6110 16785 -5990
rect 16840 -6110 16960 -5990
rect 17005 -6110 17125 -5990
rect 17170 -6110 17290 -5990
rect 17335 -6110 17455 -5990
rect 17510 -6110 17630 -5990
rect 17675 -6110 17795 -5990
rect 17840 -6110 17960 -5990
rect 18005 -6110 18125 -5990
rect 18180 -6110 18300 -5990
rect 12820 -6275 12940 -6155
rect 12985 -6275 13105 -6155
rect 13150 -6275 13270 -6155
rect 13315 -6275 13435 -6155
rect 13490 -6275 13610 -6155
rect 13655 -6275 13775 -6155
rect 13820 -6275 13940 -6155
rect 13985 -6275 14105 -6155
rect 14160 -6275 14280 -6155
rect 14325 -6275 14445 -6155
rect 14490 -6275 14610 -6155
rect 14655 -6275 14775 -6155
rect 14830 -6275 14950 -6155
rect 14995 -6275 15115 -6155
rect 15160 -6275 15280 -6155
rect 15325 -6275 15445 -6155
rect 15500 -6275 15620 -6155
rect 15665 -6275 15785 -6155
rect 15830 -6275 15950 -6155
rect 15995 -6275 16115 -6155
rect 16170 -6275 16290 -6155
rect 16335 -6275 16455 -6155
rect 16500 -6275 16620 -6155
rect 16665 -6275 16785 -6155
rect 16840 -6275 16960 -6155
rect 17005 -6275 17125 -6155
rect 17170 -6275 17290 -6155
rect 17335 -6275 17455 -6155
rect 17510 -6275 17630 -6155
rect 17675 -6275 17795 -6155
rect 17840 -6275 17960 -6155
rect 18005 -6275 18125 -6155
rect 18180 -6275 18300 -6155
rect 12820 -6440 12940 -6320
rect 12985 -6440 13105 -6320
rect 13150 -6440 13270 -6320
rect 13315 -6440 13435 -6320
rect 13490 -6440 13610 -6320
rect 13655 -6440 13775 -6320
rect 13820 -6440 13940 -6320
rect 13985 -6440 14105 -6320
rect 14160 -6440 14280 -6320
rect 14325 -6440 14445 -6320
rect 14490 -6440 14610 -6320
rect 14655 -6440 14775 -6320
rect 14830 -6440 14950 -6320
rect 14995 -6440 15115 -6320
rect 15160 -6440 15280 -6320
rect 15325 -6440 15445 -6320
rect 15500 -6440 15620 -6320
rect 15665 -6440 15785 -6320
rect 15830 -6440 15950 -6320
rect 15995 -6440 16115 -6320
rect 16170 -6440 16290 -6320
rect 16335 -6440 16455 -6320
rect 16500 -6440 16620 -6320
rect 16665 -6440 16785 -6320
rect 16840 -6440 16960 -6320
rect 17005 -6440 17125 -6320
rect 17170 -6440 17290 -6320
rect 17335 -6440 17455 -6320
rect 17510 -6440 17630 -6320
rect 17675 -6440 17795 -6320
rect 17840 -6440 17960 -6320
rect 18005 -6440 18125 -6320
rect 18180 -6440 18300 -6320
rect 12820 -6615 12940 -6495
rect 12985 -6615 13105 -6495
rect 13150 -6615 13270 -6495
rect 13315 -6615 13435 -6495
rect 13490 -6615 13610 -6495
rect 13655 -6615 13775 -6495
rect 13820 -6615 13940 -6495
rect 13985 -6615 14105 -6495
rect 14160 -6615 14280 -6495
rect 14325 -6615 14445 -6495
rect 14490 -6615 14610 -6495
rect 14655 -6615 14775 -6495
rect 14830 -6615 14950 -6495
rect 14995 -6615 15115 -6495
rect 15160 -6615 15280 -6495
rect 15325 -6615 15445 -6495
rect 15500 -6615 15620 -6495
rect 15665 -6615 15785 -6495
rect 15830 -6615 15950 -6495
rect 15995 -6615 16115 -6495
rect 16170 -6615 16290 -6495
rect 16335 -6615 16455 -6495
rect 16500 -6615 16620 -6495
rect 16665 -6615 16785 -6495
rect 16840 -6615 16960 -6495
rect 17005 -6615 17125 -6495
rect 17170 -6615 17290 -6495
rect 17335 -6615 17455 -6495
rect 17510 -6615 17630 -6495
rect 17675 -6615 17795 -6495
rect 17840 -6615 17960 -6495
rect 18005 -6615 18125 -6495
rect 18180 -6615 18300 -6495
rect 12820 -6780 12940 -6660
rect 12985 -6780 13105 -6660
rect 13150 -6780 13270 -6660
rect 13315 -6780 13435 -6660
rect 13490 -6780 13610 -6660
rect 13655 -6780 13775 -6660
rect 13820 -6780 13940 -6660
rect 13985 -6780 14105 -6660
rect 14160 -6780 14280 -6660
rect 14325 -6780 14445 -6660
rect 14490 -6780 14610 -6660
rect 14655 -6780 14775 -6660
rect 14830 -6780 14950 -6660
rect 14995 -6780 15115 -6660
rect 15160 -6780 15280 -6660
rect 15325 -6780 15445 -6660
rect 15500 -6780 15620 -6660
rect 15665 -6780 15785 -6660
rect 15830 -6780 15950 -6660
rect 15995 -6780 16115 -6660
rect 16170 -6780 16290 -6660
rect 16335 -6780 16455 -6660
rect 16500 -6780 16620 -6660
rect 16665 -6780 16785 -6660
rect 16840 -6780 16960 -6660
rect 17005 -6780 17125 -6660
rect 17170 -6780 17290 -6660
rect 17335 -6780 17455 -6660
rect 17510 -6780 17630 -6660
rect 17675 -6780 17795 -6660
rect 17840 -6780 17960 -6660
rect 18005 -6780 18125 -6660
rect 18180 -6780 18300 -6660
rect 12820 -6945 12940 -6825
rect 12985 -6945 13105 -6825
rect 13150 -6945 13270 -6825
rect 13315 -6945 13435 -6825
rect 13490 -6945 13610 -6825
rect 13655 -6945 13775 -6825
rect 13820 -6945 13940 -6825
rect 13985 -6945 14105 -6825
rect 14160 -6945 14280 -6825
rect 14325 -6945 14445 -6825
rect 14490 -6945 14610 -6825
rect 14655 -6945 14775 -6825
rect 14830 -6945 14950 -6825
rect 14995 -6945 15115 -6825
rect 15160 -6945 15280 -6825
rect 15325 -6945 15445 -6825
rect 15500 -6945 15620 -6825
rect 15665 -6945 15785 -6825
rect 15830 -6945 15950 -6825
rect 15995 -6945 16115 -6825
rect 16170 -6945 16290 -6825
rect 16335 -6945 16455 -6825
rect 16500 -6945 16620 -6825
rect 16665 -6945 16785 -6825
rect 16840 -6945 16960 -6825
rect 17005 -6945 17125 -6825
rect 17170 -6945 17290 -6825
rect 17335 -6945 17455 -6825
rect 17510 -6945 17630 -6825
rect 17675 -6945 17795 -6825
rect 17840 -6945 17960 -6825
rect 18005 -6945 18125 -6825
rect 18180 -6945 18300 -6825
rect 12820 -7110 12940 -6990
rect 12985 -7110 13105 -6990
rect 13150 -7110 13270 -6990
rect 13315 -7110 13435 -6990
rect 13490 -7110 13610 -6990
rect 13655 -7110 13775 -6990
rect 13820 -7110 13940 -6990
rect 13985 -7110 14105 -6990
rect 14160 -7110 14280 -6990
rect 14325 -7110 14445 -6990
rect 14490 -7110 14610 -6990
rect 14655 -7110 14775 -6990
rect 14830 -7110 14950 -6990
rect 14995 -7110 15115 -6990
rect 15160 -7110 15280 -6990
rect 15325 -7110 15445 -6990
rect 15500 -7110 15620 -6990
rect 15665 -7110 15785 -6990
rect 15830 -7110 15950 -6990
rect 15995 -7110 16115 -6990
rect 16170 -7110 16290 -6990
rect 16335 -7110 16455 -6990
rect 16500 -7110 16620 -6990
rect 16665 -7110 16785 -6990
rect 16840 -7110 16960 -6990
rect 17005 -7110 17125 -6990
rect 17170 -7110 17290 -6990
rect 17335 -7110 17455 -6990
rect 17510 -7110 17630 -6990
rect 17675 -7110 17795 -6990
rect 17840 -7110 17960 -6990
rect 18005 -7110 18125 -6990
rect 18180 -7110 18300 -6990
rect 12820 -7285 12940 -7165
rect 12985 -7285 13105 -7165
rect 13150 -7285 13270 -7165
rect 13315 -7285 13435 -7165
rect 13490 -7285 13610 -7165
rect 13655 -7285 13775 -7165
rect 13820 -7285 13940 -7165
rect 13985 -7285 14105 -7165
rect 14160 -7285 14280 -7165
rect 14325 -7285 14445 -7165
rect 14490 -7285 14610 -7165
rect 14655 -7285 14775 -7165
rect 14830 -7285 14950 -7165
rect 14995 -7285 15115 -7165
rect 15160 -7285 15280 -7165
rect 15325 -7285 15445 -7165
rect 15500 -7285 15620 -7165
rect 15665 -7285 15785 -7165
rect 15830 -7285 15950 -7165
rect 15995 -7285 16115 -7165
rect 16170 -7285 16290 -7165
rect 16335 -7285 16455 -7165
rect 16500 -7285 16620 -7165
rect 16665 -7285 16785 -7165
rect 16840 -7285 16960 -7165
rect 17005 -7285 17125 -7165
rect 17170 -7285 17290 -7165
rect 17335 -7285 17455 -7165
rect 17510 -7285 17630 -7165
rect 17675 -7285 17795 -7165
rect 17840 -7285 17960 -7165
rect 18005 -7285 18125 -7165
rect 18180 -7285 18300 -7165
rect 12820 -7450 12940 -7330
rect 12985 -7450 13105 -7330
rect 13150 -7450 13270 -7330
rect 13315 -7450 13435 -7330
rect 13490 -7450 13610 -7330
rect 13655 -7450 13775 -7330
rect 13820 -7450 13940 -7330
rect 13985 -7450 14105 -7330
rect 14160 -7450 14280 -7330
rect 14325 -7450 14445 -7330
rect 14490 -7450 14610 -7330
rect 14655 -7450 14775 -7330
rect 14830 -7450 14950 -7330
rect 14995 -7450 15115 -7330
rect 15160 -7450 15280 -7330
rect 15325 -7450 15445 -7330
rect 15500 -7450 15620 -7330
rect 15665 -7450 15785 -7330
rect 15830 -7450 15950 -7330
rect 15995 -7450 16115 -7330
rect 16170 -7450 16290 -7330
rect 16335 -7450 16455 -7330
rect 16500 -7450 16620 -7330
rect 16665 -7450 16785 -7330
rect 16840 -7450 16960 -7330
rect 17005 -7450 17125 -7330
rect 17170 -7450 17290 -7330
rect 17335 -7450 17455 -7330
rect 17510 -7450 17630 -7330
rect 17675 -7450 17795 -7330
rect 17840 -7450 17960 -7330
rect 18005 -7450 18125 -7330
rect 18180 -7450 18300 -7330
rect 12820 -7615 12940 -7495
rect 12985 -7615 13105 -7495
rect 13150 -7615 13270 -7495
rect 13315 -7615 13435 -7495
rect 13490 -7615 13610 -7495
rect 13655 -7615 13775 -7495
rect 13820 -7615 13940 -7495
rect 13985 -7615 14105 -7495
rect 14160 -7615 14280 -7495
rect 14325 -7615 14445 -7495
rect 14490 -7615 14610 -7495
rect 14655 -7615 14775 -7495
rect 14830 -7615 14950 -7495
rect 14995 -7615 15115 -7495
rect 15160 -7615 15280 -7495
rect 15325 -7615 15445 -7495
rect 15500 -7615 15620 -7495
rect 15665 -7615 15785 -7495
rect 15830 -7615 15950 -7495
rect 15995 -7615 16115 -7495
rect 16170 -7615 16290 -7495
rect 16335 -7615 16455 -7495
rect 16500 -7615 16620 -7495
rect 16665 -7615 16785 -7495
rect 16840 -7615 16960 -7495
rect 17005 -7615 17125 -7495
rect 17170 -7615 17290 -7495
rect 17335 -7615 17455 -7495
rect 17510 -7615 17630 -7495
rect 17675 -7615 17795 -7495
rect 17840 -7615 17960 -7495
rect 18005 -7615 18125 -7495
rect 18180 -7615 18300 -7495
rect 12820 -7780 12940 -7660
rect 12985 -7780 13105 -7660
rect 13150 -7780 13270 -7660
rect 13315 -7780 13435 -7660
rect 13490 -7780 13610 -7660
rect 13655 -7780 13775 -7660
rect 13820 -7780 13940 -7660
rect 13985 -7780 14105 -7660
rect 14160 -7780 14280 -7660
rect 14325 -7780 14445 -7660
rect 14490 -7780 14610 -7660
rect 14655 -7780 14775 -7660
rect 14830 -7780 14950 -7660
rect 14995 -7780 15115 -7660
rect 15160 -7780 15280 -7660
rect 15325 -7780 15445 -7660
rect 15500 -7780 15620 -7660
rect 15665 -7780 15785 -7660
rect 15830 -7780 15950 -7660
rect 15995 -7780 16115 -7660
rect 16170 -7780 16290 -7660
rect 16335 -7780 16455 -7660
rect 16500 -7780 16620 -7660
rect 16665 -7780 16785 -7660
rect 16840 -7780 16960 -7660
rect 17005 -7780 17125 -7660
rect 17170 -7780 17290 -7660
rect 17335 -7780 17455 -7660
rect 17510 -7780 17630 -7660
rect 17675 -7780 17795 -7660
rect 17840 -7780 17960 -7660
rect 18005 -7780 18125 -7660
rect 18180 -7780 18300 -7660
rect 12820 -7955 12940 -7835
rect 12985 -7955 13105 -7835
rect 13150 -7955 13270 -7835
rect 13315 -7955 13435 -7835
rect 13490 -7955 13610 -7835
rect 13655 -7955 13775 -7835
rect 13820 -7955 13940 -7835
rect 13985 -7955 14105 -7835
rect 14160 -7955 14280 -7835
rect 14325 -7955 14445 -7835
rect 14490 -7955 14610 -7835
rect 14655 -7955 14775 -7835
rect 14830 -7955 14950 -7835
rect 14995 -7955 15115 -7835
rect 15160 -7955 15280 -7835
rect 15325 -7955 15445 -7835
rect 15500 -7955 15620 -7835
rect 15665 -7955 15785 -7835
rect 15830 -7955 15950 -7835
rect 15995 -7955 16115 -7835
rect 16170 -7955 16290 -7835
rect 16335 -7955 16455 -7835
rect 16500 -7955 16620 -7835
rect 16665 -7955 16785 -7835
rect 16840 -7955 16960 -7835
rect 17005 -7955 17125 -7835
rect 17170 -7955 17290 -7835
rect 17335 -7955 17455 -7835
rect 17510 -7955 17630 -7835
rect 17675 -7955 17795 -7835
rect 17840 -7955 17960 -7835
rect 18005 -7955 18125 -7835
rect 18180 -7955 18300 -7835
rect 12820 -8120 12940 -8000
rect 12985 -8120 13105 -8000
rect 13150 -8120 13270 -8000
rect 13315 -8120 13435 -8000
rect 13490 -8120 13610 -8000
rect 13655 -8120 13775 -8000
rect 13820 -8120 13940 -8000
rect 13985 -8120 14105 -8000
rect 14160 -8120 14280 -8000
rect 14325 -8120 14445 -8000
rect 14490 -8120 14610 -8000
rect 14655 -8120 14775 -8000
rect 14830 -8120 14950 -8000
rect 14995 -8120 15115 -8000
rect 15160 -8120 15280 -8000
rect 15325 -8120 15445 -8000
rect 15500 -8120 15620 -8000
rect 15665 -8120 15785 -8000
rect 15830 -8120 15950 -8000
rect 15995 -8120 16115 -8000
rect 16170 -8120 16290 -8000
rect 16335 -8120 16455 -8000
rect 16500 -8120 16620 -8000
rect 16665 -8120 16785 -8000
rect 16840 -8120 16960 -8000
rect 17005 -8120 17125 -8000
rect 17170 -8120 17290 -8000
rect 17335 -8120 17455 -8000
rect 17510 -8120 17630 -8000
rect 17675 -8120 17795 -8000
rect 17840 -8120 17960 -8000
rect 18005 -8120 18125 -8000
rect 18180 -8120 18300 -8000
rect 12820 -8285 12940 -8165
rect 12985 -8285 13105 -8165
rect 13150 -8285 13270 -8165
rect 13315 -8285 13435 -8165
rect 13490 -8285 13610 -8165
rect 13655 -8285 13775 -8165
rect 13820 -8285 13940 -8165
rect 13985 -8285 14105 -8165
rect 14160 -8285 14280 -8165
rect 14325 -8285 14445 -8165
rect 14490 -8285 14610 -8165
rect 14655 -8285 14775 -8165
rect 14830 -8285 14950 -8165
rect 14995 -8285 15115 -8165
rect 15160 -8285 15280 -8165
rect 15325 -8285 15445 -8165
rect 15500 -8285 15620 -8165
rect 15665 -8285 15785 -8165
rect 15830 -8285 15950 -8165
rect 15995 -8285 16115 -8165
rect 16170 -8285 16290 -8165
rect 16335 -8285 16455 -8165
rect 16500 -8285 16620 -8165
rect 16665 -8285 16785 -8165
rect 16840 -8285 16960 -8165
rect 17005 -8285 17125 -8165
rect 17170 -8285 17290 -8165
rect 17335 -8285 17455 -8165
rect 17510 -8285 17630 -8165
rect 17675 -8285 17795 -8165
rect 17840 -8285 17960 -8165
rect 18005 -8285 18125 -8165
rect 18180 -8285 18300 -8165
rect 12820 -8450 12940 -8330
rect 12985 -8450 13105 -8330
rect 13150 -8450 13270 -8330
rect 13315 -8450 13435 -8330
rect 13490 -8450 13610 -8330
rect 13655 -8450 13775 -8330
rect 13820 -8450 13940 -8330
rect 13985 -8450 14105 -8330
rect 14160 -8450 14280 -8330
rect 14325 -8450 14445 -8330
rect 14490 -8450 14610 -8330
rect 14655 -8450 14775 -8330
rect 14830 -8450 14950 -8330
rect 14995 -8450 15115 -8330
rect 15160 -8450 15280 -8330
rect 15325 -8450 15445 -8330
rect 15500 -8450 15620 -8330
rect 15665 -8450 15785 -8330
rect 15830 -8450 15950 -8330
rect 15995 -8450 16115 -8330
rect 16170 -8450 16290 -8330
rect 16335 -8450 16455 -8330
rect 16500 -8450 16620 -8330
rect 16665 -8450 16785 -8330
rect 16840 -8450 16960 -8330
rect 17005 -8450 17125 -8330
rect 17170 -8450 17290 -8330
rect 17335 -8450 17455 -8330
rect 17510 -8450 17630 -8330
rect 17675 -8450 17795 -8330
rect 17840 -8450 17960 -8330
rect 18005 -8450 18125 -8330
rect 18180 -8450 18300 -8330
rect 12820 -8625 12940 -8505
rect 12985 -8625 13105 -8505
rect 13150 -8625 13270 -8505
rect 13315 -8625 13435 -8505
rect 13490 -8625 13610 -8505
rect 13655 -8625 13775 -8505
rect 13820 -8625 13940 -8505
rect 13985 -8625 14105 -8505
rect 14160 -8625 14280 -8505
rect 14325 -8625 14445 -8505
rect 14490 -8625 14610 -8505
rect 14655 -8625 14775 -8505
rect 14830 -8625 14950 -8505
rect 14995 -8625 15115 -8505
rect 15160 -8625 15280 -8505
rect 15325 -8625 15445 -8505
rect 15500 -8625 15620 -8505
rect 15665 -8625 15785 -8505
rect 15830 -8625 15950 -8505
rect 15995 -8625 16115 -8505
rect 16170 -8625 16290 -8505
rect 16335 -8625 16455 -8505
rect 16500 -8625 16620 -8505
rect 16665 -8625 16785 -8505
rect 16840 -8625 16960 -8505
rect 17005 -8625 17125 -8505
rect 17170 -8625 17290 -8505
rect 17335 -8625 17455 -8505
rect 17510 -8625 17630 -8505
rect 17675 -8625 17795 -8505
rect 17840 -8625 17960 -8505
rect 18005 -8625 18125 -8505
rect 18180 -8625 18300 -8505
rect 12820 -8790 12940 -8670
rect 12985 -8790 13105 -8670
rect 13150 -8790 13270 -8670
rect 13315 -8790 13435 -8670
rect 13490 -8790 13610 -8670
rect 13655 -8790 13775 -8670
rect 13820 -8790 13940 -8670
rect 13985 -8790 14105 -8670
rect 14160 -8790 14280 -8670
rect 14325 -8790 14445 -8670
rect 14490 -8790 14610 -8670
rect 14655 -8790 14775 -8670
rect 14830 -8790 14950 -8670
rect 14995 -8790 15115 -8670
rect 15160 -8790 15280 -8670
rect 15325 -8790 15445 -8670
rect 15500 -8790 15620 -8670
rect 15665 -8790 15785 -8670
rect 15830 -8790 15950 -8670
rect 15995 -8790 16115 -8670
rect 16170 -8790 16290 -8670
rect 16335 -8790 16455 -8670
rect 16500 -8790 16620 -8670
rect 16665 -8790 16785 -8670
rect 16840 -8790 16960 -8670
rect 17005 -8790 17125 -8670
rect 17170 -8790 17290 -8670
rect 17335 -8790 17455 -8670
rect 17510 -8790 17630 -8670
rect 17675 -8790 17795 -8670
rect 17840 -8790 17960 -8670
rect 18005 -8790 18125 -8670
rect 18180 -8790 18300 -8670
rect 12820 -8955 12940 -8835
rect 12985 -8955 13105 -8835
rect 13150 -8955 13270 -8835
rect 13315 -8955 13435 -8835
rect 13490 -8955 13610 -8835
rect 13655 -8955 13775 -8835
rect 13820 -8955 13940 -8835
rect 13985 -8955 14105 -8835
rect 14160 -8955 14280 -8835
rect 14325 -8955 14445 -8835
rect 14490 -8955 14610 -8835
rect 14655 -8955 14775 -8835
rect 14830 -8955 14950 -8835
rect 14995 -8955 15115 -8835
rect 15160 -8955 15280 -8835
rect 15325 -8955 15445 -8835
rect 15500 -8955 15620 -8835
rect 15665 -8955 15785 -8835
rect 15830 -8955 15950 -8835
rect 15995 -8955 16115 -8835
rect 16170 -8955 16290 -8835
rect 16335 -8955 16455 -8835
rect 16500 -8955 16620 -8835
rect 16665 -8955 16785 -8835
rect 16840 -8955 16960 -8835
rect 17005 -8955 17125 -8835
rect 17170 -8955 17290 -8835
rect 17335 -8955 17455 -8835
rect 17510 -8955 17630 -8835
rect 17675 -8955 17795 -8835
rect 17840 -8955 17960 -8835
rect 18005 -8955 18125 -8835
rect 18180 -8955 18300 -8835
rect 12820 -9120 12940 -9000
rect 12985 -9120 13105 -9000
rect 13150 -9120 13270 -9000
rect 13315 -9120 13435 -9000
rect 13490 -9120 13610 -9000
rect 13655 -9120 13775 -9000
rect 13820 -9120 13940 -9000
rect 13985 -9120 14105 -9000
rect 14160 -9120 14280 -9000
rect 14325 -9120 14445 -9000
rect 14490 -9120 14610 -9000
rect 14655 -9120 14775 -9000
rect 14830 -9120 14950 -9000
rect 14995 -9120 15115 -9000
rect 15160 -9120 15280 -9000
rect 15325 -9120 15445 -9000
rect 15500 -9120 15620 -9000
rect 15665 -9120 15785 -9000
rect 15830 -9120 15950 -9000
rect 15995 -9120 16115 -9000
rect 16170 -9120 16290 -9000
rect 16335 -9120 16455 -9000
rect 16500 -9120 16620 -9000
rect 16665 -9120 16785 -9000
rect 16840 -9120 16960 -9000
rect 17005 -9120 17125 -9000
rect 17170 -9120 17290 -9000
rect 17335 -9120 17455 -9000
rect 17510 -9120 17630 -9000
rect 17675 -9120 17795 -9000
rect 17840 -9120 17960 -9000
rect 18005 -9120 18125 -9000
rect 18180 -9120 18300 -9000
rect 12820 -9295 12940 -9175
rect 12985 -9295 13105 -9175
rect 13150 -9295 13270 -9175
rect 13315 -9295 13435 -9175
rect 13490 -9295 13610 -9175
rect 13655 -9295 13775 -9175
rect 13820 -9295 13940 -9175
rect 13985 -9295 14105 -9175
rect 14160 -9295 14280 -9175
rect 14325 -9295 14445 -9175
rect 14490 -9295 14610 -9175
rect 14655 -9295 14775 -9175
rect 14830 -9295 14950 -9175
rect 14995 -9295 15115 -9175
rect 15160 -9295 15280 -9175
rect 15325 -9295 15445 -9175
rect 15500 -9295 15620 -9175
rect 15665 -9295 15785 -9175
rect 15830 -9295 15950 -9175
rect 15995 -9295 16115 -9175
rect 16170 -9295 16290 -9175
rect 16335 -9295 16455 -9175
rect 16500 -9295 16620 -9175
rect 16665 -9295 16785 -9175
rect 16840 -9295 16960 -9175
rect 17005 -9295 17125 -9175
rect 17170 -9295 17290 -9175
rect 17335 -9295 17455 -9175
rect 17510 -9295 17630 -9175
rect 17675 -9295 17795 -9175
rect 17840 -9295 17960 -9175
rect 18005 -9295 18125 -9175
rect 18180 -9295 18300 -9175
rect 12820 -9460 12940 -9340
rect 12985 -9460 13105 -9340
rect 13150 -9460 13270 -9340
rect 13315 -9460 13435 -9340
rect 13490 -9460 13610 -9340
rect 13655 -9460 13775 -9340
rect 13820 -9460 13940 -9340
rect 13985 -9460 14105 -9340
rect 14160 -9460 14280 -9340
rect 14325 -9460 14445 -9340
rect 14490 -9460 14610 -9340
rect 14655 -9460 14775 -9340
rect 14830 -9460 14950 -9340
rect 14995 -9460 15115 -9340
rect 15160 -9460 15280 -9340
rect 15325 -9460 15445 -9340
rect 15500 -9460 15620 -9340
rect 15665 -9460 15785 -9340
rect 15830 -9460 15950 -9340
rect 15995 -9460 16115 -9340
rect 16170 -9460 16290 -9340
rect 16335 -9460 16455 -9340
rect 16500 -9460 16620 -9340
rect 16665 -9460 16785 -9340
rect 16840 -9460 16960 -9340
rect 17005 -9460 17125 -9340
rect 17170 -9460 17290 -9340
rect 17335 -9460 17455 -9340
rect 17510 -9460 17630 -9340
rect 17675 -9460 17795 -9340
rect 17840 -9460 17960 -9340
rect 18005 -9460 18125 -9340
rect 18180 -9460 18300 -9340
rect 12820 -9625 12940 -9505
rect 12985 -9625 13105 -9505
rect 13150 -9625 13270 -9505
rect 13315 -9625 13435 -9505
rect 13490 -9625 13610 -9505
rect 13655 -9625 13775 -9505
rect 13820 -9625 13940 -9505
rect 13985 -9625 14105 -9505
rect 14160 -9625 14280 -9505
rect 14325 -9625 14445 -9505
rect 14490 -9625 14610 -9505
rect 14655 -9625 14775 -9505
rect 14830 -9625 14950 -9505
rect 14995 -9625 15115 -9505
rect 15160 -9625 15280 -9505
rect 15325 -9625 15445 -9505
rect 15500 -9625 15620 -9505
rect 15665 -9625 15785 -9505
rect 15830 -9625 15950 -9505
rect 15995 -9625 16115 -9505
rect 16170 -9625 16290 -9505
rect 16335 -9625 16455 -9505
rect 16500 -9625 16620 -9505
rect 16665 -9625 16785 -9505
rect 16840 -9625 16960 -9505
rect 17005 -9625 17125 -9505
rect 17170 -9625 17290 -9505
rect 17335 -9625 17455 -9505
rect 17510 -9625 17630 -9505
rect 17675 -9625 17795 -9505
rect 17840 -9625 17960 -9505
rect 18005 -9625 18125 -9505
rect 18180 -9625 18300 -9505
rect 12820 -9790 12940 -9670
rect 12985 -9790 13105 -9670
rect 13150 -9790 13270 -9670
rect 13315 -9790 13435 -9670
rect 13490 -9790 13610 -9670
rect 13655 -9790 13775 -9670
rect 13820 -9790 13940 -9670
rect 13985 -9790 14105 -9670
rect 14160 -9790 14280 -9670
rect 14325 -9790 14445 -9670
rect 14490 -9790 14610 -9670
rect 14655 -9790 14775 -9670
rect 14830 -9790 14950 -9670
rect 14995 -9790 15115 -9670
rect 15160 -9790 15280 -9670
rect 15325 -9790 15445 -9670
rect 15500 -9790 15620 -9670
rect 15665 -9790 15785 -9670
rect 15830 -9790 15950 -9670
rect 15995 -9790 16115 -9670
rect 16170 -9790 16290 -9670
rect 16335 -9790 16455 -9670
rect 16500 -9790 16620 -9670
rect 16665 -9790 16785 -9670
rect 16840 -9790 16960 -9670
rect 17005 -9790 17125 -9670
rect 17170 -9790 17290 -9670
rect 17335 -9790 17455 -9670
rect 17510 -9790 17630 -9670
rect 17675 -9790 17795 -9670
rect 17840 -9790 17960 -9670
rect 18005 -9790 18125 -9670
rect 18180 -9790 18300 -9670
rect 18510 -4430 18630 -4310
rect 18675 -4430 18795 -4310
rect 18840 -4430 18960 -4310
rect 19005 -4430 19125 -4310
rect 19180 -4430 19300 -4310
rect 19345 -4430 19465 -4310
rect 19510 -4430 19630 -4310
rect 19675 -4430 19795 -4310
rect 19850 -4430 19970 -4310
rect 20015 -4430 20135 -4310
rect 20180 -4430 20300 -4310
rect 20345 -4430 20465 -4310
rect 20520 -4430 20640 -4310
rect 20685 -4430 20805 -4310
rect 20850 -4430 20970 -4310
rect 21015 -4430 21135 -4310
rect 21190 -4430 21310 -4310
rect 21355 -4430 21475 -4310
rect 21520 -4430 21640 -4310
rect 21685 -4430 21805 -4310
rect 21860 -4430 21980 -4310
rect 22025 -4430 22145 -4310
rect 22190 -4430 22310 -4310
rect 22355 -4430 22475 -4310
rect 22530 -4430 22650 -4310
rect 22695 -4430 22815 -4310
rect 22860 -4430 22980 -4310
rect 23025 -4430 23145 -4310
rect 23200 -4430 23320 -4310
rect 23365 -4430 23485 -4310
rect 23530 -4430 23650 -4310
rect 23695 -4430 23815 -4310
rect 23870 -4430 23990 -4310
rect 18510 -4605 18630 -4485
rect 18675 -4605 18795 -4485
rect 18840 -4605 18960 -4485
rect 19005 -4605 19125 -4485
rect 19180 -4605 19300 -4485
rect 19345 -4605 19465 -4485
rect 19510 -4605 19630 -4485
rect 19675 -4605 19795 -4485
rect 19850 -4605 19970 -4485
rect 20015 -4605 20135 -4485
rect 20180 -4605 20300 -4485
rect 20345 -4605 20465 -4485
rect 20520 -4605 20640 -4485
rect 20685 -4605 20805 -4485
rect 20850 -4605 20970 -4485
rect 21015 -4605 21135 -4485
rect 21190 -4605 21310 -4485
rect 21355 -4605 21475 -4485
rect 21520 -4605 21640 -4485
rect 21685 -4605 21805 -4485
rect 21860 -4605 21980 -4485
rect 22025 -4605 22145 -4485
rect 22190 -4605 22310 -4485
rect 22355 -4605 22475 -4485
rect 22530 -4605 22650 -4485
rect 22695 -4605 22815 -4485
rect 22860 -4605 22980 -4485
rect 23025 -4605 23145 -4485
rect 23200 -4605 23320 -4485
rect 23365 -4605 23485 -4485
rect 23530 -4605 23650 -4485
rect 23695 -4605 23815 -4485
rect 23870 -4605 23990 -4485
rect 18510 -4770 18630 -4650
rect 18675 -4770 18795 -4650
rect 18840 -4770 18960 -4650
rect 19005 -4770 19125 -4650
rect 19180 -4770 19300 -4650
rect 19345 -4770 19465 -4650
rect 19510 -4770 19630 -4650
rect 19675 -4770 19795 -4650
rect 19850 -4770 19970 -4650
rect 20015 -4770 20135 -4650
rect 20180 -4770 20300 -4650
rect 20345 -4770 20465 -4650
rect 20520 -4770 20640 -4650
rect 20685 -4770 20805 -4650
rect 20850 -4770 20970 -4650
rect 21015 -4770 21135 -4650
rect 21190 -4770 21310 -4650
rect 21355 -4770 21475 -4650
rect 21520 -4770 21640 -4650
rect 21685 -4770 21805 -4650
rect 21860 -4770 21980 -4650
rect 22025 -4770 22145 -4650
rect 22190 -4770 22310 -4650
rect 22355 -4770 22475 -4650
rect 22530 -4770 22650 -4650
rect 22695 -4770 22815 -4650
rect 22860 -4770 22980 -4650
rect 23025 -4770 23145 -4650
rect 23200 -4770 23320 -4650
rect 23365 -4770 23485 -4650
rect 23530 -4770 23650 -4650
rect 23695 -4770 23815 -4650
rect 23870 -4770 23990 -4650
rect 18510 -4935 18630 -4815
rect 18675 -4935 18795 -4815
rect 18840 -4935 18960 -4815
rect 19005 -4935 19125 -4815
rect 19180 -4935 19300 -4815
rect 19345 -4935 19465 -4815
rect 19510 -4935 19630 -4815
rect 19675 -4935 19795 -4815
rect 19850 -4935 19970 -4815
rect 20015 -4935 20135 -4815
rect 20180 -4935 20300 -4815
rect 20345 -4935 20465 -4815
rect 20520 -4935 20640 -4815
rect 20685 -4935 20805 -4815
rect 20850 -4935 20970 -4815
rect 21015 -4935 21135 -4815
rect 21190 -4935 21310 -4815
rect 21355 -4935 21475 -4815
rect 21520 -4935 21640 -4815
rect 21685 -4935 21805 -4815
rect 21860 -4935 21980 -4815
rect 22025 -4935 22145 -4815
rect 22190 -4935 22310 -4815
rect 22355 -4935 22475 -4815
rect 22530 -4935 22650 -4815
rect 22695 -4935 22815 -4815
rect 22860 -4935 22980 -4815
rect 23025 -4935 23145 -4815
rect 23200 -4935 23320 -4815
rect 23365 -4935 23485 -4815
rect 23530 -4935 23650 -4815
rect 23695 -4935 23815 -4815
rect 23870 -4935 23990 -4815
rect 18510 -5100 18630 -4980
rect 18675 -5100 18795 -4980
rect 18840 -5100 18960 -4980
rect 19005 -5100 19125 -4980
rect 19180 -5100 19300 -4980
rect 19345 -5100 19465 -4980
rect 19510 -5100 19630 -4980
rect 19675 -5100 19795 -4980
rect 19850 -5100 19970 -4980
rect 20015 -5100 20135 -4980
rect 20180 -5100 20300 -4980
rect 20345 -5100 20465 -4980
rect 20520 -5100 20640 -4980
rect 20685 -5100 20805 -4980
rect 20850 -5100 20970 -4980
rect 21015 -5100 21135 -4980
rect 21190 -5100 21310 -4980
rect 21355 -5100 21475 -4980
rect 21520 -5100 21640 -4980
rect 21685 -5100 21805 -4980
rect 21860 -5100 21980 -4980
rect 22025 -5100 22145 -4980
rect 22190 -5100 22310 -4980
rect 22355 -5100 22475 -4980
rect 22530 -5100 22650 -4980
rect 22695 -5100 22815 -4980
rect 22860 -5100 22980 -4980
rect 23025 -5100 23145 -4980
rect 23200 -5100 23320 -4980
rect 23365 -5100 23485 -4980
rect 23530 -5100 23650 -4980
rect 23695 -5100 23815 -4980
rect 23870 -5100 23990 -4980
rect 18510 -5275 18630 -5155
rect 18675 -5275 18795 -5155
rect 18840 -5275 18960 -5155
rect 19005 -5275 19125 -5155
rect 19180 -5275 19300 -5155
rect 19345 -5275 19465 -5155
rect 19510 -5275 19630 -5155
rect 19675 -5275 19795 -5155
rect 19850 -5275 19970 -5155
rect 20015 -5275 20135 -5155
rect 20180 -5275 20300 -5155
rect 20345 -5275 20465 -5155
rect 20520 -5275 20640 -5155
rect 20685 -5275 20805 -5155
rect 20850 -5275 20970 -5155
rect 21015 -5275 21135 -5155
rect 21190 -5275 21310 -5155
rect 21355 -5275 21475 -5155
rect 21520 -5275 21640 -5155
rect 21685 -5275 21805 -5155
rect 21860 -5275 21980 -5155
rect 22025 -5275 22145 -5155
rect 22190 -5275 22310 -5155
rect 22355 -5275 22475 -5155
rect 22530 -5275 22650 -5155
rect 22695 -5275 22815 -5155
rect 22860 -5275 22980 -5155
rect 23025 -5275 23145 -5155
rect 23200 -5275 23320 -5155
rect 23365 -5275 23485 -5155
rect 23530 -5275 23650 -5155
rect 23695 -5275 23815 -5155
rect 23870 -5275 23990 -5155
rect 18510 -5440 18630 -5320
rect 18675 -5440 18795 -5320
rect 18840 -5440 18960 -5320
rect 19005 -5440 19125 -5320
rect 19180 -5440 19300 -5320
rect 19345 -5440 19465 -5320
rect 19510 -5440 19630 -5320
rect 19675 -5440 19795 -5320
rect 19850 -5440 19970 -5320
rect 20015 -5440 20135 -5320
rect 20180 -5440 20300 -5320
rect 20345 -5440 20465 -5320
rect 20520 -5440 20640 -5320
rect 20685 -5440 20805 -5320
rect 20850 -5440 20970 -5320
rect 21015 -5440 21135 -5320
rect 21190 -5440 21310 -5320
rect 21355 -5440 21475 -5320
rect 21520 -5440 21640 -5320
rect 21685 -5440 21805 -5320
rect 21860 -5440 21980 -5320
rect 22025 -5440 22145 -5320
rect 22190 -5440 22310 -5320
rect 22355 -5440 22475 -5320
rect 22530 -5440 22650 -5320
rect 22695 -5440 22815 -5320
rect 22860 -5440 22980 -5320
rect 23025 -5440 23145 -5320
rect 23200 -5440 23320 -5320
rect 23365 -5440 23485 -5320
rect 23530 -5440 23650 -5320
rect 23695 -5440 23815 -5320
rect 23870 -5440 23990 -5320
rect 18510 -5605 18630 -5485
rect 18675 -5605 18795 -5485
rect 18840 -5605 18960 -5485
rect 19005 -5605 19125 -5485
rect 19180 -5605 19300 -5485
rect 19345 -5605 19465 -5485
rect 19510 -5605 19630 -5485
rect 19675 -5605 19795 -5485
rect 19850 -5605 19970 -5485
rect 20015 -5605 20135 -5485
rect 20180 -5605 20300 -5485
rect 20345 -5605 20465 -5485
rect 20520 -5605 20640 -5485
rect 20685 -5605 20805 -5485
rect 20850 -5605 20970 -5485
rect 21015 -5605 21135 -5485
rect 21190 -5605 21310 -5485
rect 21355 -5605 21475 -5485
rect 21520 -5605 21640 -5485
rect 21685 -5605 21805 -5485
rect 21860 -5605 21980 -5485
rect 22025 -5605 22145 -5485
rect 22190 -5605 22310 -5485
rect 22355 -5605 22475 -5485
rect 22530 -5605 22650 -5485
rect 22695 -5605 22815 -5485
rect 22860 -5605 22980 -5485
rect 23025 -5605 23145 -5485
rect 23200 -5605 23320 -5485
rect 23365 -5605 23485 -5485
rect 23530 -5605 23650 -5485
rect 23695 -5605 23815 -5485
rect 23870 -5605 23990 -5485
rect 18510 -5770 18630 -5650
rect 18675 -5770 18795 -5650
rect 18840 -5770 18960 -5650
rect 19005 -5770 19125 -5650
rect 19180 -5770 19300 -5650
rect 19345 -5770 19465 -5650
rect 19510 -5770 19630 -5650
rect 19675 -5770 19795 -5650
rect 19850 -5770 19970 -5650
rect 20015 -5770 20135 -5650
rect 20180 -5770 20300 -5650
rect 20345 -5770 20465 -5650
rect 20520 -5770 20640 -5650
rect 20685 -5770 20805 -5650
rect 20850 -5770 20970 -5650
rect 21015 -5770 21135 -5650
rect 21190 -5770 21310 -5650
rect 21355 -5770 21475 -5650
rect 21520 -5770 21640 -5650
rect 21685 -5770 21805 -5650
rect 21860 -5770 21980 -5650
rect 22025 -5770 22145 -5650
rect 22190 -5770 22310 -5650
rect 22355 -5770 22475 -5650
rect 22530 -5770 22650 -5650
rect 22695 -5770 22815 -5650
rect 22860 -5770 22980 -5650
rect 23025 -5770 23145 -5650
rect 23200 -5770 23320 -5650
rect 23365 -5770 23485 -5650
rect 23530 -5770 23650 -5650
rect 23695 -5770 23815 -5650
rect 23870 -5770 23990 -5650
rect 18510 -5945 18630 -5825
rect 18675 -5945 18795 -5825
rect 18840 -5945 18960 -5825
rect 19005 -5945 19125 -5825
rect 19180 -5945 19300 -5825
rect 19345 -5945 19465 -5825
rect 19510 -5945 19630 -5825
rect 19675 -5945 19795 -5825
rect 19850 -5945 19970 -5825
rect 20015 -5945 20135 -5825
rect 20180 -5945 20300 -5825
rect 20345 -5945 20465 -5825
rect 20520 -5945 20640 -5825
rect 20685 -5945 20805 -5825
rect 20850 -5945 20970 -5825
rect 21015 -5945 21135 -5825
rect 21190 -5945 21310 -5825
rect 21355 -5945 21475 -5825
rect 21520 -5945 21640 -5825
rect 21685 -5945 21805 -5825
rect 21860 -5945 21980 -5825
rect 22025 -5945 22145 -5825
rect 22190 -5945 22310 -5825
rect 22355 -5945 22475 -5825
rect 22530 -5945 22650 -5825
rect 22695 -5945 22815 -5825
rect 22860 -5945 22980 -5825
rect 23025 -5945 23145 -5825
rect 23200 -5945 23320 -5825
rect 23365 -5945 23485 -5825
rect 23530 -5945 23650 -5825
rect 23695 -5945 23815 -5825
rect 23870 -5945 23990 -5825
rect 18510 -6110 18630 -5990
rect 18675 -6110 18795 -5990
rect 18840 -6110 18960 -5990
rect 19005 -6110 19125 -5990
rect 19180 -6110 19300 -5990
rect 19345 -6110 19465 -5990
rect 19510 -6110 19630 -5990
rect 19675 -6110 19795 -5990
rect 19850 -6110 19970 -5990
rect 20015 -6110 20135 -5990
rect 20180 -6110 20300 -5990
rect 20345 -6110 20465 -5990
rect 20520 -6110 20640 -5990
rect 20685 -6110 20805 -5990
rect 20850 -6110 20970 -5990
rect 21015 -6110 21135 -5990
rect 21190 -6110 21310 -5990
rect 21355 -6110 21475 -5990
rect 21520 -6110 21640 -5990
rect 21685 -6110 21805 -5990
rect 21860 -6110 21980 -5990
rect 22025 -6110 22145 -5990
rect 22190 -6110 22310 -5990
rect 22355 -6110 22475 -5990
rect 22530 -6110 22650 -5990
rect 22695 -6110 22815 -5990
rect 22860 -6110 22980 -5990
rect 23025 -6110 23145 -5990
rect 23200 -6110 23320 -5990
rect 23365 -6110 23485 -5990
rect 23530 -6110 23650 -5990
rect 23695 -6110 23815 -5990
rect 23870 -6110 23990 -5990
rect 18510 -6275 18630 -6155
rect 18675 -6275 18795 -6155
rect 18840 -6275 18960 -6155
rect 19005 -6275 19125 -6155
rect 19180 -6275 19300 -6155
rect 19345 -6275 19465 -6155
rect 19510 -6275 19630 -6155
rect 19675 -6275 19795 -6155
rect 19850 -6275 19970 -6155
rect 20015 -6275 20135 -6155
rect 20180 -6275 20300 -6155
rect 20345 -6275 20465 -6155
rect 20520 -6275 20640 -6155
rect 20685 -6275 20805 -6155
rect 20850 -6275 20970 -6155
rect 21015 -6275 21135 -6155
rect 21190 -6275 21310 -6155
rect 21355 -6275 21475 -6155
rect 21520 -6275 21640 -6155
rect 21685 -6275 21805 -6155
rect 21860 -6275 21980 -6155
rect 22025 -6275 22145 -6155
rect 22190 -6275 22310 -6155
rect 22355 -6275 22475 -6155
rect 22530 -6275 22650 -6155
rect 22695 -6275 22815 -6155
rect 22860 -6275 22980 -6155
rect 23025 -6275 23145 -6155
rect 23200 -6275 23320 -6155
rect 23365 -6275 23485 -6155
rect 23530 -6275 23650 -6155
rect 23695 -6275 23815 -6155
rect 23870 -6275 23990 -6155
rect 18510 -6440 18630 -6320
rect 18675 -6440 18795 -6320
rect 18840 -6440 18960 -6320
rect 19005 -6440 19125 -6320
rect 19180 -6440 19300 -6320
rect 19345 -6440 19465 -6320
rect 19510 -6440 19630 -6320
rect 19675 -6440 19795 -6320
rect 19850 -6440 19970 -6320
rect 20015 -6440 20135 -6320
rect 20180 -6440 20300 -6320
rect 20345 -6440 20465 -6320
rect 20520 -6440 20640 -6320
rect 20685 -6440 20805 -6320
rect 20850 -6440 20970 -6320
rect 21015 -6440 21135 -6320
rect 21190 -6440 21310 -6320
rect 21355 -6440 21475 -6320
rect 21520 -6440 21640 -6320
rect 21685 -6440 21805 -6320
rect 21860 -6440 21980 -6320
rect 22025 -6440 22145 -6320
rect 22190 -6440 22310 -6320
rect 22355 -6440 22475 -6320
rect 22530 -6440 22650 -6320
rect 22695 -6440 22815 -6320
rect 22860 -6440 22980 -6320
rect 23025 -6440 23145 -6320
rect 23200 -6440 23320 -6320
rect 23365 -6440 23485 -6320
rect 23530 -6440 23650 -6320
rect 23695 -6440 23815 -6320
rect 23870 -6440 23990 -6320
rect 18510 -6615 18630 -6495
rect 18675 -6615 18795 -6495
rect 18840 -6615 18960 -6495
rect 19005 -6615 19125 -6495
rect 19180 -6615 19300 -6495
rect 19345 -6615 19465 -6495
rect 19510 -6615 19630 -6495
rect 19675 -6615 19795 -6495
rect 19850 -6615 19970 -6495
rect 20015 -6615 20135 -6495
rect 20180 -6615 20300 -6495
rect 20345 -6615 20465 -6495
rect 20520 -6615 20640 -6495
rect 20685 -6615 20805 -6495
rect 20850 -6615 20970 -6495
rect 21015 -6615 21135 -6495
rect 21190 -6615 21310 -6495
rect 21355 -6615 21475 -6495
rect 21520 -6615 21640 -6495
rect 21685 -6615 21805 -6495
rect 21860 -6615 21980 -6495
rect 22025 -6615 22145 -6495
rect 22190 -6615 22310 -6495
rect 22355 -6615 22475 -6495
rect 22530 -6615 22650 -6495
rect 22695 -6615 22815 -6495
rect 22860 -6615 22980 -6495
rect 23025 -6615 23145 -6495
rect 23200 -6615 23320 -6495
rect 23365 -6615 23485 -6495
rect 23530 -6615 23650 -6495
rect 23695 -6615 23815 -6495
rect 23870 -6615 23990 -6495
rect 18510 -6780 18630 -6660
rect 18675 -6780 18795 -6660
rect 18840 -6780 18960 -6660
rect 19005 -6780 19125 -6660
rect 19180 -6780 19300 -6660
rect 19345 -6780 19465 -6660
rect 19510 -6780 19630 -6660
rect 19675 -6780 19795 -6660
rect 19850 -6780 19970 -6660
rect 20015 -6780 20135 -6660
rect 20180 -6780 20300 -6660
rect 20345 -6780 20465 -6660
rect 20520 -6780 20640 -6660
rect 20685 -6780 20805 -6660
rect 20850 -6780 20970 -6660
rect 21015 -6780 21135 -6660
rect 21190 -6780 21310 -6660
rect 21355 -6780 21475 -6660
rect 21520 -6780 21640 -6660
rect 21685 -6780 21805 -6660
rect 21860 -6780 21980 -6660
rect 22025 -6780 22145 -6660
rect 22190 -6780 22310 -6660
rect 22355 -6780 22475 -6660
rect 22530 -6780 22650 -6660
rect 22695 -6780 22815 -6660
rect 22860 -6780 22980 -6660
rect 23025 -6780 23145 -6660
rect 23200 -6780 23320 -6660
rect 23365 -6780 23485 -6660
rect 23530 -6780 23650 -6660
rect 23695 -6780 23815 -6660
rect 23870 -6780 23990 -6660
rect 18510 -6945 18630 -6825
rect 18675 -6945 18795 -6825
rect 18840 -6945 18960 -6825
rect 19005 -6945 19125 -6825
rect 19180 -6945 19300 -6825
rect 19345 -6945 19465 -6825
rect 19510 -6945 19630 -6825
rect 19675 -6945 19795 -6825
rect 19850 -6945 19970 -6825
rect 20015 -6945 20135 -6825
rect 20180 -6945 20300 -6825
rect 20345 -6945 20465 -6825
rect 20520 -6945 20640 -6825
rect 20685 -6945 20805 -6825
rect 20850 -6945 20970 -6825
rect 21015 -6945 21135 -6825
rect 21190 -6945 21310 -6825
rect 21355 -6945 21475 -6825
rect 21520 -6945 21640 -6825
rect 21685 -6945 21805 -6825
rect 21860 -6945 21980 -6825
rect 22025 -6945 22145 -6825
rect 22190 -6945 22310 -6825
rect 22355 -6945 22475 -6825
rect 22530 -6945 22650 -6825
rect 22695 -6945 22815 -6825
rect 22860 -6945 22980 -6825
rect 23025 -6945 23145 -6825
rect 23200 -6945 23320 -6825
rect 23365 -6945 23485 -6825
rect 23530 -6945 23650 -6825
rect 23695 -6945 23815 -6825
rect 23870 -6945 23990 -6825
rect 18510 -7110 18630 -6990
rect 18675 -7110 18795 -6990
rect 18840 -7110 18960 -6990
rect 19005 -7110 19125 -6990
rect 19180 -7110 19300 -6990
rect 19345 -7110 19465 -6990
rect 19510 -7110 19630 -6990
rect 19675 -7110 19795 -6990
rect 19850 -7110 19970 -6990
rect 20015 -7110 20135 -6990
rect 20180 -7110 20300 -6990
rect 20345 -7110 20465 -6990
rect 20520 -7110 20640 -6990
rect 20685 -7110 20805 -6990
rect 20850 -7110 20970 -6990
rect 21015 -7110 21135 -6990
rect 21190 -7110 21310 -6990
rect 21355 -7110 21475 -6990
rect 21520 -7110 21640 -6990
rect 21685 -7110 21805 -6990
rect 21860 -7110 21980 -6990
rect 22025 -7110 22145 -6990
rect 22190 -7110 22310 -6990
rect 22355 -7110 22475 -6990
rect 22530 -7110 22650 -6990
rect 22695 -7110 22815 -6990
rect 22860 -7110 22980 -6990
rect 23025 -7110 23145 -6990
rect 23200 -7110 23320 -6990
rect 23365 -7110 23485 -6990
rect 23530 -7110 23650 -6990
rect 23695 -7110 23815 -6990
rect 23870 -7110 23990 -6990
rect 18510 -7285 18630 -7165
rect 18675 -7285 18795 -7165
rect 18840 -7285 18960 -7165
rect 19005 -7285 19125 -7165
rect 19180 -7285 19300 -7165
rect 19345 -7285 19465 -7165
rect 19510 -7285 19630 -7165
rect 19675 -7285 19795 -7165
rect 19850 -7285 19970 -7165
rect 20015 -7285 20135 -7165
rect 20180 -7285 20300 -7165
rect 20345 -7285 20465 -7165
rect 20520 -7285 20640 -7165
rect 20685 -7285 20805 -7165
rect 20850 -7285 20970 -7165
rect 21015 -7285 21135 -7165
rect 21190 -7285 21310 -7165
rect 21355 -7285 21475 -7165
rect 21520 -7285 21640 -7165
rect 21685 -7285 21805 -7165
rect 21860 -7285 21980 -7165
rect 22025 -7285 22145 -7165
rect 22190 -7285 22310 -7165
rect 22355 -7285 22475 -7165
rect 22530 -7285 22650 -7165
rect 22695 -7285 22815 -7165
rect 22860 -7285 22980 -7165
rect 23025 -7285 23145 -7165
rect 23200 -7285 23320 -7165
rect 23365 -7285 23485 -7165
rect 23530 -7285 23650 -7165
rect 23695 -7285 23815 -7165
rect 23870 -7285 23990 -7165
rect 18510 -7450 18630 -7330
rect 18675 -7450 18795 -7330
rect 18840 -7450 18960 -7330
rect 19005 -7450 19125 -7330
rect 19180 -7450 19300 -7330
rect 19345 -7450 19465 -7330
rect 19510 -7450 19630 -7330
rect 19675 -7450 19795 -7330
rect 19850 -7450 19970 -7330
rect 20015 -7450 20135 -7330
rect 20180 -7450 20300 -7330
rect 20345 -7450 20465 -7330
rect 20520 -7450 20640 -7330
rect 20685 -7450 20805 -7330
rect 20850 -7450 20970 -7330
rect 21015 -7450 21135 -7330
rect 21190 -7450 21310 -7330
rect 21355 -7450 21475 -7330
rect 21520 -7450 21640 -7330
rect 21685 -7450 21805 -7330
rect 21860 -7450 21980 -7330
rect 22025 -7450 22145 -7330
rect 22190 -7450 22310 -7330
rect 22355 -7450 22475 -7330
rect 22530 -7450 22650 -7330
rect 22695 -7450 22815 -7330
rect 22860 -7450 22980 -7330
rect 23025 -7450 23145 -7330
rect 23200 -7450 23320 -7330
rect 23365 -7450 23485 -7330
rect 23530 -7450 23650 -7330
rect 23695 -7450 23815 -7330
rect 23870 -7450 23990 -7330
rect 18510 -7615 18630 -7495
rect 18675 -7615 18795 -7495
rect 18840 -7615 18960 -7495
rect 19005 -7615 19125 -7495
rect 19180 -7615 19300 -7495
rect 19345 -7615 19465 -7495
rect 19510 -7615 19630 -7495
rect 19675 -7615 19795 -7495
rect 19850 -7615 19970 -7495
rect 20015 -7615 20135 -7495
rect 20180 -7615 20300 -7495
rect 20345 -7615 20465 -7495
rect 20520 -7615 20640 -7495
rect 20685 -7615 20805 -7495
rect 20850 -7615 20970 -7495
rect 21015 -7615 21135 -7495
rect 21190 -7615 21310 -7495
rect 21355 -7615 21475 -7495
rect 21520 -7615 21640 -7495
rect 21685 -7615 21805 -7495
rect 21860 -7615 21980 -7495
rect 22025 -7615 22145 -7495
rect 22190 -7615 22310 -7495
rect 22355 -7615 22475 -7495
rect 22530 -7615 22650 -7495
rect 22695 -7615 22815 -7495
rect 22860 -7615 22980 -7495
rect 23025 -7615 23145 -7495
rect 23200 -7615 23320 -7495
rect 23365 -7615 23485 -7495
rect 23530 -7615 23650 -7495
rect 23695 -7615 23815 -7495
rect 23870 -7615 23990 -7495
rect 18510 -7780 18630 -7660
rect 18675 -7780 18795 -7660
rect 18840 -7780 18960 -7660
rect 19005 -7780 19125 -7660
rect 19180 -7780 19300 -7660
rect 19345 -7780 19465 -7660
rect 19510 -7780 19630 -7660
rect 19675 -7780 19795 -7660
rect 19850 -7780 19970 -7660
rect 20015 -7780 20135 -7660
rect 20180 -7780 20300 -7660
rect 20345 -7780 20465 -7660
rect 20520 -7780 20640 -7660
rect 20685 -7780 20805 -7660
rect 20850 -7780 20970 -7660
rect 21015 -7780 21135 -7660
rect 21190 -7780 21310 -7660
rect 21355 -7780 21475 -7660
rect 21520 -7780 21640 -7660
rect 21685 -7780 21805 -7660
rect 21860 -7780 21980 -7660
rect 22025 -7780 22145 -7660
rect 22190 -7780 22310 -7660
rect 22355 -7780 22475 -7660
rect 22530 -7780 22650 -7660
rect 22695 -7780 22815 -7660
rect 22860 -7780 22980 -7660
rect 23025 -7780 23145 -7660
rect 23200 -7780 23320 -7660
rect 23365 -7780 23485 -7660
rect 23530 -7780 23650 -7660
rect 23695 -7780 23815 -7660
rect 23870 -7780 23990 -7660
rect 18510 -7955 18630 -7835
rect 18675 -7955 18795 -7835
rect 18840 -7955 18960 -7835
rect 19005 -7955 19125 -7835
rect 19180 -7955 19300 -7835
rect 19345 -7955 19465 -7835
rect 19510 -7955 19630 -7835
rect 19675 -7955 19795 -7835
rect 19850 -7955 19970 -7835
rect 20015 -7955 20135 -7835
rect 20180 -7955 20300 -7835
rect 20345 -7955 20465 -7835
rect 20520 -7955 20640 -7835
rect 20685 -7955 20805 -7835
rect 20850 -7955 20970 -7835
rect 21015 -7955 21135 -7835
rect 21190 -7955 21310 -7835
rect 21355 -7955 21475 -7835
rect 21520 -7955 21640 -7835
rect 21685 -7955 21805 -7835
rect 21860 -7955 21980 -7835
rect 22025 -7955 22145 -7835
rect 22190 -7955 22310 -7835
rect 22355 -7955 22475 -7835
rect 22530 -7955 22650 -7835
rect 22695 -7955 22815 -7835
rect 22860 -7955 22980 -7835
rect 23025 -7955 23145 -7835
rect 23200 -7955 23320 -7835
rect 23365 -7955 23485 -7835
rect 23530 -7955 23650 -7835
rect 23695 -7955 23815 -7835
rect 23870 -7955 23990 -7835
rect 18510 -8120 18630 -8000
rect 18675 -8120 18795 -8000
rect 18840 -8120 18960 -8000
rect 19005 -8120 19125 -8000
rect 19180 -8120 19300 -8000
rect 19345 -8120 19465 -8000
rect 19510 -8120 19630 -8000
rect 19675 -8120 19795 -8000
rect 19850 -8120 19970 -8000
rect 20015 -8120 20135 -8000
rect 20180 -8120 20300 -8000
rect 20345 -8120 20465 -8000
rect 20520 -8120 20640 -8000
rect 20685 -8120 20805 -8000
rect 20850 -8120 20970 -8000
rect 21015 -8120 21135 -8000
rect 21190 -8120 21310 -8000
rect 21355 -8120 21475 -8000
rect 21520 -8120 21640 -8000
rect 21685 -8120 21805 -8000
rect 21860 -8120 21980 -8000
rect 22025 -8120 22145 -8000
rect 22190 -8120 22310 -8000
rect 22355 -8120 22475 -8000
rect 22530 -8120 22650 -8000
rect 22695 -8120 22815 -8000
rect 22860 -8120 22980 -8000
rect 23025 -8120 23145 -8000
rect 23200 -8120 23320 -8000
rect 23365 -8120 23485 -8000
rect 23530 -8120 23650 -8000
rect 23695 -8120 23815 -8000
rect 23870 -8120 23990 -8000
rect 18510 -8285 18630 -8165
rect 18675 -8285 18795 -8165
rect 18840 -8285 18960 -8165
rect 19005 -8285 19125 -8165
rect 19180 -8285 19300 -8165
rect 19345 -8285 19465 -8165
rect 19510 -8285 19630 -8165
rect 19675 -8285 19795 -8165
rect 19850 -8285 19970 -8165
rect 20015 -8285 20135 -8165
rect 20180 -8285 20300 -8165
rect 20345 -8285 20465 -8165
rect 20520 -8285 20640 -8165
rect 20685 -8285 20805 -8165
rect 20850 -8285 20970 -8165
rect 21015 -8285 21135 -8165
rect 21190 -8285 21310 -8165
rect 21355 -8285 21475 -8165
rect 21520 -8285 21640 -8165
rect 21685 -8285 21805 -8165
rect 21860 -8285 21980 -8165
rect 22025 -8285 22145 -8165
rect 22190 -8285 22310 -8165
rect 22355 -8285 22475 -8165
rect 22530 -8285 22650 -8165
rect 22695 -8285 22815 -8165
rect 22860 -8285 22980 -8165
rect 23025 -8285 23145 -8165
rect 23200 -8285 23320 -8165
rect 23365 -8285 23485 -8165
rect 23530 -8285 23650 -8165
rect 23695 -8285 23815 -8165
rect 23870 -8285 23990 -8165
rect 18510 -8450 18630 -8330
rect 18675 -8450 18795 -8330
rect 18840 -8450 18960 -8330
rect 19005 -8450 19125 -8330
rect 19180 -8450 19300 -8330
rect 19345 -8450 19465 -8330
rect 19510 -8450 19630 -8330
rect 19675 -8450 19795 -8330
rect 19850 -8450 19970 -8330
rect 20015 -8450 20135 -8330
rect 20180 -8450 20300 -8330
rect 20345 -8450 20465 -8330
rect 20520 -8450 20640 -8330
rect 20685 -8450 20805 -8330
rect 20850 -8450 20970 -8330
rect 21015 -8450 21135 -8330
rect 21190 -8450 21310 -8330
rect 21355 -8450 21475 -8330
rect 21520 -8450 21640 -8330
rect 21685 -8450 21805 -8330
rect 21860 -8450 21980 -8330
rect 22025 -8450 22145 -8330
rect 22190 -8450 22310 -8330
rect 22355 -8450 22475 -8330
rect 22530 -8450 22650 -8330
rect 22695 -8450 22815 -8330
rect 22860 -8450 22980 -8330
rect 23025 -8450 23145 -8330
rect 23200 -8450 23320 -8330
rect 23365 -8450 23485 -8330
rect 23530 -8450 23650 -8330
rect 23695 -8450 23815 -8330
rect 23870 -8450 23990 -8330
rect 18510 -8625 18630 -8505
rect 18675 -8625 18795 -8505
rect 18840 -8625 18960 -8505
rect 19005 -8625 19125 -8505
rect 19180 -8625 19300 -8505
rect 19345 -8625 19465 -8505
rect 19510 -8625 19630 -8505
rect 19675 -8625 19795 -8505
rect 19850 -8625 19970 -8505
rect 20015 -8625 20135 -8505
rect 20180 -8625 20300 -8505
rect 20345 -8625 20465 -8505
rect 20520 -8625 20640 -8505
rect 20685 -8625 20805 -8505
rect 20850 -8625 20970 -8505
rect 21015 -8625 21135 -8505
rect 21190 -8625 21310 -8505
rect 21355 -8625 21475 -8505
rect 21520 -8625 21640 -8505
rect 21685 -8625 21805 -8505
rect 21860 -8625 21980 -8505
rect 22025 -8625 22145 -8505
rect 22190 -8625 22310 -8505
rect 22355 -8625 22475 -8505
rect 22530 -8625 22650 -8505
rect 22695 -8625 22815 -8505
rect 22860 -8625 22980 -8505
rect 23025 -8625 23145 -8505
rect 23200 -8625 23320 -8505
rect 23365 -8625 23485 -8505
rect 23530 -8625 23650 -8505
rect 23695 -8625 23815 -8505
rect 23870 -8625 23990 -8505
rect 18510 -8790 18630 -8670
rect 18675 -8790 18795 -8670
rect 18840 -8790 18960 -8670
rect 19005 -8790 19125 -8670
rect 19180 -8790 19300 -8670
rect 19345 -8790 19465 -8670
rect 19510 -8790 19630 -8670
rect 19675 -8790 19795 -8670
rect 19850 -8790 19970 -8670
rect 20015 -8790 20135 -8670
rect 20180 -8790 20300 -8670
rect 20345 -8790 20465 -8670
rect 20520 -8790 20640 -8670
rect 20685 -8790 20805 -8670
rect 20850 -8790 20970 -8670
rect 21015 -8790 21135 -8670
rect 21190 -8790 21310 -8670
rect 21355 -8790 21475 -8670
rect 21520 -8790 21640 -8670
rect 21685 -8790 21805 -8670
rect 21860 -8790 21980 -8670
rect 22025 -8790 22145 -8670
rect 22190 -8790 22310 -8670
rect 22355 -8790 22475 -8670
rect 22530 -8790 22650 -8670
rect 22695 -8790 22815 -8670
rect 22860 -8790 22980 -8670
rect 23025 -8790 23145 -8670
rect 23200 -8790 23320 -8670
rect 23365 -8790 23485 -8670
rect 23530 -8790 23650 -8670
rect 23695 -8790 23815 -8670
rect 23870 -8790 23990 -8670
rect 18510 -8955 18630 -8835
rect 18675 -8955 18795 -8835
rect 18840 -8955 18960 -8835
rect 19005 -8955 19125 -8835
rect 19180 -8955 19300 -8835
rect 19345 -8955 19465 -8835
rect 19510 -8955 19630 -8835
rect 19675 -8955 19795 -8835
rect 19850 -8955 19970 -8835
rect 20015 -8955 20135 -8835
rect 20180 -8955 20300 -8835
rect 20345 -8955 20465 -8835
rect 20520 -8955 20640 -8835
rect 20685 -8955 20805 -8835
rect 20850 -8955 20970 -8835
rect 21015 -8955 21135 -8835
rect 21190 -8955 21310 -8835
rect 21355 -8955 21475 -8835
rect 21520 -8955 21640 -8835
rect 21685 -8955 21805 -8835
rect 21860 -8955 21980 -8835
rect 22025 -8955 22145 -8835
rect 22190 -8955 22310 -8835
rect 22355 -8955 22475 -8835
rect 22530 -8955 22650 -8835
rect 22695 -8955 22815 -8835
rect 22860 -8955 22980 -8835
rect 23025 -8955 23145 -8835
rect 23200 -8955 23320 -8835
rect 23365 -8955 23485 -8835
rect 23530 -8955 23650 -8835
rect 23695 -8955 23815 -8835
rect 23870 -8955 23990 -8835
rect 18510 -9120 18630 -9000
rect 18675 -9120 18795 -9000
rect 18840 -9120 18960 -9000
rect 19005 -9120 19125 -9000
rect 19180 -9120 19300 -9000
rect 19345 -9120 19465 -9000
rect 19510 -9120 19630 -9000
rect 19675 -9120 19795 -9000
rect 19850 -9120 19970 -9000
rect 20015 -9120 20135 -9000
rect 20180 -9120 20300 -9000
rect 20345 -9120 20465 -9000
rect 20520 -9120 20640 -9000
rect 20685 -9120 20805 -9000
rect 20850 -9120 20970 -9000
rect 21015 -9120 21135 -9000
rect 21190 -9120 21310 -9000
rect 21355 -9120 21475 -9000
rect 21520 -9120 21640 -9000
rect 21685 -9120 21805 -9000
rect 21860 -9120 21980 -9000
rect 22025 -9120 22145 -9000
rect 22190 -9120 22310 -9000
rect 22355 -9120 22475 -9000
rect 22530 -9120 22650 -9000
rect 22695 -9120 22815 -9000
rect 22860 -9120 22980 -9000
rect 23025 -9120 23145 -9000
rect 23200 -9120 23320 -9000
rect 23365 -9120 23485 -9000
rect 23530 -9120 23650 -9000
rect 23695 -9120 23815 -9000
rect 23870 -9120 23990 -9000
rect 18510 -9295 18630 -9175
rect 18675 -9295 18795 -9175
rect 18840 -9295 18960 -9175
rect 19005 -9295 19125 -9175
rect 19180 -9295 19300 -9175
rect 19345 -9295 19465 -9175
rect 19510 -9295 19630 -9175
rect 19675 -9295 19795 -9175
rect 19850 -9295 19970 -9175
rect 20015 -9295 20135 -9175
rect 20180 -9295 20300 -9175
rect 20345 -9295 20465 -9175
rect 20520 -9295 20640 -9175
rect 20685 -9295 20805 -9175
rect 20850 -9295 20970 -9175
rect 21015 -9295 21135 -9175
rect 21190 -9295 21310 -9175
rect 21355 -9295 21475 -9175
rect 21520 -9295 21640 -9175
rect 21685 -9295 21805 -9175
rect 21860 -9295 21980 -9175
rect 22025 -9295 22145 -9175
rect 22190 -9295 22310 -9175
rect 22355 -9295 22475 -9175
rect 22530 -9295 22650 -9175
rect 22695 -9295 22815 -9175
rect 22860 -9295 22980 -9175
rect 23025 -9295 23145 -9175
rect 23200 -9295 23320 -9175
rect 23365 -9295 23485 -9175
rect 23530 -9295 23650 -9175
rect 23695 -9295 23815 -9175
rect 23870 -9295 23990 -9175
rect 18510 -9460 18630 -9340
rect 18675 -9460 18795 -9340
rect 18840 -9460 18960 -9340
rect 19005 -9460 19125 -9340
rect 19180 -9460 19300 -9340
rect 19345 -9460 19465 -9340
rect 19510 -9460 19630 -9340
rect 19675 -9460 19795 -9340
rect 19850 -9460 19970 -9340
rect 20015 -9460 20135 -9340
rect 20180 -9460 20300 -9340
rect 20345 -9460 20465 -9340
rect 20520 -9460 20640 -9340
rect 20685 -9460 20805 -9340
rect 20850 -9460 20970 -9340
rect 21015 -9460 21135 -9340
rect 21190 -9460 21310 -9340
rect 21355 -9460 21475 -9340
rect 21520 -9460 21640 -9340
rect 21685 -9460 21805 -9340
rect 21860 -9460 21980 -9340
rect 22025 -9460 22145 -9340
rect 22190 -9460 22310 -9340
rect 22355 -9460 22475 -9340
rect 22530 -9460 22650 -9340
rect 22695 -9460 22815 -9340
rect 22860 -9460 22980 -9340
rect 23025 -9460 23145 -9340
rect 23200 -9460 23320 -9340
rect 23365 -9460 23485 -9340
rect 23530 -9460 23650 -9340
rect 23695 -9460 23815 -9340
rect 23870 -9460 23990 -9340
rect 18510 -9625 18630 -9505
rect 18675 -9625 18795 -9505
rect 18840 -9625 18960 -9505
rect 19005 -9625 19125 -9505
rect 19180 -9625 19300 -9505
rect 19345 -9625 19465 -9505
rect 19510 -9625 19630 -9505
rect 19675 -9625 19795 -9505
rect 19850 -9625 19970 -9505
rect 20015 -9625 20135 -9505
rect 20180 -9625 20300 -9505
rect 20345 -9625 20465 -9505
rect 20520 -9625 20640 -9505
rect 20685 -9625 20805 -9505
rect 20850 -9625 20970 -9505
rect 21015 -9625 21135 -9505
rect 21190 -9625 21310 -9505
rect 21355 -9625 21475 -9505
rect 21520 -9625 21640 -9505
rect 21685 -9625 21805 -9505
rect 21860 -9625 21980 -9505
rect 22025 -9625 22145 -9505
rect 22190 -9625 22310 -9505
rect 22355 -9625 22475 -9505
rect 22530 -9625 22650 -9505
rect 22695 -9625 22815 -9505
rect 22860 -9625 22980 -9505
rect 23025 -9625 23145 -9505
rect 23200 -9625 23320 -9505
rect 23365 -9625 23485 -9505
rect 23530 -9625 23650 -9505
rect 23695 -9625 23815 -9505
rect 23870 -9625 23990 -9505
rect 18510 -9790 18630 -9670
rect 18675 -9790 18795 -9670
rect 18840 -9790 18960 -9670
rect 19005 -9790 19125 -9670
rect 19180 -9790 19300 -9670
rect 19345 -9790 19465 -9670
rect 19510 -9790 19630 -9670
rect 19675 -9790 19795 -9670
rect 19850 -9790 19970 -9670
rect 20015 -9790 20135 -9670
rect 20180 -9790 20300 -9670
rect 20345 -9790 20465 -9670
rect 20520 -9790 20640 -9670
rect 20685 -9790 20805 -9670
rect 20850 -9790 20970 -9670
rect 21015 -9790 21135 -9670
rect 21190 -9790 21310 -9670
rect 21355 -9790 21475 -9670
rect 21520 -9790 21640 -9670
rect 21685 -9790 21805 -9670
rect 21860 -9790 21980 -9670
rect 22025 -9790 22145 -9670
rect 22190 -9790 22310 -9670
rect 22355 -9790 22475 -9670
rect 22530 -9790 22650 -9670
rect 22695 -9790 22815 -9670
rect 22860 -9790 22980 -9670
rect 23025 -9790 23145 -9670
rect 23200 -9790 23320 -9670
rect 23365 -9790 23485 -9670
rect 23530 -9790 23650 -9670
rect 23695 -9790 23815 -9670
rect 23870 -9790 23990 -9670
rect 24200 -4430 24320 -4310
rect 24365 -4430 24485 -4310
rect 24530 -4430 24650 -4310
rect 24695 -4430 24815 -4310
rect 24870 -4430 24990 -4310
rect 25035 -4430 25155 -4310
rect 25200 -4430 25320 -4310
rect 25365 -4430 25485 -4310
rect 25540 -4430 25660 -4310
rect 25705 -4430 25825 -4310
rect 25870 -4430 25990 -4310
rect 26035 -4430 26155 -4310
rect 26210 -4430 26330 -4310
rect 26375 -4430 26495 -4310
rect 26540 -4430 26660 -4310
rect 26705 -4430 26825 -4310
rect 26880 -4430 27000 -4310
rect 27045 -4430 27165 -4310
rect 27210 -4430 27330 -4310
rect 27375 -4430 27495 -4310
rect 27550 -4430 27670 -4310
rect 27715 -4430 27835 -4310
rect 27880 -4430 28000 -4310
rect 28045 -4430 28165 -4310
rect 28220 -4430 28340 -4310
rect 28385 -4430 28505 -4310
rect 28550 -4430 28670 -4310
rect 28715 -4430 28835 -4310
rect 28890 -4430 29010 -4310
rect 29055 -4430 29175 -4310
rect 29220 -4430 29340 -4310
rect 29385 -4430 29505 -4310
rect 29560 -4430 29680 -4310
rect 24200 -4605 24320 -4485
rect 24365 -4605 24485 -4485
rect 24530 -4605 24650 -4485
rect 24695 -4605 24815 -4485
rect 24870 -4605 24990 -4485
rect 25035 -4605 25155 -4485
rect 25200 -4605 25320 -4485
rect 25365 -4605 25485 -4485
rect 25540 -4605 25660 -4485
rect 25705 -4605 25825 -4485
rect 25870 -4605 25990 -4485
rect 26035 -4605 26155 -4485
rect 26210 -4605 26330 -4485
rect 26375 -4605 26495 -4485
rect 26540 -4605 26660 -4485
rect 26705 -4605 26825 -4485
rect 26880 -4605 27000 -4485
rect 27045 -4605 27165 -4485
rect 27210 -4605 27330 -4485
rect 27375 -4605 27495 -4485
rect 27550 -4605 27670 -4485
rect 27715 -4605 27835 -4485
rect 27880 -4605 28000 -4485
rect 28045 -4605 28165 -4485
rect 28220 -4605 28340 -4485
rect 28385 -4605 28505 -4485
rect 28550 -4605 28670 -4485
rect 28715 -4605 28835 -4485
rect 28890 -4605 29010 -4485
rect 29055 -4605 29175 -4485
rect 29220 -4605 29340 -4485
rect 29385 -4605 29505 -4485
rect 29560 -4605 29680 -4485
rect 24200 -4770 24320 -4650
rect 24365 -4770 24485 -4650
rect 24530 -4770 24650 -4650
rect 24695 -4770 24815 -4650
rect 24870 -4770 24990 -4650
rect 25035 -4770 25155 -4650
rect 25200 -4770 25320 -4650
rect 25365 -4770 25485 -4650
rect 25540 -4770 25660 -4650
rect 25705 -4770 25825 -4650
rect 25870 -4770 25990 -4650
rect 26035 -4770 26155 -4650
rect 26210 -4770 26330 -4650
rect 26375 -4770 26495 -4650
rect 26540 -4770 26660 -4650
rect 26705 -4770 26825 -4650
rect 26880 -4770 27000 -4650
rect 27045 -4770 27165 -4650
rect 27210 -4770 27330 -4650
rect 27375 -4770 27495 -4650
rect 27550 -4770 27670 -4650
rect 27715 -4770 27835 -4650
rect 27880 -4770 28000 -4650
rect 28045 -4770 28165 -4650
rect 28220 -4770 28340 -4650
rect 28385 -4770 28505 -4650
rect 28550 -4770 28670 -4650
rect 28715 -4770 28835 -4650
rect 28890 -4770 29010 -4650
rect 29055 -4770 29175 -4650
rect 29220 -4770 29340 -4650
rect 29385 -4770 29505 -4650
rect 29560 -4770 29680 -4650
rect 24200 -4935 24320 -4815
rect 24365 -4935 24485 -4815
rect 24530 -4935 24650 -4815
rect 24695 -4935 24815 -4815
rect 24870 -4935 24990 -4815
rect 25035 -4935 25155 -4815
rect 25200 -4935 25320 -4815
rect 25365 -4935 25485 -4815
rect 25540 -4935 25660 -4815
rect 25705 -4935 25825 -4815
rect 25870 -4935 25990 -4815
rect 26035 -4935 26155 -4815
rect 26210 -4935 26330 -4815
rect 26375 -4935 26495 -4815
rect 26540 -4935 26660 -4815
rect 26705 -4935 26825 -4815
rect 26880 -4935 27000 -4815
rect 27045 -4935 27165 -4815
rect 27210 -4935 27330 -4815
rect 27375 -4935 27495 -4815
rect 27550 -4935 27670 -4815
rect 27715 -4935 27835 -4815
rect 27880 -4935 28000 -4815
rect 28045 -4935 28165 -4815
rect 28220 -4935 28340 -4815
rect 28385 -4935 28505 -4815
rect 28550 -4935 28670 -4815
rect 28715 -4935 28835 -4815
rect 28890 -4935 29010 -4815
rect 29055 -4935 29175 -4815
rect 29220 -4935 29340 -4815
rect 29385 -4935 29505 -4815
rect 29560 -4935 29680 -4815
rect 24200 -5100 24320 -4980
rect 24365 -5100 24485 -4980
rect 24530 -5100 24650 -4980
rect 24695 -5100 24815 -4980
rect 24870 -5100 24990 -4980
rect 25035 -5100 25155 -4980
rect 25200 -5100 25320 -4980
rect 25365 -5100 25485 -4980
rect 25540 -5100 25660 -4980
rect 25705 -5100 25825 -4980
rect 25870 -5100 25990 -4980
rect 26035 -5100 26155 -4980
rect 26210 -5100 26330 -4980
rect 26375 -5100 26495 -4980
rect 26540 -5100 26660 -4980
rect 26705 -5100 26825 -4980
rect 26880 -5100 27000 -4980
rect 27045 -5100 27165 -4980
rect 27210 -5100 27330 -4980
rect 27375 -5100 27495 -4980
rect 27550 -5100 27670 -4980
rect 27715 -5100 27835 -4980
rect 27880 -5100 28000 -4980
rect 28045 -5100 28165 -4980
rect 28220 -5100 28340 -4980
rect 28385 -5100 28505 -4980
rect 28550 -5100 28670 -4980
rect 28715 -5100 28835 -4980
rect 28890 -5100 29010 -4980
rect 29055 -5100 29175 -4980
rect 29220 -5100 29340 -4980
rect 29385 -5100 29505 -4980
rect 29560 -5100 29680 -4980
rect 24200 -5275 24320 -5155
rect 24365 -5275 24485 -5155
rect 24530 -5275 24650 -5155
rect 24695 -5275 24815 -5155
rect 24870 -5275 24990 -5155
rect 25035 -5275 25155 -5155
rect 25200 -5275 25320 -5155
rect 25365 -5275 25485 -5155
rect 25540 -5275 25660 -5155
rect 25705 -5275 25825 -5155
rect 25870 -5275 25990 -5155
rect 26035 -5275 26155 -5155
rect 26210 -5275 26330 -5155
rect 26375 -5275 26495 -5155
rect 26540 -5275 26660 -5155
rect 26705 -5275 26825 -5155
rect 26880 -5275 27000 -5155
rect 27045 -5275 27165 -5155
rect 27210 -5275 27330 -5155
rect 27375 -5275 27495 -5155
rect 27550 -5275 27670 -5155
rect 27715 -5275 27835 -5155
rect 27880 -5275 28000 -5155
rect 28045 -5275 28165 -5155
rect 28220 -5275 28340 -5155
rect 28385 -5275 28505 -5155
rect 28550 -5275 28670 -5155
rect 28715 -5275 28835 -5155
rect 28890 -5275 29010 -5155
rect 29055 -5275 29175 -5155
rect 29220 -5275 29340 -5155
rect 29385 -5275 29505 -5155
rect 29560 -5275 29680 -5155
rect 24200 -5440 24320 -5320
rect 24365 -5440 24485 -5320
rect 24530 -5440 24650 -5320
rect 24695 -5440 24815 -5320
rect 24870 -5440 24990 -5320
rect 25035 -5440 25155 -5320
rect 25200 -5440 25320 -5320
rect 25365 -5440 25485 -5320
rect 25540 -5440 25660 -5320
rect 25705 -5440 25825 -5320
rect 25870 -5440 25990 -5320
rect 26035 -5440 26155 -5320
rect 26210 -5440 26330 -5320
rect 26375 -5440 26495 -5320
rect 26540 -5440 26660 -5320
rect 26705 -5440 26825 -5320
rect 26880 -5440 27000 -5320
rect 27045 -5440 27165 -5320
rect 27210 -5440 27330 -5320
rect 27375 -5440 27495 -5320
rect 27550 -5440 27670 -5320
rect 27715 -5440 27835 -5320
rect 27880 -5440 28000 -5320
rect 28045 -5440 28165 -5320
rect 28220 -5440 28340 -5320
rect 28385 -5440 28505 -5320
rect 28550 -5440 28670 -5320
rect 28715 -5440 28835 -5320
rect 28890 -5440 29010 -5320
rect 29055 -5440 29175 -5320
rect 29220 -5440 29340 -5320
rect 29385 -5440 29505 -5320
rect 29560 -5440 29680 -5320
rect 24200 -5605 24320 -5485
rect 24365 -5605 24485 -5485
rect 24530 -5605 24650 -5485
rect 24695 -5605 24815 -5485
rect 24870 -5605 24990 -5485
rect 25035 -5605 25155 -5485
rect 25200 -5605 25320 -5485
rect 25365 -5605 25485 -5485
rect 25540 -5605 25660 -5485
rect 25705 -5605 25825 -5485
rect 25870 -5605 25990 -5485
rect 26035 -5605 26155 -5485
rect 26210 -5605 26330 -5485
rect 26375 -5605 26495 -5485
rect 26540 -5605 26660 -5485
rect 26705 -5605 26825 -5485
rect 26880 -5605 27000 -5485
rect 27045 -5605 27165 -5485
rect 27210 -5605 27330 -5485
rect 27375 -5605 27495 -5485
rect 27550 -5605 27670 -5485
rect 27715 -5605 27835 -5485
rect 27880 -5605 28000 -5485
rect 28045 -5605 28165 -5485
rect 28220 -5605 28340 -5485
rect 28385 -5605 28505 -5485
rect 28550 -5605 28670 -5485
rect 28715 -5605 28835 -5485
rect 28890 -5605 29010 -5485
rect 29055 -5605 29175 -5485
rect 29220 -5605 29340 -5485
rect 29385 -5605 29505 -5485
rect 29560 -5605 29680 -5485
rect 24200 -5770 24320 -5650
rect 24365 -5770 24485 -5650
rect 24530 -5770 24650 -5650
rect 24695 -5770 24815 -5650
rect 24870 -5770 24990 -5650
rect 25035 -5770 25155 -5650
rect 25200 -5770 25320 -5650
rect 25365 -5770 25485 -5650
rect 25540 -5770 25660 -5650
rect 25705 -5770 25825 -5650
rect 25870 -5770 25990 -5650
rect 26035 -5770 26155 -5650
rect 26210 -5770 26330 -5650
rect 26375 -5770 26495 -5650
rect 26540 -5770 26660 -5650
rect 26705 -5770 26825 -5650
rect 26880 -5770 27000 -5650
rect 27045 -5770 27165 -5650
rect 27210 -5770 27330 -5650
rect 27375 -5770 27495 -5650
rect 27550 -5770 27670 -5650
rect 27715 -5770 27835 -5650
rect 27880 -5770 28000 -5650
rect 28045 -5770 28165 -5650
rect 28220 -5770 28340 -5650
rect 28385 -5770 28505 -5650
rect 28550 -5770 28670 -5650
rect 28715 -5770 28835 -5650
rect 28890 -5770 29010 -5650
rect 29055 -5770 29175 -5650
rect 29220 -5770 29340 -5650
rect 29385 -5770 29505 -5650
rect 29560 -5770 29680 -5650
rect 24200 -5945 24320 -5825
rect 24365 -5945 24485 -5825
rect 24530 -5945 24650 -5825
rect 24695 -5945 24815 -5825
rect 24870 -5945 24990 -5825
rect 25035 -5945 25155 -5825
rect 25200 -5945 25320 -5825
rect 25365 -5945 25485 -5825
rect 25540 -5945 25660 -5825
rect 25705 -5945 25825 -5825
rect 25870 -5945 25990 -5825
rect 26035 -5945 26155 -5825
rect 26210 -5945 26330 -5825
rect 26375 -5945 26495 -5825
rect 26540 -5945 26660 -5825
rect 26705 -5945 26825 -5825
rect 26880 -5945 27000 -5825
rect 27045 -5945 27165 -5825
rect 27210 -5945 27330 -5825
rect 27375 -5945 27495 -5825
rect 27550 -5945 27670 -5825
rect 27715 -5945 27835 -5825
rect 27880 -5945 28000 -5825
rect 28045 -5945 28165 -5825
rect 28220 -5945 28340 -5825
rect 28385 -5945 28505 -5825
rect 28550 -5945 28670 -5825
rect 28715 -5945 28835 -5825
rect 28890 -5945 29010 -5825
rect 29055 -5945 29175 -5825
rect 29220 -5945 29340 -5825
rect 29385 -5945 29505 -5825
rect 29560 -5945 29680 -5825
rect 24200 -6110 24320 -5990
rect 24365 -6110 24485 -5990
rect 24530 -6110 24650 -5990
rect 24695 -6110 24815 -5990
rect 24870 -6110 24990 -5990
rect 25035 -6110 25155 -5990
rect 25200 -6110 25320 -5990
rect 25365 -6110 25485 -5990
rect 25540 -6110 25660 -5990
rect 25705 -6110 25825 -5990
rect 25870 -6110 25990 -5990
rect 26035 -6110 26155 -5990
rect 26210 -6110 26330 -5990
rect 26375 -6110 26495 -5990
rect 26540 -6110 26660 -5990
rect 26705 -6110 26825 -5990
rect 26880 -6110 27000 -5990
rect 27045 -6110 27165 -5990
rect 27210 -6110 27330 -5990
rect 27375 -6110 27495 -5990
rect 27550 -6110 27670 -5990
rect 27715 -6110 27835 -5990
rect 27880 -6110 28000 -5990
rect 28045 -6110 28165 -5990
rect 28220 -6110 28340 -5990
rect 28385 -6110 28505 -5990
rect 28550 -6110 28670 -5990
rect 28715 -6110 28835 -5990
rect 28890 -6110 29010 -5990
rect 29055 -6110 29175 -5990
rect 29220 -6110 29340 -5990
rect 29385 -6110 29505 -5990
rect 29560 -6110 29680 -5990
rect 24200 -6275 24320 -6155
rect 24365 -6275 24485 -6155
rect 24530 -6275 24650 -6155
rect 24695 -6275 24815 -6155
rect 24870 -6275 24990 -6155
rect 25035 -6275 25155 -6155
rect 25200 -6275 25320 -6155
rect 25365 -6275 25485 -6155
rect 25540 -6275 25660 -6155
rect 25705 -6275 25825 -6155
rect 25870 -6275 25990 -6155
rect 26035 -6275 26155 -6155
rect 26210 -6275 26330 -6155
rect 26375 -6275 26495 -6155
rect 26540 -6275 26660 -6155
rect 26705 -6275 26825 -6155
rect 26880 -6275 27000 -6155
rect 27045 -6275 27165 -6155
rect 27210 -6275 27330 -6155
rect 27375 -6275 27495 -6155
rect 27550 -6275 27670 -6155
rect 27715 -6275 27835 -6155
rect 27880 -6275 28000 -6155
rect 28045 -6275 28165 -6155
rect 28220 -6275 28340 -6155
rect 28385 -6275 28505 -6155
rect 28550 -6275 28670 -6155
rect 28715 -6275 28835 -6155
rect 28890 -6275 29010 -6155
rect 29055 -6275 29175 -6155
rect 29220 -6275 29340 -6155
rect 29385 -6275 29505 -6155
rect 29560 -6275 29680 -6155
rect 24200 -6440 24320 -6320
rect 24365 -6440 24485 -6320
rect 24530 -6440 24650 -6320
rect 24695 -6440 24815 -6320
rect 24870 -6440 24990 -6320
rect 25035 -6440 25155 -6320
rect 25200 -6440 25320 -6320
rect 25365 -6440 25485 -6320
rect 25540 -6440 25660 -6320
rect 25705 -6440 25825 -6320
rect 25870 -6440 25990 -6320
rect 26035 -6440 26155 -6320
rect 26210 -6440 26330 -6320
rect 26375 -6440 26495 -6320
rect 26540 -6440 26660 -6320
rect 26705 -6440 26825 -6320
rect 26880 -6440 27000 -6320
rect 27045 -6440 27165 -6320
rect 27210 -6440 27330 -6320
rect 27375 -6440 27495 -6320
rect 27550 -6440 27670 -6320
rect 27715 -6440 27835 -6320
rect 27880 -6440 28000 -6320
rect 28045 -6440 28165 -6320
rect 28220 -6440 28340 -6320
rect 28385 -6440 28505 -6320
rect 28550 -6440 28670 -6320
rect 28715 -6440 28835 -6320
rect 28890 -6440 29010 -6320
rect 29055 -6440 29175 -6320
rect 29220 -6440 29340 -6320
rect 29385 -6440 29505 -6320
rect 29560 -6440 29680 -6320
rect 24200 -6615 24320 -6495
rect 24365 -6615 24485 -6495
rect 24530 -6615 24650 -6495
rect 24695 -6615 24815 -6495
rect 24870 -6615 24990 -6495
rect 25035 -6615 25155 -6495
rect 25200 -6615 25320 -6495
rect 25365 -6615 25485 -6495
rect 25540 -6615 25660 -6495
rect 25705 -6615 25825 -6495
rect 25870 -6615 25990 -6495
rect 26035 -6615 26155 -6495
rect 26210 -6615 26330 -6495
rect 26375 -6615 26495 -6495
rect 26540 -6615 26660 -6495
rect 26705 -6615 26825 -6495
rect 26880 -6615 27000 -6495
rect 27045 -6615 27165 -6495
rect 27210 -6615 27330 -6495
rect 27375 -6615 27495 -6495
rect 27550 -6615 27670 -6495
rect 27715 -6615 27835 -6495
rect 27880 -6615 28000 -6495
rect 28045 -6615 28165 -6495
rect 28220 -6615 28340 -6495
rect 28385 -6615 28505 -6495
rect 28550 -6615 28670 -6495
rect 28715 -6615 28835 -6495
rect 28890 -6615 29010 -6495
rect 29055 -6615 29175 -6495
rect 29220 -6615 29340 -6495
rect 29385 -6615 29505 -6495
rect 29560 -6615 29680 -6495
rect 24200 -6780 24320 -6660
rect 24365 -6780 24485 -6660
rect 24530 -6780 24650 -6660
rect 24695 -6780 24815 -6660
rect 24870 -6780 24990 -6660
rect 25035 -6780 25155 -6660
rect 25200 -6780 25320 -6660
rect 25365 -6780 25485 -6660
rect 25540 -6780 25660 -6660
rect 25705 -6780 25825 -6660
rect 25870 -6780 25990 -6660
rect 26035 -6780 26155 -6660
rect 26210 -6780 26330 -6660
rect 26375 -6780 26495 -6660
rect 26540 -6780 26660 -6660
rect 26705 -6780 26825 -6660
rect 26880 -6780 27000 -6660
rect 27045 -6780 27165 -6660
rect 27210 -6780 27330 -6660
rect 27375 -6780 27495 -6660
rect 27550 -6780 27670 -6660
rect 27715 -6780 27835 -6660
rect 27880 -6780 28000 -6660
rect 28045 -6780 28165 -6660
rect 28220 -6780 28340 -6660
rect 28385 -6780 28505 -6660
rect 28550 -6780 28670 -6660
rect 28715 -6780 28835 -6660
rect 28890 -6780 29010 -6660
rect 29055 -6780 29175 -6660
rect 29220 -6780 29340 -6660
rect 29385 -6780 29505 -6660
rect 29560 -6780 29680 -6660
rect 24200 -6945 24320 -6825
rect 24365 -6945 24485 -6825
rect 24530 -6945 24650 -6825
rect 24695 -6945 24815 -6825
rect 24870 -6945 24990 -6825
rect 25035 -6945 25155 -6825
rect 25200 -6945 25320 -6825
rect 25365 -6945 25485 -6825
rect 25540 -6945 25660 -6825
rect 25705 -6945 25825 -6825
rect 25870 -6945 25990 -6825
rect 26035 -6945 26155 -6825
rect 26210 -6945 26330 -6825
rect 26375 -6945 26495 -6825
rect 26540 -6945 26660 -6825
rect 26705 -6945 26825 -6825
rect 26880 -6945 27000 -6825
rect 27045 -6945 27165 -6825
rect 27210 -6945 27330 -6825
rect 27375 -6945 27495 -6825
rect 27550 -6945 27670 -6825
rect 27715 -6945 27835 -6825
rect 27880 -6945 28000 -6825
rect 28045 -6945 28165 -6825
rect 28220 -6945 28340 -6825
rect 28385 -6945 28505 -6825
rect 28550 -6945 28670 -6825
rect 28715 -6945 28835 -6825
rect 28890 -6945 29010 -6825
rect 29055 -6945 29175 -6825
rect 29220 -6945 29340 -6825
rect 29385 -6945 29505 -6825
rect 29560 -6945 29680 -6825
rect 24200 -7110 24320 -6990
rect 24365 -7110 24485 -6990
rect 24530 -7110 24650 -6990
rect 24695 -7110 24815 -6990
rect 24870 -7110 24990 -6990
rect 25035 -7110 25155 -6990
rect 25200 -7110 25320 -6990
rect 25365 -7110 25485 -6990
rect 25540 -7110 25660 -6990
rect 25705 -7110 25825 -6990
rect 25870 -7110 25990 -6990
rect 26035 -7110 26155 -6990
rect 26210 -7110 26330 -6990
rect 26375 -7110 26495 -6990
rect 26540 -7110 26660 -6990
rect 26705 -7110 26825 -6990
rect 26880 -7110 27000 -6990
rect 27045 -7110 27165 -6990
rect 27210 -7110 27330 -6990
rect 27375 -7110 27495 -6990
rect 27550 -7110 27670 -6990
rect 27715 -7110 27835 -6990
rect 27880 -7110 28000 -6990
rect 28045 -7110 28165 -6990
rect 28220 -7110 28340 -6990
rect 28385 -7110 28505 -6990
rect 28550 -7110 28670 -6990
rect 28715 -7110 28835 -6990
rect 28890 -7110 29010 -6990
rect 29055 -7110 29175 -6990
rect 29220 -7110 29340 -6990
rect 29385 -7110 29505 -6990
rect 29560 -7110 29680 -6990
rect 24200 -7285 24320 -7165
rect 24365 -7285 24485 -7165
rect 24530 -7285 24650 -7165
rect 24695 -7285 24815 -7165
rect 24870 -7285 24990 -7165
rect 25035 -7285 25155 -7165
rect 25200 -7285 25320 -7165
rect 25365 -7285 25485 -7165
rect 25540 -7285 25660 -7165
rect 25705 -7285 25825 -7165
rect 25870 -7285 25990 -7165
rect 26035 -7285 26155 -7165
rect 26210 -7285 26330 -7165
rect 26375 -7285 26495 -7165
rect 26540 -7285 26660 -7165
rect 26705 -7285 26825 -7165
rect 26880 -7285 27000 -7165
rect 27045 -7285 27165 -7165
rect 27210 -7285 27330 -7165
rect 27375 -7285 27495 -7165
rect 27550 -7285 27670 -7165
rect 27715 -7285 27835 -7165
rect 27880 -7285 28000 -7165
rect 28045 -7285 28165 -7165
rect 28220 -7285 28340 -7165
rect 28385 -7285 28505 -7165
rect 28550 -7285 28670 -7165
rect 28715 -7285 28835 -7165
rect 28890 -7285 29010 -7165
rect 29055 -7285 29175 -7165
rect 29220 -7285 29340 -7165
rect 29385 -7285 29505 -7165
rect 29560 -7285 29680 -7165
rect 24200 -7450 24320 -7330
rect 24365 -7450 24485 -7330
rect 24530 -7450 24650 -7330
rect 24695 -7450 24815 -7330
rect 24870 -7450 24990 -7330
rect 25035 -7450 25155 -7330
rect 25200 -7450 25320 -7330
rect 25365 -7450 25485 -7330
rect 25540 -7450 25660 -7330
rect 25705 -7450 25825 -7330
rect 25870 -7450 25990 -7330
rect 26035 -7450 26155 -7330
rect 26210 -7450 26330 -7330
rect 26375 -7450 26495 -7330
rect 26540 -7450 26660 -7330
rect 26705 -7450 26825 -7330
rect 26880 -7450 27000 -7330
rect 27045 -7450 27165 -7330
rect 27210 -7450 27330 -7330
rect 27375 -7450 27495 -7330
rect 27550 -7450 27670 -7330
rect 27715 -7450 27835 -7330
rect 27880 -7450 28000 -7330
rect 28045 -7450 28165 -7330
rect 28220 -7450 28340 -7330
rect 28385 -7450 28505 -7330
rect 28550 -7450 28670 -7330
rect 28715 -7450 28835 -7330
rect 28890 -7450 29010 -7330
rect 29055 -7450 29175 -7330
rect 29220 -7450 29340 -7330
rect 29385 -7450 29505 -7330
rect 29560 -7450 29680 -7330
rect 24200 -7615 24320 -7495
rect 24365 -7615 24485 -7495
rect 24530 -7615 24650 -7495
rect 24695 -7615 24815 -7495
rect 24870 -7615 24990 -7495
rect 25035 -7615 25155 -7495
rect 25200 -7615 25320 -7495
rect 25365 -7615 25485 -7495
rect 25540 -7615 25660 -7495
rect 25705 -7615 25825 -7495
rect 25870 -7615 25990 -7495
rect 26035 -7615 26155 -7495
rect 26210 -7615 26330 -7495
rect 26375 -7615 26495 -7495
rect 26540 -7615 26660 -7495
rect 26705 -7615 26825 -7495
rect 26880 -7615 27000 -7495
rect 27045 -7615 27165 -7495
rect 27210 -7615 27330 -7495
rect 27375 -7615 27495 -7495
rect 27550 -7615 27670 -7495
rect 27715 -7615 27835 -7495
rect 27880 -7615 28000 -7495
rect 28045 -7615 28165 -7495
rect 28220 -7615 28340 -7495
rect 28385 -7615 28505 -7495
rect 28550 -7615 28670 -7495
rect 28715 -7615 28835 -7495
rect 28890 -7615 29010 -7495
rect 29055 -7615 29175 -7495
rect 29220 -7615 29340 -7495
rect 29385 -7615 29505 -7495
rect 29560 -7615 29680 -7495
rect 24200 -7780 24320 -7660
rect 24365 -7780 24485 -7660
rect 24530 -7780 24650 -7660
rect 24695 -7780 24815 -7660
rect 24870 -7780 24990 -7660
rect 25035 -7780 25155 -7660
rect 25200 -7780 25320 -7660
rect 25365 -7780 25485 -7660
rect 25540 -7780 25660 -7660
rect 25705 -7780 25825 -7660
rect 25870 -7780 25990 -7660
rect 26035 -7780 26155 -7660
rect 26210 -7780 26330 -7660
rect 26375 -7780 26495 -7660
rect 26540 -7780 26660 -7660
rect 26705 -7780 26825 -7660
rect 26880 -7780 27000 -7660
rect 27045 -7780 27165 -7660
rect 27210 -7780 27330 -7660
rect 27375 -7780 27495 -7660
rect 27550 -7780 27670 -7660
rect 27715 -7780 27835 -7660
rect 27880 -7780 28000 -7660
rect 28045 -7780 28165 -7660
rect 28220 -7780 28340 -7660
rect 28385 -7780 28505 -7660
rect 28550 -7780 28670 -7660
rect 28715 -7780 28835 -7660
rect 28890 -7780 29010 -7660
rect 29055 -7780 29175 -7660
rect 29220 -7780 29340 -7660
rect 29385 -7780 29505 -7660
rect 29560 -7780 29680 -7660
rect 24200 -7955 24320 -7835
rect 24365 -7955 24485 -7835
rect 24530 -7955 24650 -7835
rect 24695 -7955 24815 -7835
rect 24870 -7955 24990 -7835
rect 25035 -7955 25155 -7835
rect 25200 -7955 25320 -7835
rect 25365 -7955 25485 -7835
rect 25540 -7955 25660 -7835
rect 25705 -7955 25825 -7835
rect 25870 -7955 25990 -7835
rect 26035 -7955 26155 -7835
rect 26210 -7955 26330 -7835
rect 26375 -7955 26495 -7835
rect 26540 -7955 26660 -7835
rect 26705 -7955 26825 -7835
rect 26880 -7955 27000 -7835
rect 27045 -7955 27165 -7835
rect 27210 -7955 27330 -7835
rect 27375 -7955 27495 -7835
rect 27550 -7955 27670 -7835
rect 27715 -7955 27835 -7835
rect 27880 -7955 28000 -7835
rect 28045 -7955 28165 -7835
rect 28220 -7955 28340 -7835
rect 28385 -7955 28505 -7835
rect 28550 -7955 28670 -7835
rect 28715 -7955 28835 -7835
rect 28890 -7955 29010 -7835
rect 29055 -7955 29175 -7835
rect 29220 -7955 29340 -7835
rect 29385 -7955 29505 -7835
rect 29560 -7955 29680 -7835
rect 24200 -8120 24320 -8000
rect 24365 -8120 24485 -8000
rect 24530 -8120 24650 -8000
rect 24695 -8120 24815 -8000
rect 24870 -8120 24990 -8000
rect 25035 -8120 25155 -8000
rect 25200 -8120 25320 -8000
rect 25365 -8120 25485 -8000
rect 25540 -8120 25660 -8000
rect 25705 -8120 25825 -8000
rect 25870 -8120 25990 -8000
rect 26035 -8120 26155 -8000
rect 26210 -8120 26330 -8000
rect 26375 -8120 26495 -8000
rect 26540 -8120 26660 -8000
rect 26705 -8120 26825 -8000
rect 26880 -8120 27000 -8000
rect 27045 -8120 27165 -8000
rect 27210 -8120 27330 -8000
rect 27375 -8120 27495 -8000
rect 27550 -8120 27670 -8000
rect 27715 -8120 27835 -8000
rect 27880 -8120 28000 -8000
rect 28045 -8120 28165 -8000
rect 28220 -8120 28340 -8000
rect 28385 -8120 28505 -8000
rect 28550 -8120 28670 -8000
rect 28715 -8120 28835 -8000
rect 28890 -8120 29010 -8000
rect 29055 -8120 29175 -8000
rect 29220 -8120 29340 -8000
rect 29385 -8120 29505 -8000
rect 29560 -8120 29680 -8000
rect 24200 -8285 24320 -8165
rect 24365 -8285 24485 -8165
rect 24530 -8285 24650 -8165
rect 24695 -8285 24815 -8165
rect 24870 -8285 24990 -8165
rect 25035 -8285 25155 -8165
rect 25200 -8285 25320 -8165
rect 25365 -8285 25485 -8165
rect 25540 -8285 25660 -8165
rect 25705 -8285 25825 -8165
rect 25870 -8285 25990 -8165
rect 26035 -8285 26155 -8165
rect 26210 -8285 26330 -8165
rect 26375 -8285 26495 -8165
rect 26540 -8285 26660 -8165
rect 26705 -8285 26825 -8165
rect 26880 -8285 27000 -8165
rect 27045 -8285 27165 -8165
rect 27210 -8285 27330 -8165
rect 27375 -8285 27495 -8165
rect 27550 -8285 27670 -8165
rect 27715 -8285 27835 -8165
rect 27880 -8285 28000 -8165
rect 28045 -8285 28165 -8165
rect 28220 -8285 28340 -8165
rect 28385 -8285 28505 -8165
rect 28550 -8285 28670 -8165
rect 28715 -8285 28835 -8165
rect 28890 -8285 29010 -8165
rect 29055 -8285 29175 -8165
rect 29220 -8285 29340 -8165
rect 29385 -8285 29505 -8165
rect 29560 -8285 29680 -8165
rect 24200 -8450 24320 -8330
rect 24365 -8450 24485 -8330
rect 24530 -8450 24650 -8330
rect 24695 -8450 24815 -8330
rect 24870 -8450 24990 -8330
rect 25035 -8450 25155 -8330
rect 25200 -8450 25320 -8330
rect 25365 -8450 25485 -8330
rect 25540 -8450 25660 -8330
rect 25705 -8450 25825 -8330
rect 25870 -8450 25990 -8330
rect 26035 -8450 26155 -8330
rect 26210 -8450 26330 -8330
rect 26375 -8450 26495 -8330
rect 26540 -8450 26660 -8330
rect 26705 -8450 26825 -8330
rect 26880 -8450 27000 -8330
rect 27045 -8450 27165 -8330
rect 27210 -8450 27330 -8330
rect 27375 -8450 27495 -8330
rect 27550 -8450 27670 -8330
rect 27715 -8450 27835 -8330
rect 27880 -8450 28000 -8330
rect 28045 -8450 28165 -8330
rect 28220 -8450 28340 -8330
rect 28385 -8450 28505 -8330
rect 28550 -8450 28670 -8330
rect 28715 -8450 28835 -8330
rect 28890 -8450 29010 -8330
rect 29055 -8450 29175 -8330
rect 29220 -8450 29340 -8330
rect 29385 -8450 29505 -8330
rect 29560 -8450 29680 -8330
rect 24200 -8625 24320 -8505
rect 24365 -8625 24485 -8505
rect 24530 -8625 24650 -8505
rect 24695 -8625 24815 -8505
rect 24870 -8625 24990 -8505
rect 25035 -8625 25155 -8505
rect 25200 -8625 25320 -8505
rect 25365 -8625 25485 -8505
rect 25540 -8625 25660 -8505
rect 25705 -8625 25825 -8505
rect 25870 -8625 25990 -8505
rect 26035 -8625 26155 -8505
rect 26210 -8625 26330 -8505
rect 26375 -8625 26495 -8505
rect 26540 -8625 26660 -8505
rect 26705 -8625 26825 -8505
rect 26880 -8625 27000 -8505
rect 27045 -8625 27165 -8505
rect 27210 -8625 27330 -8505
rect 27375 -8625 27495 -8505
rect 27550 -8625 27670 -8505
rect 27715 -8625 27835 -8505
rect 27880 -8625 28000 -8505
rect 28045 -8625 28165 -8505
rect 28220 -8625 28340 -8505
rect 28385 -8625 28505 -8505
rect 28550 -8625 28670 -8505
rect 28715 -8625 28835 -8505
rect 28890 -8625 29010 -8505
rect 29055 -8625 29175 -8505
rect 29220 -8625 29340 -8505
rect 29385 -8625 29505 -8505
rect 29560 -8625 29680 -8505
rect 24200 -8790 24320 -8670
rect 24365 -8790 24485 -8670
rect 24530 -8790 24650 -8670
rect 24695 -8790 24815 -8670
rect 24870 -8790 24990 -8670
rect 25035 -8790 25155 -8670
rect 25200 -8790 25320 -8670
rect 25365 -8790 25485 -8670
rect 25540 -8790 25660 -8670
rect 25705 -8790 25825 -8670
rect 25870 -8790 25990 -8670
rect 26035 -8790 26155 -8670
rect 26210 -8790 26330 -8670
rect 26375 -8790 26495 -8670
rect 26540 -8790 26660 -8670
rect 26705 -8790 26825 -8670
rect 26880 -8790 27000 -8670
rect 27045 -8790 27165 -8670
rect 27210 -8790 27330 -8670
rect 27375 -8790 27495 -8670
rect 27550 -8790 27670 -8670
rect 27715 -8790 27835 -8670
rect 27880 -8790 28000 -8670
rect 28045 -8790 28165 -8670
rect 28220 -8790 28340 -8670
rect 28385 -8790 28505 -8670
rect 28550 -8790 28670 -8670
rect 28715 -8790 28835 -8670
rect 28890 -8790 29010 -8670
rect 29055 -8790 29175 -8670
rect 29220 -8790 29340 -8670
rect 29385 -8790 29505 -8670
rect 29560 -8790 29680 -8670
rect 24200 -8955 24320 -8835
rect 24365 -8955 24485 -8835
rect 24530 -8955 24650 -8835
rect 24695 -8955 24815 -8835
rect 24870 -8955 24990 -8835
rect 25035 -8955 25155 -8835
rect 25200 -8955 25320 -8835
rect 25365 -8955 25485 -8835
rect 25540 -8955 25660 -8835
rect 25705 -8955 25825 -8835
rect 25870 -8955 25990 -8835
rect 26035 -8955 26155 -8835
rect 26210 -8955 26330 -8835
rect 26375 -8955 26495 -8835
rect 26540 -8955 26660 -8835
rect 26705 -8955 26825 -8835
rect 26880 -8955 27000 -8835
rect 27045 -8955 27165 -8835
rect 27210 -8955 27330 -8835
rect 27375 -8955 27495 -8835
rect 27550 -8955 27670 -8835
rect 27715 -8955 27835 -8835
rect 27880 -8955 28000 -8835
rect 28045 -8955 28165 -8835
rect 28220 -8955 28340 -8835
rect 28385 -8955 28505 -8835
rect 28550 -8955 28670 -8835
rect 28715 -8955 28835 -8835
rect 28890 -8955 29010 -8835
rect 29055 -8955 29175 -8835
rect 29220 -8955 29340 -8835
rect 29385 -8955 29505 -8835
rect 29560 -8955 29680 -8835
rect 24200 -9120 24320 -9000
rect 24365 -9120 24485 -9000
rect 24530 -9120 24650 -9000
rect 24695 -9120 24815 -9000
rect 24870 -9120 24990 -9000
rect 25035 -9120 25155 -9000
rect 25200 -9120 25320 -9000
rect 25365 -9120 25485 -9000
rect 25540 -9120 25660 -9000
rect 25705 -9120 25825 -9000
rect 25870 -9120 25990 -9000
rect 26035 -9120 26155 -9000
rect 26210 -9120 26330 -9000
rect 26375 -9120 26495 -9000
rect 26540 -9120 26660 -9000
rect 26705 -9120 26825 -9000
rect 26880 -9120 27000 -9000
rect 27045 -9120 27165 -9000
rect 27210 -9120 27330 -9000
rect 27375 -9120 27495 -9000
rect 27550 -9120 27670 -9000
rect 27715 -9120 27835 -9000
rect 27880 -9120 28000 -9000
rect 28045 -9120 28165 -9000
rect 28220 -9120 28340 -9000
rect 28385 -9120 28505 -9000
rect 28550 -9120 28670 -9000
rect 28715 -9120 28835 -9000
rect 28890 -9120 29010 -9000
rect 29055 -9120 29175 -9000
rect 29220 -9120 29340 -9000
rect 29385 -9120 29505 -9000
rect 29560 -9120 29680 -9000
rect 24200 -9295 24320 -9175
rect 24365 -9295 24485 -9175
rect 24530 -9295 24650 -9175
rect 24695 -9295 24815 -9175
rect 24870 -9295 24990 -9175
rect 25035 -9295 25155 -9175
rect 25200 -9295 25320 -9175
rect 25365 -9295 25485 -9175
rect 25540 -9295 25660 -9175
rect 25705 -9295 25825 -9175
rect 25870 -9295 25990 -9175
rect 26035 -9295 26155 -9175
rect 26210 -9295 26330 -9175
rect 26375 -9295 26495 -9175
rect 26540 -9295 26660 -9175
rect 26705 -9295 26825 -9175
rect 26880 -9295 27000 -9175
rect 27045 -9295 27165 -9175
rect 27210 -9295 27330 -9175
rect 27375 -9295 27495 -9175
rect 27550 -9295 27670 -9175
rect 27715 -9295 27835 -9175
rect 27880 -9295 28000 -9175
rect 28045 -9295 28165 -9175
rect 28220 -9295 28340 -9175
rect 28385 -9295 28505 -9175
rect 28550 -9295 28670 -9175
rect 28715 -9295 28835 -9175
rect 28890 -9295 29010 -9175
rect 29055 -9295 29175 -9175
rect 29220 -9295 29340 -9175
rect 29385 -9295 29505 -9175
rect 29560 -9295 29680 -9175
rect 24200 -9460 24320 -9340
rect 24365 -9460 24485 -9340
rect 24530 -9460 24650 -9340
rect 24695 -9460 24815 -9340
rect 24870 -9460 24990 -9340
rect 25035 -9460 25155 -9340
rect 25200 -9460 25320 -9340
rect 25365 -9460 25485 -9340
rect 25540 -9460 25660 -9340
rect 25705 -9460 25825 -9340
rect 25870 -9460 25990 -9340
rect 26035 -9460 26155 -9340
rect 26210 -9460 26330 -9340
rect 26375 -9460 26495 -9340
rect 26540 -9460 26660 -9340
rect 26705 -9460 26825 -9340
rect 26880 -9460 27000 -9340
rect 27045 -9460 27165 -9340
rect 27210 -9460 27330 -9340
rect 27375 -9460 27495 -9340
rect 27550 -9460 27670 -9340
rect 27715 -9460 27835 -9340
rect 27880 -9460 28000 -9340
rect 28045 -9460 28165 -9340
rect 28220 -9460 28340 -9340
rect 28385 -9460 28505 -9340
rect 28550 -9460 28670 -9340
rect 28715 -9460 28835 -9340
rect 28890 -9460 29010 -9340
rect 29055 -9460 29175 -9340
rect 29220 -9460 29340 -9340
rect 29385 -9460 29505 -9340
rect 29560 -9460 29680 -9340
rect 24200 -9625 24320 -9505
rect 24365 -9625 24485 -9505
rect 24530 -9625 24650 -9505
rect 24695 -9625 24815 -9505
rect 24870 -9625 24990 -9505
rect 25035 -9625 25155 -9505
rect 25200 -9625 25320 -9505
rect 25365 -9625 25485 -9505
rect 25540 -9625 25660 -9505
rect 25705 -9625 25825 -9505
rect 25870 -9625 25990 -9505
rect 26035 -9625 26155 -9505
rect 26210 -9625 26330 -9505
rect 26375 -9625 26495 -9505
rect 26540 -9625 26660 -9505
rect 26705 -9625 26825 -9505
rect 26880 -9625 27000 -9505
rect 27045 -9625 27165 -9505
rect 27210 -9625 27330 -9505
rect 27375 -9625 27495 -9505
rect 27550 -9625 27670 -9505
rect 27715 -9625 27835 -9505
rect 27880 -9625 28000 -9505
rect 28045 -9625 28165 -9505
rect 28220 -9625 28340 -9505
rect 28385 -9625 28505 -9505
rect 28550 -9625 28670 -9505
rect 28715 -9625 28835 -9505
rect 28890 -9625 29010 -9505
rect 29055 -9625 29175 -9505
rect 29220 -9625 29340 -9505
rect 29385 -9625 29505 -9505
rect 29560 -9625 29680 -9505
rect 24200 -9790 24320 -9670
rect 24365 -9790 24485 -9670
rect 24530 -9790 24650 -9670
rect 24695 -9790 24815 -9670
rect 24870 -9790 24990 -9670
rect 25035 -9790 25155 -9670
rect 25200 -9790 25320 -9670
rect 25365 -9790 25485 -9670
rect 25540 -9790 25660 -9670
rect 25705 -9790 25825 -9670
rect 25870 -9790 25990 -9670
rect 26035 -9790 26155 -9670
rect 26210 -9790 26330 -9670
rect 26375 -9790 26495 -9670
rect 26540 -9790 26660 -9670
rect 26705 -9790 26825 -9670
rect 26880 -9790 27000 -9670
rect 27045 -9790 27165 -9670
rect 27210 -9790 27330 -9670
rect 27375 -9790 27495 -9670
rect 27550 -9790 27670 -9670
rect 27715 -9790 27835 -9670
rect 27880 -9790 28000 -9670
rect 28045 -9790 28165 -9670
rect 28220 -9790 28340 -9670
rect 28385 -9790 28505 -9670
rect 28550 -9790 28670 -9670
rect 28715 -9790 28835 -9670
rect 28890 -9790 29010 -9670
rect 29055 -9790 29175 -9670
rect 29220 -9790 29340 -9670
rect 29385 -9790 29505 -9670
rect 29560 -9790 29680 -9670
rect 7130 -10210 7250 -10090
rect 7305 -10210 7425 -10090
rect 7470 -10210 7590 -10090
rect 7635 -10210 7755 -10090
rect 7800 -10210 7920 -10090
rect 7975 -10210 8095 -10090
rect 8140 -10210 8260 -10090
rect 8305 -10210 8425 -10090
rect 8470 -10210 8590 -10090
rect 8645 -10210 8765 -10090
rect 8810 -10210 8930 -10090
rect 8975 -10210 9095 -10090
rect 9140 -10210 9260 -10090
rect 9315 -10210 9435 -10090
rect 9480 -10210 9600 -10090
rect 9645 -10210 9765 -10090
rect 9810 -10210 9930 -10090
rect 9985 -10210 10105 -10090
rect 10150 -10210 10270 -10090
rect 10315 -10210 10435 -10090
rect 10480 -10210 10600 -10090
rect 10655 -10210 10775 -10090
rect 10820 -10210 10940 -10090
rect 10985 -10210 11105 -10090
rect 11150 -10210 11270 -10090
rect 11325 -10210 11445 -10090
rect 11490 -10210 11610 -10090
rect 11655 -10210 11775 -10090
rect 11820 -10210 11940 -10090
rect 11995 -10210 12115 -10090
rect 12160 -10210 12280 -10090
rect 12325 -10210 12445 -10090
rect 12490 -10210 12610 -10090
rect 7130 -10375 7250 -10255
rect 7305 -10375 7425 -10255
rect 7470 -10375 7590 -10255
rect 7635 -10375 7755 -10255
rect 7800 -10375 7920 -10255
rect 7975 -10375 8095 -10255
rect 8140 -10375 8260 -10255
rect 8305 -10375 8425 -10255
rect 8470 -10375 8590 -10255
rect 8645 -10375 8765 -10255
rect 8810 -10375 8930 -10255
rect 8975 -10375 9095 -10255
rect 9140 -10375 9260 -10255
rect 9315 -10375 9435 -10255
rect 9480 -10375 9600 -10255
rect 9645 -10375 9765 -10255
rect 9810 -10375 9930 -10255
rect 9985 -10375 10105 -10255
rect 10150 -10375 10270 -10255
rect 10315 -10375 10435 -10255
rect 10480 -10375 10600 -10255
rect 10655 -10375 10775 -10255
rect 10820 -10375 10940 -10255
rect 10985 -10375 11105 -10255
rect 11150 -10375 11270 -10255
rect 11325 -10375 11445 -10255
rect 11490 -10375 11610 -10255
rect 11655 -10375 11775 -10255
rect 11820 -10375 11940 -10255
rect 11995 -10375 12115 -10255
rect 12160 -10375 12280 -10255
rect 12325 -10375 12445 -10255
rect 12490 -10375 12610 -10255
rect 7130 -10540 7250 -10420
rect 7305 -10540 7425 -10420
rect 7470 -10540 7590 -10420
rect 7635 -10540 7755 -10420
rect 7800 -10540 7920 -10420
rect 7975 -10540 8095 -10420
rect 8140 -10540 8260 -10420
rect 8305 -10540 8425 -10420
rect 8470 -10540 8590 -10420
rect 8645 -10540 8765 -10420
rect 8810 -10540 8930 -10420
rect 8975 -10540 9095 -10420
rect 9140 -10540 9260 -10420
rect 9315 -10540 9435 -10420
rect 9480 -10540 9600 -10420
rect 9645 -10540 9765 -10420
rect 9810 -10540 9930 -10420
rect 9985 -10540 10105 -10420
rect 10150 -10540 10270 -10420
rect 10315 -10540 10435 -10420
rect 10480 -10540 10600 -10420
rect 10655 -10540 10775 -10420
rect 10820 -10540 10940 -10420
rect 10985 -10540 11105 -10420
rect 11150 -10540 11270 -10420
rect 11325 -10540 11445 -10420
rect 11490 -10540 11610 -10420
rect 11655 -10540 11775 -10420
rect 11820 -10540 11940 -10420
rect 11995 -10540 12115 -10420
rect 12160 -10540 12280 -10420
rect 12325 -10540 12445 -10420
rect 12490 -10540 12610 -10420
rect 7130 -10705 7250 -10585
rect 7305 -10705 7425 -10585
rect 7470 -10705 7590 -10585
rect 7635 -10705 7755 -10585
rect 7800 -10705 7920 -10585
rect 7975 -10705 8095 -10585
rect 8140 -10705 8260 -10585
rect 8305 -10705 8425 -10585
rect 8470 -10705 8590 -10585
rect 8645 -10705 8765 -10585
rect 8810 -10705 8930 -10585
rect 8975 -10705 9095 -10585
rect 9140 -10705 9260 -10585
rect 9315 -10705 9435 -10585
rect 9480 -10705 9600 -10585
rect 9645 -10705 9765 -10585
rect 9810 -10705 9930 -10585
rect 9985 -10705 10105 -10585
rect 10150 -10705 10270 -10585
rect 10315 -10705 10435 -10585
rect 10480 -10705 10600 -10585
rect 10655 -10705 10775 -10585
rect 10820 -10705 10940 -10585
rect 10985 -10705 11105 -10585
rect 11150 -10705 11270 -10585
rect 11325 -10705 11445 -10585
rect 11490 -10705 11610 -10585
rect 11655 -10705 11775 -10585
rect 11820 -10705 11940 -10585
rect 11995 -10705 12115 -10585
rect 12160 -10705 12280 -10585
rect 12325 -10705 12445 -10585
rect 12490 -10705 12610 -10585
rect 7130 -10880 7250 -10760
rect 7305 -10880 7425 -10760
rect 7470 -10880 7590 -10760
rect 7635 -10880 7755 -10760
rect 7800 -10880 7920 -10760
rect 7975 -10880 8095 -10760
rect 8140 -10880 8260 -10760
rect 8305 -10880 8425 -10760
rect 8470 -10880 8590 -10760
rect 8645 -10880 8765 -10760
rect 8810 -10880 8930 -10760
rect 8975 -10880 9095 -10760
rect 9140 -10880 9260 -10760
rect 9315 -10880 9435 -10760
rect 9480 -10880 9600 -10760
rect 9645 -10880 9765 -10760
rect 9810 -10880 9930 -10760
rect 9985 -10880 10105 -10760
rect 10150 -10880 10270 -10760
rect 10315 -10880 10435 -10760
rect 10480 -10880 10600 -10760
rect 10655 -10880 10775 -10760
rect 10820 -10880 10940 -10760
rect 10985 -10880 11105 -10760
rect 11150 -10880 11270 -10760
rect 11325 -10880 11445 -10760
rect 11490 -10880 11610 -10760
rect 11655 -10880 11775 -10760
rect 11820 -10880 11940 -10760
rect 11995 -10880 12115 -10760
rect 12160 -10880 12280 -10760
rect 12325 -10880 12445 -10760
rect 12490 -10880 12610 -10760
rect 7130 -11045 7250 -10925
rect 7305 -11045 7425 -10925
rect 7470 -11045 7590 -10925
rect 7635 -11045 7755 -10925
rect 7800 -11045 7920 -10925
rect 7975 -11045 8095 -10925
rect 8140 -11045 8260 -10925
rect 8305 -11045 8425 -10925
rect 8470 -11045 8590 -10925
rect 8645 -11045 8765 -10925
rect 8810 -11045 8930 -10925
rect 8975 -11045 9095 -10925
rect 9140 -11045 9260 -10925
rect 9315 -11045 9435 -10925
rect 9480 -11045 9600 -10925
rect 9645 -11045 9765 -10925
rect 9810 -11045 9930 -10925
rect 9985 -11045 10105 -10925
rect 10150 -11045 10270 -10925
rect 10315 -11045 10435 -10925
rect 10480 -11045 10600 -10925
rect 10655 -11045 10775 -10925
rect 10820 -11045 10940 -10925
rect 10985 -11045 11105 -10925
rect 11150 -11045 11270 -10925
rect 11325 -11045 11445 -10925
rect 11490 -11045 11610 -10925
rect 11655 -11045 11775 -10925
rect 11820 -11045 11940 -10925
rect 11995 -11045 12115 -10925
rect 12160 -11045 12280 -10925
rect 12325 -11045 12445 -10925
rect 12490 -11045 12610 -10925
rect 7130 -11210 7250 -11090
rect 7305 -11210 7425 -11090
rect 7470 -11210 7590 -11090
rect 7635 -11210 7755 -11090
rect 7800 -11210 7920 -11090
rect 7975 -11210 8095 -11090
rect 8140 -11210 8260 -11090
rect 8305 -11210 8425 -11090
rect 8470 -11210 8590 -11090
rect 8645 -11210 8765 -11090
rect 8810 -11210 8930 -11090
rect 8975 -11210 9095 -11090
rect 9140 -11210 9260 -11090
rect 9315 -11210 9435 -11090
rect 9480 -11210 9600 -11090
rect 9645 -11210 9765 -11090
rect 9810 -11210 9930 -11090
rect 9985 -11210 10105 -11090
rect 10150 -11210 10270 -11090
rect 10315 -11210 10435 -11090
rect 10480 -11210 10600 -11090
rect 10655 -11210 10775 -11090
rect 10820 -11210 10940 -11090
rect 10985 -11210 11105 -11090
rect 11150 -11210 11270 -11090
rect 11325 -11210 11445 -11090
rect 11490 -11210 11610 -11090
rect 11655 -11210 11775 -11090
rect 11820 -11210 11940 -11090
rect 11995 -11210 12115 -11090
rect 12160 -11210 12280 -11090
rect 12325 -11210 12445 -11090
rect 12490 -11210 12610 -11090
rect 7130 -11375 7250 -11255
rect 7305 -11375 7425 -11255
rect 7470 -11375 7590 -11255
rect 7635 -11375 7755 -11255
rect 7800 -11375 7920 -11255
rect 7975 -11375 8095 -11255
rect 8140 -11375 8260 -11255
rect 8305 -11375 8425 -11255
rect 8470 -11375 8590 -11255
rect 8645 -11375 8765 -11255
rect 8810 -11375 8930 -11255
rect 8975 -11375 9095 -11255
rect 9140 -11375 9260 -11255
rect 9315 -11375 9435 -11255
rect 9480 -11375 9600 -11255
rect 9645 -11375 9765 -11255
rect 9810 -11375 9930 -11255
rect 9985 -11375 10105 -11255
rect 10150 -11375 10270 -11255
rect 10315 -11375 10435 -11255
rect 10480 -11375 10600 -11255
rect 10655 -11375 10775 -11255
rect 10820 -11375 10940 -11255
rect 10985 -11375 11105 -11255
rect 11150 -11375 11270 -11255
rect 11325 -11375 11445 -11255
rect 11490 -11375 11610 -11255
rect 11655 -11375 11775 -11255
rect 11820 -11375 11940 -11255
rect 11995 -11375 12115 -11255
rect 12160 -11375 12280 -11255
rect 12325 -11375 12445 -11255
rect 12490 -11375 12610 -11255
rect 7130 -11550 7250 -11430
rect 7305 -11550 7425 -11430
rect 7470 -11550 7590 -11430
rect 7635 -11550 7755 -11430
rect 7800 -11550 7920 -11430
rect 7975 -11550 8095 -11430
rect 8140 -11550 8260 -11430
rect 8305 -11550 8425 -11430
rect 8470 -11550 8590 -11430
rect 8645 -11550 8765 -11430
rect 8810 -11550 8930 -11430
rect 8975 -11550 9095 -11430
rect 9140 -11550 9260 -11430
rect 9315 -11550 9435 -11430
rect 9480 -11550 9600 -11430
rect 9645 -11550 9765 -11430
rect 9810 -11550 9930 -11430
rect 9985 -11550 10105 -11430
rect 10150 -11550 10270 -11430
rect 10315 -11550 10435 -11430
rect 10480 -11550 10600 -11430
rect 10655 -11550 10775 -11430
rect 10820 -11550 10940 -11430
rect 10985 -11550 11105 -11430
rect 11150 -11550 11270 -11430
rect 11325 -11550 11445 -11430
rect 11490 -11550 11610 -11430
rect 11655 -11550 11775 -11430
rect 11820 -11550 11940 -11430
rect 11995 -11550 12115 -11430
rect 12160 -11550 12280 -11430
rect 12325 -11550 12445 -11430
rect 12490 -11550 12610 -11430
rect 7130 -11715 7250 -11595
rect 7305 -11715 7425 -11595
rect 7470 -11715 7590 -11595
rect 7635 -11715 7755 -11595
rect 7800 -11715 7920 -11595
rect 7975 -11715 8095 -11595
rect 8140 -11715 8260 -11595
rect 8305 -11715 8425 -11595
rect 8470 -11715 8590 -11595
rect 8645 -11715 8765 -11595
rect 8810 -11715 8930 -11595
rect 8975 -11715 9095 -11595
rect 9140 -11715 9260 -11595
rect 9315 -11715 9435 -11595
rect 9480 -11715 9600 -11595
rect 9645 -11715 9765 -11595
rect 9810 -11715 9930 -11595
rect 9985 -11715 10105 -11595
rect 10150 -11715 10270 -11595
rect 10315 -11715 10435 -11595
rect 10480 -11715 10600 -11595
rect 10655 -11715 10775 -11595
rect 10820 -11715 10940 -11595
rect 10985 -11715 11105 -11595
rect 11150 -11715 11270 -11595
rect 11325 -11715 11445 -11595
rect 11490 -11715 11610 -11595
rect 11655 -11715 11775 -11595
rect 11820 -11715 11940 -11595
rect 11995 -11715 12115 -11595
rect 12160 -11715 12280 -11595
rect 12325 -11715 12445 -11595
rect 12490 -11715 12610 -11595
rect 7130 -11880 7250 -11760
rect 7305 -11880 7425 -11760
rect 7470 -11880 7590 -11760
rect 7635 -11880 7755 -11760
rect 7800 -11880 7920 -11760
rect 7975 -11880 8095 -11760
rect 8140 -11880 8260 -11760
rect 8305 -11880 8425 -11760
rect 8470 -11880 8590 -11760
rect 8645 -11880 8765 -11760
rect 8810 -11880 8930 -11760
rect 8975 -11880 9095 -11760
rect 9140 -11880 9260 -11760
rect 9315 -11880 9435 -11760
rect 9480 -11880 9600 -11760
rect 9645 -11880 9765 -11760
rect 9810 -11880 9930 -11760
rect 9985 -11880 10105 -11760
rect 10150 -11880 10270 -11760
rect 10315 -11880 10435 -11760
rect 10480 -11880 10600 -11760
rect 10655 -11880 10775 -11760
rect 10820 -11880 10940 -11760
rect 10985 -11880 11105 -11760
rect 11150 -11880 11270 -11760
rect 11325 -11880 11445 -11760
rect 11490 -11880 11610 -11760
rect 11655 -11880 11775 -11760
rect 11820 -11880 11940 -11760
rect 11995 -11880 12115 -11760
rect 12160 -11880 12280 -11760
rect 12325 -11880 12445 -11760
rect 12490 -11880 12610 -11760
rect 7130 -12045 7250 -11925
rect 7305 -12045 7425 -11925
rect 7470 -12045 7590 -11925
rect 7635 -12045 7755 -11925
rect 7800 -12045 7920 -11925
rect 7975 -12045 8095 -11925
rect 8140 -12045 8260 -11925
rect 8305 -12045 8425 -11925
rect 8470 -12045 8590 -11925
rect 8645 -12045 8765 -11925
rect 8810 -12045 8930 -11925
rect 8975 -12045 9095 -11925
rect 9140 -12045 9260 -11925
rect 9315 -12045 9435 -11925
rect 9480 -12045 9600 -11925
rect 9645 -12045 9765 -11925
rect 9810 -12045 9930 -11925
rect 9985 -12045 10105 -11925
rect 10150 -12045 10270 -11925
rect 10315 -12045 10435 -11925
rect 10480 -12045 10600 -11925
rect 10655 -12045 10775 -11925
rect 10820 -12045 10940 -11925
rect 10985 -12045 11105 -11925
rect 11150 -12045 11270 -11925
rect 11325 -12045 11445 -11925
rect 11490 -12045 11610 -11925
rect 11655 -12045 11775 -11925
rect 11820 -12045 11940 -11925
rect 11995 -12045 12115 -11925
rect 12160 -12045 12280 -11925
rect 12325 -12045 12445 -11925
rect 12490 -12045 12610 -11925
rect 7130 -12220 7250 -12100
rect 7305 -12220 7425 -12100
rect 7470 -12220 7590 -12100
rect 7635 -12220 7755 -12100
rect 7800 -12220 7920 -12100
rect 7975 -12220 8095 -12100
rect 8140 -12220 8260 -12100
rect 8305 -12220 8425 -12100
rect 8470 -12220 8590 -12100
rect 8645 -12220 8765 -12100
rect 8810 -12220 8930 -12100
rect 8975 -12220 9095 -12100
rect 9140 -12220 9260 -12100
rect 9315 -12220 9435 -12100
rect 9480 -12220 9600 -12100
rect 9645 -12220 9765 -12100
rect 9810 -12220 9930 -12100
rect 9985 -12220 10105 -12100
rect 10150 -12220 10270 -12100
rect 10315 -12220 10435 -12100
rect 10480 -12220 10600 -12100
rect 10655 -12220 10775 -12100
rect 10820 -12220 10940 -12100
rect 10985 -12220 11105 -12100
rect 11150 -12220 11270 -12100
rect 11325 -12220 11445 -12100
rect 11490 -12220 11610 -12100
rect 11655 -12220 11775 -12100
rect 11820 -12220 11940 -12100
rect 11995 -12220 12115 -12100
rect 12160 -12220 12280 -12100
rect 12325 -12220 12445 -12100
rect 12490 -12220 12610 -12100
rect 7130 -12385 7250 -12265
rect 7305 -12385 7425 -12265
rect 7470 -12385 7590 -12265
rect 7635 -12385 7755 -12265
rect 7800 -12385 7920 -12265
rect 7975 -12385 8095 -12265
rect 8140 -12385 8260 -12265
rect 8305 -12385 8425 -12265
rect 8470 -12385 8590 -12265
rect 8645 -12385 8765 -12265
rect 8810 -12385 8930 -12265
rect 8975 -12385 9095 -12265
rect 9140 -12385 9260 -12265
rect 9315 -12385 9435 -12265
rect 9480 -12385 9600 -12265
rect 9645 -12385 9765 -12265
rect 9810 -12385 9930 -12265
rect 9985 -12385 10105 -12265
rect 10150 -12385 10270 -12265
rect 10315 -12385 10435 -12265
rect 10480 -12385 10600 -12265
rect 10655 -12385 10775 -12265
rect 10820 -12385 10940 -12265
rect 10985 -12385 11105 -12265
rect 11150 -12385 11270 -12265
rect 11325 -12385 11445 -12265
rect 11490 -12385 11610 -12265
rect 11655 -12385 11775 -12265
rect 11820 -12385 11940 -12265
rect 11995 -12385 12115 -12265
rect 12160 -12385 12280 -12265
rect 12325 -12385 12445 -12265
rect 12490 -12385 12610 -12265
rect 7130 -12550 7250 -12430
rect 7305 -12550 7425 -12430
rect 7470 -12550 7590 -12430
rect 7635 -12550 7755 -12430
rect 7800 -12550 7920 -12430
rect 7975 -12550 8095 -12430
rect 8140 -12550 8260 -12430
rect 8305 -12550 8425 -12430
rect 8470 -12550 8590 -12430
rect 8645 -12550 8765 -12430
rect 8810 -12550 8930 -12430
rect 8975 -12550 9095 -12430
rect 9140 -12550 9260 -12430
rect 9315 -12550 9435 -12430
rect 9480 -12550 9600 -12430
rect 9645 -12550 9765 -12430
rect 9810 -12550 9930 -12430
rect 9985 -12550 10105 -12430
rect 10150 -12550 10270 -12430
rect 10315 -12550 10435 -12430
rect 10480 -12550 10600 -12430
rect 10655 -12550 10775 -12430
rect 10820 -12550 10940 -12430
rect 10985 -12550 11105 -12430
rect 11150 -12550 11270 -12430
rect 11325 -12550 11445 -12430
rect 11490 -12550 11610 -12430
rect 11655 -12550 11775 -12430
rect 11820 -12550 11940 -12430
rect 11995 -12550 12115 -12430
rect 12160 -12550 12280 -12430
rect 12325 -12550 12445 -12430
rect 12490 -12550 12610 -12430
rect 7130 -12715 7250 -12595
rect 7305 -12715 7425 -12595
rect 7470 -12715 7590 -12595
rect 7635 -12715 7755 -12595
rect 7800 -12715 7920 -12595
rect 7975 -12715 8095 -12595
rect 8140 -12715 8260 -12595
rect 8305 -12715 8425 -12595
rect 8470 -12715 8590 -12595
rect 8645 -12715 8765 -12595
rect 8810 -12715 8930 -12595
rect 8975 -12715 9095 -12595
rect 9140 -12715 9260 -12595
rect 9315 -12715 9435 -12595
rect 9480 -12715 9600 -12595
rect 9645 -12715 9765 -12595
rect 9810 -12715 9930 -12595
rect 9985 -12715 10105 -12595
rect 10150 -12715 10270 -12595
rect 10315 -12715 10435 -12595
rect 10480 -12715 10600 -12595
rect 10655 -12715 10775 -12595
rect 10820 -12715 10940 -12595
rect 10985 -12715 11105 -12595
rect 11150 -12715 11270 -12595
rect 11325 -12715 11445 -12595
rect 11490 -12715 11610 -12595
rect 11655 -12715 11775 -12595
rect 11820 -12715 11940 -12595
rect 11995 -12715 12115 -12595
rect 12160 -12715 12280 -12595
rect 12325 -12715 12445 -12595
rect 12490 -12715 12610 -12595
rect 7130 -12890 7250 -12770
rect 7305 -12890 7425 -12770
rect 7470 -12890 7590 -12770
rect 7635 -12890 7755 -12770
rect 7800 -12890 7920 -12770
rect 7975 -12890 8095 -12770
rect 8140 -12890 8260 -12770
rect 8305 -12890 8425 -12770
rect 8470 -12890 8590 -12770
rect 8645 -12890 8765 -12770
rect 8810 -12890 8930 -12770
rect 8975 -12890 9095 -12770
rect 9140 -12890 9260 -12770
rect 9315 -12890 9435 -12770
rect 9480 -12890 9600 -12770
rect 9645 -12890 9765 -12770
rect 9810 -12890 9930 -12770
rect 9985 -12890 10105 -12770
rect 10150 -12890 10270 -12770
rect 10315 -12890 10435 -12770
rect 10480 -12890 10600 -12770
rect 10655 -12890 10775 -12770
rect 10820 -12890 10940 -12770
rect 10985 -12890 11105 -12770
rect 11150 -12890 11270 -12770
rect 11325 -12890 11445 -12770
rect 11490 -12890 11610 -12770
rect 11655 -12890 11775 -12770
rect 11820 -12890 11940 -12770
rect 11995 -12890 12115 -12770
rect 12160 -12890 12280 -12770
rect 12325 -12890 12445 -12770
rect 12490 -12890 12610 -12770
rect 7130 -13055 7250 -12935
rect 7305 -13055 7425 -12935
rect 7470 -13055 7590 -12935
rect 7635 -13055 7755 -12935
rect 7800 -13055 7920 -12935
rect 7975 -13055 8095 -12935
rect 8140 -13055 8260 -12935
rect 8305 -13055 8425 -12935
rect 8470 -13055 8590 -12935
rect 8645 -13055 8765 -12935
rect 8810 -13055 8930 -12935
rect 8975 -13055 9095 -12935
rect 9140 -13055 9260 -12935
rect 9315 -13055 9435 -12935
rect 9480 -13055 9600 -12935
rect 9645 -13055 9765 -12935
rect 9810 -13055 9930 -12935
rect 9985 -13055 10105 -12935
rect 10150 -13055 10270 -12935
rect 10315 -13055 10435 -12935
rect 10480 -13055 10600 -12935
rect 10655 -13055 10775 -12935
rect 10820 -13055 10940 -12935
rect 10985 -13055 11105 -12935
rect 11150 -13055 11270 -12935
rect 11325 -13055 11445 -12935
rect 11490 -13055 11610 -12935
rect 11655 -13055 11775 -12935
rect 11820 -13055 11940 -12935
rect 11995 -13055 12115 -12935
rect 12160 -13055 12280 -12935
rect 12325 -13055 12445 -12935
rect 12490 -13055 12610 -12935
rect 7130 -13220 7250 -13100
rect 7305 -13220 7425 -13100
rect 7470 -13220 7590 -13100
rect 7635 -13220 7755 -13100
rect 7800 -13220 7920 -13100
rect 7975 -13220 8095 -13100
rect 8140 -13220 8260 -13100
rect 8305 -13220 8425 -13100
rect 8470 -13220 8590 -13100
rect 8645 -13220 8765 -13100
rect 8810 -13220 8930 -13100
rect 8975 -13220 9095 -13100
rect 9140 -13220 9260 -13100
rect 9315 -13220 9435 -13100
rect 9480 -13220 9600 -13100
rect 9645 -13220 9765 -13100
rect 9810 -13220 9930 -13100
rect 9985 -13220 10105 -13100
rect 10150 -13220 10270 -13100
rect 10315 -13220 10435 -13100
rect 10480 -13220 10600 -13100
rect 10655 -13220 10775 -13100
rect 10820 -13220 10940 -13100
rect 10985 -13220 11105 -13100
rect 11150 -13220 11270 -13100
rect 11325 -13220 11445 -13100
rect 11490 -13220 11610 -13100
rect 11655 -13220 11775 -13100
rect 11820 -13220 11940 -13100
rect 11995 -13220 12115 -13100
rect 12160 -13220 12280 -13100
rect 12325 -13220 12445 -13100
rect 12490 -13220 12610 -13100
rect 7130 -13385 7250 -13265
rect 7305 -13385 7425 -13265
rect 7470 -13385 7590 -13265
rect 7635 -13385 7755 -13265
rect 7800 -13385 7920 -13265
rect 7975 -13385 8095 -13265
rect 8140 -13385 8260 -13265
rect 8305 -13385 8425 -13265
rect 8470 -13385 8590 -13265
rect 8645 -13385 8765 -13265
rect 8810 -13385 8930 -13265
rect 8975 -13385 9095 -13265
rect 9140 -13385 9260 -13265
rect 9315 -13385 9435 -13265
rect 9480 -13385 9600 -13265
rect 9645 -13385 9765 -13265
rect 9810 -13385 9930 -13265
rect 9985 -13385 10105 -13265
rect 10150 -13385 10270 -13265
rect 10315 -13385 10435 -13265
rect 10480 -13385 10600 -13265
rect 10655 -13385 10775 -13265
rect 10820 -13385 10940 -13265
rect 10985 -13385 11105 -13265
rect 11150 -13385 11270 -13265
rect 11325 -13385 11445 -13265
rect 11490 -13385 11610 -13265
rect 11655 -13385 11775 -13265
rect 11820 -13385 11940 -13265
rect 11995 -13385 12115 -13265
rect 12160 -13385 12280 -13265
rect 12325 -13385 12445 -13265
rect 12490 -13385 12610 -13265
rect 7130 -13560 7250 -13440
rect 7305 -13560 7425 -13440
rect 7470 -13560 7590 -13440
rect 7635 -13560 7755 -13440
rect 7800 -13560 7920 -13440
rect 7975 -13560 8095 -13440
rect 8140 -13560 8260 -13440
rect 8305 -13560 8425 -13440
rect 8470 -13560 8590 -13440
rect 8645 -13560 8765 -13440
rect 8810 -13560 8930 -13440
rect 8975 -13560 9095 -13440
rect 9140 -13560 9260 -13440
rect 9315 -13560 9435 -13440
rect 9480 -13560 9600 -13440
rect 9645 -13560 9765 -13440
rect 9810 -13560 9930 -13440
rect 9985 -13560 10105 -13440
rect 10150 -13560 10270 -13440
rect 10315 -13560 10435 -13440
rect 10480 -13560 10600 -13440
rect 10655 -13560 10775 -13440
rect 10820 -13560 10940 -13440
rect 10985 -13560 11105 -13440
rect 11150 -13560 11270 -13440
rect 11325 -13560 11445 -13440
rect 11490 -13560 11610 -13440
rect 11655 -13560 11775 -13440
rect 11820 -13560 11940 -13440
rect 11995 -13560 12115 -13440
rect 12160 -13560 12280 -13440
rect 12325 -13560 12445 -13440
rect 12490 -13560 12610 -13440
rect 7130 -13725 7250 -13605
rect 7305 -13725 7425 -13605
rect 7470 -13725 7590 -13605
rect 7635 -13725 7755 -13605
rect 7800 -13725 7920 -13605
rect 7975 -13725 8095 -13605
rect 8140 -13725 8260 -13605
rect 8305 -13725 8425 -13605
rect 8470 -13725 8590 -13605
rect 8645 -13725 8765 -13605
rect 8810 -13725 8930 -13605
rect 8975 -13725 9095 -13605
rect 9140 -13725 9260 -13605
rect 9315 -13725 9435 -13605
rect 9480 -13725 9600 -13605
rect 9645 -13725 9765 -13605
rect 9810 -13725 9930 -13605
rect 9985 -13725 10105 -13605
rect 10150 -13725 10270 -13605
rect 10315 -13725 10435 -13605
rect 10480 -13725 10600 -13605
rect 10655 -13725 10775 -13605
rect 10820 -13725 10940 -13605
rect 10985 -13725 11105 -13605
rect 11150 -13725 11270 -13605
rect 11325 -13725 11445 -13605
rect 11490 -13725 11610 -13605
rect 11655 -13725 11775 -13605
rect 11820 -13725 11940 -13605
rect 11995 -13725 12115 -13605
rect 12160 -13725 12280 -13605
rect 12325 -13725 12445 -13605
rect 12490 -13725 12610 -13605
rect 7130 -13890 7250 -13770
rect 7305 -13890 7425 -13770
rect 7470 -13890 7590 -13770
rect 7635 -13890 7755 -13770
rect 7800 -13890 7920 -13770
rect 7975 -13890 8095 -13770
rect 8140 -13890 8260 -13770
rect 8305 -13890 8425 -13770
rect 8470 -13890 8590 -13770
rect 8645 -13890 8765 -13770
rect 8810 -13890 8930 -13770
rect 8975 -13890 9095 -13770
rect 9140 -13890 9260 -13770
rect 9315 -13890 9435 -13770
rect 9480 -13890 9600 -13770
rect 9645 -13890 9765 -13770
rect 9810 -13890 9930 -13770
rect 9985 -13890 10105 -13770
rect 10150 -13890 10270 -13770
rect 10315 -13890 10435 -13770
rect 10480 -13890 10600 -13770
rect 10655 -13890 10775 -13770
rect 10820 -13890 10940 -13770
rect 10985 -13890 11105 -13770
rect 11150 -13890 11270 -13770
rect 11325 -13890 11445 -13770
rect 11490 -13890 11610 -13770
rect 11655 -13890 11775 -13770
rect 11820 -13890 11940 -13770
rect 11995 -13890 12115 -13770
rect 12160 -13890 12280 -13770
rect 12325 -13890 12445 -13770
rect 12490 -13890 12610 -13770
rect 7130 -14055 7250 -13935
rect 7305 -14055 7425 -13935
rect 7470 -14055 7590 -13935
rect 7635 -14055 7755 -13935
rect 7800 -14055 7920 -13935
rect 7975 -14055 8095 -13935
rect 8140 -14055 8260 -13935
rect 8305 -14055 8425 -13935
rect 8470 -14055 8590 -13935
rect 8645 -14055 8765 -13935
rect 8810 -14055 8930 -13935
rect 8975 -14055 9095 -13935
rect 9140 -14055 9260 -13935
rect 9315 -14055 9435 -13935
rect 9480 -14055 9600 -13935
rect 9645 -14055 9765 -13935
rect 9810 -14055 9930 -13935
rect 9985 -14055 10105 -13935
rect 10150 -14055 10270 -13935
rect 10315 -14055 10435 -13935
rect 10480 -14055 10600 -13935
rect 10655 -14055 10775 -13935
rect 10820 -14055 10940 -13935
rect 10985 -14055 11105 -13935
rect 11150 -14055 11270 -13935
rect 11325 -14055 11445 -13935
rect 11490 -14055 11610 -13935
rect 11655 -14055 11775 -13935
rect 11820 -14055 11940 -13935
rect 11995 -14055 12115 -13935
rect 12160 -14055 12280 -13935
rect 12325 -14055 12445 -13935
rect 12490 -14055 12610 -13935
rect 7130 -14230 7250 -14110
rect 7305 -14230 7425 -14110
rect 7470 -14230 7590 -14110
rect 7635 -14230 7755 -14110
rect 7800 -14230 7920 -14110
rect 7975 -14230 8095 -14110
rect 8140 -14230 8260 -14110
rect 8305 -14230 8425 -14110
rect 8470 -14230 8590 -14110
rect 8645 -14230 8765 -14110
rect 8810 -14230 8930 -14110
rect 8975 -14230 9095 -14110
rect 9140 -14230 9260 -14110
rect 9315 -14230 9435 -14110
rect 9480 -14230 9600 -14110
rect 9645 -14230 9765 -14110
rect 9810 -14230 9930 -14110
rect 9985 -14230 10105 -14110
rect 10150 -14230 10270 -14110
rect 10315 -14230 10435 -14110
rect 10480 -14230 10600 -14110
rect 10655 -14230 10775 -14110
rect 10820 -14230 10940 -14110
rect 10985 -14230 11105 -14110
rect 11150 -14230 11270 -14110
rect 11325 -14230 11445 -14110
rect 11490 -14230 11610 -14110
rect 11655 -14230 11775 -14110
rect 11820 -14230 11940 -14110
rect 11995 -14230 12115 -14110
rect 12160 -14230 12280 -14110
rect 12325 -14230 12445 -14110
rect 12490 -14230 12610 -14110
rect 7130 -14395 7250 -14275
rect 7305 -14395 7425 -14275
rect 7470 -14395 7590 -14275
rect 7635 -14395 7755 -14275
rect 7800 -14395 7920 -14275
rect 7975 -14395 8095 -14275
rect 8140 -14395 8260 -14275
rect 8305 -14395 8425 -14275
rect 8470 -14395 8590 -14275
rect 8645 -14395 8765 -14275
rect 8810 -14395 8930 -14275
rect 8975 -14395 9095 -14275
rect 9140 -14395 9260 -14275
rect 9315 -14395 9435 -14275
rect 9480 -14395 9600 -14275
rect 9645 -14395 9765 -14275
rect 9810 -14395 9930 -14275
rect 9985 -14395 10105 -14275
rect 10150 -14395 10270 -14275
rect 10315 -14395 10435 -14275
rect 10480 -14395 10600 -14275
rect 10655 -14395 10775 -14275
rect 10820 -14395 10940 -14275
rect 10985 -14395 11105 -14275
rect 11150 -14395 11270 -14275
rect 11325 -14395 11445 -14275
rect 11490 -14395 11610 -14275
rect 11655 -14395 11775 -14275
rect 11820 -14395 11940 -14275
rect 11995 -14395 12115 -14275
rect 12160 -14395 12280 -14275
rect 12325 -14395 12445 -14275
rect 12490 -14395 12610 -14275
rect 7130 -14560 7250 -14440
rect 7305 -14560 7425 -14440
rect 7470 -14560 7590 -14440
rect 7635 -14560 7755 -14440
rect 7800 -14560 7920 -14440
rect 7975 -14560 8095 -14440
rect 8140 -14560 8260 -14440
rect 8305 -14560 8425 -14440
rect 8470 -14560 8590 -14440
rect 8645 -14560 8765 -14440
rect 8810 -14560 8930 -14440
rect 8975 -14560 9095 -14440
rect 9140 -14560 9260 -14440
rect 9315 -14560 9435 -14440
rect 9480 -14560 9600 -14440
rect 9645 -14560 9765 -14440
rect 9810 -14560 9930 -14440
rect 9985 -14560 10105 -14440
rect 10150 -14560 10270 -14440
rect 10315 -14560 10435 -14440
rect 10480 -14560 10600 -14440
rect 10655 -14560 10775 -14440
rect 10820 -14560 10940 -14440
rect 10985 -14560 11105 -14440
rect 11150 -14560 11270 -14440
rect 11325 -14560 11445 -14440
rect 11490 -14560 11610 -14440
rect 11655 -14560 11775 -14440
rect 11820 -14560 11940 -14440
rect 11995 -14560 12115 -14440
rect 12160 -14560 12280 -14440
rect 12325 -14560 12445 -14440
rect 12490 -14560 12610 -14440
rect 7130 -14725 7250 -14605
rect 7305 -14725 7425 -14605
rect 7470 -14725 7590 -14605
rect 7635 -14725 7755 -14605
rect 7800 -14725 7920 -14605
rect 7975 -14725 8095 -14605
rect 8140 -14725 8260 -14605
rect 8305 -14725 8425 -14605
rect 8470 -14725 8590 -14605
rect 8645 -14725 8765 -14605
rect 8810 -14725 8930 -14605
rect 8975 -14725 9095 -14605
rect 9140 -14725 9260 -14605
rect 9315 -14725 9435 -14605
rect 9480 -14725 9600 -14605
rect 9645 -14725 9765 -14605
rect 9810 -14725 9930 -14605
rect 9985 -14725 10105 -14605
rect 10150 -14725 10270 -14605
rect 10315 -14725 10435 -14605
rect 10480 -14725 10600 -14605
rect 10655 -14725 10775 -14605
rect 10820 -14725 10940 -14605
rect 10985 -14725 11105 -14605
rect 11150 -14725 11270 -14605
rect 11325 -14725 11445 -14605
rect 11490 -14725 11610 -14605
rect 11655 -14725 11775 -14605
rect 11820 -14725 11940 -14605
rect 11995 -14725 12115 -14605
rect 12160 -14725 12280 -14605
rect 12325 -14725 12445 -14605
rect 12490 -14725 12610 -14605
rect 7130 -14900 7250 -14780
rect 7305 -14900 7425 -14780
rect 7470 -14900 7590 -14780
rect 7635 -14900 7755 -14780
rect 7800 -14900 7920 -14780
rect 7975 -14900 8095 -14780
rect 8140 -14900 8260 -14780
rect 8305 -14900 8425 -14780
rect 8470 -14900 8590 -14780
rect 8645 -14900 8765 -14780
rect 8810 -14900 8930 -14780
rect 8975 -14900 9095 -14780
rect 9140 -14900 9260 -14780
rect 9315 -14900 9435 -14780
rect 9480 -14900 9600 -14780
rect 9645 -14900 9765 -14780
rect 9810 -14900 9930 -14780
rect 9985 -14900 10105 -14780
rect 10150 -14900 10270 -14780
rect 10315 -14900 10435 -14780
rect 10480 -14900 10600 -14780
rect 10655 -14900 10775 -14780
rect 10820 -14900 10940 -14780
rect 10985 -14900 11105 -14780
rect 11150 -14900 11270 -14780
rect 11325 -14900 11445 -14780
rect 11490 -14900 11610 -14780
rect 11655 -14900 11775 -14780
rect 11820 -14900 11940 -14780
rect 11995 -14900 12115 -14780
rect 12160 -14900 12280 -14780
rect 12325 -14900 12445 -14780
rect 12490 -14900 12610 -14780
rect 7130 -15065 7250 -14945
rect 7305 -15065 7425 -14945
rect 7470 -15065 7590 -14945
rect 7635 -15065 7755 -14945
rect 7800 -15065 7920 -14945
rect 7975 -15065 8095 -14945
rect 8140 -15065 8260 -14945
rect 8305 -15065 8425 -14945
rect 8470 -15065 8590 -14945
rect 8645 -15065 8765 -14945
rect 8810 -15065 8930 -14945
rect 8975 -15065 9095 -14945
rect 9140 -15065 9260 -14945
rect 9315 -15065 9435 -14945
rect 9480 -15065 9600 -14945
rect 9645 -15065 9765 -14945
rect 9810 -15065 9930 -14945
rect 9985 -15065 10105 -14945
rect 10150 -15065 10270 -14945
rect 10315 -15065 10435 -14945
rect 10480 -15065 10600 -14945
rect 10655 -15065 10775 -14945
rect 10820 -15065 10940 -14945
rect 10985 -15065 11105 -14945
rect 11150 -15065 11270 -14945
rect 11325 -15065 11445 -14945
rect 11490 -15065 11610 -14945
rect 11655 -15065 11775 -14945
rect 11820 -15065 11940 -14945
rect 11995 -15065 12115 -14945
rect 12160 -15065 12280 -14945
rect 12325 -15065 12445 -14945
rect 12490 -15065 12610 -14945
rect 7130 -15230 7250 -15110
rect 7305 -15230 7425 -15110
rect 7470 -15230 7590 -15110
rect 7635 -15230 7755 -15110
rect 7800 -15230 7920 -15110
rect 7975 -15230 8095 -15110
rect 8140 -15230 8260 -15110
rect 8305 -15230 8425 -15110
rect 8470 -15230 8590 -15110
rect 8645 -15230 8765 -15110
rect 8810 -15230 8930 -15110
rect 8975 -15230 9095 -15110
rect 9140 -15230 9260 -15110
rect 9315 -15230 9435 -15110
rect 9480 -15230 9600 -15110
rect 9645 -15230 9765 -15110
rect 9810 -15230 9930 -15110
rect 9985 -15230 10105 -15110
rect 10150 -15230 10270 -15110
rect 10315 -15230 10435 -15110
rect 10480 -15230 10600 -15110
rect 10655 -15230 10775 -15110
rect 10820 -15230 10940 -15110
rect 10985 -15230 11105 -15110
rect 11150 -15230 11270 -15110
rect 11325 -15230 11445 -15110
rect 11490 -15230 11610 -15110
rect 11655 -15230 11775 -15110
rect 11820 -15230 11940 -15110
rect 11995 -15230 12115 -15110
rect 12160 -15230 12280 -15110
rect 12325 -15230 12445 -15110
rect 12490 -15230 12610 -15110
rect 7130 -15395 7250 -15275
rect 7305 -15395 7425 -15275
rect 7470 -15395 7590 -15275
rect 7635 -15395 7755 -15275
rect 7800 -15395 7920 -15275
rect 7975 -15395 8095 -15275
rect 8140 -15395 8260 -15275
rect 8305 -15395 8425 -15275
rect 8470 -15395 8590 -15275
rect 8645 -15395 8765 -15275
rect 8810 -15395 8930 -15275
rect 8975 -15395 9095 -15275
rect 9140 -15395 9260 -15275
rect 9315 -15395 9435 -15275
rect 9480 -15395 9600 -15275
rect 9645 -15395 9765 -15275
rect 9810 -15395 9930 -15275
rect 9985 -15395 10105 -15275
rect 10150 -15395 10270 -15275
rect 10315 -15395 10435 -15275
rect 10480 -15395 10600 -15275
rect 10655 -15395 10775 -15275
rect 10820 -15395 10940 -15275
rect 10985 -15395 11105 -15275
rect 11150 -15395 11270 -15275
rect 11325 -15395 11445 -15275
rect 11490 -15395 11610 -15275
rect 11655 -15395 11775 -15275
rect 11820 -15395 11940 -15275
rect 11995 -15395 12115 -15275
rect 12160 -15395 12280 -15275
rect 12325 -15395 12445 -15275
rect 12490 -15395 12610 -15275
rect 7130 -15570 7250 -15450
rect 7305 -15570 7425 -15450
rect 7470 -15570 7590 -15450
rect 7635 -15570 7755 -15450
rect 7800 -15570 7920 -15450
rect 7975 -15570 8095 -15450
rect 8140 -15570 8260 -15450
rect 8305 -15570 8425 -15450
rect 8470 -15570 8590 -15450
rect 8645 -15570 8765 -15450
rect 8810 -15570 8930 -15450
rect 8975 -15570 9095 -15450
rect 9140 -15570 9260 -15450
rect 9315 -15570 9435 -15450
rect 9480 -15570 9600 -15450
rect 9645 -15570 9765 -15450
rect 9810 -15570 9930 -15450
rect 9985 -15570 10105 -15450
rect 10150 -15570 10270 -15450
rect 10315 -15570 10435 -15450
rect 10480 -15570 10600 -15450
rect 10655 -15570 10775 -15450
rect 10820 -15570 10940 -15450
rect 10985 -15570 11105 -15450
rect 11150 -15570 11270 -15450
rect 11325 -15570 11445 -15450
rect 11490 -15570 11610 -15450
rect 11655 -15570 11775 -15450
rect 11820 -15570 11940 -15450
rect 11995 -15570 12115 -15450
rect 12160 -15570 12280 -15450
rect 12325 -15570 12445 -15450
rect 12490 -15570 12610 -15450
rect 12820 -10210 12940 -10090
rect 12995 -10210 13115 -10090
rect 13160 -10210 13280 -10090
rect 13325 -10210 13445 -10090
rect 13490 -10210 13610 -10090
rect 13665 -10210 13785 -10090
rect 13830 -10210 13950 -10090
rect 13995 -10210 14115 -10090
rect 14160 -10210 14280 -10090
rect 14335 -10210 14455 -10090
rect 14500 -10210 14620 -10090
rect 14665 -10210 14785 -10090
rect 14830 -10210 14950 -10090
rect 15005 -10210 15125 -10090
rect 15170 -10210 15290 -10090
rect 15335 -10210 15455 -10090
rect 15500 -10210 15620 -10090
rect 15675 -10210 15795 -10090
rect 15840 -10210 15960 -10090
rect 16005 -10210 16125 -10090
rect 16170 -10210 16290 -10090
rect 16345 -10210 16465 -10090
rect 16510 -10210 16630 -10090
rect 16675 -10210 16795 -10090
rect 16840 -10210 16960 -10090
rect 17015 -10210 17135 -10090
rect 17180 -10210 17300 -10090
rect 17345 -10210 17465 -10090
rect 17510 -10210 17630 -10090
rect 17685 -10210 17805 -10090
rect 17850 -10210 17970 -10090
rect 18015 -10210 18135 -10090
rect 18180 -10210 18300 -10090
rect 12820 -10375 12940 -10255
rect 12995 -10375 13115 -10255
rect 13160 -10375 13280 -10255
rect 13325 -10375 13445 -10255
rect 13490 -10375 13610 -10255
rect 13665 -10375 13785 -10255
rect 13830 -10375 13950 -10255
rect 13995 -10375 14115 -10255
rect 14160 -10375 14280 -10255
rect 14335 -10375 14455 -10255
rect 14500 -10375 14620 -10255
rect 14665 -10375 14785 -10255
rect 14830 -10375 14950 -10255
rect 15005 -10375 15125 -10255
rect 15170 -10375 15290 -10255
rect 15335 -10375 15455 -10255
rect 15500 -10375 15620 -10255
rect 15675 -10375 15795 -10255
rect 15840 -10375 15960 -10255
rect 16005 -10375 16125 -10255
rect 16170 -10375 16290 -10255
rect 16345 -10375 16465 -10255
rect 16510 -10375 16630 -10255
rect 16675 -10375 16795 -10255
rect 16840 -10375 16960 -10255
rect 17015 -10375 17135 -10255
rect 17180 -10375 17300 -10255
rect 17345 -10375 17465 -10255
rect 17510 -10375 17630 -10255
rect 17685 -10375 17805 -10255
rect 17850 -10375 17970 -10255
rect 18015 -10375 18135 -10255
rect 18180 -10375 18300 -10255
rect 12820 -10540 12940 -10420
rect 12995 -10540 13115 -10420
rect 13160 -10540 13280 -10420
rect 13325 -10540 13445 -10420
rect 13490 -10540 13610 -10420
rect 13665 -10540 13785 -10420
rect 13830 -10540 13950 -10420
rect 13995 -10540 14115 -10420
rect 14160 -10540 14280 -10420
rect 14335 -10540 14455 -10420
rect 14500 -10540 14620 -10420
rect 14665 -10540 14785 -10420
rect 14830 -10540 14950 -10420
rect 15005 -10540 15125 -10420
rect 15170 -10540 15290 -10420
rect 15335 -10540 15455 -10420
rect 15500 -10540 15620 -10420
rect 15675 -10540 15795 -10420
rect 15840 -10540 15960 -10420
rect 16005 -10540 16125 -10420
rect 16170 -10540 16290 -10420
rect 16345 -10540 16465 -10420
rect 16510 -10540 16630 -10420
rect 16675 -10540 16795 -10420
rect 16840 -10540 16960 -10420
rect 17015 -10540 17135 -10420
rect 17180 -10540 17300 -10420
rect 17345 -10540 17465 -10420
rect 17510 -10540 17630 -10420
rect 17685 -10540 17805 -10420
rect 17850 -10540 17970 -10420
rect 18015 -10540 18135 -10420
rect 18180 -10540 18300 -10420
rect 12820 -10705 12940 -10585
rect 12995 -10705 13115 -10585
rect 13160 -10705 13280 -10585
rect 13325 -10705 13445 -10585
rect 13490 -10705 13610 -10585
rect 13665 -10705 13785 -10585
rect 13830 -10705 13950 -10585
rect 13995 -10705 14115 -10585
rect 14160 -10705 14280 -10585
rect 14335 -10705 14455 -10585
rect 14500 -10705 14620 -10585
rect 14665 -10705 14785 -10585
rect 14830 -10705 14950 -10585
rect 15005 -10705 15125 -10585
rect 15170 -10705 15290 -10585
rect 15335 -10705 15455 -10585
rect 15500 -10705 15620 -10585
rect 15675 -10705 15795 -10585
rect 15840 -10705 15960 -10585
rect 16005 -10705 16125 -10585
rect 16170 -10705 16290 -10585
rect 16345 -10705 16465 -10585
rect 16510 -10705 16630 -10585
rect 16675 -10705 16795 -10585
rect 16840 -10705 16960 -10585
rect 17015 -10705 17135 -10585
rect 17180 -10705 17300 -10585
rect 17345 -10705 17465 -10585
rect 17510 -10705 17630 -10585
rect 17685 -10705 17805 -10585
rect 17850 -10705 17970 -10585
rect 18015 -10705 18135 -10585
rect 18180 -10705 18300 -10585
rect 12820 -10880 12940 -10760
rect 12995 -10880 13115 -10760
rect 13160 -10880 13280 -10760
rect 13325 -10880 13445 -10760
rect 13490 -10880 13610 -10760
rect 13665 -10880 13785 -10760
rect 13830 -10880 13950 -10760
rect 13995 -10880 14115 -10760
rect 14160 -10880 14280 -10760
rect 14335 -10880 14455 -10760
rect 14500 -10880 14620 -10760
rect 14665 -10880 14785 -10760
rect 14830 -10880 14950 -10760
rect 15005 -10880 15125 -10760
rect 15170 -10880 15290 -10760
rect 15335 -10880 15455 -10760
rect 15500 -10880 15620 -10760
rect 15675 -10880 15795 -10760
rect 15840 -10880 15960 -10760
rect 16005 -10880 16125 -10760
rect 16170 -10880 16290 -10760
rect 16345 -10880 16465 -10760
rect 16510 -10880 16630 -10760
rect 16675 -10880 16795 -10760
rect 16840 -10880 16960 -10760
rect 17015 -10880 17135 -10760
rect 17180 -10880 17300 -10760
rect 17345 -10880 17465 -10760
rect 17510 -10880 17630 -10760
rect 17685 -10880 17805 -10760
rect 17850 -10880 17970 -10760
rect 18015 -10880 18135 -10760
rect 18180 -10880 18300 -10760
rect 12820 -11045 12940 -10925
rect 12995 -11045 13115 -10925
rect 13160 -11045 13280 -10925
rect 13325 -11045 13445 -10925
rect 13490 -11045 13610 -10925
rect 13665 -11045 13785 -10925
rect 13830 -11045 13950 -10925
rect 13995 -11045 14115 -10925
rect 14160 -11045 14280 -10925
rect 14335 -11045 14455 -10925
rect 14500 -11045 14620 -10925
rect 14665 -11045 14785 -10925
rect 14830 -11045 14950 -10925
rect 15005 -11045 15125 -10925
rect 15170 -11045 15290 -10925
rect 15335 -11045 15455 -10925
rect 15500 -11045 15620 -10925
rect 15675 -11045 15795 -10925
rect 15840 -11045 15960 -10925
rect 16005 -11045 16125 -10925
rect 16170 -11045 16290 -10925
rect 16345 -11045 16465 -10925
rect 16510 -11045 16630 -10925
rect 16675 -11045 16795 -10925
rect 16840 -11045 16960 -10925
rect 17015 -11045 17135 -10925
rect 17180 -11045 17300 -10925
rect 17345 -11045 17465 -10925
rect 17510 -11045 17630 -10925
rect 17685 -11045 17805 -10925
rect 17850 -11045 17970 -10925
rect 18015 -11045 18135 -10925
rect 18180 -11045 18300 -10925
rect 12820 -11210 12940 -11090
rect 12995 -11210 13115 -11090
rect 13160 -11210 13280 -11090
rect 13325 -11210 13445 -11090
rect 13490 -11210 13610 -11090
rect 13665 -11210 13785 -11090
rect 13830 -11210 13950 -11090
rect 13995 -11210 14115 -11090
rect 14160 -11210 14280 -11090
rect 14335 -11210 14455 -11090
rect 14500 -11210 14620 -11090
rect 14665 -11210 14785 -11090
rect 14830 -11210 14950 -11090
rect 15005 -11210 15125 -11090
rect 15170 -11210 15290 -11090
rect 15335 -11210 15455 -11090
rect 15500 -11210 15620 -11090
rect 15675 -11210 15795 -11090
rect 15840 -11210 15960 -11090
rect 16005 -11210 16125 -11090
rect 16170 -11210 16290 -11090
rect 16345 -11210 16465 -11090
rect 16510 -11210 16630 -11090
rect 16675 -11210 16795 -11090
rect 16840 -11210 16960 -11090
rect 17015 -11210 17135 -11090
rect 17180 -11210 17300 -11090
rect 17345 -11210 17465 -11090
rect 17510 -11210 17630 -11090
rect 17685 -11210 17805 -11090
rect 17850 -11210 17970 -11090
rect 18015 -11210 18135 -11090
rect 18180 -11210 18300 -11090
rect 12820 -11375 12940 -11255
rect 12995 -11375 13115 -11255
rect 13160 -11375 13280 -11255
rect 13325 -11375 13445 -11255
rect 13490 -11375 13610 -11255
rect 13665 -11375 13785 -11255
rect 13830 -11375 13950 -11255
rect 13995 -11375 14115 -11255
rect 14160 -11375 14280 -11255
rect 14335 -11375 14455 -11255
rect 14500 -11375 14620 -11255
rect 14665 -11375 14785 -11255
rect 14830 -11375 14950 -11255
rect 15005 -11375 15125 -11255
rect 15170 -11375 15290 -11255
rect 15335 -11375 15455 -11255
rect 15500 -11375 15620 -11255
rect 15675 -11375 15795 -11255
rect 15840 -11375 15960 -11255
rect 16005 -11375 16125 -11255
rect 16170 -11375 16290 -11255
rect 16345 -11375 16465 -11255
rect 16510 -11375 16630 -11255
rect 16675 -11375 16795 -11255
rect 16840 -11375 16960 -11255
rect 17015 -11375 17135 -11255
rect 17180 -11375 17300 -11255
rect 17345 -11375 17465 -11255
rect 17510 -11375 17630 -11255
rect 17685 -11375 17805 -11255
rect 17850 -11375 17970 -11255
rect 18015 -11375 18135 -11255
rect 18180 -11375 18300 -11255
rect 12820 -11550 12940 -11430
rect 12995 -11550 13115 -11430
rect 13160 -11550 13280 -11430
rect 13325 -11550 13445 -11430
rect 13490 -11550 13610 -11430
rect 13665 -11550 13785 -11430
rect 13830 -11550 13950 -11430
rect 13995 -11550 14115 -11430
rect 14160 -11550 14280 -11430
rect 14335 -11550 14455 -11430
rect 14500 -11550 14620 -11430
rect 14665 -11550 14785 -11430
rect 14830 -11550 14950 -11430
rect 15005 -11550 15125 -11430
rect 15170 -11550 15290 -11430
rect 15335 -11550 15455 -11430
rect 15500 -11550 15620 -11430
rect 15675 -11550 15795 -11430
rect 15840 -11550 15960 -11430
rect 16005 -11550 16125 -11430
rect 16170 -11550 16290 -11430
rect 16345 -11550 16465 -11430
rect 16510 -11550 16630 -11430
rect 16675 -11550 16795 -11430
rect 16840 -11550 16960 -11430
rect 17015 -11550 17135 -11430
rect 17180 -11550 17300 -11430
rect 17345 -11550 17465 -11430
rect 17510 -11550 17630 -11430
rect 17685 -11550 17805 -11430
rect 17850 -11550 17970 -11430
rect 18015 -11550 18135 -11430
rect 18180 -11550 18300 -11430
rect 12820 -11715 12940 -11595
rect 12995 -11715 13115 -11595
rect 13160 -11715 13280 -11595
rect 13325 -11715 13445 -11595
rect 13490 -11715 13610 -11595
rect 13665 -11715 13785 -11595
rect 13830 -11715 13950 -11595
rect 13995 -11715 14115 -11595
rect 14160 -11715 14280 -11595
rect 14335 -11715 14455 -11595
rect 14500 -11715 14620 -11595
rect 14665 -11715 14785 -11595
rect 14830 -11715 14950 -11595
rect 15005 -11715 15125 -11595
rect 15170 -11715 15290 -11595
rect 15335 -11715 15455 -11595
rect 15500 -11715 15620 -11595
rect 15675 -11715 15795 -11595
rect 15840 -11715 15960 -11595
rect 16005 -11715 16125 -11595
rect 16170 -11715 16290 -11595
rect 16345 -11715 16465 -11595
rect 16510 -11715 16630 -11595
rect 16675 -11715 16795 -11595
rect 16840 -11715 16960 -11595
rect 17015 -11715 17135 -11595
rect 17180 -11715 17300 -11595
rect 17345 -11715 17465 -11595
rect 17510 -11715 17630 -11595
rect 17685 -11715 17805 -11595
rect 17850 -11715 17970 -11595
rect 18015 -11715 18135 -11595
rect 18180 -11715 18300 -11595
rect 12820 -11880 12940 -11760
rect 12995 -11880 13115 -11760
rect 13160 -11880 13280 -11760
rect 13325 -11880 13445 -11760
rect 13490 -11880 13610 -11760
rect 13665 -11880 13785 -11760
rect 13830 -11880 13950 -11760
rect 13995 -11880 14115 -11760
rect 14160 -11880 14280 -11760
rect 14335 -11880 14455 -11760
rect 14500 -11880 14620 -11760
rect 14665 -11880 14785 -11760
rect 14830 -11880 14950 -11760
rect 15005 -11880 15125 -11760
rect 15170 -11880 15290 -11760
rect 15335 -11880 15455 -11760
rect 15500 -11880 15620 -11760
rect 15675 -11880 15795 -11760
rect 15840 -11880 15960 -11760
rect 16005 -11880 16125 -11760
rect 16170 -11880 16290 -11760
rect 16345 -11880 16465 -11760
rect 16510 -11880 16630 -11760
rect 16675 -11880 16795 -11760
rect 16840 -11880 16960 -11760
rect 17015 -11880 17135 -11760
rect 17180 -11880 17300 -11760
rect 17345 -11880 17465 -11760
rect 17510 -11880 17630 -11760
rect 17685 -11880 17805 -11760
rect 17850 -11880 17970 -11760
rect 18015 -11880 18135 -11760
rect 18180 -11880 18300 -11760
rect 12820 -12045 12940 -11925
rect 12995 -12045 13115 -11925
rect 13160 -12045 13280 -11925
rect 13325 -12045 13445 -11925
rect 13490 -12045 13610 -11925
rect 13665 -12045 13785 -11925
rect 13830 -12045 13950 -11925
rect 13995 -12045 14115 -11925
rect 14160 -12045 14280 -11925
rect 14335 -12045 14455 -11925
rect 14500 -12045 14620 -11925
rect 14665 -12045 14785 -11925
rect 14830 -12045 14950 -11925
rect 15005 -12045 15125 -11925
rect 15170 -12045 15290 -11925
rect 15335 -12045 15455 -11925
rect 15500 -12045 15620 -11925
rect 15675 -12045 15795 -11925
rect 15840 -12045 15960 -11925
rect 16005 -12045 16125 -11925
rect 16170 -12045 16290 -11925
rect 16345 -12045 16465 -11925
rect 16510 -12045 16630 -11925
rect 16675 -12045 16795 -11925
rect 16840 -12045 16960 -11925
rect 17015 -12045 17135 -11925
rect 17180 -12045 17300 -11925
rect 17345 -12045 17465 -11925
rect 17510 -12045 17630 -11925
rect 17685 -12045 17805 -11925
rect 17850 -12045 17970 -11925
rect 18015 -12045 18135 -11925
rect 18180 -12045 18300 -11925
rect 12820 -12220 12940 -12100
rect 12995 -12220 13115 -12100
rect 13160 -12220 13280 -12100
rect 13325 -12220 13445 -12100
rect 13490 -12220 13610 -12100
rect 13665 -12220 13785 -12100
rect 13830 -12220 13950 -12100
rect 13995 -12220 14115 -12100
rect 14160 -12220 14280 -12100
rect 14335 -12220 14455 -12100
rect 14500 -12220 14620 -12100
rect 14665 -12220 14785 -12100
rect 14830 -12220 14950 -12100
rect 15005 -12220 15125 -12100
rect 15170 -12220 15290 -12100
rect 15335 -12220 15455 -12100
rect 15500 -12220 15620 -12100
rect 15675 -12220 15795 -12100
rect 15840 -12220 15960 -12100
rect 16005 -12220 16125 -12100
rect 16170 -12220 16290 -12100
rect 16345 -12220 16465 -12100
rect 16510 -12220 16630 -12100
rect 16675 -12220 16795 -12100
rect 16840 -12220 16960 -12100
rect 17015 -12220 17135 -12100
rect 17180 -12220 17300 -12100
rect 17345 -12220 17465 -12100
rect 17510 -12220 17630 -12100
rect 17685 -12220 17805 -12100
rect 17850 -12220 17970 -12100
rect 18015 -12220 18135 -12100
rect 18180 -12220 18300 -12100
rect 12820 -12385 12940 -12265
rect 12995 -12385 13115 -12265
rect 13160 -12385 13280 -12265
rect 13325 -12385 13445 -12265
rect 13490 -12385 13610 -12265
rect 13665 -12385 13785 -12265
rect 13830 -12385 13950 -12265
rect 13995 -12385 14115 -12265
rect 14160 -12385 14280 -12265
rect 14335 -12385 14455 -12265
rect 14500 -12385 14620 -12265
rect 14665 -12385 14785 -12265
rect 14830 -12385 14950 -12265
rect 15005 -12385 15125 -12265
rect 15170 -12385 15290 -12265
rect 15335 -12385 15455 -12265
rect 15500 -12385 15620 -12265
rect 15675 -12385 15795 -12265
rect 15840 -12385 15960 -12265
rect 16005 -12385 16125 -12265
rect 16170 -12385 16290 -12265
rect 16345 -12385 16465 -12265
rect 16510 -12385 16630 -12265
rect 16675 -12385 16795 -12265
rect 16840 -12385 16960 -12265
rect 17015 -12385 17135 -12265
rect 17180 -12385 17300 -12265
rect 17345 -12385 17465 -12265
rect 17510 -12385 17630 -12265
rect 17685 -12385 17805 -12265
rect 17850 -12385 17970 -12265
rect 18015 -12385 18135 -12265
rect 18180 -12385 18300 -12265
rect 12820 -12550 12940 -12430
rect 12995 -12550 13115 -12430
rect 13160 -12550 13280 -12430
rect 13325 -12550 13445 -12430
rect 13490 -12550 13610 -12430
rect 13665 -12550 13785 -12430
rect 13830 -12550 13950 -12430
rect 13995 -12550 14115 -12430
rect 14160 -12550 14280 -12430
rect 14335 -12550 14455 -12430
rect 14500 -12550 14620 -12430
rect 14665 -12550 14785 -12430
rect 14830 -12550 14950 -12430
rect 15005 -12550 15125 -12430
rect 15170 -12550 15290 -12430
rect 15335 -12550 15455 -12430
rect 15500 -12550 15620 -12430
rect 15675 -12550 15795 -12430
rect 15840 -12550 15960 -12430
rect 16005 -12550 16125 -12430
rect 16170 -12550 16290 -12430
rect 16345 -12550 16465 -12430
rect 16510 -12550 16630 -12430
rect 16675 -12550 16795 -12430
rect 16840 -12550 16960 -12430
rect 17015 -12550 17135 -12430
rect 17180 -12550 17300 -12430
rect 17345 -12550 17465 -12430
rect 17510 -12550 17630 -12430
rect 17685 -12550 17805 -12430
rect 17850 -12550 17970 -12430
rect 18015 -12550 18135 -12430
rect 18180 -12550 18300 -12430
rect 12820 -12715 12940 -12595
rect 12995 -12715 13115 -12595
rect 13160 -12715 13280 -12595
rect 13325 -12715 13445 -12595
rect 13490 -12715 13610 -12595
rect 13665 -12715 13785 -12595
rect 13830 -12715 13950 -12595
rect 13995 -12715 14115 -12595
rect 14160 -12715 14280 -12595
rect 14335 -12715 14455 -12595
rect 14500 -12715 14620 -12595
rect 14665 -12715 14785 -12595
rect 14830 -12715 14950 -12595
rect 15005 -12715 15125 -12595
rect 15170 -12715 15290 -12595
rect 15335 -12715 15455 -12595
rect 15500 -12715 15620 -12595
rect 15675 -12715 15795 -12595
rect 15840 -12715 15960 -12595
rect 16005 -12715 16125 -12595
rect 16170 -12715 16290 -12595
rect 16345 -12715 16465 -12595
rect 16510 -12715 16630 -12595
rect 16675 -12715 16795 -12595
rect 16840 -12715 16960 -12595
rect 17015 -12715 17135 -12595
rect 17180 -12715 17300 -12595
rect 17345 -12715 17465 -12595
rect 17510 -12715 17630 -12595
rect 17685 -12715 17805 -12595
rect 17850 -12715 17970 -12595
rect 18015 -12715 18135 -12595
rect 18180 -12715 18300 -12595
rect 12820 -12890 12940 -12770
rect 12995 -12890 13115 -12770
rect 13160 -12890 13280 -12770
rect 13325 -12890 13445 -12770
rect 13490 -12890 13610 -12770
rect 13665 -12890 13785 -12770
rect 13830 -12890 13950 -12770
rect 13995 -12890 14115 -12770
rect 14160 -12890 14280 -12770
rect 14335 -12890 14455 -12770
rect 14500 -12890 14620 -12770
rect 14665 -12890 14785 -12770
rect 14830 -12890 14950 -12770
rect 15005 -12890 15125 -12770
rect 15170 -12890 15290 -12770
rect 15335 -12890 15455 -12770
rect 15500 -12890 15620 -12770
rect 15675 -12890 15795 -12770
rect 15840 -12890 15960 -12770
rect 16005 -12890 16125 -12770
rect 16170 -12890 16290 -12770
rect 16345 -12890 16465 -12770
rect 16510 -12890 16630 -12770
rect 16675 -12890 16795 -12770
rect 16840 -12890 16960 -12770
rect 17015 -12890 17135 -12770
rect 17180 -12890 17300 -12770
rect 17345 -12890 17465 -12770
rect 17510 -12890 17630 -12770
rect 17685 -12890 17805 -12770
rect 17850 -12890 17970 -12770
rect 18015 -12890 18135 -12770
rect 18180 -12890 18300 -12770
rect 12820 -13055 12940 -12935
rect 12995 -13055 13115 -12935
rect 13160 -13055 13280 -12935
rect 13325 -13055 13445 -12935
rect 13490 -13055 13610 -12935
rect 13665 -13055 13785 -12935
rect 13830 -13055 13950 -12935
rect 13995 -13055 14115 -12935
rect 14160 -13055 14280 -12935
rect 14335 -13055 14455 -12935
rect 14500 -13055 14620 -12935
rect 14665 -13055 14785 -12935
rect 14830 -13055 14950 -12935
rect 15005 -13055 15125 -12935
rect 15170 -13055 15290 -12935
rect 15335 -13055 15455 -12935
rect 15500 -13055 15620 -12935
rect 15675 -13055 15795 -12935
rect 15840 -13055 15960 -12935
rect 16005 -13055 16125 -12935
rect 16170 -13055 16290 -12935
rect 16345 -13055 16465 -12935
rect 16510 -13055 16630 -12935
rect 16675 -13055 16795 -12935
rect 16840 -13055 16960 -12935
rect 17015 -13055 17135 -12935
rect 17180 -13055 17300 -12935
rect 17345 -13055 17465 -12935
rect 17510 -13055 17630 -12935
rect 17685 -13055 17805 -12935
rect 17850 -13055 17970 -12935
rect 18015 -13055 18135 -12935
rect 18180 -13055 18300 -12935
rect 12820 -13220 12940 -13100
rect 12995 -13220 13115 -13100
rect 13160 -13220 13280 -13100
rect 13325 -13220 13445 -13100
rect 13490 -13220 13610 -13100
rect 13665 -13220 13785 -13100
rect 13830 -13220 13950 -13100
rect 13995 -13220 14115 -13100
rect 14160 -13220 14280 -13100
rect 14335 -13220 14455 -13100
rect 14500 -13220 14620 -13100
rect 14665 -13220 14785 -13100
rect 14830 -13220 14950 -13100
rect 15005 -13220 15125 -13100
rect 15170 -13220 15290 -13100
rect 15335 -13220 15455 -13100
rect 15500 -13220 15620 -13100
rect 15675 -13220 15795 -13100
rect 15840 -13220 15960 -13100
rect 16005 -13220 16125 -13100
rect 16170 -13220 16290 -13100
rect 16345 -13220 16465 -13100
rect 16510 -13220 16630 -13100
rect 16675 -13220 16795 -13100
rect 16840 -13220 16960 -13100
rect 17015 -13220 17135 -13100
rect 17180 -13220 17300 -13100
rect 17345 -13220 17465 -13100
rect 17510 -13220 17630 -13100
rect 17685 -13220 17805 -13100
rect 17850 -13220 17970 -13100
rect 18015 -13220 18135 -13100
rect 18180 -13220 18300 -13100
rect 12820 -13385 12940 -13265
rect 12995 -13385 13115 -13265
rect 13160 -13385 13280 -13265
rect 13325 -13385 13445 -13265
rect 13490 -13385 13610 -13265
rect 13665 -13385 13785 -13265
rect 13830 -13385 13950 -13265
rect 13995 -13385 14115 -13265
rect 14160 -13385 14280 -13265
rect 14335 -13385 14455 -13265
rect 14500 -13385 14620 -13265
rect 14665 -13385 14785 -13265
rect 14830 -13385 14950 -13265
rect 15005 -13385 15125 -13265
rect 15170 -13385 15290 -13265
rect 15335 -13385 15455 -13265
rect 15500 -13385 15620 -13265
rect 15675 -13385 15795 -13265
rect 15840 -13385 15960 -13265
rect 16005 -13385 16125 -13265
rect 16170 -13385 16290 -13265
rect 16345 -13385 16465 -13265
rect 16510 -13385 16630 -13265
rect 16675 -13385 16795 -13265
rect 16840 -13385 16960 -13265
rect 17015 -13385 17135 -13265
rect 17180 -13385 17300 -13265
rect 17345 -13385 17465 -13265
rect 17510 -13385 17630 -13265
rect 17685 -13385 17805 -13265
rect 17850 -13385 17970 -13265
rect 18015 -13385 18135 -13265
rect 18180 -13385 18300 -13265
rect 12820 -13560 12940 -13440
rect 12995 -13560 13115 -13440
rect 13160 -13560 13280 -13440
rect 13325 -13560 13445 -13440
rect 13490 -13560 13610 -13440
rect 13665 -13560 13785 -13440
rect 13830 -13560 13950 -13440
rect 13995 -13560 14115 -13440
rect 14160 -13560 14280 -13440
rect 14335 -13560 14455 -13440
rect 14500 -13560 14620 -13440
rect 14665 -13560 14785 -13440
rect 14830 -13560 14950 -13440
rect 15005 -13560 15125 -13440
rect 15170 -13560 15290 -13440
rect 15335 -13560 15455 -13440
rect 15500 -13560 15620 -13440
rect 15675 -13560 15795 -13440
rect 15840 -13560 15960 -13440
rect 16005 -13560 16125 -13440
rect 16170 -13560 16290 -13440
rect 16345 -13560 16465 -13440
rect 16510 -13560 16630 -13440
rect 16675 -13560 16795 -13440
rect 16840 -13560 16960 -13440
rect 17015 -13560 17135 -13440
rect 17180 -13560 17300 -13440
rect 17345 -13560 17465 -13440
rect 17510 -13560 17630 -13440
rect 17685 -13560 17805 -13440
rect 17850 -13560 17970 -13440
rect 18015 -13560 18135 -13440
rect 18180 -13560 18300 -13440
rect 12820 -13725 12940 -13605
rect 12995 -13725 13115 -13605
rect 13160 -13725 13280 -13605
rect 13325 -13725 13445 -13605
rect 13490 -13725 13610 -13605
rect 13665 -13725 13785 -13605
rect 13830 -13725 13950 -13605
rect 13995 -13725 14115 -13605
rect 14160 -13725 14280 -13605
rect 14335 -13725 14455 -13605
rect 14500 -13725 14620 -13605
rect 14665 -13725 14785 -13605
rect 14830 -13725 14950 -13605
rect 15005 -13725 15125 -13605
rect 15170 -13725 15290 -13605
rect 15335 -13725 15455 -13605
rect 15500 -13725 15620 -13605
rect 15675 -13725 15795 -13605
rect 15840 -13725 15960 -13605
rect 16005 -13725 16125 -13605
rect 16170 -13725 16290 -13605
rect 16345 -13725 16465 -13605
rect 16510 -13725 16630 -13605
rect 16675 -13725 16795 -13605
rect 16840 -13725 16960 -13605
rect 17015 -13725 17135 -13605
rect 17180 -13725 17300 -13605
rect 17345 -13725 17465 -13605
rect 17510 -13725 17630 -13605
rect 17685 -13725 17805 -13605
rect 17850 -13725 17970 -13605
rect 18015 -13725 18135 -13605
rect 18180 -13725 18300 -13605
rect 12820 -13890 12940 -13770
rect 12995 -13890 13115 -13770
rect 13160 -13890 13280 -13770
rect 13325 -13890 13445 -13770
rect 13490 -13890 13610 -13770
rect 13665 -13890 13785 -13770
rect 13830 -13890 13950 -13770
rect 13995 -13890 14115 -13770
rect 14160 -13890 14280 -13770
rect 14335 -13890 14455 -13770
rect 14500 -13890 14620 -13770
rect 14665 -13890 14785 -13770
rect 14830 -13890 14950 -13770
rect 15005 -13890 15125 -13770
rect 15170 -13890 15290 -13770
rect 15335 -13890 15455 -13770
rect 15500 -13890 15620 -13770
rect 15675 -13890 15795 -13770
rect 15840 -13890 15960 -13770
rect 16005 -13890 16125 -13770
rect 16170 -13890 16290 -13770
rect 16345 -13890 16465 -13770
rect 16510 -13890 16630 -13770
rect 16675 -13890 16795 -13770
rect 16840 -13890 16960 -13770
rect 17015 -13890 17135 -13770
rect 17180 -13890 17300 -13770
rect 17345 -13890 17465 -13770
rect 17510 -13890 17630 -13770
rect 17685 -13890 17805 -13770
rect 17850 -13890 17970 -13770
rect 18015 -13890 18135 -13770
rect 18180 -13890 18300 -13770
rect 12820 -14055 12940 -13935
rect 12995 -14055 13115 -13935
rect 13160 -14055 13280 -13935
rect 13325 -14055 13445 -13935
rect 13490 -14055 13610 -13935
rect 13665 -14055 13785 -13935
rect 13830 -14055 13950 -13935
rect 13995 -14055 14115 -13935
rect 14160 -14055 14280 -13935
rect 14335 -14055 14455 -13935
rect 14500 -14055 14620 -13935
rect 14665 -14055 14785 -13935
rect 14830 -14055 14950 -13935
rect 15005 -14055 15125 -13935
rect 15170 -14055 15290 -13935
rect 15335 -14055 15455 -13935
rect 15500 -14055 15620 -13935
rect 15675 -14055 15795 -13935
rect 15840 -14055 15960 -13935
rect 16005 -14055 16125 -13935
rect 16170 -14055 16290 -13935
rect 16345 -14055 16465 -13935
rect 16510 -14055 16630 -13935
rect 16675 -14055 16795 -13935
rect 16840 -14055 16960 -13935
rect 17015 -14055 17135 -13935
rect 17180 -14055 17300 -13935
rect 17345 -14055 17465 -13935
rect 17510 -14055 17630 -13935
rect 17685 -14055 17805 -13935
rect 17850 -14055 17970 -13935
rect 18015 -14055 18135 -13935
rect 18180 -14055 18300 -13935
rect 12820 -14230 12940 -14110
rect 12995 -14230 13115 -14110
rect 13160 -14230 13280 -14110
rect 13325 -14230 13445 -14110
rect 13490 -14230 13610 -14110
rect 13665 -14230 13785 -14110
rect 13830 -14230 13950 -14110
rect 13995 -14230 14115 -14110
rect 14160 -14230 14280 -14110
rect 14335 -14230 14455 -14110
rect 14500 -14230 14620 -14110
rect 14665 -14230 14785 -14110
rect 14830 -14230 14950 -14110
rect 15005 -14230 15125 -14110
rect 15170 -14230 15290 -14110
rect 15335 -14230 15455 -14110
rect 15500 -14230 15620 -14110
rect 15675 -14230 15795 -14110
rect 15840 -14230 15960 -14110
rect 16005 -14230 16125 -14110
rect 16170 -14230 16290 -14110
rect 16345 -14230 16465 -14110
rect 16510 -14230 16630 -14110
rect 16675 -14230 16795 -14110
rect 16840 -14230 16960 -14110
rect 17015 -14230 17135 -14110
rect 17180 -14230 17300 -14110
rect 17345 -14230 17465 -14110
rect 17510 -14230 17630 -14110
rect 17685 -14230 17805 -14110
rect 17850 -14230 17970 -14110
rect 18015 -14230 18135 -14110
rect 18180 -14230 18300 -14110
rect 12820 -14395 12940 -14275
rect 12995 -14395 13115 -14275
rect 13160 -14395 13280 -14275
rect 13325 -14395 13445 -14275
rect 13490 -14395 13610 -14275
rect 13665 -14395 13785 -14275
rect 13830 -14395 13950 -14275
rect 13995 -14395 14115 -14275
rect 14160 -14395 14280 -14275
rect 14335 -14395 14455 -14275
rect 14500 -14395 14620 -14275
rect 14665 -14395 14785 -14275
rect 14830 -14395 14950 -14275
rect 15005 -14395 15125 -14275
rect 15170 -14395 15290 -14275
rect 15335 -14395 15455 -14275
rect 15500 -14395 15620 -14275
rect 15675 -14395 15795 -14275
rect 15840 -14395 15960 -14275
rect 16005 -14395 16125 -14275
rect 16170 -14395 16290 -14275
rect 16345 -14395 16465 -14275
rect 16510 -14395 16630 -14275
rect 16675 -14395 16795 -14275
rect 16840 -14395 16960 -14275
rect 17015 -14395 17135 -14275
rect 17180 -14395 17300 -14275
rect 17345 -14395 17465 -14275
rect 17510 -14395 17630 -14275
rect 17685 -14395 17805 -14275
rect 17850 -14395 17970 -14275
rect 18015 -14395 18135 -14275
rect 18180 -14395 18300 -14275
rect 12820 -14560 12940 -14440
rect 12995 -14560 13115 -14440
rect 13160 -14560 13280 -14440
rect 13325 -14560 13445 -14440
rect 13490 -14560 13610 -14440
rect 13665 -14560 13785 -14440
rect 13830 -14560 13950 -14440
rect 13995 -14560 14115 -14440
rect 14160 -14560 14280 -14440
rect 14335 -14560 14455 -14440
rect 14500 -14560 14620 -14440
rect 14665 -14560 14785 -14440
rect 14830 -14560 14950 -14440
rect 15005 -14560 15125 -14440
rect 15170 -14560 15290 -14440
rect 15335 -14560 15455 -14440
rect 15500 -14560 15620 -14440
rect 15675 -14560 15795 -14440
rect 15840 -14560 15960 -14440
rect 16005 -14560 16125 -14440
rect 16170 -14560 16290 -14440
rect 16345 -14560 16465 -14440
rect 16510 -14560 16630 -14440
rect 16675 -14560 16795 -14440
rect 16840 -14560 16960 -14440
rect 17015 -14560 17135 -14440
rect 17180 -14560 17300 -14440
rect 17345 -14560 17465 -14440
rect 17510 -14560 17630 -14440
rect 17685 -14560 17805 -14440
rect 17850 -14560 17970 -14440
rect 18015 -14560 18135 -14440
rect 18180 -14560 18300 -14440
rect 12820 -14725 12940 -14605
rect 12995 -14725 13115 -14605
rect 13160 -14725 13280 -14605
rect 13325 -14725 13445 -14605
rect 13490 -14725 13610 -14605
rect 13665 -14725 13785 -14605
rect 13830 -14725 13950 -14605
rect 13995 -14725 14115 -14605
rect 14160 -14725 14280 -14605
rect 14335 -14725 14455 -14605
rect 14500 -14725 14620 -14605
rect 14665 -14725 14785 -14605
rect 14830 -14725 14950 -14605
rect 15005 -14725 15125 -14605
rect 15170 -14725 15290 -14605
rect 15335 -14725 15455 -14605
rect 15500 -14725 15620 -14605
rect 15675 -14725 15795 -14605
rect 15840 -14725 15960 -14605
rect 16005 -14725 16125 -14605
rect 16170 -14725 16290 -14605
rect 16345 -14725 16465 -14605
rect 16510 -14725 16630 -14605
rect 16675 -14725 16795 -14605
rect 16840 -14725 16960 -14605
rect 17015 -14725 17135 -14605
rect 17180 -14725 17300 -14605
rect 17345 -14725 17465 -14605
rect 17510 -14725 17630 -14605
rect 17685 -14725 17805 -14605
rect 17850 -14725 17970 -14605
rect 18015 -14725 18135 -14605
rect 18180 -14725 18300 -14605
rect 12820 -14900 12940 -14780
rect 12995 -14900 13115 -14780
rect 13160 -14900 13280 -14780
rect 13325 -14900 13445 -14780
rect 13490 -14900 13610 -14780
rect 13665 -14900 13785 -14780
rect 13830 -14900 13950 -14780
rect 13995 -14900 14115 -14780
rect 14160 -14900 14280 -14780
rect 14335 -14900 14455 -14780
rect 14500 -14900 14620 -14780
rect 14665 -14900 14785 -14780
rect 14830 -14900 14950 -14780
rect 15005 -14900 15125 -14780
rect 15170 -14900 15290 -14780
rect 15335 -14900 15455 -14780
rect 15500 -14900 15620 -14780
rect 15675 -14900 15795 -14780
rect 15840 -14900 15960 -14780
rect 16005 -14900 16125 -14780
rect 16170 -14900 16290 -14780
rect 16345 -14900 16465 -14780
rect 16510 -14900 16630 -14780
rect 16675 -14900 16795 -14780
rect 16840 -14900 16960 -14780
rect 17015 -14900 17135 -14780
rect 17180 -14900 17300 -14780
rect 17345 -14900 17465 -14780
rect 17510 -14900 17630 -14780
rect 17685 -14900 17805 -14780
rect 17850 -14900 17970 -14780
rect 18015 -14900 18135 -14780
rect 18180 -14900 18300 -14780
rect 12820 -15065 12940 -14945
rect 12995 -15065 13115 -14945
rect 13160 -15065 13280 -14945
rect 13325 -15065 13445 -14945
rect 13490 -15065 13610 -14945
rect 13665 -15065 13785 -14945
rect 13830 -15065 13950 -14945
rect 13995 -15065 14115 -14945
rect 14160 -15065 14280 -14945
rect 14335 -15065 14455 -14945
rect 14500 -15065 14620 -14945
rect 14665 -15065 14785 -14945
rect 14830 -15065 14950 -14945
rect 15005 -15065 15125 -14945
rect 15170 -15065 15290 -14945
rect 15335 -15065 15455 -14945
rect 15500 -15065 15620 -14945
rect 15675 -15065 15795 -14945
rect 15840 -15065 15960 -14945
rect 16005 -15065 16125 -14945
rect 16170 -15065 16290 -14945
rect 16345 -15065 16465 -14945
rect 16510 -15065 16630 -14945
rect 16675 -15065 16795 -14945
rect 16840 -15065 16960 -14945
rect 17015 -15065 17135 -14945
rect 17180 -15065 17300 -14945
rect 17345 -15065 17465 -14945
rect 17510 -15065 17630 -14945
rect 17685 -15065 17805 -14945
rect 17850 -15065 17970 -14945
rect 18015 -15065 18135 -14945
rect 18180 -15065 18300 -14945
rect 12820 -15230 12940 -15110
rect 12995 -15230 13115 -15110
rect 13160 -15230 13280 -15110
rect 13325 -15230 13445 -15110
rect 13490 -15230 13610 -15110
rect 13665 -15230 13785 -15110
rect 13830 -15230 13950 -15110
rect 13995 -15230 14115 -15110
rect 14160 -15230 14280 -15110
rect 14335 -15230 14455 -15110
rect 14500 -15230 14620 -15110
rect 14665 -15230 14785 -15110
rect 14830 -15230 14950 -15110
rect 15005 -15230 15125 -15110
rect 15170 -15230 15290 -15110
rect 15335 -15230 15455 -15110
rect 15500 -15230 15620 -15110
rect 15675 -15230 15795 -15110
rect 15840 -15230 15960 -15110
rect 16005 -15230 16125 -15110
rect 16170 -15230 16290 -15110
rect 16345 -15230 16465 -15110
rect 16510 -15230 16630 -15110
rect 16675 -15230 16795 -15110
rect 16840 -15230 16960 -15110
rect 17015 -15230 17135 -15110
rect 17180 -15230 17300 -15110
rect 17345 -15230 17465 -15110
rect 17510 -15230 17630 -15110
rect 17685 -15230 17805 -15110
rect 17850 -15230 17970 -15110
rect 18015 -15230 18135 -15110
rect 18180 -15230 18300 -15110
rect 12820 -15395 12940 -15275
rect 12995 -15395 13115 -15275
rect 13160 -15395 13280 -15275
rect 13325 -15395 13445 -15275
rect 13490 -15395 13610 -15275
rect 13665 -15395 13785 -15275
rect 13830 -15395 13950 -15275
rect 13995 -15395 14115 -15275
rect 14160 -15395 14280 -15275
rect 14335 -15395 14455 -15275
rect 14500 -15395 14620 -15275
rect 14665 -15395 14785 -15275
rect 14830 -15395 14950 -15275
rect 15005 -15395 15125 -15275
rect 15170 -15395 15290 -15275
rect 15335 -15395 15455 -15275
rect 15500 -15395 15620 -15275
rect 15675 -15395 15795 -15275
rect 15840 -15395 15960 -15275
rect 16005 -15395 16125 -15275
rect 16170 -15395 16290 -15275
rect 16345 -15395 16465 -15275
rect 16510 -15395 16630 -15275
rect 16675 -15395 16795 -15275
rect 16840 -15395 16960 -15275
rect 17015 -15395 17135 -15275
rect 17180 -15395 17300 -15275
rect 17345 -15395 17465 -15275
rect 17510 -15395 17630 -15275
rect 17685 -15395 17805 -15275
rect 17850 -15395 17970 -15275
rect 18015 -15395 18135 -15275
rect 18180 -15395 18300 -15275
rect 12820 -15570 12940 -15450
rect 12995 -15570 13115 -15450
rect 13160 -15570 13280 -15450
rect 13325 -15570 13445 -15450
rect 13490 -15570 13610 -15450
rect 13665 -15570 13785 -15450
rect 13830 -15570 13950 -15450
rect 13995 -15570 14115 -15450
rect 14160 -15570 14280 -15450
rect 14335 -15570 14455 -15450
rect 14500 -15570 14620 -15450
rect 14665 -15570 14785 -15450
rect 14830 -15570 14950 -15450
rect 15005 -15570 15125 -15450
rect 15170 -15570 15290 -15450
rect 15335 -15570 15455 -15450
rect 15500 -15570 15620 -15450
rect 15675 -15570 15795 -15450
rect 15840 -15570 15960 -15450
rect 16005 -15570 16125 -15450
rect 16170 -15570 16290 -15450
rect 16345 -15570 16465 -15450
rect 16510 -15570 16630 -15450
rect 16675 -15570 16795 -15450
rect 16840 -15570 16960 -15450
rect 17015 -15570 17135 -15450
rect 17180 -15570 17300 -15450
rect 17345 -15570 17465 -15450
rect 17510 -15570 17630 -15450
rect 17685 -15570 17805 -15450
rect 17850 -15570 17970 -15450
rect 18015 -15570 18135 -15450
rect 18180 -15570 18300 -15450
rect 18510 -10210 18630 -10090
rect 18685 -10210 18805 -10090
rect 18850 -10210 18970 -10090
rect 19015 -10210 19135 -10090
rect 19180 -10210 19300 -10090
rect 19355 -10210 19475 -10090
rect 19520 -10210 19640 -10090
rect 19685 -10210 19805 -10090
rect 19850 -10210 19970 -10090
rect 20025 -10210 20145 -10090
rect 20190 -10210 20310 -10090
rect 20355 -10210 20475 -10090
rect 20520 -10210 20640 -10090
rect 20695 -10210 20815 -10090
rect 20860 -10210 20980 -10090
rect 21025 -10210 21145 -10090
rect 21190 -10210 21310 -10090
rect 21365 -10210 21485 -10090
rect 21530 -10210 21650 -10090
rect 21695 -10210 21815 -10090
rect 21860 -10210 21980 -10090
rect 22035 -10210 22155 -10090
rect 22200 -10210 22320 -10090
rect 22365 -10210 22485 -10090
rect 22530 -10210 22650 -10090
rect 22705 -10210 22825 -10090
rect 22870 -10210 22990 -10090
rect 23035 -10210 23155 -10090
rect 23200 -10210 23320 -10090
rect 23375 -10210 23495 -10090
rect 23540 -10210 23660 -10090
rect 23705 -10210 23825 -10090
rect 23870 -10210 23990 -10090
rect 18510 -10375 18630 -10255
rect 18685 -10375 18805 -10255
rect 18850 -10375 18970 -10255
rect 19015 -10375 19135 -10255
rect 19180 -10375 19300 -10255
rect 19355 -10375 19475 -10255
rect 19520 -10375 19640 -10255
rect 19685 -10375 19805 -10255
rect 19850 -10375 19970 -10255
rect 20025 -10375 20145 -10255
rect 20190 -10375 20310 -10255
rect 20355 -10375 20475 -10255
rect 20520 -10375 20640 -10255
rect 20695 -10375 20815 -10255
rect 20860 -10375 20980 -10255
rect 21025 -10375 21145 -10255
rect 21190 -10375 21310 -10255
rect 21365 -10375 21485 -10255
rect 21530 -10375 21650 -10255
rect 21695 -10375 21815 -10255
rect 21860 -10375 21980 -10255
rect 22035 -10375 22155 -10255
rect 22200 -10375 22320 -10255
rect 22365 -10375 22485 -10255
rect 22530 -10375 22650 -10255
rect 22705 -10375 22825 -10255
rect 22870 -10375 22990 -10255
rect 23035 -10375 23155 -10255
rect 23200 -10375 23320 -10255
rect 23375 -10375 23495 -10255
rect 23540 -10375 23660 -10255
rect 23705 -10375 23825 -10255
rect 23870 -10375 23990 -10255
rect 18510 -10540 18630 -10420
rect 18685 -10540 18805 -10420
rect 18850 -10540 18970 -10420
rect 19015 -10540 19135 -10420
rect 19180 -10540 19300 -10420
rect 19355 -10540 19475 -10420
rect 19520 -10540 19640 -10420
rect 19685 -10540 19805 -10420
rect 19850 -10540 19970 -10420
rect 20025 -10540 20145 -10420
rect 20190 -10540 20310 -10420
rect 20355 -10540 20475 -10420
rect 20520 -10540 20640 -10420
rect 20695 -10540 20815 -10420
rect 20860 -10540 20980 -10420
rect 21025 -10540 21145 -10420
rect 21190 -10540 21310 -10420
rect 21365 -10540 21485 -10420
rect 21530 -10540 21650 -10420
rect 21695 -10540 21815 -10420
rect 21860 -10540 21980 -10420
rect 22035 -10540 22155 -10420
rect 22200 -10540 22320 -10420
rect 22365 -10540 22485 -10420
rect 22530 -10540 22650 -10420
rect 22705 -10540 22825 -10420
rect 22870 -10540 22990 -10420
rect 23035 -10540 23155 -10420
rect 23200 -10540 23320 -10420
rect 23375 -10540 23495 -10420
rect 23540 -10540 23660 -10420
rect 23705 -10540 23825 -10420
rect 23870 -10540 23990 -10420
rect 18510 -10705 18630 -10585
rect 18685 -10705 18805 -10585
rect 18850 -10705 18970 -10585
rect 19015 -10705 19135 -10585
rect 19180 -10705 19300 -10585
rect 19355 -10705 19475 -10585
rect 19520 -10705 19640 -10585
rect 19685 -10705 19805 -10585
rect 19850 -10705 19970 -10585
rect 20025 -10705 20145 -10585
rect 20190 -10705 20310 -10585
rect 20355 -10705 20475 -10585
rect 20520 -10705 20640 -10585
rect 20695 -10705 20815 -10585
rect 20860 -10705 20980 -10585
rect 21025 -10705 21145 -10585
rect 21190 -10705 21310 -10585
rect 21365 -10705 21485 -10585
rect 21530 -10705 21650 -10585
rect 21695 -10705 21815 -10585
rect 21860 -10705 21980 -10585
rect 22035 -10705 22155 -10585
rect 22200 -10705 22320 -10585
rect 22365 -10705 22485 -10585
rect 22530 -10705 22650 -10585
rect 22705 -10705 22825 -10585
rect 22870 -10705 22990 -10585
rect 23035 -10705 23155 -10585
rect 23200 -10705 23320 -10585
rect 23375 -10705 23495 -10585
rect 23540 -10705 23660 -10585
rect 23705 -10705 23825 -10585
rect 23870 -10705 23990 -10585
rect 18510 -10880 18630 -10760
rect 18685 -10880 18805 -10760
rect 18850 -10880 18970 -10760
rect 19015 -10880 19135 -10760
rect 19180 -10880 19300 -10760
rect 19355 -10880 19475 -10760
rect 19520 -10880 19640 -10760
rect 19685 -10880 19805 -10760
rect 19850 -10880 19970 -10760
rect 20025 -10880 20145 -10760
rect 20190 -10880 20310 -10760
rect 20355 -10880 20475 -10760
rect 20520 -10880 20640 -10760
rect 20695 -10880 20815 -10760
rect 20860 -10880 20980 -10760
rect 21025 -10880 21145 -10760
rect 21190 -10880 21310 -10760
rect 21365 -10880 21485 -10760
rect 21530 -10880 21650 -10760
rect 21695 -10880 21815 -10760
rect 21860 -10880 21980 -10760
rect 22035 -10880 22155 -10760
rect 22200 -10880 22320 -10760
rect 22365 -10880 22485 -10760
rect 22530 -10880 22650 -10760
rect 22705 -10880 22825 -10760
rect 22870 -10880 22990 -10760
rect 23035 -10880 23155 -10760
rect 23200 -10880 23320 -10760
rect 23375 -10880 23495 -10760
rect 23540 -10880 23660 -10760
rect 23705 -10880 23825 -10760
rect 23870 -10880 23990 -10760
rect 18510 -11045 18630 -10925
rect 18685 -11045 18805 -10925
rect 18850 -11045 18970 -10925
rect 19015 -11045 19135 -10925
rect 19180 -11045 19300 -10925
rect 19355 -11045 19475 -10925
rect 19520 -11045 19640 -10925
rect 19685 -11045 19805 -10925
rect 19850 -11045 19970 -10925
rect 20025 -11045 20145 -10925
rect 20190 -11045 20310 -10925
rect 20355 -11045 20475 -10925
rect 20520 -11045 20640 -10925
rect 20695 -11045 20815 -10925
rect 20860 -11045 20980 -10925
rect 21025 -11045 21145 -10925
rect 21190 -11045 21310 -10925
rect 21365 -11045 21485 -10925
rect 21530 -11045 21650 -10925
rect 21695 -11045 21815 -10925
rect 21860 -11045 21980 -10925
rect 22035 -11045 22155 -10925
rect 22200 -11045 22320 -10925
rect 22365 -11045 22485 -10925
rect 22530 -11045 22650 -10925
rect 22705 -11045 22825 -10925
rect 22870 -11045 22990 -10925
rect 23035 -11045 23155 -10925
rect 23200 -11045 23320 -10925
rect 23375 -11045 23495 -10925
rect 23540 -11045 23660 -10925
rect 23705 -11045 23825 -10925
rect 23870 -11045 23990 -10925
rect 18510 -11210 18630 -11090
rect 18685 -11210 18805 -11090
rect 18850 -11210 18970 -11090
rect 19015 -11210 19135 -11090
rect 19180 -11210 19300 -11090
rect 19355 -11210 19475 -11090
rect 19520 -11210 19640 -11090
rect 19685 -11210 19805 -11090
rect 19850 -11210 19970 -11090
rect 20025 -11210 20145 -11090
rect 20190 -11210 20310 -11090
rect 20355 -11210 20475 -11090
rect 20520 -11210 20640 -11090
rect 20695 -11210 20815 -11090
rect 20860 -11210 20980 -11090
rect 21025 -11210 21145 -11090
rect 21190 -11210 21310 -11090
rect 21365 -11210 21485 -11090
rect 21530 -11210 21650 -11090
rect 21695 -11210 21815 -11090
rect 21860 -11210 21980 -11090
rect 22035 -11210 22155 -11090
rect 22200 -11210 22320 -11090
rect 22365 -11210 22485 -11090
rect 22530 -11210 22650 -11090
rect 22705 -11210 22825 -11090
rect 22870 -11210 22990 -11090
rect 23035 -11210 23155 -11090
rect 23200 -11210 23320 -11090
rect 23375 -11210 23495 -11090
rect 23540 -11210 23660 -11090
rect 23705 -11210 23825 -11090
rect 23870 -11210 23990 -11090
rect 18510 -11375 18630 -11255
rect 18685 -11375 18805 -11255
rect 18850 -11375 18970 -11255
rect 19015 -11375 19135 -11255
rect 19180 -11375 19300 -11255
rect 19355 -11375 19475 -11255
rect 19520 -11375 19640 -11255
rect 19685 -11375 19805 -11255
rect 19850 -11375 19970 -11255
rect 20025 -11375 20145 -11255
rect 20190 -11375 20310 -11255
rect 20355 -11375 20475 -11255
rect 20520 -11375 20640 -11255
rect 20695 -11375 20815 -11255
rect 20860 -11375 20980 -11255
rect 21025 -11375 21145 -11255
rect 21190 -11375 21310 -11255
rect 21365 -11375 21485 -11255
rect 21530 -11375 21650 -11255
rect 21695 -11375 21815 -11255
rect 21860 -11375 21980 -11255
rect 22035 -11375 22155 -11255
rect 22200 -11375 22320 -11255
rect 22365 -11375 22485 -11255
rect 22530 -11375 22650 -11255
rect 22705 -11375 22825 -11255
rect 22870 -11375 22990 -11255
rect 23035 -11375 23155 -11255
rect 23200 -11375 23320 -11255
rect 23375 -11375 23495 -11255
rect 23540 -11375 23660 -11255
rect 23705 -11375 23825 -11255
rect 23870 -11375 23990 -11255
rect 18510 -11550 18630 -11430
rect 18685 -11550 18805 -11430
rect 18850 -11550 18970 -11430
rect 19015 -11550 19135 -11430
rect 19180 -11550 19300 -11430
rect 19355 -11550 19475 -11430
rect 19520 -11550 19640 -11430
rect 19685 -11550 19805 -11430
rect 19850 -11550 19970 -11430
rect 20025 -11550 20145 -11430
rect 20190 -11550 20310 -11430
rect 20355 -11550 20475 -11430
rect 20520 -11550 20640 -11430
rect 20695 -11550 20815 -11430
rect 20860 -11550 20980 -11430
rect 21025 -11550 21145 -11430
rect 21190 -11550 21310 -11430
rect 21365 -11550 21485 -11430
rect 21530 -11550 21650 -11430
rect 21695 -11550 21815 -11430
rect 21860 -11550 21980 -11430
rect 22035 -11550 22155 -11430
rect 22200 -11550 22320 -11430
rect 22365 -11550 22485 -11430
rect 22530 -11550 22650 -11430
rect 22705 -11550 22825 -11430
rect 22870 -11550 22990 -11430
rect 23035 -11550 23155 -11430
rect 23200 -11550 23320 -11430
rect 23375 -11550 23495 -11430
rect 23540 -11550 23660 -11430
rect 23705 -11550 23825 -11430
rect 23870 -11550 23990 -11430
rect 18510 -11715 18630 -11595
rect 18685 -11715 18805 -11595
rect 18850 -11715 18970 -11595
rect 19015 -11715 19135 -11595
rect 19180 -11715 19300 -11595
rect 19355 -11715 19475 -11595
rect 19520 -11715 19640 -11595
rect 19685 -11715 19805 -11595
rect 19850 -11715 19970 -11595
rect 20025 -11715 20145 -11595
rect 20190 -11715 20310 -11595
rect 20355 -11715 20475 -11595
rect 20520 -11715 20640 -11595
rect 20695 -11715 20815 -11595
rect 20860 -11715 20980 -11595
rect 21025 -11715 21145 -11595
rect 21190 -11715 21310 -11595
rect 21365 -11715 21485 -11595
rect 21530 -11715 21650 -11595
rect 21695 -11715 21815 -11595
rect 21860 -11715 21980 -11595
rect 22035 -11715 22155 -11595
rect 22200 -11715 22320 -11595
rect 22365 -11715 22485 -11595
rect 22530 -11715 22650 -11595
rect 22705 -11715 22825 -11595
rect 22870 -11715 22990 -11595
rect 23035 -11715 23155 -11595
rect 23200 -11715 23320 -11595
rect 23375 -11715 23495 -11595
rect 23540 -11715 23660 -11595
rect 23705 -11715 23825 -11595
rect 23870 -11715 23990 -11595
rect 18510 -11880 18630 -11760
rect 18685 -11880 18805 -11760
rect 18850 -11880 18970 -11760
rect 19015 -11880 19135 -11760
rect 19180 -11880 19300 -11760
rect 19355 -11880 19475 -11760
rect 19520 -11880 19640 -11760
rect 19685 -11880 19805 -11760
rect 19850 -11880 19970 -11760
rect 20025 -11880 20145 -11760
rect 20190 -11880 20310 -11760
rect 20355 -11880 20475 -11760
rect 20520 -11880 20640 -11760
rect 20695 -11880 20815 -11760
rect 20860 -11880 20980 -11760
rect 21025 -11880 21145 -11760
rect 21190 -11880 21310 -11760
rect 21365 -11880 21485 -11760
rect 21530 -11880 21650 -11760
rect 21695 -11880 21815 -11760
rect 21860 -11880 21980 -11760
rect 22035 -11880 22155 -11760
rect 22200 -11880 22320 -11760
rect 22365 -11880 22485 -11760
rect 22530 -11880 22650 -11760
rect 22705 -11880 22825 -11760
rect 22870 -11880 22990 -11760
rect 23035 -11880 23155 -11760
rect 23200 -11880 23320 -11760
rect 23375 -11880 23495 -11760
rect 23540 -11880 23660 -11760
rect 23705 -11880 23825 -11760
rect 23870 -11880 23990 -11760
rect 18510 -12045 18630 -11925
rect 18685 -12045 18805 -11925
rect 18850 -12045 18970 -11925
rect 19015 -12045 19135 -11925
rect 19180 -12045 19300 -11925
rect 19355 -12045 19475 -11925
rect 19520 -12045 19640 -11925
rect 19685 -12045 19805 -11925
rect 19850 -12045 19970 -11925
rect 20025 -12045 20145 -11925
rect 20190 -12045 20310 -11925
rect 20355 -12045 20475 -11925
rect 20520 -12045 20640 -11925
rect 20695 -12045 20815 -11925
rect 20860 -12045 20980 -11925
rect 21025 -12045 21145 -11925
rect 21190 -12045 21310 -11925
rect 21365 -12045 21485 -11925
rect 21530 -12045 21650 -11925
rect 21695 -12045 21815 -11925
rect 21860 -12045 21980 -11925
rect 22035 -12045 22155 -11925
rect 22200 -12045 22320 -11925
rect 22365 -12045 22485 -11925
rect 22530 -12045 22650 -11925
rect 22705 -12045 22825 -11925
rect 22870 -12045 22990 -11925
rect 23035 -12045 23155 -11925
rect 23200 -12045 23320 -11925
rect 23375 -12045 23495 -11925
rect 23540 -12045 23660 -11925
rect 23705 -12045 23825 -11925
rect 23870 -12045 23990 -11925
rect 18510 -12220 18630 -12100
rect 18685 -12220 18805 -12100
rect 18850 -12220 18970 -12100
rect 19015 -12220 19135 -12100
rect 19180 -12220 19300 -12100
rect 19355 -12220 19475 -12100
rect 19520 -12220 19640 -12100
rect 19685 -12220 19805 -12100
rect 19850 -12220 19970 -12100
rect 20025 -12220 20145 -12100
rect 20190 -12220 20310 -12100
rect 20355 -12220 20475 -12100
rect 20520 -12220 20640 -12100
rect 20695 -12220 20815 -12100
rect 20860 -12220 20980 -12100
rect 21025 -12220 21145 -12100
rect 21190 -12220 21310 -12100
rect 21365 -12220 21485 -12100
rect 21530 -12220 21650 -12100
rect 21695 -12220 21815 -12100
rect 21860 -12220 21980 -12100
rect 22035 -12220 22155 -12100
rect 22200 -12220 22320 -12100
rect 22365 -12220 22485 -12100
rect 22530 -12220 22650 -12100
rect 22705 -12220 22825 -12100
rect 22870 -12220 22990 -12100
rect 23035 -12220 23155 -12100
rect 23200 -12220 23320 -12100
rect 23375 -12220 23495 -12100
rect 23540 -12220 23660 -12100
rect 23705 -12220 23825 -12100
rect 23870 -12220 23990 -12100
rect 18510 -12385 18630 -12265
rect 18685 -12385 18805 -12265
rect 18850 -12385 18970 -12265
rect 19015 -12385 19135 -12265
rect 19180 -12385 19300 -12265
rect 19355 -12385 19475 -12265
rect 19520 -12385 19640 -12265
rect 19685 -12385 19805 -12265
rect 19850 -12385 19970 -12265
rect 20025 -12385 20145 -12265
rect 20190 -12385 20310 -12265
rect 20355 -12385 20475 -12265
rect 20520 -12385 20640 -12265
rect 20695 -12385 20815 -12265
rect 20860 -12385 20980 -12265
rect 21025 -12385 21145 -12265
rect 21190 -12385 21310 -12265
rect 21365 -12385 21485 -12265
rect 21530 -12385 21650 -12265
rect 21695 -12385 21815 -12265
rect 21860 -12385 21980 -12265
rect 22035 -12385 22155 -12265
rect 22200 -12385 22320 -12265
rect 22365 -12385 22485 -12265
rect 22530 -12385 22650 -12265
rect 22705 -12385 22825 -12265
rect 22870 -12385 22990 -12265
rect 23035 -12385 23155 -12265
rect 23200 -12385 23320 -12265
rect 23375 -12385 23495 -12265
rect 23540 -12385 23660 -12265
rect 23705 -12385 23825 -12265
rect 23870 -12385 23990 -12265
rect 18510 -12550 18630 -12430
rect 18685 -12550 18805 -12430
rect 18850 -12550 18970 -12430
rect 19015 -12550 19135 -12430
rect 19180 -12550 19300 -12430
rect 19355 -12550 19475 -12430
rect 19520 -12550 19640 -12430
rect 19685 -12550 19805 -12430
rect 19850 -12550 19970 -12430
rect 20025 -12550 20145 -12430
rect 20190 -12550 20310 -12430
rect 20355 -12550 20475 -12430
rect 20520 -12550 20640 -12430
rect 20695 -12550 20815 -12430
rect 20860 -12550 20980 -12430
rect 21025 -12550 21145 -12430
rect 21190 -12550 21310 -12430
rect 21365 -12550 21485 -12430
rect 21530 -12550 21650 -12430
rect 21695 -12550 21815 -12430
rect 21860 -12550 21980 -12430
rect 22035 -12550 22155 -12430
rect 22200 -12550 22320 -12430
rect 22365 -12550 22485 -12430
rect 22530 -12550 22650 -12430
rect 22705 -12550 22825 -12430
rect 22870 -12550 22990 -12430
rect 23035 -12550 23155 -12430
rect 23200 -12550 23320 -12430
rect 23375 -12550 23495 -12430
rect 23540 -12550 23660 -12430
rect 23705 -12550 23825 -12430
rect 23870 -12550 23990 -12430
rect 18510 -12715 18630 -12595
rect 18685 -12715 18805 -12595
rect 18850 -12715 18970 -12595
rect 19015 -12715 19135 -12595
rect 19180 -12715 19300 -12595
rect 19355 -12715 19475 -12595
rect 19520 -12715 19640 -12595
rect 19685 -12715 19805 -12595
rect 19850 -12715 19970 -12595
rect 20025 -12715 20145 -12595
rect 20190 -12715 20310 -12595
rect 20355 -12715 20475 -12595
rect 20520 -12715 20640 -12595
rect 20695 -12715 20815 -12595
rect 20860 -12715 20980 -12595
rect 21025 -12715 21145 -12595
rect 21190 -12715 21310 -12595
rect 21365 -12715 21485 -12595
rect 21530 -12715 21650 -12595
rect 21695 -12715 21815 -12595
rect 21860 -12715 21980 -12595
rect 22035 -12715 22155 -12595
rect 22200 -12715 22320 -12595
rect 22365 -12715 22485 -12595
rect 22530 -12715 22650 -12595
rect 22705 -12715 22825 -12595
rect 22870 -12715 22990 -12595
rect 23035 -12715 23155 -12595
rect 23200 -12715 23320 -12595
rect 23375 -12715 23495 -12595
rect 23540 -12715 23660 -12595
rect 23705 -12715 23825 -12595
rect 23870 -12715 23990 -12595
rect 18510 -12890 18630 -12770
rect 18685 -12890 18805 -12770
rect 18850 -12890 18970 -12770
rect 19015 -12890 19135 -12770
rect 19180 -12890 19300 -12770
rect 19355 -12890 19475 -12770
rect 19520 -12890 19640 -12770
rect 19685 -12890 19805 -12770
rect 19850 -12890 19970 -12770
rect 20025 -12890 20145 -12770
rect 20190 -12890 20310 -12770
rect 20355 -12890 20475 -12770
rect 20520 -12890 20640 -12770
rect 20695 -12890 20815 -12770
rect 20860 -12890 20980 -12770
rect 21025 -12890 21145 -12770
rect 21190 -12890 21310 -12770
rect 21365 -12890 21485 -12770
rect 21530 -12890 21650 -12770
rect 21695 -12890 21815 -12770
rect 21860 -12890 21980 -12770
rect 22035 -12890 22155 -12770
rect 22200 -12890 22320 -12770
rect 22365 -12890 22485 -12770
rect 22530 -12890 22650 -12770
rect 22705 -12890 22825 -12770
rect 22870 -12890 22990 -12770
rect 23035 -12890 23155 -12770
rect 23200 -12890 23320 -12770
rect 23375 -12890 23495 -12770
rect 23540 -12890 23660 -12770
rect 23705 -12890 23825 -12770
rect 23870 -12890 23990 -12770
rect 18510 -13055 18630 -12935
rect 18685 -13055 18805 -12935
rect 18850 -13055 18970 -12935
rect 19015 -13055 19135 -12935
rect 19180 -13055 19300 -12935
rect 19355 -13055 19475 -12935
rect 19520 -13055 19640 -12935
rect 19685 -13055 19805 -12935
rect 19850 -13055 19970 -12935
rect 20025 -13055 20145 -12935
rect 20190 -13055 20310 -12935
rect 20355 -13055 20475 -12935
rect 20520 -13055 20640 -12935
rect 20695 -13055 20815 -12935
rect 20860 -13055 20980 -12935
rect 21025 -13055 21145 -12935
rect 21190 -13055 21310 -12935
rect 21365 -13055 21485 -12935
rect 21530 -13055 21650 -12935
rect 21695 -13055 21815 -12935
rect 21860 -13055 21980 -12935
rect 22035 -13055 22155 -12935
rect 22200 -13055 22320 -12935
rect 22365 -13055 22485 -12935
rect 22530 -13055 22650 -12935
rect 22705 -13055 22825 -12935
rect 22870 -13055 22990 -12935
rect 23035 -13055 23155 -12935
rect 23200 -13055 23320 -12935
rect 23375 -13055 23495 -12935
rect 23540 -13055 23660 -12935
rect 23705 -13055 23825 -12935
rect 23870 -13055 23990 -12935
rect 18510 -13220 18630 -13100
rect 18685 -13220 18805 -13100
rect 18850 -13220 18970 -13100
rect 19015 -13220 19135 -13100
rect 19180 -13220 19300 -13100
rect 19355 -13220 19475 -13100
rect 19520 -13220 19640 -13100
rect 19685 -13220 19805 -13100
rect 19850 -13220 19970 -13100
rect 20025 -13220 20145 -13100
rect 20190 -13220 20310 -13100
rect 20355 -13220 20475 -13100
rect 20520 -13220 20640 -13100
rect 20695 -13220 20815 -13100
rect 20860 -13220 20980 -13100
rect 21025 -13220 21145 -13100
rect 21190 -13220 21310 -13100
rect 21365 -13220 21485 -13100
rect 21530 -13220 21650 -13100
rect 21695 -13220 21815 -13100
rect 21860 -13220 21980 -13100
rect 22035 -13220 22155 -13100
rect 22200 -13220 22320 -13100
rect 22365 -13220 22485 -13100
rect 22530 -13220 22650 -13100
rect 22705 -13220 22825 -13100
rect 22870 -13220 22990 -13100
rect 23035 -13220 23155 -13100
rect 23200 -13220 23320 -13100
rect 23375 -13220 23495 -13100
rect 23540 -13220 23660 -13100
rect 23705 -13220 23825 -13100
rect 23870 -13220 23990 -13100
rect 18510 -13385 18630 -13265
rect 18685 -13385 18805 -13265
rect 18850 -13385 18970 -13265
rect 19015 -13385 19135 -13265
rect 19180 -13385 19300 -13265
rect 19355 -13385 19475 -13265
rect 19520 -13385 19640 -13265
rect 19685 -13385 19805 -13265
rect 19850 -13385 19970 -13265
rect 20025 -13385 20145 -13265
rect 20190 -13385 20310 -13265
rect 20355 -13385 20475 -13265
rect 20520 -13385 20640 -13265
rect 20695 -13385 20815 -13265
rect 20860 -13385 20980 -13265
rect 21025 -13385 21145 -13265
rect 21190 -13385 21310 -13265
rect 21365 -13385 21485 -13265
rect 21530 -13385 21650 -13265
rect 21695 -13385 21815 -13265
rect 21860 -13385 21980 -13265
rect 22035 -13385 22155 -13265
rect 22200 -13385 22320 -13265
rect 22365 -13385 22485 -13265
rect 22530 -13385 22650 -13265
rect 22705 -13385 22825 -13265
rect 22870 -13385 22990 -13265
rect 23035 -13385 23155 -13265
rect 23200 -13385 23320 -13265
rect 23375 -13385 23495 -13265
rect 23540 -13385 23660 -13265
rect 23705 -13385 23825 -13265
rect 23870 -13385 23990 -13265
rect 18510 -13560 18630 -13440
rect 18685 -13560 18805 -13440
rect 18850 -13560 18970 -13440
rect 19015 -13560 19135 -13440
rect 19180 -13560 19300 -13440
rect 19355 -13560 19475 -13440
rect 19520 -13560 19640 -13440
rect 19685 -13560 19805 -13440
rect 19850 -13560 19970 -13440
rect 20025 -13560 20145 -13440
rect 20190 -13560 20310 -13440
rect 20355 -13560 20475 -13440
rect 20520 -13560 20640 -13440
rect 20695 -13560 20815 -13440
rect 20860 -13560 20980 -13440
rect 21025 -13560 21145 -13440
rect 21190 -13560 21310 -13440
rect 21365 -13560 21485 -13440
rect 21530 -13560 21650 -13440
rect 21695 -13560 21815 -13440
rect 21860 -13560 21980 -13440
rect 22035 -13560 22155 -13440
rect 22200 -13560 22320 -13440
rect 22365 -13560 22485 -13440
rect 22530 -13560 22650 -13440
rect 22705 -13560 22825 -13440
rect 22870 -13560 22990 -13440
rect 23035 -13560 23155 -13440
rect 23200 -13560 23320 -13440
rect 23375 -13560 23495 -13440
rect 23540 -13560 23660 -13440
rect 23705 -13560 23825 -13440
rect 23870 -13560 23990 -13440
rect 18510 -13725 18630 -13605
rect 18685 -13725 18805 -13605
rect 18850 -13725 18970 -13605
rect 19015 -13725 19135 -13605
rect 19180 -13725 19300 -13605
rect 19355 -13725 19475 -13605
rect 19520 -13725 19640 -13605
rect 19685 -13725 19805 -13605
rect 19850 -13725 19970 -13605
rect 20025 -13725 20145 -13605
rect 20190 -13725 20310 -13605
rect 20355 -13725 20475 -13605
rect 20520 -13725 20640 -13605
rect 20695 -13725 20815 -13605
rect 20860 -13725 20980 -13605
rect 21025 -13725 21145 -13605
rect 21190 -13725 21310 -13605
rect 21365 -13725 21485 -13605
rect 21530 -13725 21650 -13605
rect 21695 -13725 21815 -13605
rect 21860 -13725 21980 -13605
rect 22035 -13725 22155 -13605
rect 22200 -13725 22320 -13605
rect 22365 -13725 22485 -13605
rect 22530 -13725 22650 -13605
rect 22705 -13725 22825 -13605
rect 22870 -13725 22990 -13605
rect 23035 -13725 23155 -13605
rect 23200 -13725 23320 -13605
rect 23375 -13725 23495 -13605
rect 23540 -13725 23660 -13605
rect 23705 -13725 23825 -13605
rect 23870 -13725 23990 -13605
rect 18510 -13890 18630 -13770
rect 18685 -13890 18805 -13770
rect 18850 -13890 18970 -13770
rect 19015 -13890 19135 -13770
rect 19180 -13890 19300 -13770
rect 19355 -13890 19475 -13770
rect 19520 -13890 19640 -13770
rect 19685 -13890 19805 -13770
rect 19850 -13890 19970 -13770
rect 20025 -13890 20145 -13770
rect 20190 -13890 20310 -13770
rect 20355 -13890 20475 -13770
rect 20520 -13890 20640 -13770
rect 20695 -13890 20815 -13770
rect 20860 -13890 20980 -13770
rect 21025 -13890 21145 -13770
rect 21190 -13890 21310 -13770
rect 21365 -13890 21485 -13770
rect 21530 -13890 21650 -13770
rect 21695 -13890 21815 -13770
rect 21860 -13890 21980 -13770
rect 22035 -13890 22155 -13770
rect 22200 -13890 22320 -13770
rect 22365 -13890 22485 -13770
rect 22530 -13890 22650 -13770
rect 22705 -13890 22825 -13770
rect 22870 -13890 22990 -13770
rect 23035 -13890 23155 -13770
rect 23200 -13890 23320 -13770
rect 23375 -13890 23495 -13770
rect 23540 -13890 23660 -13770
rect 23705 -13890 23825 -13770
rect 23870 -13890 23990 -13770
rect 18510 -14055 18630 -13935
rect 18685 -14055 18805 -13935
rect 18850 -14055 18970 -13935
rect 19015 -14055 19135 -13935
rect 19180 -14055 19300 -13935
rect 19355 -14055 19475 -13935
rect 19520 -14055 19640 -13935
rect 19685 -14055 19805 -13935
rect 19850 -14055 19970 -13935
rect 20025 -14055 20145 -13935
rect 20190 -14055 20310 -13935
rect 20355 -14055 20475 -13935
rect 20520 -14055 20640 -13935
rect 20695 -14055 20815 -13935
rect 20860 -14055 20980 -13935
rect 21025 -14055 21145 -13935
rect 21190 -14055 21310 -13935
rect 21365 -14055 21485 -13935
rect 21530 -14055 21650 -13935
rect 21695 -14055 21815 -13935
rect 21860 -14055 21980 -13935
rect 22035 -14055 22155 -13935
rect 22200 -14055 22320 -13935
rect 22365 -14055 22485 -13935
rect 22530 -14055 22650 -13935
rect 22705 -14055 22825 -13935
rect 22870 -14055 22990 -13935
rect 23035 -14055 23155 -13935
rect 23200 -14055 23320 -13935
rect 23375 -14055 23495 -13935
rect 23540 -14055 23660 -13935
rect 23705 -14055 23825 -13935
rect 23870 -14055 23990 -13935
rect 18510 -14230 18630 -14110
rect 18685 -14230 18805 -14110
rect 18850 -14230 18970 -14110
rect 19015 -14230 19135 -14110
rect 19180 -14230 19300 -14110
rect 19355 -14230 19475 -14110
rect 19520 -14230 19640 -14110
rect 19685 -14230 19805 -14110
rect 19850 -14230 19970 -14110
rect 20025 -14230 20145 -14110
rect 20190 -14230 20310 -14110
rect 20355 -14230 20475 -14110
rect 20520 -14230 20640 -14110
rect 20695 -14230 20815 -14110
rect 20860 -14230 20980 -14110
rect 21025 -14230 21145 -14110
rect 21190 -14230 21310 -14110
rect 21365 -14230 21485 -14110
rect 21530 -14230 21650 -14110
rect 21695 -14230 21815 -14110
rect 21860 -14230 21980 -14110
rect 22035 -14230 22155 -14110
rect 22200 -14230 22320 -14110
rect 22365 -14230 22485 -14110
rect 22530 -14230 22650 -14110
rect 22705 -14230 22825 -14110
rect 22870 -14230 22990 -14110
rect 23035 -14230 23155 -14110
rect 23200 -14230 23320 -14110
rect 23375 -14230 23495 -14110
rect 23540 -14230 23660 -14110
rect 23705 -14230 23825 -14110
rect 23870 -14230 23990 -14110
rect 18510 -14395 18630 -14275
rect 18685 -14395 18805 -14275
rect 18850 -14395 18970 -14275
rect 19015 -14395 19135 -14275
rect 19180 -14395 19300 -14275
rect 19355 -14395 19475 -14275
rect 19520 -14395 19640 -14275
rect 19685 -14395 19805 -14275
rect 19850 -14395 19970 -14275
rect 20025 -14395 20145 -14275
rect 20190 -14395 20310 -14275
rect 20355 -14395 20475 -14275
rect 20520 -14395 20640 -14275
rect 20695 -14395 20815 -14275
rect 20860 -14395 20980 -14275
rect 21025 -14395 21145 -14275
rect 21190 -14395 21310 -14275
rect 21365 -14395 21485 -14275
rect 21530 -14395 21650 -14275
rect 21695 -14395 21815 -14275
rect 21860 -14395 21980 -14275
rect 22035 -14395 22155 -14275
rect 22200 -14395 22320 -14275
rect 22365 -14395 22485 -14275
rect 22530 -14395 22650 -14275
rect 22705 -14395 22825 -14275
rect 22870 -14395 22990 -14275
rect 23035 -14395 23155 -14275
rect 23200 -14395 23320 -14275
rect 23375 -14395 23495 -14275
rect 23540 -14395 23660 -14275
rect 23705 -14395 23825 -14275
rect 23870 -14395 23990 -14275
rect 18510 -14560 18630 -14440
rect 18685 -14560 18805 -14440
rect 18850 -14560 18970 -14440
rect 19015 -14560 19135 -14440
rect 19180 -14560 19300 -14440
rect 19355 -14560 19475 -14440
rect 19520 -14560 19640 -14440
rect 19685 -14560 19805 -14440
rect 19850 -14560 19970 -14440
rect 20025 -14560 20145 -14440
rect 20190 -14560 20310 -14440
rect 20355 -14560 20475 -14440
rect 20520 -14560 20640 -14440
rect 20695 -14560 20815 -14440
rect 20860 -14560 20980 -14440
rect 21025 -14560 21145 -14440
rect 21190 -14560 21310 -14440
rect 21365 -14560 21485 -14440
rect 21530 -14560 21650 -14440
rect 21695 -14560 21815 -14440
rect 21860 -14560 21980 -14440
rect 22035 -14560 22155 -14440
rect 22200 -14560 22320 -14440
rect 22365 -14560 22485 -14440
rect 22530 -14560 22650 -14440
rect 22705 -14560 22825 -14440
rect 22870 -14560 22990 -14440
rect 23035 -14560 23155 -14440
rect 23200 -14560 23320 -14440
rect 23375 -14560 23495 -14440
rect 23540 -14560 23660 -14440
rect 23705 -14560 23825 -14440
rect 23870 -14560 23990 -14440
rect 18510 -14725 18630 -14605
rect 18685 -14725 18805 -14605
rect 18850 -14725 18970 -14605
rect 19015 -14725 19135 -14605
rect 19180 -14725 19300 -14605
rect 19355 -14725 19475 -14605
rect 19520 -14725 19640 -14605
rect 19685 -14725 19805 -14605
rect 19850 -14725 19970 -14605
rect 20025 -14725 20145 -14605
rect 20190 -14725 20310 -14605
rect 20355 -14725 20475 -14605
rect 20520 -14725 20640 -14605
rect 20695 -14725 20815 -14605
rect 20860 -14725 20980 -14605
rect 21025 -14725 21145 -14605
rect 21190 -14725 21310 -14605
rect 21365 -14725 21485 -14605
rect 21530 -14725 21650 -14605
rect 21695 -14725 21815 -14605
rect 21860 -14725 21980 -14605
rect 22035 -14725 22155 -14605
rect 22200 -14725 22320 -14605
rect 22365 -14725 22485 -14605
rect 22530 -14725 22650 -14605
rect 22705 -14725 22825 -14605
rect 22870 -14725 22990 -14605
rect 23035 -14725 23155 -14605
rect 23200 -14725 23320 -14605
rect 23375 -14725 23495 -14605
rect 23540 -14725 23660 -14605
rect 23705 -14725 23825 -14605
rect 23870 -14725 23990 -14605
rect 18510 -14900 18630 -14780
rect 18685 -14900 18805 -14780
rect 18850 -14900 18970 -14780
rect 19015 -14900 19135 -14780
rect 19180 -14900 19300 -14780
rect 19355 -14900 19475 -14780
rect 19520 -14900 19640 -14780
rect 19685 -14900 19805 -14780
rect 19850 -14900 19970 -14780
rect 20025 -14900 20145 -14780
rect 20190 -14900 20310 -14780
rect 20355 -14900 20475 -14780
rect 20520 -14900 20640 -14780
rect 20695 -14900 20815 -14780
rect 20860 -14900 20980 -14780
rect 21025 -14900 21145 -14780
rect 21190 -14900 21310 -14780
rect 21365 -14900 21485 -14780
rect 21530 -14900 21650 -14780
rect 21695 -14900 21815 -14780
rect 21860 -14900 21980 -14780
rect 22035 -14900 22155 -14780
rect 22200 -14900 22320 -14780
rect 22365 -14900 22485 -14780
rect 22530 -14900 22650 -14780
rect 22705 -14900 22825 -14780
rect 22870 -14900 22990 -14780
rect 23035 -14900 23155 -14780
rect 23200 -14900 23320 -14780
rect 23375 -14900 23495 -14780
rect 23540 -14900 23660 -14780
rect 23705 -14900 23825 -14780
rect 23870 -14900 23990 -14780
rect 18510 -15065 18630 -14945
rect 18685 -15065 18805 -14945
rect 18850 -15065 18970 -14945
rect 19015 -15065 19135 -14945
rect 19180 -15065 19300 -14945
rect 19355 -15065 19475 -14945
rect 19520 -15065 19640 -14945
rect 19685 -15065 19805 -14945
rect 19850 -15065 19970 -14945
rect 20025 -15065 20145 -14945
rect 20190 -15065 20310 -14945
rect 20355 -15065 20475 -14945
rect 20520 -15065 20640 -14945
rect 20695 -15065 20815 -14945
rect 20860 -15065 20980 -14945
rect 21025 -15065 21145 -14945
rect 21190 -15065 21310 -14945
rect 21365 -15065 21485 -14945
rect 21530 -15065 21650 -14945
rect 21695 -15065 21815 -14945
rect 21860 -15065 21980 -14945
rect 22035 -15065 22155 -14945
rect 22200 -15065 22320 -14945
rect 22365 -15065 22485 -14945
rect 22530 -15065 22650 -14945
rect 22705 -15065 22825 -14945
rect 22870 -15065 22990 -14945
rect 23035 -15065 23155 -14945
rect 23200 -15065 23320 -14945
rect 23375 -15065 23495 -14945
rect 23540 -15065 23660 -14945
rect 23705 -15065 23825 -14945
rect 23870 -15065 23990 -14945
rect 18510 -15230 18630 -15110
rect 18685 -15230 18805 -15110
rect 18850 -15230 18970 -15110
rect 19015 -15230 19135 -15110
rect 19180 -15230 19300 -15110
rect 19355 -15230 19475 -15110
rect 19520 -15230 19640 -15110
rect 19685 -15230 19805 -15110
rect 19850 -15230 19970 -15110
rect 20025 -15230 20145 -15110
rect 20190 -15230 20310 -15110
rect 20355 -15230 20475 -15110
rect 20520 -15230 20640 -15110
rect 20695 -15230 20815 -15110
rect 20860 -15230 20980 -15110
rect 21025 -15230 21145 -15110
rect 21190 -15230 21310 -15110
rect 21365 -15230 21485 -15110
rect 21530 -15230 21650 -15110
rect 21695 -15230 21815 -15110
rect 21860 -15230 21980 -15110
rect 22035 -15230 22155 -15110
rect 22200 -15230 22320 -15110
rect 22365 -15230 22485 -15110
rect 22530 -15230 22650 -15110
rect 22705 -15230 22825 -15110
rect 22870 -15230 22990 -15110
rect 23035 -15230 23155 -15110
rect 23200 -15230 23320 -15110
rect 23375 -15230 23495 -15110
rect 23540 -15230 23660 -15110
rect 23705 -15230 23825 -15110
rect 23870 -15230 23990 -15110
rect 18510 -15395 18630 -15275
rect 18685 -15395 18805 -15275
rect 18850 -15395 18970 -15275
rect 19015 -15395 19135 -15275
rect 19180 -15395 19300 -15275
rect 19355 -15395 19475 -15275
rect 19520 -15395 19640 -15275
rect 19685 -15395 19805 -15275
rect 19850 -15395 19970 -15275
rect 20025 -15395 20145 -15275
rect 20190 -15395 20310 -15275
rect 20355 -15395 20475 -15275
rect 20520 -15395 20640 -15275
rect 20695 -15395 20815 -15275
rect 20860 -15395 20980 -15275
rect 21025 -15395 21145 -15275
rect 21190 -15395 21310 -15275
rect 21365 -15395 21485 -15275
rect 21530 -15395 21650 -15275
rect 21695 -15395 21815 -15275
rect 21860 -15395 21980 -15275
rect 22035 -15395 22155 -15275
rect 22200 -15395 22320 -15275
rect 22365 -15395 22485 -15275
rect 22530 -15395 22650 -15275
rect 22705 -15395 22825 -15275
rect 22870 -15395 22990 -15275
rect 23035 -15395 23155 -15275
rect 23200 -15395 23320 -15275
rect 23375 -15395 23495 -15275
rect 23540 -15395 23660 -15275
rect 23705 -15395 23825 -15275
rect 23870 -15395 23990 -15275
rect 18510 -15570 18630 -15450
rect 18685 -15570 18805 -15450
rect 18850 -15570 18970 -15450
rect 19015 -15570 19135 -15450
rect 19180 -15570 19300 -15450
rect 19355 -15570 19475 -15450
rect 19520 -15570 19640 -15450
rect 19685 -15570 19805 -15450
rect 19850 -15570 19970 -15450
rect 20025 -15570 20145 -15450
rect 20190 -15570 20310 -15450
rect 20355 -15570 20475 -15450
rect 20520 -15570 20640 -15450
rect 20695 -15570 20815 -15450
rect 20860 -15570 20980 -15450
rect 21025 -15570 21145 -15450
rect 21190 -15570 21310 -15450
rect 21365 -15570 21485 -15450
rect 21530 -15570 21650 -15450
rect 21695 -15570 21815 -15450
rect 21860 -15570 21980 -15450
rect 22035 -15570 22155 -15450
rect 22200 -15570 22320 -15450
rect 22365 -15570 22485 -15450
rect 22530 -15570 22650 -15450
rect 22705 -15570 22825 -15450
rect 22870 -15570 22990 -15450
rect 23035 -15570 23155 -15450
rect 23200 -15570 23320 -15450
rect 23375 -15570 23495 -15450
rect 23540 -15570 23660 -15450
rect 23705 -15570 23825 -15450
rect 23870 -15570 23990 -15450
rect 24200 -10210 24320 -10090
rect 24375 -10210 24495 -10090
rect 24540 -10210 24660 -10090
rect 24705 -10210 24825 -10090
rect 24870 -10210 24990 -10090
rect 25045 -10210 25165 -10090
rect 25210 -10210 25330 -10090
rect 25375 -10210 25495 -10090
rect 25540 -10210 25660 -10090
rect 25715 -10210 25835 -10090
rect 25880 -10210 26000 -10090
rect 26045 -10210 26165 -10090
rect 26210 -10210 26330 -10090
rect 26385 -10210 26505 -10090
rect 26550 -10210 26670 -10090
rect 26715 -10210 26835 -10090
rect 26880 -10210 27000 -10090
rect 27055 -10210 27175 -10090
rect 27220 -10210 27340 -10090
rect 27385 -10210 27505 -10090
rect 27550 -10210 27670 -10090
rect 27725 -10210 27845 -10090
rect 27890 -10210 28010 -10090
rect 28055 -10210 28175 -10090
rect 28220 -10210 28340 -10090
rect 28395 -10210 28515 -10090
rect 28560 -10210 28680 -10090
rect 28725 -10210 28845 -10090
rect 28890 -10210 29010 -10090
rect 29065 -10210 29185 -10090
rect 29230 -10210 29350 -10090
rect 29395 -10210 29515 -10090
rect 29560 -10210 29680 -10090
rect 24200 -10375 24320 -10255
rect 24375 -10375 24495 -10255
rect 24540 -10375 24660 -10255
rect 24705 -10375 24825 -10255
rect 24870 -10375 24990 -10255
rect 25045 -10375 25165 -10255
rect 25210 -10375 25330 -10255
rect 25375 -10375 25495 -10255
rect 25540 -10375 25660 -10255
rect 25715 -10375 25835 -10255
rect 25880 -10375 26000 -10255
rect 26045 -10375 26165 -10255
rect 26210 -10375 26330 -10255
rect 26385 -10375 26505 -10255
rect 26550 -10375 26670 -10255
rect 26715 -10375 26835 -10255
rect 26880 -10375 27000 -10255
rect 27055 -10375 27175 -10255
rect 27220 -10375 27340 -10255
rect 27385 -10375 27505 -10255
rect 27550 -10375 27670 -10255
rect 27725 -10375 27845 -10255
rect 27890 -10375 28010 -10255
rect 28055 -10375 28175 -10255
rect 28220 -10375 28340 -10255
rect 28395 -10375 28515 -10255
rect 28560 -10375 28680 -10255
rect 28725 -10375 28845 -10255
rect 28890 -10375 29010 -10255
rect 29065 -10375 29185 -10255
rect 29230 -10375 29350 -10255
rect 29395 -10375 29515 -10255
rect 29560 -10375 29680 -10255
rect 24200 -10540 24320 -10420
rect 24375 -10540 24495 -10420
rect 24540 -10540 24660 -10420
rect 24705 -10540 24825 -10420
rect 24870 -10540 24990 -10420
rect 25045 -10540 25165 -10420
rect 25210 -10540 25330 -10420
rect 25375 -10540 25495 -10420
rect 25540 -10540 25660 -10420
rect 25715 -10540 25835 -10420
rect 25880 -10540 26000 -10420
rect 26045 -10540 26165 -10420
rect 26210 -10540 26330 -10420
rect 26385 -10540 26505 -10420
rect 26550 -10540 26670 -10420
rect 26715 -10540 26835 -10420
rect 26880 -10540 27000 -10420
rect 27055 -10540 27175 -10420
rect 27220 -10540 27340 -10420
rect 27385 -10540 27505 -10420
rect 27550 -10540 27670 -10420
rect 27725 -10540 27845 -10420
rect 27890 -10540 28010 -10420
rect 28055 -10540 28175 -10420
rect 28220 -10540 28340 -10420
rect 28395 -10540 28515 -10420
rect 28560 -10540 28680 -10420
rect 28725 -10540 28845 -10420
rect 28890 -10540 29010 -10420
rect 29065 -10540 29185 -10420
rect 29230 -10540 29350 -10420
rect 29395 -10540 29515 -10420
rect 29560 -10540 29680 -10420
rect 24200 -10705 24320 -10585
rect 24375 -10705 24495 -10585
rect 24540 -10705 24660 -10585
rect 24705 -10705 24825 -10585
rect 24870 -10705 24990 -10585
rect 25045 -10705 25165 -10585
rect 25210 -10705 25330 -10585
rect 25375 -10705 25495 -10585
rect 25540 -10705 25660 -10585
rect 25715 -10705 25835 -10585
rect 25880 -10705 26000 -10585
rect 26045 -10705 26165 -10585
rect 26210 -10705 26330 -10585
rect 26385 -10705 26505 -10585
rect 26550 -10705 26670 -10585
rect 26715 -10705 26835 -10585
rect 26880 -10705 27000 -10585
rect 27055 -10705 27175 -10585
rect 27220 -10705 27340 -10585
rect 27385 -10705 27505 -10585
rect 27550 -10705 27670 -10585
rect 27725 -10705 27845 -10585
rect 27890 -10705 28010 -10585
rect 28055 -10705 28175 -10585
rect 28220 -10705 28340 -10585
rect 28395 -10705 28515 -10585
rect 28560 -10705 28680 -10585
rect 28725 -10705 28845 -10585
rect 28890 -10705 29010 -10585
rect 29065 -10705 29185 -10585
rect 29230 -10705 29350 -10585
rect 29395 -10705 29515 -10585
rect 29560 -10705 29680 -10585
rect 24200 -10880 24320 -10760
rect 24375 -10880 24495 -10760
rect 24540 -10880 24660 -10760
rect 24705 -10880 24825 -10760
rect 24870 -10880 24990 -10760
rect 25045 -10880 25165 -10760
rect 25210 -10880 25330 -10760
rect 25375 -10880 25495 -10760
rect 25540 -10880 25660 -10760
rect 25715 -10880 25835 -10760
rect 25880 -10880 26000 -10760
rect 26045 -10880 26165 -10760
rect 26210 -10880 26330 -10760
rect 26385 -10880 26505 -10760
rect 26550 -10880 26670 -10760
rect 26715 -10880 26835 -10760
rect 26880 -10880 27000 -10760
rect 27055 -10880 27175 -10760
rect 27220 -10880 27340 -10760
rect 27385 -10880 27505 -10760
rect 27550 -10880 27670 -10760
rect 27725 -10880 27845 -10760
rect 27890 -10880 28010 -10760
rect 28055 -10880 28175 -10760
rect 28220 -10880 28340 -10760
rect 28395 -10880 28515 -10760
rect 28560 -10880 28680 -10760
rect 28725 -10880 28845 -10760
rect 28890 -10880 29010 -10760
rect 29065 -10880 29185 -10760
rect 29230 -10880 29350 -10760
rect 29395 -10880 29515 -10760
rect 29560 -10880 29680 -10760
rect 24200 -11045 24320 -10925
rect 24375 -11045 24495 -10925
rect 24540 -11045 24660 -10925
rect 24705 -11045 24825 -10925
rect 24870 -11045 24990 -10925
rect 25045 -11045 25165 -10925
rect 25210 -11045 25330 -10925
rect 25375 -11045 25495 -10925
rect 25540 -11045 25660 -10925
rect 25715 -11045 25835 -10925
rect 25880 -11045 26000 -10925
rect 26045 -11045 26165 -10925
rect 26210 -11045 26330 -10925
rect 26385 -11045 26505 -10925
rect 26550 -11045 26670 -10925
rect 26715 -11045 26835 -10925
rect 26880 -11045 27000 -10925
rect 27055 -11045 27175 -10925
rect 27220 -11045 27340 -10925
rect 27385 -11045 27505 -10925
rect 27550 -11045 27670 -10925
rect 27725 -11045 27845 -10925
rect 27890 -11045 28010 -10925
rect 28055 -11045 28175 -10925
rect 28220 -11045 28340 -10925
rect 28395 -11045 28515 -10925
rect 28560 -11045 28680 -10925
rect 28725 -11045 28845 -10925
rect 28890 -11045 29010 -10925
rect 29065 -11045 29185 -10925
rect 29230 -11045 29350 -10925
rect 29395 -11045 29515 -10925
rect 29560 -11045 29680 -10925
rect 24200 -11210 24320 -11090
rect 24375 -11210 24495 -11090
rect 24540 -11210 24660 -11090
rect 24705 -11210 24825 -11090
rect 24870 -11210 24990 -11090
rect 25045 -11210 25165 -11090
rect 25210 -11210 25330 -11090
rect 25375 -11210 25495 -11090
rect 25540 -11210 25660 -11090
rect 25715 -11210 25835 -11090
rect 25880 -11210 26000 -11090
rect 26045 -11210 26165 -11090
rect 26210 -11210 26330 -11090
rect 26385 -11210 26505 -11090
rect 26550 -11210 26670 -11090
rect 26715 -11210 26835 -11090
rect 26880 -11210 27000 -11090
rect 27055 -11210 27175 -11090
rect 27220 -11210 27340 -11090
rect 27385 -11210 27505 -11090
rect 27550 -11210 27670 -11090
rect 27725 -11210 27845 -11090
rect 27890 -11210 28010 -11090
rect 28055 -11210 28175 -11090
rect 28220 -11210 28340 -11090
rect 28395 -11210 28515 -11090
rect 28560 -11210 28680 -11090
rect 28725 -11210 28845 -11090
rect 28890 -11210 29010 -11090
rect 29065 -11210 29185 -11090
rect 29230 -11210 29350 -11090
rect 29395 -11210 29515 -11090
rect 29560 -11210 29680 -11090
rect 24200 -11375 24320 -11255
rect 24375 -11375 24495 -11255
rect 24540 -11375 24660 -11255
rect 24705 -11375 24825 -11255
rect 24870 -11375 24990 -11255
rect 25045 -11375 25165 -11255
rect 25210 -11375 25330 -11255
rect 25375 -11375 25495 -11255
rect 25540 -11375 25660 -11255
rect 25715 -11375 25835 -11255
rect 25880 -11375 26000 -11255
rect 26045 -11375 26165 -11255
rect 26210 -11375 26330 -11255
rect 26385 -11375 26505 -11255
rect 26550 -11375 26670 -11255
rect 26715 -11375 26835 -11255
rect 26880 -11375 27000 -11255
rect 27055 -11375 27175 -11255
rect 27220 -11375 27340 -11255
rect 27385 -11375 27505 -11255
rect 27550 -11375 27670 -11255
rect 27725 -11375 27845 -11255
rect 27890 -11375 28010 -11255
rect 28055 -11375 28175 -11255
rect 28220 -11375 28340 -11255
rect 28395 -11375 28515 -11255
rect 28560 -11375 28680 -11255
rect 28725 -11375 28845 -11255
rect 28890 -11375 29010 -11255
rect 29065 -11375 29185 -11255
rect 29230 -11375 29350 -11255
rect 29395 -11375 29515 -11255
rect 29560 -11375 29680 -11255
rect 24200 -11550 24320 -11430
rect 24375 -11550 24495 -11430
rect 24540 -11550 24660 -11430
rect 24705 -11550 24825 -11430
rect 24870 -11550 24990 -11430
rect 25045 -11550 25165 -11430
rect 25210 -11550 25330 -11430
rect 25375 -11550 25495 -11430
rect 25540 -11550 25660 -11430
rect 25715 -11550 25835 -11430
rect 25880 -11550 26000 -11430
rect 26045 -11550 26165 -11430
rect 26210 -11550 26330 -11430
rect 26385 -11550 26505 -11430
rect 26550 -11550 26670 -11430
rect 26715 -11550 26835 -11430
rect 26880 -11550 27000 -11430
rect 27055 -11550 27175 -11430
rect 27220 -11550 27340 -11430
rect 27385 -11550 27505 -11430
rect 27550 -11550 27670 -11430
rect 27725 -11550 27845 -11430
rect 27890 -11550 28010 -11430
rect 28055 -11550 28175 -11430
rect 28220 -11550 28340 -11430
rect 28395 -11550 28515 -11430
rect 28560 -11550 28680 -11430
rect 28725 -11550 28845 -11430
rect 28890 -11550 29010 -11430
rect 29065 -11550 29185 -11430
rect 29230 -11550 29350 -11430
rect 29395 -11550 29515 -11430
rect 29560 -11550 29680 -11430
rect 24200 -11715 24320 -11595
rect 24375 -11715 24495 -11595
rect 24540 -11715 24660 -11595
rect 24705 -11715 24825 -11595
rect 24870 -11715 24990 -11595
rect 25045 -11715 25165 -11595
rect 25210 -11715 25330 -11595
rect 25375 -11715 25495 -11595
rect 25540 -11715 25660 -11595
rect 25715 -11715 25835 -11595
rect 25880 -11715 26000 -11595
rect 26045 -11715 26165 -11595
rect 26210 -11715 26330 -11595
rect 26385 -11715 26505 -11595
rect 26550 -11715 26670 -11595
rect 26715 -11715 26835 -11595
rect 26880 -11715 27000 -11595
rect 27055 -11715 27175 -11595
rect 27220 -11715 27340 -11595
rect 27385 -11715 27505 -11595
rect 27550 -11715 27670 -11595
rect 27725 -11715 27845 -11595
rect 27890 -11715 28010 -11595
rect 28055 -11715 28175 -11595
rect 28220 -11715 28340 -11595
rect 28395 -11715 28515 -11595
rect 28560 -11715 28680 -11595
rect 28725 -11715 28845 -11595
rect 28890 -11715 29010 -11595
rect 29065 -11715 29185 -11595
rect 29230 -11715 29350 -11595
rect 29395 -11715 29515 -11595
rect 29560 -11715 29680 -11595
rect 24200 -11880 24320 -11760
rect 24375 -11880 24495 -11760
rect 24540 -11880 24660 -11760
rect 24705 -11880 24825 -11760
rect 24870 -11880 24990 -11760
rect 25045 -11880 25165 -11760
rect 25210 -11880 25330 -11760
rect 25375 -11880 25495 -11760
rect 25540 -11880 25660 -11760
rect 25715 -11880 25835 -11760
rect 25880 -11880 26000 -11760
rect 26045 -11880 26165 -11760
rect 26210 -11880 26330 -11760
rect 26385 -11880 26505 -11760
rect 26550 -11880 26670 -11760
rect 26715 -11880 26835 -11760
rect 26880 -11880 27000 -11760
rect 27055 -11880 27175 -11760
rect 27220 -11880 27340 -11760
rect 27385 -11880 27505 -11760
rect 27550 -11880 27670 -11760
rect 27725 -11880 27845 -11760
rect 27890 -11880 28010 -11760
rect 28055 -11880 28175 -11760
rect 28220 -11880 28340 -11760
rect 28395 -11880 28515 -11760
rect 28560 -11880 28680 -11760
rect 28725 -11880 28845 -11760
rect 28890 -11880 29010 -11760
rect 29065 -11880 29185 -11760
rect 29230 -11880 29350 -11760
rect 29395 -11880 29515 -11760
rect 29560 -11880 29680 -11760
rect 24200 -12045 24320 -11925
rect 24375 -12045 24495 -11925
rect 24540 -12045 24660 -11925
rect 24705 -12045 24825 -11925
rect 24870 -12045 24990 -11925
rect 25045 -12045 25165 -11925
rect 25210 -12045 25330 -11925
rect 25375 -12045 25495 -11925
rect 25540 -12045 25660 -11925
rect 25715 -12045 25835 -11925
rect 25880 -12045 26000 -11925
rect 26045 -12045 26165 -11925
rect 26210 -12045 26330 -11925
rect 26385 -12045 26505 -11925
rect 26550 -12045 26670 -11925
rect 26715 -12045 26835 -11925
rect 26880 -12045 27000 -11925
rect 27055 -12045 27175 -11925
rect 27220 -12045 27340 -11925
rect 27385 -12045 27505 -11925
rect 27550 -12045 27670 -11925
rect 27725 -12045 27845 -11925
rect 27890 -12045 28010 -11925
rect 28055 -12045 28175 -11925
rect 28220 -12045 28340 -11925
rect 28395 -12045 28515 -11925
rect 28560 -12045 28680 -11925
rect 28725 -12045 28845 -11925
rect 28890 -12045 29010 -11925
rect 29065 -12045 29185 -11925
rect 29230 -12045 29350 -11925
rect 29395 -12045 29515 -11925
rect 29560 -12045 29680 -11925
rect 24200 -12220 24320 -12100
rect 24375 -12220 24495 -12100
rect 24540 -12220 24660 -12100
rect 24705 -12220 24825 -12100
rect 24870 -12220 24990 -12100
rect 25045 -12220 25165 -12100
rect 25210 -12220 25330 -12100
rect 25375 -12220 25495 -12100
rect 25540 -12220 25660 -12100
rect 25715 -12220 25835 -12100
rect 25880 -12220 26000 -12100
rect 26045 -12220 26165 -12100
rect 26210 -12220 26330 -12100
rect 26385 -12220 26505 -12100
rect 26550 -12220 26670 -12100
rect 26715 -12220 26835 -12100
rect 26880 -12220 27000 -12100
rect 27055 -12220 27175 -12100
rect 27220 -12220 27340 -12100
rect 27385 -12220 27505 -12100
rect 27550 -12220 27670 -12100
rect 27725 -12220 27845 -12100
rect 27890 -12220 28010 -12100
rect 28055 -12220 28175 -12100
rect 28220 -12220 28340 -12100
rect 28395 -12220 28515 -12100
rect 28560 -12220 28680 -12100
rect 28725 -12220 28845 -12100
rect 28890 -12220 29010 -12100
rect 29065 -12220 29185 -12100
rect 29230 -12220 29350 -12100
rect 29395 -12220 29515 -12100
rect 29560 -12220 29680 -12100
rect 24200 -12385 24320 -12265
rect 24375 -12385 24495 -12265
rect 24540 -12385 24660 -12265
rect 24705 -12385 24825 -12265
rect 24870 -12385 24990 -12265
rect 25045 -12385 25165 -12265
rect 25210 -12385 25330 -12265
rect 25375 -12385 25495 -12265
rect 25540 -12385 25660 -12265
rect 25715 -12385 25835 -12265
rect 25880 -12385 26000 -12265
rect 26045 -12385 26165 -12265
rect 26210 -12385 26330 -12265
rect 26385 -12385 26505 -12265
rect 26550 -12385 26670 -12265
rect 26715 -12385 26835 -12265
rect 26880 -12385 27000 -12265
rect 27055 -12385 27175 -12265
rect 27220 -12385 27340 -12265
rect 27385 -12385 27505 -12265
rect 27550 -12385 27670 -12265
rect 27725 -12385 27845 -12265
rect 27890 -12385 28010 -12265
rect 28055 -12385 28175 -12265
rect 28220 -12385 28340 -12265
rect 28395 -12385 28515 -12265
rect 28560 -12385 28680 -12265
rect 28725 -12385 28845 -12265
rect 28890 -12385 29010 -12265
rect 29065 -12385 29185 -12265
rect 29230 -12385 29350 -12265
rect 29395 -12385 29515 -12265
rect 29560 -12385 29680 -12265
rect 24200 -12550 24320 -12430
rect 24375 -12550 24495 -12430
rect 24540 -12550 24660 -12430
rect 24705 -12550 24825 -12430
rect 24870 -12550 24990 -12430
rect 25045 -12550 25165 -12430
rect 25210 -12550 25330 -12430
rect 25375 -12550 25495 -12430
rect 25540 -12550 25660 -12430
rect 25715 -12550 25835 -12430
rect 25880 -12550 26000 -12430
rect 26045 -12550 26165 -12430
rect 26210 -12550 26330 -12430
rect 26385 -12550 26505 -12430
rect 26550 -12550 26670 -12430
rect 26715 -12550 26835 -12430
rect 26880 -12550 27000 -12430
rect 27055 -12550 27175 -12430
rect 27220 -12550 27340 -12430
rect 27385 -12550 27505 -12430
rect 27550 -12550 27670 -12430
rect 27725 -12550 27845 -12430
rect 27890 -12550 28010 -12430
rect 28055 -12550 28175 -12430
rect 28220 -12550 28340 -12430
rect 28395 -12550 28515 -12430
rect 28560 -12550 28680 -12430
rect 28725 -12550 28845 -12430
rect 28890 -12550 29010 -12430
rect 29065 -12550 29185 -12430
rect 29230 -12550 29350 -12430
rect 29395 -12550 29515 -12430
rect 29560 -12550 29680 -12430
rect 24200 -12715 24320 -12595
rect 24375 -12715 24495 -12595
rect 24540 -12715 24660 -12595
rect 24705 -12715 24825 -12595
rect 24870 -12715 24990 -12595
rect 25045 -12715 25165 -12595
rect 25210 -12715 25330 -12595
rect 25375 -12715 25495 -12595
rect 25540 -12715 25660 -12595
rect 25715 -12715 25835 -12595
rect 25880 -12715 26000 -12595
rect 26045 -12715 26165 -12595
rect 26210 -12715 26330 -12595
rect 26385 -12715 26505 -12595
rect 26550 -12715 26670 -12595
rect 26715 -12715 26835 -12595
rect 26880 -12715 27000 -12595
rect 27055 -12715 27175 -12595
rect 27220 -12715 27340 -12595
rect 27385 -12715 27505 -12595
rect 27550 -12715 27670 -12595
rect 27725 -12715 27845 -12595
rect 27890 -12715 28010 -12595
rect 28055 -12715 28175 -12595
rect 28220 -12715 28340 -12595
rect 28395 -12715 28515 -12595
rect 28560 -12715 28680 -12595
rect 28725 -12715 28845 -12595
rect 28890 -12715 29010 -12595
rect 29065 -12715 29185 -12595
rect 29230 -12715 29350 -12595
rect 29395 -12715 29515 -12595
rect 29560 -12715 29680 -12595
rect 24200 -12890 24320 -12770
rect 24375 -12890 24495 -12770
rect 24540 -12890 24660 -12770
rect 24705 -12890 24825 -12770
rect 24870 -12890 24990 -12770
rect 25045 -12890 25165 -12770
rect 25210 -12890 25330 -12770
rect 25375 -12890 25495 -12770
rect 25540 -12890 25660 -12770
rect 25715 -12890 25835 -12770
rect 25880 -12890 26000 -12770
rect 26045 -12890 26165 -12770
rect 26210 -12890 26330 -12770
rect 26385 -12890 26505 -12770
rect 26550 -12890 26670 -12770
rect 26715 -12890 26835 -12770
rect 26880 -12890 27000 -12770
rect 27055 -12890 27175 -12770
rect 27220 -12890 27340 -12770
rect 27385 -12890 27505 -12770
rect 27550 -12890 27670 -12770
rect 27725 -12890 27845 -12770
rect 27890 -12890 28010 -12770
rect 28055 -12890 28175 -12770
rect 28220 -12890 28340 -12770
rect 28395 -12890 28515 -12770
rect 28560 -12890 28680 -12770
rect 28725 -12890 28845 -12770
rect 28890 -12890 29010 -12770
rect 29065 -12890 29185 -12770
rect 29230 -12890 29350 -12770
rect 29395 -12890 29515 -12770
rect 29560 -12890 29680 -12770
rect 24200 -13055 24320 -12935
rect 24375 -13055 24495 -12935
rect 24540 -13055 24660 -12935
rect 24705 -13055 24825 -12935
rect 24870 -13055 24990 -12935
rect 25045 -13055 25165 -12935
rect 25210 -13055 25330 -12935
rect 25375 -13055 25495 -12935
rect 25540 -13055 25660 -12935
rect 25715 -13055 25835 -12935
rect 25880 -13055 26000 -12935
rect 26045 -13055 26165 -12935
rect 26210 -13055 26330 -12935
rect 26385 -13055 26505 -12935
rect 26550 -13055 26670 -12935
rect 26715 -13055 26835 -12935
rect 26880 -13055 27000 -12935
rect 27055 -13055 27175 -12935
rect 27220 -13055 27340 -12935
rect 27385 -13055 27505 -12935
rect 27550 -13055 27670 -12935
rect 27725 -13055 27845 -12935
rect 27890 -13055 28010 -12935
rect 28055 -13055 28175 -12935
rect 28220 -13055 28340 -12935
rect 28395 -13055 28515 -12935
rect 28560 -13055 28680 -12935
rect 28725 -13055 28845 -12935
rect 28890 -13055 29010 -12935
rect 29065 -13055 29185 -12935
rect 29230 -13055 29350 -12935
rect 29395 -13055 29515 -12935
rect 29560 -13055 29680 -12935
rect 24200 -13220 24320 -13100
rect 24375 -13220 24495 -13100
rect 24540 -13220 24660 -13100
rect 24705 -13220 24825 -13100
rect 24870 -13220 24990 -13100
rect 25045 -13220 25165 -13100
rect 25210 -13220 25330 -13100
rect 25375 -13220 25495 -13100
rect 25540 -13220 25660 -13100
rect 25715 -13220 25835 -13100
rect 25880 -13220 26000 -13100
rect 26045 -13220 26165 -13100
rect 26210 -13220 26330 -13100
rect 26385 -13220 26505 -13100
rect 26550 -13220 26670 -13100
rect 26715 -13220 26835 -13100
rect 26880 -13220 27000 -13100
rect 27055 -13220 27175 -13100
rect 27220 -13220 27340 -13100
rect 27385 -13220 27505 -13100
rect 27550 -13220 27670 -13100
rect 27725 -13220 27845 -13100
rect 27890 -13220 28010 -13100
rect 28055 -13220 28175 -13100
rect 28220 -13220 28340 -13100
rect 28395 -13220 28515 -13100
rect 28560 -13220 28680 -13100
rect 28725 -13220 28845 -13100
rect 28890 -13220 29010 -13100
rect 29065 -13220 29185 -13100
rect 29230 -13220 29350 -13100
rect 29395 -13220 29515 -13100
rect 29560 -13220 29680 -13100
rect 24200 -13385 24320 -13265
rect 24375 -13385 24495 -13265
rect 24540 -13385 24660 -13265
rect 24705 -13385 24825 -13265
rect 24870 -13385 24990 -13265
rect 25045 -13385 25165 -13265
rect 25210 -13385 25330 -13265
rect 25375 -13385 25495 -13265
rect 25540 -13385 25660 -13265
rect 25715 -13385 25835 -13265
rect 25880 -13385 26000 -13265
rect 26045 -13385 26165 -13265
rect 26210 -13385 26330 -13265
rect 26385 -13385 26505 -13265
rect 26550 -13385 26670 -13265
rect 26715 -13385 26835 -13265
rect 26880 -13385 27000 -13265
rect 27055 -13385 27175 -13265
rect 27220 -13385 27340 -13265
rect 27385 -13385 27505 -13265
rect 27550 -13385 27670 -13265
rect 27725 -13385 27845 -13265
rect 27890 -13385 28010 -13265
rect 28055 -13385 28175 -13265
rect 28220 -13385 28340 -13265
rect 28395 -13385 28515 -13265
rect 28560 -13385 28680 -13265
rect 28725 -13385 28845 -13265
rect 28890 -13385 29010 -13265
rect 29065 -13385 29185 -13265
rect 29230 -13385 29350 -13265
rect 29395 -13385 29515 -13265
rect 29560 -13385 29680 -13265
rect 24200 -13560 24320 -13440
rect 24375 -13560 24495 -13440
rect 24540 -13560 24660 -13440
rect 24705 -13560 24825 -13440
rect 24870 -13560 24990 -13440
rect 25045 -13560 25165 -13440
rect 25210 -13560 25330 -13440
rect 25375 -13560 25495 -13440
rect 25540 -13560 25660 -13440
rect 25715 -13560 25835 -13440
rect 25880 -13560 26000 -13440
rect 26045 -13560 26165 -13440
rect 26210 -13560 26330 -13440
rect 26385 -13560 26505 -13440
rect 26550 -13560 26670 -13440
rect 26715 -13560 26835 -13440
rect 26880 -13560 27000 -13440
rect 27055 -13560 27175 -13440
rect 27220 -13560 27340 -13440
rect 27385 -13560 27505 -13440
rect 27550 -13560 27670 -13440
rect 27725 -13560 27845 -13440
rect 27890 -13560 28010 -13440
rect 28055 -13560 28175 -13440
rect 28220 -13560 28340 -13440
rect 28395 -13560 28515 -13440
rect 28560 -13560 28680 -13440
rect 28725 -13560 28845 -13440
rect 28890 -13560 29010 -13440
rect 29065 -13560 29185 -13440
rect 29230 -13560 29350 -13440
rect 29395 -13560 29515 -13440
rect 29560 -13560 29680 -13440
rect 24200 -13725 24320 -13605
rect 24375 -13725 24495 -13605
rect 24540 -13725 24660 -13605
rect 24705 -13725 24825 -13605
rect 24870 -13725 24990 -13605
rect 25045 -13725 25165 -13605
rect 25210 -13725 25330 -13605
rect 25375 -13725 25495 -13605
rect 25540 -13725 25660 -13605
rect 25715 -13725 25835 -13605
rect 25880 -13725 26000 -13605
rect 26045 -13725 26165 -13605
rect 26210 -13725 26330 -13605
rect 26385 -13725 26505 -13605
rect 26550 -13725 26670 -13605
rect 26715 -13725 26835 -13605
rect 26880 -13725 27000 -13605
rect 27055 -13725 27175 -13605
rect 27220 -13725 27340 -13605
rect 27385 -13725 27505 -13605
rect 27550 -13725 27670 -13605
rect 27725 -13725 27845 -13605
rect 27890 -13725 28010 -13605
rect 28055 -13725 28175 -13605
rect 28220 -13725 28340 -13605
rect 28395 -13725 28515 -13605
rect 28560 -13725 28680 -13605
rect 28725 -13725 28845 -13605
rect 28890 -13725 29010 -13605
rect 29065 -13725 29185 -13605
rect 29230 -13725 29350 -13605
rect 29395 -13725 29515 -13605
rect 29560 -13725 29680 -13605
rect 24200 -13890 24320 -13770
rect 24375 -13890 24495 -13770
rect 24540 -13890 24660 -13770
rect 24705 -13890 24825 -13770
rect 24870 -13890 24990 -13770
rect 25045 -13890 25165 -13770
rect 25210 -13890 25330 -13770
rect 25375 -13890 25495 -13770
rect 25540 -13890 25660 -13770
rect 25715 -13890 25835 -13770
rect 25880 -13890 26000 -13770
rect 26045 -13890 26165 -13770
rect 26210 -13890 26330 -13770
rect 26385 -13890 26505 -13770
rect 26550 -13890 26670 -13770
rect 26715 -13890 26835 -13770
rect 26880 -13890 27000 -13770
rect 27055 -13890 27175 -13770
rect 27220 -13890 27340 -13770
rect 27385 -13890 27505 -13770
rect 27550 -13890 27670 -13770
rect 27725 -13890 27845 -13770
rect 27890 -13890 28010 -13770
rect 28055 -13890 28175 -13770
rect 28220 -13890 28340 -13770
rect 28395 -13890 28515 -13770
rect 28560 -13890 28680 -13770
rect 28725 -13890 28845 -13770
rect 28890 -13890 29010 -13770
rect 29065 -13890 29185 -13770
rect 29230 -13890 29350 -13770
rect 29395 -13890 29515 -13770
rect 29560 -13890 29680 -13770
rect 24200 -14055 24320 -13935
rect 24375 -14055 24495 -13935
rect 24540 -14055 24660 -13935
rect 24705 -14055 24825 -13935
rect 24870 -14055 24990 -13935
rect 25045 -14055 25165 -13935
rect 25210 -14055 25330 -13935
rect 25375 -14055 25495 -13935
rect 25540 -14055 25660 -13935
rect 25715 -14055 25835 -13935
rect 25880 -14055 26000 -13935
rect 26045 -14055 26165 -13935
rect 26210 -14055 26330 -13935
rect 26385 -14055 26505 -13935
rect 26550 -14055 26670 -13935
rect 26715 -14055 26835 -13935
rect 26880 -14055 27000 -13935
rect 27055 -14055 27175 -13935
rect 27220 -14055 27340 -13935
rect 27385 -14055 27505 -13935
rect 27550 -14055 27670 -13935
rect 27725 -14055 27845 -13935
rect 27890 -14055 28010 -13935
rect 28055 -14055 28175 -13935
rect 28220 -14055 28340 -13935
rect 28395 -14055 28515 -13935
rect 28560 -14055 28680 -13935
rect 28725 -14055 28845 -13935
rect 28890 -14055 29010 -13935
rect 29065 -14055 29185 -13935
rect 29230 -14055 29350 -13935
rect 29395 -14055 29515 -13935
rect 29560 -14055 29680 -13935
rect 24200 -14230 24320 -14110
rect 24375 -14230 24495 -14110
rect 24540 -14230 24660 -14110
rect 24705 -14230 24825 -14110
rect 24870 -14230 24990 -14110
rect 25045 -14230 25165 -14110
rect 25210 -14230 25330 -14110
rect 25375 -14230 25495 -14110
rect 25540 -14230 25660 -14110
rect 25715 -14230 25835 -14110
rect 25880 -14230 26000 -14110
rect 26045 -14230 26165 -14110
rect 26210 -14230 26330 -14110
rect 26385 -14230 26505 -14110
rect 26550 -14230 26670 -14110
rect 26715 -14230 26835 -14110
rect 26880 -14230 27000 -14110
rect 27055 -14230 27175 -14110
rect 27220 -14230 27340 -14110
rect 27385 -14230 27505 -14110
rect 27550 -14230 27670 -14110
rect 27725 -14230 27845 -14110
rect 27890 -14230 28010 -14110
rect 28055 -14230 28175 -14110
rect 28220 -14230 28340 -14110
rect 28395 -14230 28515 -14110
rect 28560 -14230 28680 -14110
rect 28725 -14230 28845 -14110
rect 28890 -14230 29010 -14110
rect 29065 -14230 29185 -14110
rect 29230 -14230 29350 -14110
rect 29395 -14230 29515 -14110
rect 29560 -14230 29680 -14110
rect 24200 -14395 24320 -14275
rect 24375 -14395 24495 -14275
rect 24540 -14395 24660 -14275
rect 24705 -14395 24825 -14275
rect 24870 -14395 24990 -14275
rect 25045 -14395 25165 -14275
rect 25210 -14395 25330 -14275
rect 25375 -14395 25495 -14275
rect 25540 -14395 25660 -14275
rect 25715 -14395 25835 -14275
rect 25880 -14395 26000 -14275
rect 26045 -14395 26165 -14275
rect 26210 -14395 26330 -14275
rect 26385 -14395 26505 -14275
rect 26550 -14395 26670 -14275
rect 26715 -14395 26835 -14275
rect 26880 -14395 27000 -14275
rect 27055 -14395 27175 -14275
rect 27220 -14395 27340 -14275
rect 27385 -14395 27505 -14275
rect 27550 -14395 27670 -14275
rect 27725 -14395 27845 -14275
rect 27890 -14395 28010 -14275
rect 28055 -14395 28175 -14275
rect 28220 -14395 28340 -14275
rect 28395 -14395 28515 -14275
rect 28560 -14395 28680 -14275
rect 28725 -14395 28845 -14275
rect 28890 -14395 29010 -14275
rect 29065 -14395 29185 -14275
rect 29230 -14395 29350 -14275
rect 29395 -14395 29515 -14275
rect 29560 -14395 29680 -14275
rect 24200 -14560 24320 -14440
rect 24375 -14560 24495 -14440
rect 24540 -14560 24660 -14440
rect 24705 -14560 24825 -14440
rect 24870 -14560 24990 -14440
rect 25045 -14560 25165 -14440
rect 25210 -14560 25330 -14440
rect 25375 -14560 25495 -14440
rect 25540 -14560 25660 -14440
rect 25715 -14560 25835 -14440
rect 25880 -14560 26000 -14440
rect 26045 -14560 26165 -14440
rect 26210 -14560 26330 -14440
rect 26385 -14560 26505 -14440
rect 26550 -14560 26670 -14440
rect 26715 -14560 26835 -14440
rect 26880 -14560 27000 -14440
rect 27055 -14560 27175 -14440
rect 27220 -14560 27340 -14440
rect 27385 -14560 27505 -14440
rect 27550 -14560 27670 -14440
rect 27725 -14560 27845 -14440
rect 27890 -14560 28010 -14440
rect 28055 -14560 28175 -14440
rect 28220 -14560 28340 -14440
rect 28395 -14560 28515 -14440
rect 28560 -14560 28680 -14440
rect 28725 -14560 28845 -14440
rect 28890 -14560 29010 -14440
rect 29065 -14560 29185 -14440
rect 29230 -14560 29350 -14440
rect 29395 -14560 29515 -14440
rect 29560 -14560 29680 -14440
rect 24200 -14725 24320 -14605
rect 24375 -14725 24495 -14605
rect 24540 -14725 24660 -14605
rect 24705 -14725 24825 -14605
rect 24870 -14725 24990 -14605
rect 25045 -14725 25165 -14605
rect 25210 -14725 25330 -14605
rect 25375 -14725 25495 -14605
rect 25540 -14725 25660 -14605
rect 25715 -14725 25835 -14605
rect 25880 -14725 26000 -14605
rect 26045 -14725 26165 -14605
rect 26210 -14725 26330 -14605
rect 26385 -14725 26505 -14605
rect 26550 -14725 26670 -14605
rect 26715 -14725 26835 -14605
rect 26880 -14725 27000 -14605
rect 27055 -14725 27175 -14605
rect 27220 -14725 27340 -14605
rect 27385 -14725 27505 -14605
rect 27550 -14725 27670 -14605
rect 27725 -14725 27845 -14605
rect 27890 -14725 28010 -14605
rect 28055 -14725 28175 -14605
rect 28220 -14725 28340 -14605
rect 28395 -14725 28515 -14605
rect 28560 -14725 28680 -14605
rect 28725 -14725 28845 -14605
rect 28890 -14725 29010 -14605
rect 29065 -14725 29185 -14605
rect 29230 -14725 29350 -14605
rect 29395 -14725 29515 -14605
rect 29560 -14725 29680 -14605
rect 24200 -14900 24320 -14780
rect 24375 -14900 24495 -14780
rect 24540 -14900 24660 -14780
rect 24705 -14900 24825 -14780
rect 24870 -14900 24990 -14780
rect 25045 -14900 25165 -14780
rect 25210 -14900 25330 -14780
rect 25375 -14900 25495 -14780
rect 25540 -14900 25660 -14780
rect 25715 -14900 25835 -14780
rect 25880 -14900 26000 -14780
rect 26045 -14900 26165 -14780
rect 26210 -14900 26330 -14780
rect 26385 -14900 26505 -14780
rect 26550 -14900 26670 -14780
rect 26715 -14900 26835 -14780
rect 26880 -14900 27000 -14780
rect 27055 -14900 27175 -14780
rect 27220 -14900 27340 -14780
rect 27385 -14900 27505 -14780
rect 27550 -14900 27670 -14780
rect 27725 -14900 27845 -14780
rect 27890 -14900 28010 -14780
rect 28055 -14900 28175 -14780
rect 28220 -14900 28340 -14780
rect 28395 -14900 28515 -14780
rect 28560 -14900 28680 -14780
rect 28725 -14900 28845 -14780
rect 28890 -14900 29010 -14780
rect 29065 -14900 29185 -14780
rect 29230 -14900 29350 -14780
rect 29395 -14900 29515 -14780
rect 29560 -14900 29680 -14780
rect 24200 -15065 24320 -14945
rect 24375 -15065 24495 -14945
rect 24540 -15065 24660 -14945
rect 24705 -15065 24825 -14945
rect 24870 -15065 24990 -14945
rect 25045 -15065 25165 -14945
rect 25210 -15065 25330 -14945
rect 25375 -15065 25495 -14945
rect 25540 -15065 25660 -14945
rect 25715 -15065 25835 -14945
rect 25880 -15065 26000 -14945
rect 26045 -15065 26165 -14945
rect 26210 -15065 26330 -14945
rect 26385 -15065 26505 -14945
rect 26550 -15065 26670 -14945
rect 26715 -15065 26835 -14945
rect 26880 -15065 27000 -14945
rect 27055 -15065 27175 -14945
rect 27220 -15065 27340 -14945
rect 27385 -15065 27505 -14945
rect 27550 -15065 27670 -14945
rect 27725 -15065 27845 -14945
rect 27890 -15065 28010 -14945
rect 28055 -15065 28175 -14945
rect 28220 -15065 28340 -14945
rect 28395 -15065 28515 -14945
rect 28560 -15065 28680 -14945
rect 28725 -15065 28845 -14945
rect 28890 -15065 29010 -14945
rect 29065 -15065 29185 -14945
rect 29230 -15065 29350 -14945
rect 29395 -15065 29515 -14945
rect 29560 -15065 29680 -14945
rect 24200 -15230 24320 -15110
rect 24375 -15230 24495 -15110
rect 24540 -15230 24660 -15110
rect 24705 -15230 24825 -15110
rect 24870 -15230 24990 -15110
rect 25045 -15230 25165 -15110
rect 25210 -15230 25330 -15110
rect 25375 -15230 25495 -15110
rect 25540 -15230 25660 -15110
rect 25715 -15230 25835 -15110
rect 25880 -15230 26000 -15110
rect 26045 -15230 26165 -15110
rect 26210 -15230 26330 -15110
rect 26385 -15230 26505 -15110
rect 26550 -15230 26670 -15110
rect 26715 -15230 26835 -15110
rect 26880 -15230 27000 -15110
rect 27055 -15230 27175 -15110
rect 27220 -15230 27340 -15110
rect 27385 -15230 27505 -15110
rect 27550 -15230 27670 -15110
rect 27725 -15230 27845 -15110
rect 27890 -15230 28010 -15110
rect 28055 -15230 28175 -15110
rect 28220 -15230 28340 -15110
rect 28395 -15230 28515 -15110
rect 28560 -15230 28680 -15110
rect 28725 -15230 28845 -15110
rect 28890 -15230 29010 -15110
rect 29065 -15230 29185 -15110
rect 29230 -15230 29350 -15110
rect 29395 -15230 29515 -15110
rect 29560 -15230 29680 -15110
rect 24200 -15395 24320 -15275
rect 24375 -15395 24495 -15275
rect 24540 -15395 24660 -15275
rect 24705 -15395 24825 -15275
rect 24870 -15395 24990 -15275
rect 25045 -15395 25165 -15275
rect 25210 -15395 25330 -15275
rect 25375 -15395 25495 -15275
rect 25540 -15395 25660 -15275
rect 25715 -15395 25835 -15275
rect 25880 -15395 26000 -15275
rect 26045 -15395 26165 -15275
rect 26210 -15395 26330 -15275
rect 26385 -15395 26505 -15275
rect 26550 -15395 26670 -15275
rect 26715 -15395 26835 -15275
rect 26880 -15395 27000 -15275
rect 27055 -15395 27175 -15275
rect 27220 -15395 27340 -15275
rect 27385 -15395 27505 -15275
rect 27550 -15395 27670 -15275
rect 27725 -15395 27845 -15275
rect 27890 -15395 28010 -15275
rect 28055 -15395 28175 -15275
rect 28220 -15395 28340 -15275
rect 28395 -15395 28515 -15275
rect 28560 -15395 28680 -15275
rect 28725 -15395 28845 -15275
rect 28890 -15395 29010 -15275
rect 29065 -15395 29185 -15275
rect 29230 -15395 29350 -15275
rect 29395 -15395 29515 -15275
rect 29560 -15395 29680 -15275
rect 24200 -15570 24320 -15450
rect 24375 -15570 24495 -15450
rect 24540 -15570 24660 -15450
rect 24705 -15570 24825 -15450
rect 24870 -15570 24990 -15450
rect 25045 -15570 25165 -15450
rect 25210 -15570 25330 -15450
rect 25375 -15570 25495 -15450
rect 25540 -15570 25660 -15450
rect 25715 -15570 25835 -15450
rect 25880 -15570 26000 -15450
rect 26045 -15570 26165 -15450
rect 26210 -15570 26330 -15450
rect 26385 -15570 26505 -15450
rect 26550 -15570 26670 -15450
rect 26715 -15570 26835 -15450
rect 26880 -15570 27000 -15450
rect 27055 -15570 27175 -15450
rect 27220 -15570 27340 -15450
rect 27385 -15570 27505 -15450
rect 27550 -15570 27670 -15450
rect 27725 -15570 27845 -15450
rect 27890 -15570 28010 -15450
rect 28055 -15570 28175 -15450
rect 28220 -15570 28340 -15450
rect 28395 -15570 28515 -15450
rect 28560 -15570 28680 -15450
rect 28725 -15570 28845 -15450
rect 28890 -15570 29010 -15450
rect 29065 -15570 29185 -15450
rect 29230 -15570 29350 -15450
rect 29395 -15570 29515 -15450
rect 29560 -15570 29680 -15450
<< metal5 >>
rect 7105 7160 12635 7185
rect 7105 7040 7130 7160
rect 7250 7040 7295 7160
rect 7415 7040 7460 7160
rect 7580 7040 7625 7160
rect 7745 7040 7800 7160
rect 7920 7040 7965 7160
rect 8085 7040 8130 7160
rect 8250 7040 8295 7160
rect 8415 7040 8470 7160
rect 8590 7040 8635 7160
rect 8755 7040 8800 7160
rect 8920 7040 8965 7160
rect 9085 7040 9140 7160
rect 9260 7040 9305 7160
rect 9425 7040 9470 7160
rect 9590 7040 9635 7160
rect 9755 7040 9810 7160
rect 9930 7040 9975 7160
rect 10095 7040 10140 7160
rect 10260 7040 10305 7160
rect 10425 7040 10480 7160
rect 10600 7040 10645 7160
rect 10765 7040 10810 7160
rect 10930 7040 10975 7160
rect 11095 7040 11150 7160
rect 11270 7040 11315 7160
rect 11435 7040 11480 7160
rect 11600 7040 11645 7160
rect 11765 7040 11820 7160
rect 11940 7040 11985 7160
rect 12105 7040 12150 7160
rect 12270 7040 12315 7160
rect 12435 7040 12490 7160
rect 12610 7040 12635 7160
rect 7105 6985 12635 7040
rect 7105 6865 7130 6985
rect 7250 6865 7295 6985
rect 7415 6865 7460 6985
rect 7580 6865 7625 6985
rect 7745 6865 7800 6985
rect 7920 6865 7965 6985
rect 8085 6865 8130 6985
rect 8250 6865 8295 6985
rect 8415 6865 8470 6985
rect 8590 6865 8635 6985
rect 8755 6865 8800 6985
rect 8920 6865 8965 6985
rect 9085 6865 9140 6985
rect 9260 6865 9305 6985
rect 9425 6865 9470 6985
rect 9590 6865 9635 6985
rect 9755 6865 9810 6985
rect 9930 6865 9975 6985
rect 10095 6865 10140 6985
rect 10260 6865 10305 6985
rect 10425 6865 10480 6985
rect 10600 6865 10645 6985
rect 10765 6865 10810 6985
rect 10930 6865 10975 6985
rect 11095 6865 11150 6985
rect 11270 6865 11315 6985
rect 11435 6865 11480 6985
rect 11600 6865 11645 6985
rect 11765 6865 11820 6985
rect 11940 6865 11985 6985
rect 12105 6865 12150 6985
rect 12270 6865 12315 6985
rect 12435 6865 12490 6985
rect 12610 6865 12635 6985
rect 7105 6820 12635 6865
rect 7105 6700 7130 6820
rect 7250 6700 7295 6820
rect 7415 6700 7460 6820
rect 7580 6700 7625 6820
rect 7745 6700 7800 6820
rect 7920 6700 7965 6820
rect 8085 6700 8130 6820
rect 8250 6700 8295 6820
rect 8415 6700 8470 6820
rect 8590 6700 8635 6820
rect 8755 6700 8800 6820
rect 8920 6700 8965 6820
rect 9085 6700 9140 6820
rect 9260 6700 9305 6820
rect 9425 6700 9470 6820
rect 9590 6700 9635 6820
rect 9755 6700 9810 6820
rect 9930 6700 9975 6820
rect 10095 6700 10140 6820
rect 10260 6700 10305 6820
rect 10425 6700 10480 6820
rect 10600 6700 10645 6820
rect 10765 6700 10810 6820
rect 10930 6700 10975 6820
rect 11095 6700 11150 6820
rect 11270 6700 11315 6820
rect 11435 6700 11480 6820
rect 11600 6700 11645 6820
rect 11765 6700 11820 6820
rect 11940 6700 11985 6820
rect 12105 6700 12150 6820
rect 12270 6700 12315 6820
rect 12435 6700 12490 6820
rect 12610 6700 12635 6820
rect 7105 6655 12635 6700
rect 7105 6535 7130 6655
rect 7250 6535 7295 6655
rect 7415 6535 7460 6655
rect 7580 6535 7625 6655
rect 7745 6535 7800 6655
rect 7920 6535 7965 6655
rect 8085 6535 8130 6655
rect 8250 6535 8295 6655
rect 8415 6535 8470 6655
rect 8590 6535 8635 6655
rect 8755 6535 8800 6655
rect 8920 6535 8965 6655
rect 9085 6535 9140 6655
rect 9260 6535 9305 6655
rect 9425 6535 9470 6655
rect 9590 6535 9635 6655
rect 9755 6535 9810 6655
rect 9930 6535 9975 6655
rect 10095 6535 10140 6655
rect 10260 6535 10305 6655
rect 10425 6535 10480 6655
rect 10600 6535 10645 6655
rect 10765 6535 10810 6655
rect 10930 6535 10975 6655
rect 11095 6535 11150 6655
rect 11270 6535 11315 6655
rect 11435 6535 11480 6655
rect 11600 6535 11645 6655
rect 11765 6535 11820 6655
rect 11940 6535 11985 6655
rect 12105 6535 12150 6655
rect 12270 6535 12315 6655
rect 12435 6535 12490 6655
rect 12610 6535 12635 6655
rect 7105 6490 12635 6535
rect 7105 6370 7130 6490
rect 7250 6370 7295 6490
rect 7415 6370 7460 6490
rect 7580 6370 7625 6490
rect 7745 6370 7800 6490
rect 7920 6370 7965 6490
rect 8085 6370 8130 6490
rect 8250 6370 8295 6490
rect 8415 6370 8470 6490
rect 8590 6370 8635 6490
rect 8755 6370 8800 6490
rect 8920 6370 8965 6490
rect 9085 6370 9140 6490
rect 9260 6370 9305 6490
rect 9425 6370 9470 6490
rect 9590 6370 9635 6490
rect 9755 6370 9810 6490
rect 9930 6370 9975 6490
rect 10095 6370 10140 6490
rect 10260 6370 10305 6490
rect 10425 6370 10480 6490
rect 10600 6370 10645 6490
rect 10765 6370 10810 6490
rect 10930 6370 10975 6490
rect 11095 6370 11150 6490
rect 11270 6370 11315 6490
rect 11435 6370 11480 6490
rect 11600 6370 11645 6490
rect 11765 6370 11820 6490
rect 11940 6370 11985 6490
rect 12105 6370 12150 6490
rect 12270 6370 12315 6490
rect 12435 6370 12490 6490
rect 12610 6370 12635 6490
rect 7105 6315 12635 6370
rect 7105 6195 7130 6315
rect 7250 6195 7295 6315
rect 7415 6195 7460 6315
rect 7580 6195 7625 6315
rect 7745 6195 7800 6315
rect 7920 6195 7965 6315
rect 8085 6195 8130 6315
rect 8250 6195 8295 6315
rect 8415 6195 8470 6315
rect 8590 6195 8635 6315
rect 8755 6195 8800 6315
rect 8920 6195 8965 6315
rect 9085 6195 9140 6315
rect 9260 6195 9305 6315
rect 9425 6195 9470 6315
rect 9590 6195 9635 6315
rect 9755 6195 9810 6315
rect 9930 6195 9975 6315
rect 10095 6195 10140 6315
rect 10260 6195 10305 6315
rect 10425 6195 10480 6315
rect 10600 6195 10645 6315
rect 10765 6195 10810 6315
rect 10930 6195 10975 6315
rect 11095 6195 11150 6315
rect 11270 6195 11315 6315
rect 11435 6195 11480 6315
rect 11600 6195 11645 6315
rect 11765 6195 11820 6315
rect 11940 6195 11985 6315
rect 12105 6195 12150 6315
rect 12270 6195 12315 6315
rect 12435 6195 12490 6315
rect 12610 6195 12635 6315
rect 7105 6150 12635 6195
rect 7105 6030 7130 6150
rect 7250 6030 7295 6150
rect 7415 6030 7460 6150
rect 7580 6030 7625 6150
rect 7745 6030 7800 6150
rect 7920 6030 7965 6150
rect 8085 6030 8130 6150
rect 8250 6030 8295 6150
rect 8415 6030 8470 6150
rect 8590 6030 8635 6150
rect 8755 6030 8800 6150
rect 8920 6030 8965 6150
rect 9085 6030 9140 6150
rect 9260 6030 9305 6150
rect 9425 6030 9470 6150
rect 9590 6030 9635 6150
rect 9755 6030 9810 6150
rect 9930 6030 9975 6150
rect 10095 6030 10140 6150
rect 10260 6030 10305 6150
rect 10425 6030 10480 6150
rect 10600 6030 10645 6150
rect 10765 6030 10810 6150
rect 10930 6030 10975 6150
rect 11095 6030 11150 6150
rect 11270 6030 11315 6150
rect 11435 6030 11480 6150
rect 11600 6030 11645 6150
rect 11765 6030 11820 6150
rect 11940 6030 11985 6150
rect 12105 6030 12150 6150
rect 12270 6030 12315 6150
rect 12435 6030 12490 6150
rect 12610 6030 12635 6150
rect 7105 5985 12635 6030
rect 7105 5865 7130 5985
rect 7250 5865 7295 5985
rect 7415 5865 7460 5985
rect 7580 5865 7625 5985
rect 7745 5865 7800 5985
rect 7920 5865 7965 5985
rect 8085 5865 8130 5985
rect 8250 5865 8295 5985
rect 8415 5865 8470 5985
rect 8590 5865 8635 5985
rect 8755 5865 8800 5985
rect 8920 5865 8965 5985
rect 9085 5865 9140 5985
rect 9260 5865 9305 5985
rect 9425 5865 9470 5985
rect 9590 5865 9635 5985
rect 9755 5865 9810 5985
rect 9930 5865 9975 5985
rect 10095 5865 10140 5985
rect 10260 5865 10305 5985
rect 10425 5865 10480 5985
rect 10600 5865 10645 5985
rect 10765 5865 10810 5985
rect 10930 5865 10975 5985
rect 11095 5865 11150 5985
rect 11270 5865 11315 5985
rect 11435 5865 11480 5985
rect 11600 5865 11645 5985
rect 11765 5865 11820 5985
rect 11940 5865 11985 5985
rect 12105 5865 12150 5985
rect 12270 5865 12315 5985
rect 12435 5865 12490 5985
rect 12610 5865 12635 5985
rect 7105 5820 12635 5865
rect 7105 5700 7130 5820
rect 7250 5700 7295 5820
rect 7415 5700 7460 5820
rect 7580 5700 7625 5820
rect 7745 5700 7800 5820
rect 7920 5700 7965 5820
rect 8085 5700 8130 5820
rect 8250 5700 8295 5820
rect 8415 5700 8470 5820
rect 8590 5700 8635 5820
rect 8755 5700 8800 5820
rect 8920 5700 8965 5820
rect 9085 5700 9140 5820
rect 9260 5700 9305 5820
rect 9425 5700 9470 5820
rect 9590 5700 9635 5820
rect 9755 5700 9810 5820
rect 9930 5700 9975 5820
rect 10095 5700 10140 5820
rect 10260 5700 10305 5820
rect 10425 5700 10480 5820
rect 10600 5700 10645 5820
rect 10765 5700 10810 5820
rect 10930 5700 10975 5820
rect 11095 5700 11150 5820
rect 11270 5700 11315 5820
rect 11435 5700 11480 5820
rect 11600 5700 11645 5820
rect 11765 5700 11820 5820
rect 11940 5700 11985 5820
rect 12105 5700 12150 5820
rect 12270 5700 12315 5820
rect 12435 5700 12490 5820
rect 12610 5700 12635 5820
rect 7105 5645 12635 5700
rect 7105 5525 7130 5645
rect 7250 5525 7295 5645
rect 7415 5525 7460 5645
rect 7580 5525 7625 5645
rect 7745 5525 7800 5645
rect 7920 5525 7965 5645
rect 8085 5525 8130 5645
rect 8250 5525 8295 5645
rect 8415 5525 8470 5645
rect 8590 5525 8635 5645
rect 8755 5525 8800 5645
rect 8920 5525 8965 5645
rect 9085 5525 9140 5645
rect 9260 5525 9305 5645
rect 9425 5525 9470 5645
rect 9590 5525 9635 5645
rect 9755 5525 9810 5645
rect 9930 5525 9975 5645
rect 10095 5525 10140 5645
rect 10260 5525 10305 5645
rect 10425 5525 10480 5645
rect 10600 5525 10645 5645
rect 10765 5525 10810 5645
rect 10930 5525 10975 5645
rect 11095 5525 11150 5645
rect 11270 5525 11315 5645
rect 11435 5525 11480 5645
rect 11600 5525 11645 5645
rect 11765 5525 11820 5645
rect 11940 5525 11985 5645
rect 12105 5525 12150 5645
rect 12270 5525 12315 5645
rect 12435 5525 12490 5645
rect 12610 5525 12635 5645
rect 7105 5480 12635 5525
rect 7105 5360 7130 5480
rect 7250 5360 7295 5480
rect 7415 5360 7460 5480
rect 7580 5360 7625 5480
rect 7745 5360 7800 5480
rect 7920 5360 7965 5480
rect 8085 5360 8130 5480
rect 8250 5360 8295 5480
rect 8415 5360 8470 5480
rect 8590 5360 8635 5480
rect 8755 5360 8800 5480
rect 8920 5360 8965 5480
rect 9085 5360 9140 5480
rect 9260 5360 9305 5480
rect 9425 5360 9470 5480
rect 9590 5360 9635 5480
rect 9755 5360 9810 5480
rect 9930 5360 9975 5480
rect 10095 5360 10140 5480
rect 10260 5360 10305 5480
rect 10425 5360 10480 5480
rect 10600 5360 10645 5480
rect 10765 5360 10810 5480
rect 10930 5360 10975 5480
rect 11095 5360 11150 5480
rect 11270 5360 11315 5480
rect 11435 5360 11480 5480
rect 11600 5360 11645 5480
rect 11765 5360 11820 5480
rect 11940 5360 11985 5480
rect 12105 5360 12150 5480
rect 12270 5360 12315 5480
rect 12435 5360 12490 5480
rect 12610 5360 12635 5480
rect 7105 5315 12635 5360
rect 7105 5195 7130 5315
rect 7250 5195 7295 5315
rect 7415 5195 7460 5315
rect 7580 5195 7625 5315
rect 7745 5195 7800 5315
rect 7920 5195 7965 5315
rect 8085 5195 8130 5315
rect 8250 5195 8295 5315
rect 8415 5195 8470 5315
rect 8590 5195 8635 5315
rect 8755 5195 8800 5315
rect 8920 5195 8965 5315
rect 9085 5195 9140 5315
rect 9260 5195 9305 5315
rect 9425 5195 9470 5315
rect 9590 5195 9635 5315
rect 9755 5195 9810 5315
rect 9930 5195 9975 5315
rect 10095 5195 10140 5315
rect 10260 5195 10305 5315
rect 10425 5195 10480 5315
rect 10600 5195 10645 5315
rect 10765 5195 10810 5315
rect 10930 5195 10975 5315
rect 11095 5195 11150 5315
rect 11270 5195 11315 5315
rect 11435 5195 11480 5315
rect 11600 5195 11645 5315
rect 11765 5195 11820 5315
rect 11940 5195 11985 5315
rect 12105 5195 12150 5315
rect 12270 5195 12315 5315
rect 12435 5195 12490 5315
rect 12610 5195 12635 5315
rect 7105 5150 12635 5195
rect 7105 5030 7130 5150
rect 7250 5030 7295 5150
rect 7415 5030 7460 5150
rect 7580 5030 7625 5150
rect 7745 5030 7800 5150
rect 7920 5030 7965 5150
rect 8085 5030 8130 5150
rect 8250 5030 8295 5150
rect 8415 5030 8470 5150
rect 8590 5030 8635 5150
rect 8755 5030 8800 5150
rect 8920 5030 8965 5150
rect 9085 5030 9140 5150
rect 9260 5030 9305 5150
rect 9425 5030 9470 5150
rect 9590 5030 9635 5150
rect 9755 5030 9810 5150
rect 9930 5030 9975 5150
rect 10095 5030 10140 5150
rect 10260 5030 10305 5150
rect 10425 5030 10480 5150
rect 10600 5030 10645 5150
rect 10765 5030 10810 5150
rect 10930 5030 10975 5150
rect 11095 5030 11150 5150
rect 11270 5030 11315 5150
rect 11435 5030 11480 5150
rect 11600 5030 11645 5150
rect 11765 5030 11820 5150
rect 11940 5030 11985 5150
rect 12105 5030 12150 5150
rect 12270 5030 12315 5150
rect 12435 5030 12490 5150
rect 12610 5030 12635 5150
rect 7105 4975 12635 5030
rect 7105 4855 7130 4975
rect 7250 4855 7295 4975
rect 7415 4855 7460 4975
rect 7580 4855 7625 4975
rect 7745 4855 7800 4975
rect 7920 4855 7965 4975
rect 8085 4855 8130 4975
rect 8250 4855 8295 4975
rect 8415 4855 8470 4975
rect 8590 4855 8635 4975
rect 8755 4855 8800 4975
rect 8920 4855 8965 4975
rect 9085 4855 9140 4975
rect 9260 4855 9305 4975
rect 9425 4855 9470 4975
rect 9590 4855 9635 4975
rect 9755 4855 9810 4975
rect 9930 4855 9975 4975
rect 10095 4855 10140 4975
rect 10260 4855 10305 4975
rect 10425 4855 10480 4975
rect 10600 4855 10645 4975
rect 10765 4855 10810 4975
rect 10930 4855 10975 4975
rect 11095 4855 11150 4975
rect 11270 4855 11315 4975
rect 11435 4855 11480 4975
rect 11600 4855 11645 4975
rect 11765 4855 11820 4975
rect 11940 4855 11985 4975
rect 12105 4855 12150 4975
rect 12270 4855 12315 4975
rect 12435 4855 12490 4975
rect 12610 4855 12635 4975
rect 7105 4810 12635 4855
rect 7105 4690 7130 4810
rect 7250 4690 7295 4810
rect 7415 4690 7460 4810
rect 7580 4690 7625 4810
rect 7745 4690 7800 4810
rect 7920 4690 7965 4810
rect 8085 4690 8130 4810
rect 8250 4690 8295 4810
rect 8415 4690 8470 4810
rect 8590 4690 8635 4810
rect 8755 4690 8800 4810
rect 8920 4690 8965 4810
rect 9085 4690 9140 4810
rect 9260 4690 9305 4810
rect 9425 4690 9470 4810
rect 9590 4690 9635 4810
rect 9755 4690 9810 4810
rect 9930 4690 9975 4810
rect 10095 4690 10140 4810
rect 10260 4690 10305 4810
rect 10425 4690 10480 4810
rect 10600 4690 10645 4810
rect 10765 4690 10810 4810
rect 10930 4690 10975 4810
rect 11095 4690 11150 4810
rect 11270 4690 11315 4810
rect 11435 4690 11480 4810
rect 11600 4690 11645 4810
rect 11765 4690 11820 4810
rect 11940 4690 11985 4810
rect 12105 4690 12150 4810
rect 12270 4690 12315 4810
rect 12435 4690 12490 4810
rect 12610 4690 12635 4810
rect 7105 4645 12635 4690
rect 7105 4525 7130 4645
rect 7250 4525 7295 4645
rect 7415 4525 7460 4645
rect 7580 4525 7625 4645
rect 7745 4525 7800 4645
rect 7920 4525 7965 4645
rect 8085 4525 8130 4645
rect 8250 4525 8295 4645
rect 8415 4525 8470 4645
rect 8590 4525 8635 4645
rect 8755 4525 8800 4645
rect 8920 4525 8965 4645
rect 9085 4525 9140 4645
rect 9260 4525 9305 4645
rect 9425 4525 9470 4645
rect 9590 4525 9635 4645
rect 9755 4525 9810 4645
rect 9930 4525 9975 4645
rect 10095 4525 10140 4645
rect 10260 4525 10305 4645
rect 10425 4525 10480 4645
rect 10600 4525 10645 4645
rect 10765 4525 10810 4645
rect 10930 4525 10975 4645
rect 11095 4525 11150 4645
rect 11270 4525 11315 4645
rect 11435 4525 11480 4645
rect 11600 4525 11645 4645
rect 11765 4525 11820 4645
rect 11940 4525 11985 4645
rect 12105 4525 12150 4645
rect 12270 4525 12315 4645
rect 12435 4525 12490 4645
rect 12610 4525 12635 4645
rect 7105 4480 12635 4525
rect 7105 4360 7130 4480
rect 7250 4360 7295 4480
rect 7415 4360 7460 4480
rect 7580 4360 7625 4480
rect 7745 4360 7800 4480
rect 7920 4360 7965 4480
rect 8085 4360 8130 4480
rect 8250 4360 8295 4480
rect 8415 4360 8470 4480
rect 8590 4360 8635 4480
rect 8755 4360 8800 4480
rect 8920 4360 8965 4480
rect 9085 4360 9140 4480
rect 9260 4360 9305 4480
rect 9425 4360 9470 4480
rect 9590 4360 9635 4480
rect 9755 4360 9810 4480
rect 9930 4360 9975 4480
rect 10095 4360 10140 4480
rect 10260 4360 10305 4480
rect 10425 4360 10480 4480
rect 10600 4360 10645 4480
rect 10765 4360 10810 4480
rect 10930 4360 10975 4480
rect 11095 4360 11150 4480
rect 11270 4360 11315 4480
rect 11435 4360 11480 4480
rect 11600 4360 11645 4480
rect 11765 4360 11820 4480
rect 11940 4360 11985 4480
rect 12105 4360 12150 4480
rect 12270 4360 12315 4480
rect 12435 4360 12490 4480
rect 12610 4360 12635 4480
rect 7105 4305 12635 4360
rect 7105 4185 7130 4305
rect 7250 4185 7295 4305
rect 7415 4185 7460 4305
rect 7580 4185 7625 4305
rect 7745 4185 7800 4305
rect 7920 4185 7965 4305
rect 8085 4185 8130 4305
rect 8250 4185 8295 4305
rect 8415 4185 8470 4305
rect 8590 4185 8635 4305
rect 8755 4185 8800 4305
rect 8920 4185 8965 4305
rect 9085 4185 9140 4305
rect 9260 4185 9305 4305
rect 9425 4185 9470 4305
rect 9590 4185 9635 4305
rect 9755 4185 9810 4305
rect 9930 4185 9975 4305
rect 10095 4185 10140 4305
rect 10260 4185 10305 4305
rect 10425 4185 10480 4305
rect 10600 4185 10645 4305
rect 10765 4185 10810 4305
rect 10930 4185 10975 4305
rect 11095 4185 11150 4305
rect 11270 4185 11315 4305
rect 11435 4185 11480 4305
rect 11600 4185 11645 4305
rect 11765 4185 11820 4305
rect 11940 4185 11985 4305
rect 12105 4185 12150 4305
rect 12270 4185 12315 4305
rect 12435 4185 12490 4305
rect 12610 4185 12635 4305
rect 7105 4140 12635 4185
rect 7105 4020 7130 4140
rect 7250 4020 7295 4140
rect 7415 4020 7460 4140
rect 7580 4020 7625 4140
rect 7745 4020 7800 4140
rect 7920 4020 7965 4140
rect 8085 4020 8130 4140
rect 8250 4020 8295 4140
rect 8415 4020 8470 4140
rect 8590 4020 8635 4140
rect 8755 4020 8800 4140
rect 8920 4020 8965 4140
rect 9085 4020 9140 4140
rect 9260 4020 9305 4140
rect 9425 4020 9470 4140
rect 9590 4020 9635 4140
rect 9755 4020 9810 4140
rect 9930 4020 9975 4140
rect 10095 4020 10140 4140
rect 10260 4020 10305 4140
rect 10425 4020 10480 4140
rect 10600 4020 10645 4140
rect 10765 4020 10810 4140
rect 10930 4020 10975 4140
rect 11095 4020 11150 4140
rect 11270 4020 11315 4140
rect 11435 4020 11480 4140
rect 11600 4020 11645 4140
rect 11765 4020 11820 4140
rect 11940 4020 11985 4140
rect 12105 4020 12150 4140
rect 12270 4020 12315 4140
rect 12435 4020 12490 4140
rect 12610 4020 12635 4140
rect 7105 3975 12635 4020
rect 7105 3855 7130 3975
rect 7250 3855 7295 3975
rect 7415 3855 7460 3975
rect 7580 3855 7625 3975
rect 7745 3855 7800 3975
rect 7920 3855 7965 3975
rect 8085 3855 8130 3975
rect 8250 3855 8295 3975
rect 8415 3855 8470 3975
rect 8590 3855 8635 3975
rect 8755 3855 8800 3975
rect 8920 3855 8965 3975
rect 9085 3855 9140 3975
rect 9260 3855 9305 3975
rect 9425 3855 9470 3975
rect 9590 3855 9635 3975
rect 9755 3855 9810 3975
rect 9930 3855 9975 3975
rect 10095 3855 10140 3975
rect 10260 3855 10305 3975
rect 10425 3855 10480 3975
rect 10600 3855 10645 3975
rect 10765 3855 10810 3975
rect 10930 3855 10975 3975
rect 11095 3855 11150 3975
rect 11270 3855 11315 3975
rect 11435 3855 11480 3975
rect 11600 3855 11645 3975
rect 11765 3855 11820 3975
rect 11940 3855 11985 3975
rect 12105 3855 12150 3975
rect 12270 3855 12315 3975
rect 12435 3855 12490 3975
rect 12610 3855 12635 3975
rect 7105 3810 12635 3855
rect 7105 3690 7130 3810
rect 7250 3690 7295 3810
rect 7415 3690 7460 3810
rect 7580 3690 7625 3810
rect 7745 3690 7800 3810
rect 7920 3690 7965 3810
rect 8085 3690 8130 3810
rect 8250 3690 8295 3810
rect 8415 3690 8470 3810
rect 8590 3690 8635 3810
rect 8755 3690 8800 3810
rect 8920 3690 8965 3810
rect 9085 3690 9140 3810
rect 9260 3690 9305 3810
rect 9425 3690 9470 3810
rect 9590 3690 9635 3810
rect 9755 3690 9810 3810
rect 9930 3690 9975 3810
rect 10095 3690 10140 3810
rect 10260 3690 10305 3810
rect 10425 3690 10480 3810
rect 10600 3690 10645 3810
rect 10765 3690 10810 3810
rect 10930 3690 10975 3810
rect 11095 3690 11150 3810
rect 11270 3690 11315 3810
rect 11435 3690 11480 3810
rect 11600 3690 11645 3810
rect 11765 3690 11820 3810
rect 11940 3690 11985 3810
rect 12105 3690 12150 3810
rect 12270 3690 12315 3810
rect 12435 3690 12490 3810
rect 12610 3690 12635 3810
rect 7105 3635 12635 3690
rect 7105 3515 7130 3635
rect 7250 3515 7295 3635
rect 7415 3515 7460 3635
rect 7580 3515 7625 3635
rect 7745 3515 7800 3635
rect 7920 3515 7965 3635
rect 8085 3515 8130 3635
rect 8250 3515 8295 3635
rect 8415 3515 8470 3635
rect 8590 3515 8635 3635
rect 8755 3515 8800 3635
rect 8920 3515 8965 3635
rect 9085 3515 9140 3635
rect 9260 3515 9305 3635
rect 9425 3515 9470 3635
rect 9590 3515 9635 3635
rect 9755 3515 9810 3635
rect 9930 3515 9975 3635
rect 10095 3515 10140 3635
rect 10260 3515 10305 3635
rect 10425 3515 10480 3635
rect 10600 3515 10645 3635
rect 10765 3515 10810 3635
rect 10930 3515 10975 3635
rect 11095 3515 11150 3635
rect 11270 3515 11315 3635
rect 11435 3515 11480 3635
rect 11600 3515 11645 3635
rect 11765 3515 11820 3635
rect 11940 3515 11985 3635
rect 12105 3515 12150 3635
rect 12270 3515 12315 3635
rect 12435 3515 12490 3635
rect 12610 3515 12635 3635
rect 7105 3470 12635 3515
rect 7105 3350 7130 3470
rect 7250 3350 7295 3470
rect 7415 3350 7460 3470
rect 7580 3350 7625 3470
rect 7745 3350 7800 3470
rect 7920 3350 7965 3470
rect 8085 3350 8130 3470
rect 8250 3350 8295 3470
rect 8415 3350 8470 3470
rect 8590 3350 8635 3470
rect 8755 3350 8800 3470
rect 8920 3350 8965 3470
rect 9085 3350 9140 3470
rect 9260 3350 9305 3470
rect 9425 3350 9470 3470
rect 9590 3350 9635 3470
rect 9755 3350 9810 3470
rect 9930 3350 9975 3470
rect 10095 3350 10140 3470
rect 10260 3350 10305 3470
rect 10425 3350 10480 3470
rect 10600 3350 10645 3470
rect 10765 3350 10810 3470
rect 10930 3350 10975 3470
rect 11095 3350 11150 3470
rect 11270 3350 11315 3470
rect 11435 3350 11480 3470
rect 11600 3350 11645 3470
rect 11765 3350 11820 3470
rect 11940 3350 11985 3470
rect 12105 3350 12150 3470
rect 12270 3350 12315 3470
rect 12435 3350 12490 3470
rect 12610 3350 12635 3470
rect 7105 3305 12635 3350
rect 7105 3185 7130 3305
rect 7250 3185 7295 3305
rect 7415 3185 7460 3305
rect 7580 3185 7625 3305
rect 7745 3185 7800 3305
rect 7920 3185 7965 3305
rect 8085 3185 8130 3305
rect 8250 3185 8295 3305
rect 8415 3185 8470 3305
rect 8590 3185 8635 3305
rect 8755 3185 8800 3305
rect 8920 3185 8965 3305
rect 9085 3185 9140 3305
rect 9260 3185 9305 3305
rect 9425 3185 9470 3305
rect 9590 3185 9635 3305
rect 9755 3185 9810 3305
rect 9930 3185 9975 3305
rect 10095 3185 10140 3305
rect 10260 3185 10305 3305
rect 10425 3185 10480 3305
rect 10600 3185 10645 3305
rect 10765 3185 10810 3305
rect 10930 3185 10975 3305
rect 11095 3185 11150 3305
rect 11270 3185 11315 3305
rect 11435 3185 11480 3305
rect 11600 3185 11645 3305
rect 11765 3185 11820 3305
rect 11940 3185 11985 3305
rect 12105 3185 12150 3305
rect 12270 3185 12315 3305
rect 12435 3185 12490 3305
rect 12610 3185 12635 3305
rect 7105 3140 12635 3185
rect 7105 3020 7130 3140
rect 7250 3020 7295 3140
rect 7415 3020 7460 3140
rect 7580 3020 7625 3140
rect 7745 3020 7800 3140
rect 7920 3020 7965 3140
rect 8085 3020 8130 3140
rect 8250 3020 8295 3140
rect 8415 3020 8470 3140
rect 8590 3020 8635 3140
rect 8755 3020 8800 3140
rect 8920 3020 8965 3140
rect 9085 3020 9140 3140
rect 9260 3020 9305 3140
rect 9425 3020 9470 3140
rect 9590 3020 9635 3140
rect 9755 3020 9810 3140
rect 9930 3020 9975 3140
rect 10095 3020 10140 3140
rect 10260 3020 10305 3140
rect 10425 3020 10480 3140
rect 10600 3020 10645 3140
rect 10765 3020 10810 3140
rect 10930 3020 10975 3140
rect 11095 3020 11150 3140
rect 11270 3020 11315 3140
rect 11435 3020 11480 3140
rect 11600 3020 11645 3140
rect 11765 3020 11820 3140
rect 11940 3020 11985 3140
rect 12105 3020 12150 3140
rect 12270 3020 12315 3140
rect 12435 3020 12490 3140
rect 12610 3020 12635 3140
rect 7105 2965 12635 3020
rect 7105 2845 7130 2965
rect 7250 2845 7295 2965
rect 7415 2845 7460 2965
rect 7580 2845 7625 2965
rect 7745 2845 7800 2965
rect 7920 2845 7965 2965
rect 8085 2845 8130 2965
rect 8250 2845 8295 2965
rect 8415 2845 8470 2965
rect 8590 2845 8635 2965
rect 8755 2845 8800 2965
rect 8920 2845 8965 2965
rect 9085 2845 9140 2965
rect 9260 2845 9305 2965
rect 9425 2845 9470 2965
rect 9590 2845 9635 2965
rect 9755 2845 9810 2965
rect 9930 2845 9975 2965
rect 10095 2845 10140 2965
rect 10260 2845 10305 2965
rect 10425 2845 10480 2965
rect 10600 2845 10645 2965
rect 10765 2845 10810 2965
rect 10930 2845 10975 2965
rect 11095 2845 11150 2965
rect 11270 2845 11315 2965
rect 11435 2845 11480 2965
rect 11600 2845 11645 2965
rect 11765 2845 11820 2965
rect 11940 2845 11985 2965
rect 12105 2845 12150 2965
rect 12270 2845 12315 2965
rect 12435 2845 12490 2965
rect 12610 2845 12635 2965
rect 7105 2800 12635 2845
rect 7105 2680 7130 2800
rect 7250 2680 7295 2800
rect 7415 2680 7460 2800
rect 7580 2680 7625 2800
rect 7745 2680 7800 2800
rect 7920 2680 7965 2800
rect 8085 2680 8130 2800
rect 8250 2680 8295 2800
rect 8415 2680 8470 2800
rect 8590 2680 8635 2800
rect 8755 2680 8800 2800
rect 8920 2680 8965 2800
rect 9085 2680 9140 2800
rect 9260 2680 9305 2800
rect 9425 2680 9470 2800
rect 9590 2680 9635 2800
rect 9755 2680 9810 2800
rect 9930 2680 9975 2800
rect 10095 2680 10140 2800
rect 10260 2680 10305 2800
rect 10425 2680 10480 2800
rect 10600 2680 10645 2800
rect 10765 2680 10810 2800
rect 10930 2680 10975 2800
rect 11095 2680 11150 2800
rect 11270 2680 11315 2800
rect 11435 2680 11480 2800
rect 11600 2680 11645 2800
rect 11765 2680 11820 2800
rect 11940 2680 11985 2800
rect 12105 2680 12150 2800
rect 12270 2680 12315 2800
rect 12435 2680 12490 2800
rect 12610 2680 12635 2800
rect 7105 2635 12635 2680
rect 7105 2515 7130 2635
rect 7250 2515 7295 2635
rect 7415 2515 7460 2635
rect 7580 2515 7625 2635
rect 7745 2515 7800 2635
rect 7920 2515 7965 2635
rect 8085 2515 8130 2635
rect 8250 2515 8295 2635
rect 8415 2515 8470 2635
rect 8590 2515 8635 2635
rect 8755 2515 8800 2635
rect 8920 2515 8965 2635
rect 9085 2515 9140 2635
rect 9260 2515 9305 2635
rect 9425 2515 9470 2635
rect 9590 2515 9635 2635
rect 9755 2515 9810 2635
rect 9930 2515 9975 2635
rect 10095 2515 10140 2635
rect 10260 2515 10305 2635
rect 10425 2515 10480 2635
rect 10600 2515 10645 2635
rect 10765 2515 10810 2635
rect 10930 2515 10975 2635
rect 11095 2515 11150 2635
rect 11270 2515 11315 2635
rect 11435 2515 11480 2635
rect 11600 2515 11645 2635
rect 11765 2515 11820 2635
rect 11940 2515 11985 2635
rect 12105 2515 12150 2635
rect 12270 2515 12315 2635
rect 12435 2515 12490 2635
rect 12610 2515 12635 2635
rect 7105 2470 12635 2515
rect 7105 2350 7130 2470
rect 7250 2350 7295 2470
rect 7415 2350 7460 2470
rect 7580 2350 7625 2470
rect 7745 2350 7800 2470
rect 7920 2350 7965 2470
rect 8085 2350 8130 2470
rect 8250 2350 8295 2470
rect 8415 2350 8470 2470
rect 8590 2350 8635 2470
rect 8755 2350 8800 2470
rect 8920 2350 8965 2470
rect 9085 2350 9140 2470
rect 9260 2350 9305 2470
rect 9425 2350 9470 2470
rect 9590 2350 9635 2470
rect 9755 2350 9810 2470
rect 9930 2350 9975 2470
rect 10095 2350 10140 2470
rect 10260 2350 10305 2470
rect 10425 2350 10480 2470
rect 10600 2350 10645 2470
rect 10765 2350 10810 2470
rect 10930 2350 10975 2470
rect 11095 2350 11150 2470
rect 11270 2350 11315 2470
rect 11435 2350 11480 2470
rect 11600 2350 11645 2470
rect 11765 2350 11820 2470
rect 11940 2350 11985 2470
rect 12105 2350 12150 2470
rect 12270 2350 12315 2470
rect 12435 2350 12490 2470
rect 12610 2350 12635 2470
rect 7105 2295 12635 2350
rect 7105 2175 7130 2295
rect 7250 2175 7295 2295
rect 7415 2175 7460 2295
rect 7580 2175 7625 2295
rect 7745 2175 7800 2295
rect 7920 2175 7965 2295
rect 8085 2175 8130 2295
rect 8250 2175 8295 2295
rect 8415 2175 8470 2295
rect 8590 2175 8635 2295
rect 8755 2175 8800 2295
rect 8920 2175 8965 2295
rect 9085 2175 9140 2295
rect 9260 2175 9305 2295
rect 9425 2175 9470 2295
rect 9590 2175 9635 2295
rect 9755 2175 9810 2295
rect 9930 2175 9975 2295
rect 10095 2175 10140 2295
rect 10260 2175 10305 2295
rect 10425 2175 10480 2295
rect 10600 2175 10645 2295
rect 10765 2175 10810 2295
rect 10930 2175 10975 2295
rect 11095 2175 11150 2295
rect 11270 2175 11315 2295
rect 11435 2175 11480 2295
rect 11600 2175 11645 2295
rect 11765 2175 11820 2295
rect 11940 2175 11985 2295
rect 12105 2175 12150 2295
rect 12270 2175 12315 2295
rect 12435 2175 12490 2295
rect 12610 2175 12635 2295
rect 7105 2130 12635 2175
rect 7105 2010 7130 2130
rect 7250 2010 7295 2130
rect 7415 2010 7460 2130
rect 7580 2010 7625 2130
rect 7745 2010 7800 2130
rect 7920 2010 7965 2130
rect 8085 2010 8130 2130
rect 8250 2010 8295 2130
rect 8415 2010 8470 2130
rect 8590 2010 8635 2130
rect 8755 2010 8800 2130
rect 8920 2010 8965 2130
rect 9085 2010 9140 2130
rect 9260 2010 9305 2130
rect 9425 2010 9470 2130
rect 9590 2010 9635 2130
rect 9755 2010 9810 2130
rect 9930 2010 9975 2130
rect 10095 2010 10140 2130
rect 10260 2010 10305 2130
rect 10425 2010 10480 2130
rect 10600 2010 10645 2130
rect 10765 2010 10810 2130
rect 10930 2010 10975 2130
rect 11095 2010 11150 2130
rect 11270 2010 11315 2130
rect 11435 2010 11480 2130
rect 11600 2010 11645 2130
rect 11765 2010 11820 2130
rect 11940 2010 11985 2130
rect 12105 2010 12150 2130
rect 12270 2010 12315 2130
rect 12435 2010 12490 2130
rect 12610 2010 12635 2130
rect 7105 1965 12635 2010
rect 7105 1845 7130 1965
rect 7250 1845 7295 1965
rect 7415 1845 7460 1965
rect 7580 1845 7625 1965
rect 7745 1845 7800 1965
rect 7920 1845 7965 1965
rect 8085 1845 8130 1965
rect 8250 1845 8295 1965
rect 8415 1845 8470 1965
rect 8590 1845 8635 1965
rect 8755 1845 8800 1965
rect 8920 1845 8965 1965
rect 9085 1845 9140 1965
rect 9260 1845 9305 1965
rect 9425 1845 9470 1965
rect 9590 1845 9635 1965
rect 9755 1845 9810 1965
rect 9930 1845 9975 1965
rect 10095 1845 10140 1965
rect 10260 1845 10305 1965
rect 10425 1845 10480 1965
rect 10600 1845 10645 1965
rect 10765 1845 10810 1965
rect 10930 1845 10975 1965
rect 11095 1845 11150 1965
rect 11270 1845 11315 1965
rect 11435 1845 11480 1965
rect 11600 1845 11645 1965
rect 11765 1845 11820 1965
rect 11940 1845 11985 1965
rect 12105 1845 12150 1965
rect 12270 1845 12315 1965
rect 12435 1845 12490 1965
rect 12610 1845 12635 1965
rect 7105 1800 12635 1845
rect 7105 1680 7130 1800
rect 7250 1680 7295 1800
rect 7415 1680 7460 1800
rect 7580 1680 7625 1800
rect 7745 1680 7800 1800
rect 7920 1680 7965 1800
rect 8085 1680 8130 1800
rect 8250 1680 8295 1800
rect 8415 1680 8470 1800
rect 8590 1680 8635 1800
rect 8755 1680 8800 1800
rect 8920 1680 8965 1800
rect 9085 1680 9140 1800
rect 9260 1680 9305 1800
rect 9425 1680 9470 1800
rect 9590 1680 9635 1800
rect 9755 1680 9810 1800
rect 9930 1680 9975 1800
rect 10095 1680 10140 1800
rect 10260 1680 10305 1800
rect 10425 1680 10480 1800
rect 10600 1680 10645 1800
rect 10765 1680 10810 1800
rect 10930 1680 10975 1800
rect 11095 1680 11150 1800
rect 11270 1680 11315 1800
rect 11435 1680 11480 1800
rect 11600 1680 11645 1800
rect 11765 1680 11820 1800
rect 11940 1680 11985 1800
rect 12105 1680 12150 1800
rect 12270 1680 12315 1800
rect 12435 1680 12490 1800
rect 12610 1680 12635 1800
rect 7105 1610 12635 1680
rect 12795 7160 18325 7185
rect 12795 7040 12820 7160
rect 12940 7040 12985 7160
rect 13105 7040 13150 7160
rect 13270 7040 13315 7160
rect 13435 7040 13490 7160
rect 13610 7040 13655 7160
rect 13775 7040 13820 7160
rect 13940 7040 13985 7160
rect 14105 7040 14160 7160
rect 14280 7040 14325 7160
rect 14445 7040 14490 7160
rect 14610 7040 14655 7160
rect 14775 7040 14830 7160
rect 14950 7040 14995 7160
rect 15115 7040 15160 7160
rect 15280 7040 15325 7160
rect 15445 7040 15500 7160
rect 15620 7040 15665 7160
rect 15785 7040 15830 7160
rect 15950 7040 15995 7160
rect 16115 7040 16170 7160
rect 16290 7040 16335 7160
rect 16455 7040 16500 7160
rect 16620 7040 16665 7160
rect 16785 7040 16840 7160
rect 16960 7040 17005 7160
rect 17125 7040 17170 7160
rect 17290 7040 17335 7160
rect 17455 7040 17510 7160
rect 17630 7040 17675 7160
rect 17795 7040 17840 7160
rect 17960 7040 18005 7160
rect 18125 7040 18180 7160
rect 18300 7040 18325 7160
rect 12795 6985 18325 7040
rect 12795 6865 12820 6985
rect 12940 6865 12985 6985
rect 13105 6865 13150 6985
rect 13270 6865 13315 6985
rect 13435 6865 13490 6985
rect 13610 6865 13655 6985
rect 13775 6865 13820 6985
rect 13940 6865 13985 6985
rect 14105 6865 14160 6985
rect 14280 6865 14325 6985
rect 14445 6865 14490 6985
rect 14610 6865 14655 6985
rect 14775 6865 14830 6985
rect 14950 6865 14995 6985
rect 15115 6865 15160 6985
rect 15280 6865 15325 6985
rect 15445 6865 15500 6985
rect 15620 6865 15665 6985
rect 15785 6865 15830 6985
rect 15950 6865 15995 6985
rect 16115 6865 16170 6985
rect 16290 6865 16335 6985
rect 16455 6865 16500 6985
rect 16620 6865 16665 6985
rect 16785 6865 16840 6985
rect 16960 6865 17005 6985
rect 17125 6865 17170 6985
rect 17290 6865 17335 6985
rect 17455 6865 17510 6985
rect 17630 6865 17675 6985
rect 17795 6865 17840 6985
rect 17960 6865 18005 6985
rect 18125 6865 18180 6985
rect 18300 6865 18325 6985
rect 12795 6820 18325 6865
rect 12795 6700 12820 6820
rect 12940 6700 12985 6820
rect 13105 6700 13150 6820
rect 13270 6700 13315 6820
rect 13435 6700 13490 6820
rect 13610 6700 13655 6820
rect 13775 6700 13820 6820
rect 13940 6700 13985 6820
rect 14105 6700 14160 6820
rect 14280 6700 14325 6820
rect 14445 6700 14490 6820
rect 14610 6700 14655 6820
rect 14775 6700 14830 6820
rect 14950 6700 14995 6820
rect 15115 6700 15160 6820
rect 15280 6700 15325 6820
rect 15445 6700 15500 6820
rect 15620 6700 15665 6820
rect 15785 6700 15830 6820
rect 15950 6700 15995 6820
rect 16115 6700 16170 6820
rect 16290 6700 16335 6820
rect 16455 6700 16500 6820
rect 16620 6700 16665 6820
rect 16785 6700 16840 6820
rect 16960 6700 17005 6820
rect 17125 6700 17170 6820
rect 17290 6700 17335 6820
rect 17455 6700 17510 6820
rect 17630 6700 17675 6820
rect 17795 6700 17840 6820
rect 17960 6700 18005 6820
rect 18125 6700 18180 6820
rect 18300 6700 18325 6820
rect 12795 6655 18325 6700
rect 12795 6535 12820 6655
rect 12940 6535 12985 6655
rect 13105 6535 13150 6655
rect 13270 6535 13315 6655
rect 13435 6535 13490 6655
rect 13610 6535 13655 6655
rect 13775 6535 13820 6655
rect 13940 6535 13985 6655
rect 14105 6535 14160 6655
rect 14280 6535 14325 6655
rect 14445 6535 14490 6655
rect 14610 6535 14655 6655
rect 14775 6535 14830 6655
rect 14950 6535 14995 6655
rect 15115 6535 15160 6655
rect 15280 6535 15325 6655
rect 15445 6535 15500 6655
rect 15620 6535 15665 6655
rect 15785 6535 15830 6655
rect 15950 6535 15995 6655
rect 16115 6535 16170 6655
rect 16290 6535 16335 6655
rect 16455 6535 16500 6655
rect 16620 6535 16665 6655
rect 16785 6535 16840 6655
rect 16960 6535 17005 6655
rect 17125 6535 17170 6655
rect 17290 6535 17335 6655
rect 17455 6535 17510 6655
rect 17630 6535 17675 6655
rect 17795 6535 17840 6655
rect 17960 6535 18005 6655
rect 18125 6535 18180 6655
rect 18300 6535 18325 6655
rect 12795 6490 18325 6535
rect 12795 6370 12820 6490
rect 12940 6370 12985 6490
rect 13105 6370 13150 6490
rect 13270 6370 13315 6490
rect 13435 6370 13490 6490
rect 13610 6370 13655 6490
rect 13775 6370 13820 6490
rect 13940 6370 13985 6490
rect 14105 6370 14160 6490
rect 14280 6370 14325 6490
rect 14445 6370 14490 6490
rect 14610 6370 14655 6490
rect 14775 6370 14830 6490
rect 14950 6370 14995 6490
rect 15115 6370 15160 6490
rect 15280 6370 15325 6490
rect 15445 6370 15500 6490
rect 15620 6370 15665 6490
rect 15785 6370 15830 6490
rect 15950 6370 15995 6490
rect 16115 6370 16170 6490
rect 16290 6370 16335 6490
rect 16455 6370 16500 6490
rect 16620 6370 16665 6490
rect 16785 6370 16840 6490
rect 16960 6370 17005 6490
rect 17125 6370 17170 6490
rect 17290 6370 17335 6490
rect 17455 6370 17510 6490
rect 17630 6370 17675 6490
rect 17795 6370 17840 6490
rect 17960 6370 18005 6490
rect 18125 6370 18180 6490
rect 18300 6370 18325 6490
rect 12795 6315 18325 6370
rect 12795 6195 12820 6315
rect 12940 6195 12985 6315
rect 13105 6195 13150 6315
rect 13270 6195 13315 6315
rect 13435 6195 13490 6315
rect 13610 6195 13655 6315
rect 13775 6195 13820 6315
rect 13940 6195 13985 6315
rect 14105 6195 14160 6315
rect 14280 6195 14325 6315
rect 14445 6195 14490 6315
rect 14610 6195 14655 6315
rect 14775 6195 14830 6315
rect 14950 6195 14995 6315
rect 15115 6195 15160 6315
rect 15280 6195 15325 6315
rect 15445 6195 15500 6315
rect 15620 6195 15665 6315
rect 15785 6195 15830 6315
rect 15950 6195 15995 6315
rect 16115 6195 16170 6315
rect 16290 6195 16335 6315
rect 16455 6195 16500 6315
rect 16620 6195 16665 6315
rect 16785 6195 16840 6315
rect 16960 6195 17005 6315
rect 17125 6195 17170 6315
rect 17290 6195 17335 6315
rect 17455 6195 17510 6315
rect 17630 6195 17675 6315
rect 17795 6195 17840 6315
rect 17960 6195 18005 6315
rect 18125 6195 18180 6315
rect 18300 6195 18325 6315
rect 12795 6150 18325 6195
rect 12795 6030 12820 6150
rect 12940 6030 12985 6150
rect 13105 6030 13150 6150
rect 13270 6030 13315 6150
rect 13435 6030 13490 6150
rect 13610 6030 13655 6150
rect 13775 6030 13820 6150
rect 13940 6030 13985 6150
rect 14105 6030 14160 6150
rect 14280 6030 14325 6150
rect 14445 6030 14490 6150
rect 14610 6030 14655 6150
rect 14775 6030 14830 6150
rect 14950 6030 14995 6150
rect 15115 6030 15160 6150
rect 15280 6030 15325 6150
rect 15445 6030 15500 6150
rect 15620 6030 15665 6150
rect 15785 6030 15830 6150
rect 15950 6030 15995 6150
rect 16115 6030 16170 6150
rect 16290 6030 16335 6150
rect 16455 6030 16500 6150
rect 16620 6030 16665 6150
rect 16785 6030 16840 6150
rect 16960 6030 17005 6150
rect 17125 6030 17170 6150
rect 17290 6030 17335 6150
rect 17455 6030 17510 6150
rect 17630 6030 17675 6150
rect 17795 6030 17840 6150
rect 17960 6030 18005 6150
rect 18125 6030 18180 6150
rect 18300 6030 18325 6150
rect 12795 5985 18325 6030
rect 12795 5865 12820 5985
rect 12940 5865 12985 5985
rect 13105 5865 13150 5985
rect 13270 5865 13315 5985
rect 13435 5865 13490 5985
rect 13610 5865 13655 5985
rect 13775 5865 13820 5985
rect 13940 5865 13985 5985
rect 14105 5865 14160 5985
rect 14280 5865 14325 5985
rect 14445 5865 14490 5985
rect 14610 5865 14655 5985
rect 14775 5865 14830 5985
rect 14950 5865 14995 5985
rect 15115 5865 15160 5985
rect 15280 5865 15325 5985
rect 15445 5865 15500 5985
rect 15620 5865 15665 5985
rect 15785 5865 15830 5985
rect 15950 5865 15995 5985
rect 16115 5865 16170 5985
rect 16290 5865 16335 5985
rect 16455 5865 16500 5985
rect 16620 5865 16665 5985
rect 16785 5865 16840 5985
rect 16960 5865 17005 5985
rect 17125 5865 17170 5985
rect 17290 5865 17335 5985
rect 17455 5865 17510 5985
rect 17630 5865 17675 5985
rect 17795 5865 17840 5985
rect 17960 5865 18005 5985
rect 18125 5865 18180 5985
rect 18300 5865 18325 5985
rect 12795 5820 18325 5865
rect 12795 5700 12820 5820
rect 12940 5700 12985 5820
rect 13105 5700 13150 5820
rect 13270 5700 13315 5820
rect 13435 5700 13490 5820
rect 13610 5700 13655 5820
rect 13775 5700 13820 5820
rect 13940 5700 13985 5820
rect 14105 5700 14160 5820
rect 14280 5700 14325 5820
rect 14445 5700 14490 5820
rect 14610 5700 14655 5820
rect 14775 5700 14830 5820
rect 14950 5700 14995 5820
rect 15115 5700 15160 5820
rect 15280 5700 15325 5820
rect 15445 5700 15500 5820
rect 15620 5700 15665 5820
rect 15785 5700 15830 5820
rect 15950 5700 15995 5820
rect 16115 5700 16170 5820
rect 16290 5700 16335 5820
rect 16455 5700 16500 5820
rect 16620 5700 16665 5820
rect 16785 5700 16840 5820
rect 16960 5700 17005 5820
rect 17125 5700 17170 5820
rect 17290 5700 17335 5820
rect 17455 5700 17510 5820
rect 17630 5700 17675 5820
rect 17795 5700 17840 5820
rect 17960 5700 18005 5820
rect 18125 5700 18180 5820
rect 18300 5700 18325 5820
rect 12795 5645 18325 5700
rect 12795 5525 12820 5645
rect 12940 5525 12985 5645
rect 13105 5525 13150 5645
rect 13270 5525 13315 5645
rect 13435 5525 13490 5645
rect 13610 5525 13655 5645
rect 13775 5525 13820 5645
rect 13940 5525 13985 5645
rect 14105 5525 14160 5645
rect 14280 5525 14325 5645
rect 14445 5525 14490 5645
rect 14610 5525 14655 5645
rect 14775 5525 14830 5645
rect 14950 5525 14995 5645
rect 15115 5525 15160 5645
rect 15280 5525 15325 5645
rect 15445 5525 15500 5645
rect 15620 5525 15665 5645
rect 15785 5525 15830 5645
rect 15950 5525 15995 5645
rect 16115 5525 16170 5645
rect 16290 5525 16335 5645
rect 16455 5525 16500 5645
rect 16620 5525 16665 5645
rect 16785 5525 16840 5645
rect 16960 5525 17005 5645
rect 17125 5525 17170 5645
rect 17290 5525 17335 5645
rect 17455 5525 17510 5645
rect 17630 5525 17675 5645
rect 17795 5525 17840 5645
rect 17960 5525 18005 5645
rect 18125 5525 18180 5645
rect 18300 5525 18325 5645
rect 12795 5480 18325 5525
rect 12795 5360 12820 5480
rect 12940 5360 12985 5480
rect 13105 5360 13150 5480
rect 13270 5360 13315 5480
rect 13435 5360 13490 5480
rect 13610 5360 13655 5480
rect 13775 5360 13820 5480
rect 13940 5360 13985 5480
rect 14105 5360 14160 5480
rect 14280 5360 14325 5480
rect 14445 5360 14490 5480
rect 14610 5360 14655 5480
rect 14775 5360 14830 5480
rect 14950 5360 14995 5480
rect 15115 5360 15160 5480
rect 15280 5360 15325 5480
rect 15445 5360 15500 5480
rect 15620 5360 15665 5480
rect 15785 5360 15830 5480
rect 15950 5360 15995 5480
rect 16115 5360 16170 5480
rect 16290 5360 16335 5480
rect 16455 5360 16500 5480
rect 16620 5360 16665 5480
rect 16785 5360 16840 5480
rect 16960 5360 17005 5480
rect 17125 5360 17170 5480
rect 17290 5360 17335 5480
rect 17455 5360 17510 5480
rect 17630 5360 17675 5480
rect 17795 5360 17840 5480
rect 17960 5360 18005 5480
rect 18125 5360 18180 5480
rect 18300 5360 18325 5480
rect 12795 5315 18325 5360
rect 12795 5195 12820 5315
rect 12940 5195 12985 5315
rect 13105 5195 13150 5315
rect 13270 5195 13315 5315
rect 13435 5195 13490 5315
rect 13610 5195 13655 5315
rect 13775 5195 13820 5315
rect 13940 5195 13985 5315
rect 14105 5195 14160 5315
rect 14280 5195 14325 5315
rect 14445 5195 14490 5315
rect 14610 5195 14655 5315
rect 14775 5195 14830 5315
rect 14950 5195 14995 5315
rect 15115 5195 15160 5315
rect 15280 5195 15325 5315
rect 15445 5195 15500 5315
rect 15620 5195 15665 5315
rect 15785 5195 15830 5315
rect 15950 5195 15995 5315
rect 16115 5195 16170 5315
rect 16290 5195 16335 5315
rect 16455 5195 16500 5315
rect 16620 5195 16665 5315
rect 16785 5195 16840 5315
rect 16960 5195 17005 5315
rect 17125 5195 17170 5315
rect 17290 5195 17335 5315
rect 17455 5195 17510 5315
rect 17630 5195 17675 5315
rect 17795 5195 17840 5315
rect 17960 5195 18005 5315
rect 18125 5195 18180 5315
rect 18300 5195 18325 5315
rect 12795 5150 18325 5195
rect 12795 5030 12820 5150
rect 12940 5030 12985 5150
rect 13105 5030 13150 5150
rect 13270 5030 13315 5150
rect 13435 5030 13490 5150
rect 13610 5030 13655 5150
rect 13775 5030 13820 5150
rect 13940 5030 13985 5150
rect 14105 5030 14160 5150
rect 14280 5030 14325 5150
rect 14445 5030 14490 5150
rect 14610 5030 14655 5150
rect 14775 5030 14830 5150
rect 14950 5030 14995 5150
rect 15115 5030 15160 5150
rect 15280 5030 15325 5150
rect 15445 5030 15500 5150
rect 15620 5030 15665 5150
rect 15785 5030 15830 5150
rect 15950 5030 15995 5150
rect 16115 5030 16170 5150
rect 16290 5030 16335 5150
rect 16455 5030 16500 5150
rect 16620 5030 16665 5150
rect 16785 5030 16840 5150
rect 16960 5030 17005 5150
rect 17125 5030 17170 5150
rect 17290 5030 17335 5150
rect 17455 5030 17510 5150
rect 17630 5030 17675 5150
rect 17795 5030 17840 5150
rect 17960 5030 18005 5150
rect 18125 5030 18180 5150
rect 18300 5030 18325 5150
rect 12795 4975 18325 5030
rect 12795 4855 12820 4975
rect 12940 4855 12985 4975
rect 13105 4855 13150 4975
rect 13270 4855 13315 4975
rect 13435 4855 13490 4975
rect 13610 4855 13655 4975
rect 13775 4855 13820 4975
rect 13940 4855 13985 4975
rect 14105 4855 14160 4975
rect 14280 4855 14325 4975
rect 14445 4855 14490 4975
rect 14610 4855 14655 4975
rect 14775 4855 14830 4975
rect 14950 4855 14995 4975
rect 15115 4855 15160 4975
rect 15280 4855 15325 4975
rect 15445 4855 15500 4975
rect 15620 4855 15665 4975
rect 15785 4855 15830 4975
rect 15950 4855 15995 4975
rect 16115 4855 16170 4975
rect 16290 4855 16335 4975
rect 16455 4855 16500 4975
rect 16620 4855 16665 4975
rect 16785 4855 16840 4975
rect 16960 4855 17005 4975
rect 17125 4855 17170 4975
rect 17290 4855 17335 4975
rect 17455 4855 17510 4975
rect 17630 4855 17675 4975
rect 17795 4855 17840 4975
rect 17960 4855 18005 4975
rect 18125 4855 18180 4975
rect 18300 4855 18325 4975
rect 12795 4810 18325 4855
rect 12795 4690 12820 4810
rect 12940 4690 12985 4810
rect 13105 4690 13150 4810
rect 13270 4690 13315 4810
rect 13435 4690 13490 4810
rect 13610 4690 13655 4810
rect 13775 4690 13820 4810
rect 13940 4690 13985 4810
rect 14105 4690 14160 4810
rect 14280 4690 14325 4810
rect 14445 4690 14490 4810
rect 14610 4690 14655 4810
rect 14775 4690 14830 4810
rect 14950 4690 14995 4810
rect 15115 4690 15160 4810
rect 15280 4690 15325 4810
rect 15445 4690 15500 4810
rect 15620 4690 15665 4810
rect 15785 4690 15830 4810
rect 15950 4690 15995 4810
rect 16115 4690 16170 4810
rect 16290 4690 16335 4810
rect 16455 4690 16500 4810
rect 16620 4690 16665 4810
rect 16785 4690 16840 4810
rect 16960 4690 17005 4810
rect 17125 4690 17170 4810
rect 17290 4690 17335 4810
rect 17455 4690 17510 4810
rect 17630 4690 17675 4810
rect 17795 4690 17840 4810
rect 17960 4690 18005 4810
rect 18125 4690 18180 4810
rect 18300 4690 18325 4810
rect 12795 4645 18325 4690
rect 12795 4525 12820 4645
rect 12940 4525 12985 4645
rect 13105 4525 13150 4645
rect 13270 4525 13315 4645
rect 13435 4525 13490 4645
rect 13610 4525 13655 4645
rect 13775 4525 13820 4645
rect 13940 4525 13985 4645
rect 14105 4525 14160 4645
rect 14280 4525 14325 4645
rect 14445 4525 14490 4645
rect 14610 4525 14655 4645
rect 14775 4525 14830 4645
rect 14950 4525 14995 4645
rect 15115 4525 15160 4645
rect 15280 4525 15325 4645
rect 15445 4525 15500 4645
rect 15620 4525 15665 4645
rect 15785 4525 15830 4645
rect 15950 4525 15995 4645
rect 16115 4525 16170 4645
rect 16290 4525 16335 4645
rect 16455 4525 16500 4645
rect 16620 4525 16665 4645
rect 16785 4525 16840 4645
rect 16960 4525 17005 4645
rect 17125 4525 17170 4645
rect 17290 4525 17335 4645
rect 17455 4525 17510 4645
rect 17630 4525 17675 4645
rect 17795 4525 17840 4645
rect 17960 4525 18005 4645
rect 18125 4525 18180 4645
rect 18300 4525 18325 4645
rect 12795 4480 18325 4525
rect 12795 4360 12820 4480
rect 12940 4360 12985 4480
rect 13105 4360 13150 4480
rect 13270 4360 13315 4480
rect 13435 4360 13490 4480
rect 13610 4360 13655 4480
rect 13775 4360 13820 4480
rect 13940 4360 13985 4480
rect 14105 4360 14160 4480
rect 14280 4360 14325 4480
rect 14445 4360 14490 4480
rect 14610 4360 14655 4480
rect 14775 4360 14830 4480
rect 14950 4360 14995 4480
rect 15115 4360 15160 4480
rect 15280 4360 15325 4480
rect 15445 4360 15500 4480
rect 15620 4360 15665 4480
rect 15785 4360 15830 4480
rect 15950 4360 15995 4480
rect 16115 4360 16170 4480
rect 16290 4360 16335 4480
rect 16455 4360 16500 4480
rect 16620 4360 16665 4480
rect 16785 4360 16840 4480
rect 16960 4360 17005 4480
rect 17125 4360 17170 4480
rect 17290 4360 17335 4480
rect 17455 4360 17510 4480
rect 17630 4360 17675 4480
rect 17795 4360 17840 4480
rect 17960 4360 18005 4480
rect 18125 4360 18180 4480
rect 18300 4360 18325 4480
rect 12795 4305 18325 4360
rect 12795 4185 12820 4305
rect 12940 4185 12985 4305
rect 13105 4185 13150 4305
rect 13270 4185 13315 4305
rect 13435 4185 13490 4305
rect 13610 4185 13655 4305
rect 13775 4185 13820 4305
rect 13940 4185 13985 4305
rect 14105 4185 14160 4305
rect 14280 4185 14325 4305
rect 14445 4185 14490 4305
rect 14610 4185 14655 4305
rect 14775 4185 14830 4305
rect 14950 4185 14995 4305
rect 15115 4185 15160 4305
rect 15280 4185 15325 4305
rect 15445 4185 15500 4305
rect 15620 4185 15665 4305
rect 15785 4185 15830 4305
rect 15950 4185 15995 4305
rect 16115 4185 16170 4305
rect 16290 4185 16335 4305
rect 16455 4185 16500 4305
rect 16620 4185 16665 4305
rect 16785 4185 16840 4305
rect 16960 4185 17005 4305
rect 17125 4185 17170 4305
rect 17290 4185 17335 4305
rect 17455 4185 17510 4305
rect 17630 4185 17675 4305
rect 17795 4185 17840 4305
rect 17960 4185 18005 4305
rect 18125 4185 18180 4305
rect 18300 4185 18325 4305
rect 12795 4140 18325 4185
rect 12795 4020 12820 4140
rect 12940 4020 12985 4140
rect 13105 4020 13150 4140
rect 13270 4020 13315 4140
rect 13435 4020 13490 4140
rect 13610 4020 13655 4140
rect 13775 4020 13820 4140
rect 13940 4020 13985 4140
rect 14105 4020 14160 4140
rect 14280 4020 14325 4140
rect 14445 4020 14490 4140
rect 14610 4020 14655 4140
rect 14775 4020 14830 4140
rect 14950 4020 14995 4140
rect 15115 4020 15160 4140
rect 15280 4020 15325 4140
rect 15445 4020 15500 4140
rect 15620 4020 15665 4140
rect 15785 4020 15830 4140
rect 15950 4020 15995 4140
rect 16115 4020 16170 4140
rect 16290 4020 16335 4140
rect 16455 4020 16500 4140
rect 16620 4020 16665 4140
rect 16785 4020 16840 4140
rect 16960 4020 17005 4140
rect 17125 4020 17170 4140
rect 17290 4020 17335 4140
rect 17455 4020 17510 4140
rect 17630 4020 17675 4140
rect 17795 4020 17840 4140
rect 17960 4020 18005 4140
rect 18125 4020 18180 4140
rect 18300 4020 18325 4140
rect 12795 3975 18325 4020
rect 12795 3855 12820 3975
rect 12940 3855 12985 3975
rect 13105 3855 13150 3975
rect 13270 3855 13315 3975
rect 13435 3855 13490 3975
rect 13610 3855 13655 3975
rect 13775 3855 13820 3975
rect 13940 3855 13985 3975
rect 14105 3855 14160 3975
rect 14280 3855 14325 3975
rect 14445 3855 14490 3975
rect 14610 3855 14655 3975
rect 14775 3855 14830 3975
rect 14950 3855 14995 3975
rect 15115 3855 15160 3975
rect 15280 3855 15325 3975
rect 15445 3855 15500 3975
rect 15620 3855 15665 3975
rect 15785 3855 15830 3975
rect 15950 3855 15995 3975
rect 16115 3855 16170 3975
rect 16290 3855 16335 3975
rect 16455 3855 16500 3975
rect 16620 3855 16665 3975
rect 16785 3855 16840 3975
rect 16960 3855 17005 3975
rect 17125 3855 17170 3975
rect 17290 3855 17335 3975
rect 17455 3855 17510 3975
rect 17630 3855 17675 3975
rect 17795 3855 17840 3975
rect 17960 3855 18005 3975
rect 18125 3855 18180 3975
rect 18300 3855 18325 3975
rect 12795 3810 18325 3855
rect 12795 3690 12820 3810
rect 12940 3690 12985 3810
rect 13105 3690 13150 3810
rect 13270 3690 13315 3810
rect 13435 3690 13490 3810
rect 13610 3690 13655 3810
rect 13775 3690 13820 3810
rect 13940 3690 13985 3810
rect 14105 3690 14160 3810
rect 14280 3690 14325 3810
rect 14445 3690 14490 3810
rect 14610 3690 14655 3810
rect 14775 3690 14830 3810
rect 14950 3690 14995 3810
rect 15115 3690 15160 3810
rect 15280 3690 15325 3810
rect 15445 3690 15500 3810
rect 15620 3690 15665 3810
rect 15785 3690 15830 3810
rect 15950 3690 15995 3810
rect 16115 3690 16170 3810
rect 16290 3690 16335 3810
rect 16455 3690 16500 3810
rect 16620 3690 16665 3810
rect 16785 3690 16840 3810
rect 16960 3690 17005 3810
rect 17125 3690 17170 3810
rect 17290 3690 17335 3810
rect 17455 3690 17510 3810
rect 17630 3690 17675 3810
rect 17795 3690 17840 3810
rect 17960 3690 18005 3810
rect 18125 3690 18180 3810
rect 18300 3690 18325 3810
rect 12795 3635 18325 3690
rect 12795 3515 12820 3635
rect 12940 3515 12985 3635
rect 13105 3515 13150 3635
rect 13270 3515 13315 3635
rect 13435 3515 13490 3635
rect 13610 3515 13655 3635
rect 13775 3515 13820 3635
rect 13940 3515 13985 3635
rect 14105 3515 14160 3635
rect 14280 3515 14325 3635
rect 14445 3515 14490 3635
rect 14610 3515 14655 3635
rect 14775 3515 14830 3635
rect 14950 3515 14995 3635
rect 15115 3515 15160 3635
rect 15280 3515 15325 3635
rect 15445 3515 15500 3635
rect 15620 3515 15665 3635
rect 15785 3515 15830 3635
rect 15950 3515 15995 3635
rect 16115 3515 16170 3635
rect 16290 3515 16335 3635
rect 16455 3515 16500 3635
rect 16620 3515 16665 3635
rect 16785 3515 16840 3635
rect 16960 3515 17005 3635
rect 17125 3515 17170 3635
rect 17290 3515 17335 3635
rect 17455 3515 17510 3635
rect 17630 3515 17675 3635
rect 17795 3515 17840 3635
rect 17960 3515 18005 3635
rect 18125 3515 18180 3635
rect 18300 3515 18325 3635
rect 12795 3470 18325 3515
rect 12795 3350 12820 3470
rect 12940 3350 12985 3470
rect 13105 3350 13150 3470
rect 13270 3350 13315 3470
rect 13435 3350 13490 3470
rect 13610 3350 13655 3470
rect 13775 3350 13820 3470
rect 13940 3350 13985 3470
rect 14105 3350 14160 3470
rect 14280 3350 14325 3470
rect 14445 3350 14490 3470
rect 14610 3350 14655 3470
rect 14775 3350 14830 3470
rect 14950 3350 14995 3470
rect 15115 3350 15160 3470
rect 15280 3350 15325 3470
rect 15445 3350 15500 3470
rect 15620 3350 15665 3470
rect 15785 3350 15830 3470
rect 15950 3350 15995 3470
rect 16115 3350 16170 3470
rect 16290 3350 16335 3470
rect 16455 3350 16500 3470
rect 16620 3350 16665 3470
rect 16785 3350 16840 3470
rect 16960 3350 17005 3470
rect 17125 3350 17170 3470
rect 17290 3350 17335 3470
rect 17455 3350 17510 3470
rect 17630 3350 17675 3470
rect 17795 3350 17840 3470
rect 17960 3350 18005 3470
rect 18125 3350 18180 3470
rect 18300 3350 18325 3470
rect 12795 3305 18325 3350
rect 12795 3185 12820 3305
rect 12940 3185 12985 3305
rect 13105 3185 13150 3305
rect 13270 3185 13315 3305
rect 13435 3185 13490 3305
rect 13610 3185 13655 3305
rect 13775 3185 13820 3305
rect 13940 3185 13985 3305
rect 14105 3185 14160 3305
rect 14280 3185 14325 3305
rect 14445 3185 14490 3305
rect 14610 3185 14655 3305
rect 14775 3185 14830 3305
rect 14950 3185 14995 3305
rect 15115 3185 15160 3305
rect 15280 3185 15325 3305
rect 15445 3185 15500 3305
rect 15620 3185 15665 3305
rect 15785 3185 15830 3305
rect 15950 3185 15995 3305
rect 16115 3185 16170 3305
rect 16290 3185 16335 3305
rect 16455 3185 16500 3305
rect 16620 3185 16665 3305
rect 16785 3185 16840 3305
rect 16960 3185 17005 3305
rect 17125 3185 17170 3305
rect 17290 3185 17335 3305
rect 17455 3185 17510 3305
rect 17630 3185 17675 3305
rect 17795 3185 17840 3305
rect 17960 3185 18005 3305
rect 18125 3185 18180 3305
rect 18300 3185 18325 3305
rect 12795 3140 18325 3185
rect 12795 3020 12820 3140
rect 12940 3020 12985 3140
rect 13105 3020 13150 3140
rect 13270 3020 13315 3140
rect 13435 3020 13490 3140
rect 13610 3020 13655 3140
rect 13775 3020 13820 3140
rect 13940 3020 13985 3140
rect 14105 3020 14160 3140
rect 14280 3020 14325 3140
rect 14445 3020 14490 3140
rect 14610 3020 14655 3140
rect 14775 3020 14830 3140
rect 14950 3020 14995 3140
rect 15115 3020 15160 3140
rect 15280 3020 15325 3140
rect 15445 3020 15500 3140
rect 15620 3020 15665 3140
rect 15785 3020 15830 3140
rect 15950 3020 15995 3140
rect 16115 3020 16170 3140
rect 16290 3020 16335 3140
rect 16455 3020 16500 3140
rect 16620 3020 16665 3140
rect 16785 3020 16840 3140
rect 16960 3020 17005 3140
rect 17125 3020 17170 3140
rect 17290 3020 17335 3140
rect 17455 3020 17510 3140
rect 17630 3020 17675 3140
rect 17795 3020 17840 3140
rect 17960 3020 18005 3140
rect 18125 3020 18180 3140
rect 18300 3020 18325 3140
rect 12795 2965 18325 3020
rect 12795 2845 12820 2965
rect 12940 2845 12985 2965
rect 13105 2845 13150 2965
rect 13270 2845 13315 2965
rect 13435 2845 13490 2965
rect 13610 2845 13655 2965
rect 13775 2845 13820 2965
rect 13940 2845 13985 2965
rect 14105 2845 14160 2965
rect 14280 2845 14325 2965
rect 14445 2845 14490 2965
rect 14610 2845 14655 2965
rect 14775 2845 14830 2965
rect 14950 2845 14995 2965
rect 15115 2845 15160 2965
rect 15280 2845 15325 2965
rect 15445 2845 15500 2965
rect 15620 2845 15665 2965
rect 15785 2845 15830 2965
rect 15950 2845 15995 2965
rect 16115 2845 16170 2965
rect 16290 2845 16335 2965
rect 16455 2845 16500 2965
rect 16620 2845 16665 2965
rect 16785 2845 16840 2965
rect 16960 2845 17005 2965
rect 17125 2845 17170 2965
rect 17290 2845 17335 2965
rect 17455 2845 17510 2965
rect 17630 2845 17675 2965
rect 17795 2845 17840 2965
rect 17960 2845 18005 2965
rect 18125 2845 18180 2965
rect 18300 2845 18325 2965
rect 12795 2800 18325 2845
rect 12795 2680 12820 2800
rect 12940 2680 12985 2800
rect 13105 2680 13150 2800
rect 13270 2680 13315 2800
rect 13435 2680 13490 2800
rect 13610 2680 13655 2800
rect 13775 2680 13820 2800
rect 13940 2680 13985 2800
rect 14105 2680 14160 2800
rect 14280 2680 14325 2800
rect 14445 2680 14490 2800
rect 14610 2680 14655 2800
rect 14775 2680 14830 2800
rect 14950 2680 14995 2800
rect 15115 2680 15160 2800
rect 15280 2680 15325 2800
rect 15445 2680 15500 2800
rect 15620 2680 15665 2800
rect 15785 2680 15830 2800
rect 15950 2680 15995 2800
rect 16115 2680 16170 2800
rect 16290 2680 16335 2800
rect 16455 2680 16500 2800
rect 16620 2680 16665 2800
rect 16785 2680 16840 2800
rect 16960 2680 17005 2800
rect 17125 2680 17170 2800
rect 17290 2680 17335 2800
rect 17455 2680 17510 2800
rect 17630 2680 17675 2800
rect 17795 2680 17840 2800
rect 17960 2680 18005 2800
rect 18125 2680 18180 2800
rect 18300 2680 18325 2800
rect 12795 2635 18325 2680
rect 12795 2515 12820 2635
rect 12940 2515 12985 2635
rect 13105 2515 13150 2635
rect 13270 2515 13315 2635
rect 13435 2515 13490 2635
rect 13610 2515 13655 2635
rect 13775 2515 13820 2635
rect 13940 2515 13985 2635
rect 14105 2515 14160 2635
rect 14280 2515 14325 2635
rect 14445 2515 14490 2635
rect 14610 2515 14655 2635
rect 14775 2515 14830 2635
rect 14950 2515 14995 2635
rect 15115 2515 15160 2635
rect 15280 2515 15325 2635
rect 15445 2515 15500 2635
rect 15620 2515 15665 2635
rect 15785 2515 15830 2635
rect 15950 2515 15995 2635
rect 16115 2515 16170 2635
rect 16290 2515 16335 2635
rect 16455 2515 16500 2635
rect 16620 2515 16665 2635
rect 16785 2515 16840 2635
rect 16960 2515 17005 2635
rect 17125 2515 17170 2635
rect 17290 2515 17335 2635
rect 17455 2515 17510 2635
rect 17630 2515 17675 2635
rect 17795 2515 17840 2635
rect 17960 2515 18005 2635
rect 18125 2515 18180 2635
rect 18300 2515 18325 2635
rect 12795 2470 18325 2515
rect 12795 2350 12820 2470
rect 12940 2350 12985 2470
rect 13105 2350 13150 2470
rect 13270 2350 13315 2470
rect 13435 2350 13490 2470
rect 13610 2350 13655 2470
rect 13775 2350 13820 2470
rect 13940 2350 13985 2470
rect 14105 2350 14160 2470
rect 14280 2350 14325 2470
rect 14445 2350 14490 2470
rect 14610 2350 14655 2470
rect 14775 2350 14830 2470
rect 14950 2350 14995 2470
rect 15115 2350 15160 2470
rect 15280 2350 15325 2470
rect 15445 2350 15500 2470
rect 15620 2350 15665 2470
rect 15785 2350 15830 2470
rect 15950 2350 15995 2470
rect 16115 2350 16170 2470
rect 16290 2350 16335 2470
rect 16455 2350 16500 2470
rect 16620 2350 16665 2470
rect 16785 2350 16840 2470
rect 16960 2350 17005 2470
rect 17125 2350 17170 2470
rect 17290 2350 17335 2470
rect 17455 2350 17510 2470
rect 17630 2350 17675 2470
rect 17795 2350 17840 2470
rect 17960 2350 18005 2470
rect 18125 2350 18180 2470
rect 18300 2350 18325 2470
rect 12795 2295 18325 2350
rect 12795 2175 12820 2295
rect 12940 2175 12985 2295
rect 13105 2175 13150 2295
rect 13270 2175 13315 2295
rect 13435 2175 13490 2295
rect 13610 2175 13655 2295
rect 13775 2175 13820 2295
rect 13940 2175 13985 2295
rect 14105 2175 14160 2295
rect 14280 2175 14325 2295
rect 14445 2175 14490 2295
rect 14610 2175 14655 2295
rect 14775 2175 14830 2295
rect 14950 2175 14995 2295
rect 15115 2175 15160 2295
rect 15280 2175 15325 2295
rect 15445 2175 15500 2295
rect 15620 2175 15665 2295
rect 15785 2175 15830 2295
rect 15950 2175 15995 2295
rect 16115 2175 16170 2295
rect 16290 2175 16335 2295
rect 16455 2175 16500 2295
rect 16620 2175 16665 2295
rect 16785 2175 16840 2295
rect 16960 2175 17005 2295
rect 17125 2175 17170 2295
rect 17290 2175 17335 2295
rect 17455 2175 17510 2295
rect 17630 2175 17675 2295
rect 17795 2175 17840 2295
rect 17960 2175 18005 2295
rect 18125 2175 18180 2295
rect 18300 2175 18325 2295
rect 12795 2130 18325 2175
rect 12795 2010 12820 2130
rect 12940 2010 12985 2130
rect 13105 2010 13150 2130
rect 13270 2010 13315 2130
rect 13435 2010 13490 2130
rect 13610 2010 13655 2130
rect 13775 2010 13820 2130
rect 13940 2010 13985 2130
rect 14105 2010 14160 2130
rect 14280 2010 14325 2130
rect 14445 2010 14490 2130
rect 14610 2010 14655 2130
rect 14775 2010 14830 2130
rect 14950 2010 14995 2130
rect 15115 2010 15160 2130
rect 15280 2010 15325 2130
rect 15445 2010 15500 2130
rect 15620 2010 15665 2130
rect 15785 2010 15830 2130
rect 15950 2010 15995 2130
rect 16115 2010 16170 2130
rect 16290 2010 16335 2130
rect 16455 2010 16500 2130
rect 16620 2010 16665 2130
rect 16785 2010 16840 2130
rect 16960 2010 17005 2130
rect 17125 2010 17170 2130
rect 17290 2010 17335 2130
rect 17455 2010 17510 2130
rect 17630 2010 17675 2130
rect 17795 2010 17840 2130
rect 17960 2010 18005 2130
rect 18125 2010 18180 2130
rect 18300 2010 18325 2130
rect 12795 1965 18325 2010
rect 12795 1845 12820 1965
rect 12940 1845 12985 1965
rect 13105 1845 13150 1965
rect 13270 1845 13315 1965
rect 13435 1845 13490 1965
rect 13610 1845 13655 1965
rect 13775 1845 13820 1965
rect 13940 1845 13985 1965
rect 14105 1845 14160 1965
rect 14280 1845 14325 1965
rect 14445 1845 14490 1965
rect 14610 1845 14655 1965
rect 14775 1845 14830 1965
rect 14950 1845 14995 1965
rect 15115 1845 15160 1965
rect 15280 1845 15325 1965
rect 15445 1845 15500 1965
rect 15620 1845 15665 1965
rect 15785 1845 15830 1965
rect 15950 1845 15995 1965
rect 16115 1845 16170 1965
rect 16290 1845 16335 1965
rect 16455 1845 16500 1965
rect 16620 1845 16665 1965
rect 16785 1845 16840 1965
rect 16960 1845 17005 1965
rect 17125 1845 17170 1965
rect 17290 1845 17335 1965
rect 17455 1845 17510 1965
rect 17630 1845 17675 1965
rect 17795 1845 17840 1965
rect 17960 1845 18005 1965
rect 18125 1845 18180 1965
rect 18300 1845 18325 1965
rect 12795 1800 18325 1845
rect 12795 1680 12820 1800
rect 12940 1680 12985 1800
rect 13105 1680 13150 1800
rect 13270 1680 13315 1800
rect 13435 1680 13490 1800
rect 13610 1680 13655 1800
rect 13775 1680 13820 1800
rect 13940 1680 13985 1800
rect 14105 1680 14160 1800
rect 14280 1680 14325 1800
rect 14445 1680 14490 1800
rect 14610 1680 14655 1800
rect 14775 1680 14830 1800
rect 14950 1680 14995 1800
rect 15115 1680 15160 1800
rect 15280 1680 15325 1800
rect 15445 1680 15500 1800
rect 15620 1680 15665 1800
rect 15785 1680 15830 1800
rect 15950 1680 15995 1800
rect 16115 1680 16170 1800
rect 16290 1680 16335 1800
rect 16455 1680 16500 1800
rect 16620 1680 16665 1800
rect 16785 1680 16840 1800
rect 16960 1680 17005 1800
rect 17125 1680 17170 1800
rect 17290 1680 17335 1800
rect 17455 1680 17510 1800
rect 17630 1680 17675 1800
rect 17795 1680 17840 1800
rect 17960 1680 18005 1800
rect 18125 1680 18180 1800
rect 18300 1680 18325 1800
rect 12795 1610 18325 1680
rect 18485 7160 24015 7185
rect 18485 7040 18510 7160
rect 18630 7040 18675 7160
rect 18795 7040 18840 7160
rect 18960 7040 19005 7160
rect 19125 7040 19180 7160
rect 19300 7040 19345 7160
rect 19465 7040 19510 7160
rect 19630 7040 19675 7160
rect 19795 7040 19850 7160
rect 19970 7040 20015 7160
rect 20135 7040 20180 7160
rect 20300 7040 20345 7160
rect 20465 7040 20520 7160
rect 20640 7040 20685 7160
rect 20805 7040 20850 7160
rect 20970 7040 21015 7160
rect 21135 7040 21190 7160
rect 21310 7040 21355 7160
rect 21475 7040 21520 7160
rect 21640 7040 21685 7160
rect 21805 7040 21860 7160
rect 21980 7040 22025 7160
rect 22145 7040 22190 7160
rect 22310 7040 22355 7160
rect 22475 7040 22530 7160
rect 22650 7040 22695 7160
rect 22815 7040 22860 7160
rect 22980 7040 23025 7160
rect 23145 7040 23200 7160
rect 23320 7040 23365 7160
rect 23485 7040 23530 7160
rect 23650 7040 23695 7160
rect 23815 7040 23870 7160
rect 23990 7040 24015 7160
rect 18485 6985 24015 7040
rect 18485 6865 18510 6985
rect 18630 6865 18675 6985
rect 18795 6865 18840 6985
rect 18960 6865 19005 6985
rect 19125 6865 19180 6985
rect 19300 6865 19345 6985
rect 19465 6865 19510 6985
rect 19630 6865 19675 6985
rect 19795 6865 19850 6985
rect 19970 6865 20015 6985
rect 20135 6865 20180 6985
rect 20300 6865 20345 6985
rect 20465 6865 20520 6985
rect 20640 6865 20685 6985
rect 20805 6865 20850 6985
rect 20970 6865 21015 6985
rect 21135 6865 21190 6985
rect 21310 6865 21355 6985
rect 21475 6865 21520 6985
rect 21640 6865 21685 6985
rect 21805 6865 21860 6985
rect 21980 6865 22025 6985
rect 22145 6865 22190 6985
rect 22310 6865 22355 6985
rect 22475 6865 22530 6985
rect 22650 6865 22695 6985
rect 22815 6865 22860 6985
rect 22980 6865 23025 6985
rect 23145 6865 23200 6985
rect 23320 6865 23365 6985
rect 23485 6865 23530 6985
rect 23650 6865 23695 6985
rect 23815 6865 23870 6985
rect 23990 6865 24015 6985
rect 18485 6820 24015 6865
rect 18485 6700 18510 6820
rect 18630 6700 18675 6820
rect 18795 6700 18840 6820
rect 18960 6700 19005 6820
rect 19125 6700 19180 6820
rect 19300 6700 19345 6820
rect 19465 6700 19510 6820
rect 19630 6700 19675 6820
rect 19795 6700 19850 6820
rect 19970 6700 20015 6820
rect 20135 6700 20180 6820
rect 20300 6700 20345 6820
rect 20465 6700 20520 6820
rect 20640 6700 20685 6820
rect 20805 6700 20850 6820
rect 20970 6700 21015 6820
rect 21135 6700 21190 6820
rect 21310 6700 21355 6820
rect 21475 6700 21520 6820
rect 21640 6700 21685 6820
rect 21805 6700 21860 6820
rect 21980 6700 22025 6820
rect 22145 6700 22190 6820
rect 22310 6700 22355 6820
rect 22475 6700 22530 6820
rect 22650 6700 22695 6820
rect 22815 6700 22860 6820
rect 22980 6700 23025 6820
rect 23145 6700 23200 6820
rect 23320 6700 23365 6820
rect 23485 6700 23530 6820
rect 23650 6700 23695 6820
rect 23815 6700 23870 6820
rect 23990 6700 24015 6820
rect 18485 6655 24015 6700
rect 18485 6535 18510 6655
rect 18630 6535 18675 6655
rect 18795 6535 18840 6655
rect 18960 6535 19005 6655
rect 19125 6535 19180 6655
rect 19300 6535 19345 6655
rect 19465 6535 19510 6655
rect 19630 6535 19675 6655
rect 19795 6535 19850 6655
rect 19970 6535 20015 6655
rect 20135 6535 20180 6655
rect 20300 6535 20345 6655
rect 20465 6535 20520 6655
rect 20640 6535 20685 6655
rect 20805 6535 20850 6655
rect 20970 6535 21015 6655
rect 21135 6535 21190 6655
rect 21310 6535 21355 6655
rect 21475 6535 21520 6655
rect 21640 6535 21685 6655
rect 21805 6535 21860 6655
rect 21980 6535 22025 6655
rect 22145 6535 22190 6655
rect 22310 6535 22355 6655
rect 22475 6535 22530 6655
rect 22650 6535 22695 6655
rect 22815 6535 22860 6655
rect 22980 6535 23025 6655
rect 23145 6535 23200 6655
rect 23320 6535 23365 6655
rect 23485 6535 23530 6655
rect 23650 6535 23695 6655
rect 23815 6535 23870 6655
rect 23990 6535 24015 6655
rect 18485 6490 24015 6535
rect 18485 6370 18510 6490
rect 18630 6370 18675 6490
rect 18795 6370 18840 6490
rect 18960 6370 19005 6490
rect 19125 6370 19180 6490
rect 19300 6370 19345 6490
rect 19465 6370 19510 6490
rect 19630 6370 19675 6490
rect 19795 6370 19850 6490
rect 19970 6370 20015 6490
rect 20135 6370 20180 6490
rect 20300 6370 20345 6490
rect 20465 6370 20520 6490
rect 20640 6370 20685 6490
rect 20805 6370 20850 6490
rect 20970 6370 21015 6490
rect 21135 6370 21190 6490
rect 21310 6370 21355 6490
rect 21475 6370 21520 6490
rect 21640 6370 21685 6490
rect 21805 6370 21860 6490
rect 21980 6370 22025 6490
rect 22145 6370 22190 6490
rect 22310 6370 22355 6490
rect 22475 6370 22530 6490
rect 22650 6370 22695 6490
rect 22815 6370 22860 6490
rect 22980 6370 23025 6490
rect 23145 6370 23200 6490
rect 23320 6370 23365 6490
rect 23485 6370 23530 6490
rect 23650 6370 23695 6490
rect 23815 6370 23870 6490
rect 23990 6370 24015 6490
rect 18485 6315 24015 6370
rect 18485 6195 18510 6315
rect 18630 6195 18675 6315
rect 18795 6195 18840 6315
rect 18960 6195 19005 6315
rect 19125 6195 19180 6315
rect 19300 6195 19345 6315
rect 19465 6195 19510 6315
rect 19630 6195 19675 6315
rect 19795 6195 19850 6315
rect 19970 6195 20015 6315
rect 20135 6195 20180 6315
rect 20300 6195 20345 6315
rect 20465 6195 20520 6315
rect 20640 6195 20685 6315
rect 20805 6195 20850 6315
rect 20970 6195 21015 6315
rect 21135 6195 21190 6315
rect 21310 6195 21355 6315
rect 21475 6195 21520 6315
rect 21640 6195 21685 6315
rect 21805 6195 21860 6315
rect 21980 6195 22025 6315
rect 22145 6195 22190 6315
rect 22310 6195 22355 6315
rect 22475 6195 22530 6315
rect 22650 6195 22695 6315
rect 22815 6195 22860 6315
rect 22980 6195 23025 6315
rect 23145 6195 23200 6315
rect 23320 6195 23365 6315
rect 23485 6195 23530 6315
rect 23650 6195 23695 6315
rect 23815 6195 23870 6315
rect 23990 6195 24015 6315
rect 18485 6150 24015 6195
rect 18485 6030 18510 6150
rect 18630 6030 18675 6150
rect 18795 6030 18840 6150
rect 18960 6030 19005 6150
rect 19125 6030 19180 6150
rect 19300 6030 19345 6150
rect 19465 6030 19510 6150
rect 19630 6030 19675 6150
rect 19795 6030 19850 6150
rect 19970 6030 20015 6150
rect 20135 6030 20180 6150
rect 20300 6030 20345 6150
rect 20465 6030 20520 6150
rect 20640 6030 20685 6150
rect 20805 6030 20850 6150
rect 20970 6030 21015 6150
rect 21135 6030 21190 6150
rect 21310 6030 21355 6150
rect 21475 6030 21520 6150
rect 21640 6030 21685 6150
rect 21805 6030 21860 6150
rect 21980 6030 22025 6150
rect 22145 6030 22190 6150
rect 22310 6030 22355 6150
rect 22475 6030 22530 6150
rect 22650 6030 22695 6150
rect 22815 6030 22860 6150
rect 22980 6030 23025 6150
rect 23145 6030 23200 6150
rect 23320 6030 23365 6150
rect 23485 6030 23530 6150
rect 23650 6030 23695 6150
rect 23815 6030 23870 6150
rect 23990 6030 24015 6150
rect 18485 5985 24015 6030
rect 18485 5865 18510 5985
rect 18630 5865 18675 5985
rect 18795 5865 18840 5985
rect 18960 5865 19005 5985
rect 19125 5865 19180 5985
rect 19300 5865 19345 5985
rect 19465 5865 19510 5985
rect 19630 5865 19675 5985
rect 19795 5865 19850 5985
rect 19970 5865 20015 5985
rect 20135 5865 20180 5985
rect 20300 5865 20345 5985
rect 20465 5865 20520 5985
rect 20640 5865 20685 5985
rect 20805 5865 20850 5985
rect 20970 5865 21015 5985
rect 21135 5865 21190 5985
rect 21310 5865 21355 5985
rect 21475 5865 21520 5985
rect 21640 5865 21685 5985
rect 21805 5865 21860 5985
rect 21980 5865 22025 5985
rect 22145 5865 22190 5985
rect 22310 5865 22355 5985
rect 22475 5865 22530 5985
rect 22650 5865 22695 5985
rect 22815 5865 22860 5985
rect 22980 5865 23025 5985
rect 23145 5865 23200 5985
rect 23320 5865 23365 5985
rect 23485 5865 23530 5985
rect 23650 5865 23695 5985
rect 23815 5865 23870 5985
rect 23990 5865 24015 5985
rect 18485 5820 24015 5865
rect 18485 5700 18510 5820
rect 18630 5700 18675 5820
rect 18795 5700 18840 5820
rect 18960 5700 19005 5820
rect 19125 5700 19180 5820
rect 19300 5700 19345 5820
rect 19465 5700 19510 5820
rect 19630 5700 19675 5820
rect 19795 5700 19850 5820
rect 19970 5700 20015 5820
rect 20135 5700 20180 5820
rect 20300 5700 20345 5820
rect 20465 5700 20520 5820
rect 20640 5700 20685 5820
rect 20805 5700 20850 5820
rect 20970 5700 21015 5820
rect 21135 5700 21190 5820
rect 21310 5700 21355 5820
rect 21475 5700 21520 5820
rect 21640 5700 21685 5820
rect 21805 5700 21860 5820
rect 21980 5700 22025 5820
rect 22145 5700 22190 5820
rect 22310 5700 22355 5820
rect 22475 5700 22530 5820
rect 22650 5700 22695 5820
rect 22815 5700 22860 5820
rect 22980 5700 23025 5820
rect 23145 5700 23200 5820
rect 23320 5700 23365 5820
rect 23485 5700 23530 5820
rect 23650 5700 23695 5820
rect 23815 5700 23870 5820
rect 23990 5700 24015 5820
rect 18485 5645 24015 5700
rect 18485 5525 18510 5645
rect 18630 5525 18675 5645
rect 18795 5525 18840 5645
rect 18960 5525 19005 5645
rect 19125 5525 19180 5645
rect 19300 5525 19345 5645
rect 19465 5525 19510 5645
rect 19630 5525 19675 5645
rect 19795 5525 19850 5645
rect 19970 5525 20015 5645
rect 20135 5525 20180 5645
rect 20300 5525 20345 5645
rect 20465 5525 20520 5645
rect 20640 5525 20685 5645
rect 20805 5525 20850 5645
rect 20970 5525 21015 5645
rect 21135 5525 21190 5645
rect 21310 5525 21355 5645
rect 21475 5525 21520 5645
rect 21640 5525 21685 5645
rect 21805 5525 21860 5645
rect 21980 5525 22025 5645
rect 22145 5525 22190 5645
rect 22310 5525 22355 5645
rect 22475 5525 22530 5645
rect 22650 5525 22695 5645
rect 22815 5525 22860 5645
rect 22980 5525 23025 5645
rect 23145 5525 23200 5645
rect 23320 5525 23365 5645
rect 23485 5525 23530 5645
rect 23650 5525 23695 5645
rect 23815 5525 23870 5645
rect 23990 5525 24015 5645
rect 18485 5480 24015 5525
rect 18485 5360 18510 5480
rect 18630 5360 18675 5480
rect 18795 5360 18840 5480
rect 18960 5360 19005 5480
rect 19125 5360 19180 5480
rect 19300 5360 19345 5480
rect 19465 5360 19510 5480
rect 19630 5360 19675 5480
rect 19795 5360 19850 5480
rect 19970 5360 20015 5480
rect 20135 5360 20180 5480
rect 20300 5360 20345 5480
rect 20465 5360 20520 5480
rect 20640 5360 20685 5480
rect 20805 5360 20850 5480
rect 20970 5360 21015 5480
rect 21135 5360 21190 5480
rect 21310 5360 21355 5480
rect 21475 5360 21520 5480
rect 21640 5360 21685 5480
rect 21805 5360 21860 5480
rect 21980 5360 22025 5480
rect 22145 5360 22190 5480
rect 22310 5360 22355 5480
rect 22475 5360 22530 5480
rect 22650 5360 22695 5480
rect 22815 5360 22860 5480
rect 22980 5360 23025 5480
rect 23145 5360 23200 5480
rect 23320 5360 23365 5480
rect 23485 5360 23530 5480
rect 23650 5360 23695 5480
rect 23815 5360 23870 5480
rect 23990 5360 24015 5480
rect 18485 5315 24015 5360
rect 18485 5195 18510 5315
rect 18630 5195 18675 5315
rect 18795 5195 18840 5315
rect 18960 5195 19005 5315
rect 19125 5195 19180 5315
rect 19300 5195 19345 5315
rect 19465 5195 19510 5315
rect 19630 5195 19675 5315
rect 19795 5195 19850 5315
rect 19970 5195 20015 5315
rect 20135 5195 20180 5315
rect 20300 5195 20345 5315
rect 20465 5195 20520 5315
rect 20640 5195 20685 5315
rect 20805 5195 20850 5315
rect 20970 5195 21015 5315
rect 21135 5195 21190 5315
rect 21310 5195 21355 5315
rect 21475 5195 21520 5315
rect 21640 5195 21685 5315
rect 21805 5195 21860 5315
rect 21980 5195 22025 5315
rect 22145 5195 22190 5315
rect 22310 5195 22355 5315
rect 22475 5195 22530 5315
rect 22650 5195 22695 5315
rect 22815 5195 22860 5315
rect 22980 5195 23025 5315
rect 23145 5195 23200 5315
rect 23320 5195 23365 5315
rect 23485 5195 23530 5315
rect 23650 5195 23695 5315
rect 23815 5195 23870 5315
rect 23990 5195 24015 5315
rect 18485 5150 24015 5195
rect 18485 5030 18510 5150
rect 18630 5030 18675 5150
rect 18795 5030 18840 5150
rect 18960 5030 19005 5150
rect 19125 5030 19180 5150
rect 19300 5030 19345 5150
rect 19465 5030 19510 5150
rect 19630 5030 19675 5150
rect 19795 5030 19850 5150
rect 19970 5030 20015 5150
rect 20135 5030 20180 5150
rect 20300 5030 20345 5150
rect 20465 5030 20520 5150
rect 20640 5030 20685 5150
rect 20805 5030 20850 5150
rect 20970 5030 21015 5150
rect 21135 5030 21190 5150
rect 21310 5030 21355 5150
rect 21475 5030 21520 5150
rect 21640 5030 21685 5150
rect 21805 5030 21860 5150
rect 21980 5030 22025 5150
rect 22145 5030 22190 5150
rect 22310 5030 22355 5150
rect 22475 5030 22530 5150
rect 22650 5030 22695 5150
rect 22815 5030 22860 5150
rect 22980 5030 23025 5150
rect 23145 5030 23200 5150
rect 23320 5030 23365 5150
rect 23485 5030 23530 5150
rect 23650 5030 23695 5150
rect 23815 5030 23870 5150
rect 23990 5030 24015 5150
rect 18485 4975 24015 5030
rect 18485 4855 18510 4975
rect 18630 4855 18675 4975
rect 18795 4855 18840 4975
rect 18960 4855 19005 4975
rect 19125 4855 19180 4975
rect 19300 4855 19345 4975
rect 19465 4855 19510 4975
rect 19630 4855 19675 4975
rect 19795 4855 19850 4975
rect 19970 4855 20015 4975
rect 20135 4855 20180 4975
rect 20300 4855 20345 4975
rect 20465 4855 20520 4975
rect 20640 4855 20685 4975
rect 20805 4855 20850 4975
rect 20970 4855 21015 4975
rect 21135 4855 21190 4975
rect 21310 4855 21355 4975
rect 21475 4855 21520 4975
rect 21640 4855 21685 4975
rect 21805 4855 21860 4975
rect 21980 4855 22025 4975
rect 22145 4855 22190 4975
rect 22310 4855 22355 4975
rect 22475 4855 22530 4975
rect 22650 4855 22695 4975
rect 22815 4855 22860 4975
rect 22980 4855 23025 4975
rect 23145 4855 23200 4975
rect 23320 4855 23365 4975
rect 23485 4855 23530 4975
rect 23650 4855 23695 4975
rect 23815 4855 23870 4975
rect 23990 4855 24015 4975
rect 18485 4810 24015 4855
rect 18485 4690 18510 4810
rect 18630 4690 18675 4810
rect 18795 4690 18840 4810
rect 18960 4690 19005 4810
rect 19125 4690 19180 4810
rect 19300 4690 19345 4810
rect 19465 4690 19510 4810
rect 19630 4690 19675 4810
rect 19795 4690 19850 4810
rect 19970 4690 20015 4810
rect 20135 4690 20180 4810
rect 20300 4690 20345 4810
rect 20465 4690 20520 4810
rect 20640 4690 20685 4810
rect 20805 4690 20850 4810
rect 20970 4690 21015 4810
rect 21135 4690 21190 4810
rect 21310 4690 21355 4810
rect 21475 4690 21520 4810
rect 21640 4690 21685 4810
rect 21805 4690 21860 4810
rect 21980 4690 22025 4810
rect 22145 4690 22190 4810
rect 22310 4690 22355 4810
rect 22475 4690 22530 4810
rect 22650 4690 22695 4810
rect 22815 4690 22860 4810
rect 22980 4690 23025 4810
rect 23145 4690 23200 4810
rect 23320 4690 23365 4810
rect 23485 4690 23530 4810
rect 23650 4690 23695 4810
rect 23815 4690 23870 4810
rect 23990 4690 24015 4810
rect 18485 4645 24015 4690
rect 18485 4525 18510 4645
rect 18630 4525 18675 4645
rect 18795 4525 18840 4645
rect 18960 4525 19005 4645
rect 19125 4525 19180 4645
rect 19300 4525 19345 4645
rect 19465 4525 19510 4645
rect 19630 4525 19675 4645
rect 19795 4525 19850 4645
rect 19970 4525 20015 4645
rect 20135 4525 20180 4645
rect 20300 4525 20345 4645
rect 20465 4525 20520 4645
rect 20640 4525 20685 4645
rect 20805 4525 20850 4645
rect 20970 4525 21015 4645
rect 21135 4525 21190 4645
rect 21310 4525 21355 4645
rect 21475 4525 21520 4645
rect 21640 4525 21685 4645
rect 21805 4525 21860 4645
rect 21980 4525 22025 4645
rect 22145 4525 22190 4645
rect 22310 4525 22355 4645
rect 22475 4525 22530 4645
rect 22650 4525 22695 4645
rect 22815 4525 22860 4645
rect 22980 4525 23025 4645
rect 23145 4525 23200 4645
rect 23320 4525 23365 4645
rect 23485 4525 23530 4645
rect 23650 4525 23695 4645
rect 23815 4525 23870 4645
rect 23990 4525 24015 4645
rect 18485 4480 24015 4525
rect 18485 4360 18510 4480
rect 18630 4360 18675 4480
rect 18795 4360 18840 4480
rect 18960 4360 19005 4480
rect 19125 4360 19180 4480
rect 19300 4360 19345 4480
rect 19465 4360 19510 4480
rect 19630 4360 19675 4480
rect 19795 4360 19850 4480
rect 19970 4360 20015 4480
rect 20135 4360 20180 4480
rect 20300 4360 20345 4480
rect 20465 4360 20520 4480
rect 20640 4360 20685 4480
rect 20805 4360 20850 4480
rect 20970 4360 21015 4480
rect 21135 4360 21190 4480
rect 21310 4360 21355 4480
rect 21475 4360 21520 4480
rect 21640 4360 21685 4480
rect 21805 4360 21860 4480
rect 21980 4360 22025 4480
rect 22145 4360 22190 4480
rect 22310 4360 22355 4480
rect 22475 4360 22530 4480
rect 22650 4360 22695 4480
rect 22815 4360 22860 4480
rect 22980 4360 23025 4480
rect 23145 4360 23200 4480
rect 23320 4360 23365 4480
rect 23485 4360 23530 4480
rect 23650 4360 23695 4480
rect 23815 4360 23870 4480
rect 23990 4360 24015 4480
rect 18485 4305 24015 4360
rect 18485 4185 18510 4305
rect 18630 4185 18675 4305
rect 18795 4185 18840 4305
rect 18960 4185 19005 4305
rect 19125 4185 19180 4305
rect 19300 4185 19345 4305
rect 19465 4185 19510 4305
rect 19630 4185 19675 4305
rect 19795 4185 19850 4305
rect 19970 4185 20015 4305
rect 20135 4185 20180 4305
rect 20300 4185 20345 4305
rect 20465 4185 20520 4305
rect 20640 4185 20685 4305
rect 20805 4185 20850 4305
rect 20970 4185 21015 4305
rect 21135 4185 21190 4305
rect 21310 4185 21355 4305
rect 21475 4185 21520 4305
rect 21640 4185 21685 4305
rect 21805 4185 21860 4305
rect 21980 4185 22025 4305
rect 22145 4185 22190 4305
rect 22310 4185 22355 4305
rect 22475 4185 22530 4305
rect 22650 4185 22695 4305
rect 22815 4185 22860 4305
rect 22980 4185 23025 4305
rect 23145 4185 23200 4305
rect 23320 4185 23365 4305
rect 23485 4185 23530 4305
rect 23650 4185 23695 4305
rect 23815 4185 23870 4305
rect 23990 4185 24015 4305
rect 18485 4140 24015 4185
rect 18485 4020 18510 4140
rect 18630 4020 18675 4140
rect 18795 4020 18840 4140
rect 18960 4020 19005 4140
rect 19125 4020 19180 4140
rect 19300 4020 19345 4140
rect 19465 4020 19510 4140
rect 19630 4020 19675 4140
rect 19795 4020 19850 4140
rect 19970 4020 20015 4140
rect 20135 4020 20180 4140
rect 20300 4020 20345 4140
rect 20465 4020 20520 4140
rect 20640 4020 20685 4140
rect 20805 4020 20850 4140
rect 20970 4020 21015 4140
rect 21135 4020 21190 4140
rect 21310 4020 21355 4140
rect 21475 4020 21520 4140
rect 21640 4020 21685 4140
rect 21805 4020 21860 4140
rect 21980 4020 22025 4140
rect 22145 4020 22190 4140
rect 22310 4020 22355 4140
rect 22475 4020 22530 4140
rect 22650 4020 22695 4140
rect 22815 4020 22860 4140
rect 22980 4020 23025 4140
rect 23145 4020 23200 4140
rect 23320 4020 23365 4140
rect 23485 4020 23530 4140
rect 23650 4020 23695 4140
rect 23815 4020 23870 4140
rect 23990 4020 24015 4140
rect 18485 3975 24015 4020
rect 18485 3855 18510 3975
rect 18630 3855 18675 3975
rect 18795 3855 18840 3975
rect 18960 3855 19005 3975
rect 19125 3855 19180 3975
rect 19300 3855 19345 3975
rect 19465 3855 19510 3975
rect 19630 3855 19675 3975
rect 19795 3855 19850 3975
rect 19970 3855 20015 3975
rect 20135 3855 20180 3975
rect 20300 3855 20345 3975
rect 20465 3855 20520 3975
rect 20640 3855 20685 3975
rect 20805 3855 20850 3975
rect 20970 3855 21015 3975
rect 21135 3855 21190 3975
rect 21310 3855 21355 3975
rect 21475 3855 21520 3975
rect 21640 3855 21685 3975
rect 21805 3855 21860 3975
rect 21980 3855 22025 3975
rect 22145 3855 22190 3975
rect 22310 3855 22355 3975
rect 22475 3855 22530 3975
rect 22650 3855 22695 3975
rect 22815 3855 22860 3975
rect 22980 3855 23025 3975
rect 23145 3855 23200 3975
rect 23320 3855 23365 3975
rect 23485 3855 23530 3975
rect 23650 3855 23695 3975
rect 23815 3855 23870 3975
rect 23990 3855 24015 3975
rect 18485 3810 24015 3855
rect 18485 3690 18510 3810
rect 18630 3690 18675 3810
rect 18795 3690 18840 3810
rect 18960 3690 19005 3810
rect 19125 3690 19180 3810
rect 19300 3690 19345 3810
rect 19465 3690 19510 3810
rect 19630 3690 19675 3810
rect 19795 3690 19850 3810
rect 19970 3690 20015 3810
rect 20135 3690 20180 3810
rect 20300 3690 20345 3810
rect 20465 3690 20520 3810
rect 20640 3690 20685 3810
rect 20805 3690 20850 3810
rect 20970 3690 21015 3810
rect 21135 3690 21190 3810
rect 21310 3690 21355 3810
rect 21475 3690 21520 3810
rect 21640 3690 21685 3810
rect 21805 3690 21860 3810
rect 21980 3690 22025 3810
rect 22145 3690 22190 3810
rect 22310 3690 22355 3810
rect 22475 3690 22530 3810
rect 22650 3690 22695 3810
rect 22815 3690 22860 3810
rect 22980 3690 23025 3810
rect 23145 3690 23200 3810
rect 23320 3690 23365 3810
rect 23485 3690 23530 3810
rect 23650 3690 23695 3810
rect 23815 3690 23870 3810
rect 23990 3690 24015 3810
rect 18485 3635 24015 3690
rect 18485 3515 18510 3635
rect 18630 3515 18675 3635
rect 18795 3515 18840 3635
rect 18960 3515 19005 3635
rect 19125 3515 19180 3635
rect 19300 3515 19345 3635
rect 19465 3515 19510 3635
rect 19630 3515 19675 3635
rect 19795 3515 19850 3635
rect 19970 3515 20015 3635
rect 20135 3515 20180 3635
rect 20300 3515 20345 3635
rect 20465 3515 20520 3635
rect 20640 3515 20685 3635
rect 20805 3515 20850 3635
rect 20970 3515 21015 3635
rect 21135 3515 21190 3635
rect 21310 3515 21355 3635
rect 21475 3515 21520 3635
rect 21640 3515 21685 3635
rect 21805 3515 21860 3635
rect 21980 3515 22025 3635
rect 22145 3515 22190 3635
rect 22310 3515 22355 3635
rect 22475 3515 22530 3635
rect 22650 3515 22695 3635
rect 22815 3515 22860 3635
rect 22980 3515 23025 3635
rect 23145 3515 23200 3635
rect 23320 3515 23365 3635
rect 23485 3515 23530 3635
rect 23650 3515 23695 3635
rect 23815 3515 23870 3635
rect 23990 3515 24015 3635
rect 18485 3470 24015 3515
rect 18485 3350 18510 3470
rect 18630 3350 18675 3470
rect 18795 3350 18840 3470
rect 18960 3350 19005 3470
rect 19125 3350 19180 3470
rect 19300 3350 19345 3470
rect 19465 3350 19510 3470
rect 19630 3350 19675 3470
rect 19795 3350 19850 3470
rect 19970 3350 20015 3470
rect 20135 3350 20180 3470
rect 20300 3350 20345 3470
rect 20465 3350 20520 3470
rect 20640 3350 20685 3470
rect 20805 3350 20850 3470
rect 20970 3350 21015 3470
rect 21135 3350 21190 3470
rect 21310 3350 21355 3470
rect 21475 3350 21520 3470
rect 21640 3350 21685 3470
rect 21805 3350 21860 3470
rect 21980 3350 22025 3470
rect 22145 3350 22190 3470
rect 22310 3350 22355 3470
rect 22475 3350 22530 3470
rect 22650 3350 22695 3470
rect 22815 3350 22860 3470
rect 22980 3350 23025 3470
rect 23145 3350 23200 3470
rect 23320 3350 23365 3470
rect 23485 3350 23530 3470
rect 23650 3350 23695 3470
rect 23815 3350 23870 3470
rect 23990 3350 24015 3470
rect 18485 3305 24015 3350
rect 18485 3185 18510 3305
rect 18630 3185 18675 3305
rect 18795 3185 18840 3305
rect 18960 3185 19005 3305
rect 19125 3185 19180 3305
rect 19300 3185 19345 3305
rect 19465 3185 19510 3305
rect 19630 3185 19675 3305
rect 19795 3185 19850 3305
rect 19970 3185 20015 3305
rect 20135 3185 20180 3305
rect 20300 3185 20345 3305
rect 20465 3185 20520 3305
rect 20640 3185 20685 3305
rect 20805 3185 20850 3305
rect 20970 3185 21015 3305
rect 21135 3185 21190 3305
rect 21310 3185 21355 3305
rect 21475 3185 21520 3305
rect 21640 3185 21685 3305
rect 21805 3185 21860 3305
rect 21980 3185 22025 3305
rect 22145 3185 22190 3305
rect 22310 3185 22355 3305
rect 22475 3185 22530 3305
rect 22650 3185 22695 3305
rect 22815 3185 22860 3305
rect 22980 3185 23025 3305
rect 23145 3185 23200 3305
rect 23320 3185 23365 3305
rect 23485 3185 23530 3305
rect 23650 3185 23695 3305
rect 23815 3185 23870 3305
rect 23990 3185 24015 3305
rect 18485 3140 24015 3185
rect 18485 3020 18510 3140
rect 18630 3020 18675 3140
rect 18795 3020 18840 3140
rect 18960 3020 19005 3140
rect 19125 3020 19180 3140
rect 19300 3020 19345 3140
rect 19465 3020 19510 3140
rect 19630 3020 19675 3140
rect 19795 3020 19850 3140
rect 19970 3020 20015 3140
rect 20135 3020 20180 3140
rect 20300 3020 20345 3140
rect 20465 3020 20520 3140
rect 20640 3020 20685 3140
rect 20805 3020 20850 3140
rect 20970 3020 21015 3140
rect 21135 3020 21190 3140
rect 21310 3020 21355 3140
rect 21475 3020 21520 3140
rect 21640 3020 21685 3140
rect 21805 3020 21860 3140
rect 21980 3020 22025 3140
rect 22145 3020 22190 3140
rect 22310 3020 22355 3140
rect 22475 3020 22530 3140
rect 22650 3020 22695 3140
rect 22815 3020 22860 3140
rect 22980 3020 23025 3140
rect 23145 3020 23200 3140
rect 23320 3020 23365 3140
rect 23485 3020 23530 3140
rect 23650 3020 23695 3140
rect 23815 3020 23870 3140
rect 23990 3020 24015 3140
rect 18485 2965 24015 3020
rect 18485 2845 18510 2965
rect 18630 2845 18675 2965
rect 18795 2845 18840 2965
rect 18960 2845 19005 2965
rect 19125 2845 19180 2965
rect 19300 2845 19345 2965
rect 19465 2845 19510 2965
rect 19630 2845 19675 2965
rect 19795 2845 19850 2965
rect 19970 2845 20015 2965
rect 20135 2845 20180 2965
rect 20300 2845 20345 2965
rect 20465 2845 20520 2965
rect 20640 2845 20685 2965
rect 20805 2845 20850 2965
rect 20970 2845 21015 2965
rect 21135 2845 21190 2965
rect 21310 2845 21355 2965
rect 21475 2845 21520 2965
rect 21640 2845 21685 2965
rect 21805 2845 21860 2965
rect 21980 2845 22025 2965
rect 22145 2845 22190 2965
rect 22310 2845 22355 2965
rect 22475 2845 22530 2965
rect 22650 2845 22695 2965
rect 22815 2845 22860 2965
rect 22980 2845 23025 2965
rect 23145 2845 23200 2965
rect 23320 2845 23365 2965
rect 23485 2845 23530 2965
rect 23650 2845 23695 2965
rect 23815 2845 23870 2965
rect 23990 2845 24015 2965
rect 18485 2800 24015 2845
rect 18485 2680 18510 2800
rect 18630 2680 18675 2800
rect 18795 2680 18840 2800
rect 18960 2680 19005 2800
rect 19125 2680 19180 2800
rect 19300 2680 19345 2800
rect 19465 2680 19510 2800
rect 19630 2680 19675 2800
rect 19795 2680 19850 2800
rect 19970 2680 20015 2800
rect 20135 2680 20180 2800
rect 20300 2680 20345 2800
rect 20465 2680 20520 2800
rect 20640 2680 20685 2800
rect 20805 2680 20850 2800
rect 20970 2680 21015 2800
rect 21135 2680 21190 2800
rect 21310 2680 21355 2800
rect 21475 2680 21520 2800
rect 21640 2680 21685 2800
rect 21805 2680 21860 2800
rect 21980 2680 22025 2800
rect 22145 2680 22190 2800
rect 22310 2680 22355 2800
rect 22475 2680 22530 2800
rect 22650 2680 22695 2800
rect 22815 2680 22860 2800
rect 22980 2680 23025 2800
rect 23145 2680 23200 2800
rect 23320 2680 23365 2800
rect 23485 2680 23530 2800
rect 23650 2680 23695 2800
rect 23815 2680 23870 2800
rect 23990 2680 24015 2800
rect 18485 2635 24015 2680
rect 18485 2515 18510 2635
rect 18630 2515 18675 2635
rect 18795 2515 18840 2635
rect 18960 2515 19005 2635
rect 19125 2515 19180 2635
rect 19300 2515 19345 2635
rect 19465 2515 19510 2635
rect 19630 2515 19675 2635
rect 19795 2515 19850 2635
rect 19970 2515 20015 2635
rect 20135 2515 20180 2635
rect 20300 2515 20345 2635
rect 20465 2515 20520 2635
rect 20640 2515 20685 2635
rect 20805 2515 20850 2635
rect 20970 2515 21015 2635
rect 21135 2515 21190 2635
rect 21310 2515 21355 2635
rect 21475 2515 21520 2635
rect 21640 2515 21685 2635
rect 21805 2515 21860 2635
rect 21980 2515 22025 2635
rect 22145 2515 22190 2635
rect 22310 2515 22355 2635
rect 22475 2515 22530 2635
rect 22650 2515 22695 2635
rect 22815 2515 22860 2635
rect 22980 2515 23025 2635
rect 23145 2515 23200 2635
rect 23320 2515 23365 2635
rect 23485 2515 23530 2635
rect 23650 2515 23695 2635
rect 23815 2515 23870 2635
rect 23990 2515 24015 2635
rect 18485 2470 24015 2515
rect 18485 2350 18510 2470
rect 18630 2350 18675 2470
rect 18795 2350 18840 2470
rect 18960 2350 19005 2470
rect 19125 2350 19180 2470
rect 19300 2350 19345 2470
rect 19465 2350 19510 2470
rect 19630 2350 19675 2470
rect 19795 2350 19850 2470
rect 19970 2350 20015 2470
rect 20135 2350 20180 2470
rect 20300 2350 20345 2470
rect 20465 2350 20520 2470
rect 20640 2350 20685 2470
rect 20805 2350 20850 2470
rect 20970 2350 21015 2470
rect 21135 2350 21190 2470
rect 21310 2350 21355 2470
rect 21475 2350 21520 2470
rect 21640 2350 21685 2470
rect 21805 2350 21860 2470
rect 21980 2350 22025 2470
rect 22145 2350 22190 2470
rect 22310 2350 22355 2470
rect 22475 2350 22530 2470
rect 22650 2350 22695 2470
rect 22815 2350 22860 2470
rect 22980 2350 23025 2470
rect 23145 2350 23200 2470
rect 23320 2350 23365 2470
rect 23485 2350 23530 2470
rect 23650 2350 23695 2470
rect 23815 2350 23870 2470
rect 23990 2350 24015 2470
rect 18485 2295 24015 2350
rect 18485 2175 18510 2295
rect 18630 2175 18675 2295
rect 18795 2175 18840 2295
rect 18960 2175 19005 2295
rect 19125 2175 19180 2295
rect 19300 2175 19345 2295
rect 19465 2175 19510 2295
rect 19630 2175 19675 2295
rect 19795 2175 19850 2295
rect 19970 2175 20015 2295
rect 20135 2175 20180 2295
rect 20300 2175 20345 2295
rect 20465 2175 20520 2295
rect 20640 2175 20685 2295
rect 20805 2175 20850 2295
rect 20970 2175 21015 2295
rect 21135 2175 21190 2295
rect 21310 2175 21355 2295
rect 21475 2175 21520 2295
rect 21640 2175 21685 2295
rect 21805 2175 21860 2295
rect 21980 2175 22025 2295
rect 22145 2175 22190 2295
rect 22310 2175 22355 2295
rect 22475 2175 22530 2295
rect 22650 2175 22695 2295
rect 22815 2175 22860 2295
rect 22980 2175 23025 2295
rect 23145 2175 23200 2295
rect 23320 2175 23365 2295
rect 23485 2175 23530 2295
rect 23650 2175 23695 2295
rect 23815 2175 23870 2295
rect 23990 2175 24015 2295
rect 18485 2130 24015 2175
rect 18485 2010 18510 2130
rect 18630 2010 18675 2130
rect 18795 2010 18840 2130
rect 18960 2010 19005 2130
rect 19125 2010 19180 2130
rect 19300 2010 19345 2130
rect 19465 2010 19510 2130
rect 19630 2010 19675 2130
rect 19795 2010 19850 2130
rect 19970 2010 20015 2130
rect 20135 2010 20180 2130
rect 20300 2010 20345 2130
rect 20465 2010 20520 2130
rect 20640 2010 20685 2130
rect 20805 2010 20850 2130
rect 20970 2010 21015 2130
rect 21135 2010 21190 2130
rect 21310 2010 21355 2130
rect 21475 2010 21520 2130
rect 21640 2010 21685 2130
rect 21805 2010 21860 2130
rect 21980 2010 22025 2130
rect 22145 2010 22190 2130
rect 22310 2010 22355 2130
rect 22475 2010 22530 2130
rect 22650 2010 22695 2130
rect 22815 2010 22860 2130
rect 22980 2010 23025 2130
rect 23145 2010 23200 2130
rect 23320 2010 23365 2130
rect 23485 2010 23530 2130
rect 23650 2010 23695 2130
rect 23815 2010 23870 2130
rect 23990 2010 24015 2130
rect 18485 1965 24015 2010
rect 18485 1845 18510 1965
rect 18630 1845 18675 1965
rect 18795 1845 18840 1965
rect 18960 1845 19005 1965
rect 19125 1845 19180 1965
rect 19300 1845 19345 1965
rect 19465 1845 19510 1965
rect 19630 1845 19675 1965
rect 19795 1845 19850 1965
rect 19970 1845 20015 1965
rect 20135 1845 20180 1965
rect 20300 1845 20345 1965
rect 20465 1845 20520 1965
rect 20640 1845 20685 1965
rect 20805 1845 20850 1965
rect 20970 1845 21015 1965
rect 21135 1845 21190 1965
rect 21310 1845 21355 1965
rect 21475 1845 21520 1965
rect 21640 1845 21685 1965
rect 21805 1845 21860 1965
rect 21980 1845 22025 1965
rect 22145 1845 22190 1965
rect 22310 1845 22355 1965
rect 22475 1845 22530 1965
rect 22650 1845 22695 1965
rect 22815 1845 22860 1965
rect 22980 1845 23025 1965
rect 23145 1845 23200 1965
rect 23320 1845 23365 1965
rect 23485 1845 23530 1965
rect 23650 1845 23695 1965
rect 23815 1845 23870 1965
rect 23990 1845 24015 1965
rect 18485 1800 24015 1845
rect 18485 1680 18510 1800
rect 18630 1680 18675 1800
rect 18795 1680 18840 1800
rect 18960 1680 19005 1800
rect 19125 1680 19180 1800
rect 19300 1680 19345 1800
rect 19465 1680 19510 1800
rect 19630 1680 19675 1800
rect 19795 1680 19850 1800
rect 19970 1680 20015 1800
rect 20135 1680 20180 1800
rect 20300 1680 20345 1800
rect 20465 1680 20520 1800
rect 20640 1680 20685 1800
rect 20805 1680 20850 1800
rect 20970 1680 21015 1800
rect 21135 1680 21190 1800
rect 21310 1680 21355 1800
rect 21475 1680 21520 1800
rect 21640 1680 21685 1800
rect 21805 1680 21860 1800
rect 21980 1680 22025 1800
rect 22145 1680 22190 1800
rect 22310 1680 22355 1800
rect 22475 1680 22530 1800
rect 22650 1680 22695 1800
rect 22815 1680 22860 1800
rect 22980 1680 23025 1800
rect 23145 1680 23200 1800
rect 23320 1680 23365 1800
rect 23485 1680 23530 1800
rect 23650 1680 23695 1800
rect 23815 1680 23870 1800
rect 23990 1680 24015 1800
rect 18485 1610 24015 1680
rect 24175 7160 29705 7185
rect 24175 7040 24200 7160
rect 24320 7040 24365 7160
rect 24485 7040 24530 7160
rect 24650 7040 24695 7160
rect 24815 7040 24870 7160
rect 24990 7040 25035 7160
rect 25155 7040 25200 7160
rect 25320 7040 25365 7160
rect 25485 7040 25540 7160
rect 25660 7040 25705 7160
rect 25825 7040 25870 7160
rect 25990 7040 26035 7160
rect 26155 7040 26210 7160
rect 26330 7040 26375 7160
rect 26495 7040 26540 7160
rect 26660 7040 26705 7160
rect 26825 7040 26880 7160
rect 27000 7040 27045 7160
rect 27165 7040 27210 7160
rect 27330 7040 27375 7160
rect 27495 7040 27550 7160
rect 27670 7040 27715 7160
rect 27835 7040 27880 7160
rect 28000 7040 28045 7160
rect 28165 7040 28220 7160
rect 28340 7040 28385 7160
rect 28505 7040 28550 7160
rect 28670 7040 28715 7160
rect 28835 7040 28890 7160
rect 29010 7040 29055 7160
rect 29175 7040 29220 7160
rect 29340 7040 29385 7160
rect 29505 7040 29560 7160
rect 29680 7040 29705 7160
rect 24175 6985 29705 7040
rect 24175 6865 24200 6985
rect 24320 6865 24365 6985
rect 24485 6865 24530 6985
rect 24650 6865 24695 6985
rect 24815 6865 24870 6985
rect 24990 6865 25035 6985
rect 25155 6865 25200 6985
rect 25320 6865 25365 6985
rect 25485 6865 25540 6985
rect 25660 6865 25705 6985
rect 25825 6865 25870 6985
rect 25990 6865 26035 6985
rect 26155 6865 26210 6985
rect 26330 6865 26375 6985
rect 26495 6865 26540 6985
rect 26660 6865 26705 6985
rect 26825 6865 26880 6985
rect 27000 6865 27045 6985
rect 27165 6865 27210 6985
rect 27330 6865 27375 6985
rect 27495 6865 27550 6985
rect 27670 6865 27715 6985
rect 27835 6865 27880 6985
rect 28000 6865 28045 6985
rect 28165 6865 28220 6985
rect 28340 6865 28385 6985
rect 28505 6865 28550 6985
rect 28670 6865 28715 6985
rect 28835 6865 28890 6985
rect 29010 6865 29055 6985
rect 29175 6865 29220 6985
rect 29340 6865 29385 6985
rect 29505 6865 29560 6985
rect 29680 6865 29705 6985
rect 24175 6820 29705 6865
rect 24175 6700 24200 6820
rect 24320 6700 24365 6820
rect 24485 6700 24530 6820
rect 24650 6700 24695 6820
rect 24815 6700 24870 6820
rect 24990 6700 25035 6820
rect 25155 6700 25200 6820
rect 25320 6700 25365 6820
rect 25485 6700 25540 6820
rect 25660 6700 25705 6820
rect 25825 6700 25870 6820
rect 25990 6700 26035 6820
rect 26155 6700 26210 6820
rect 26330 6700 26375 6820
rect 26495 6700 26540 6820
rect 26660 6700 26705 6820
rect 26825 6700 26880 6820
rect 27000 6700 27045 6820
rect 27165 6700 27210 6820
rect 27330 6700 27375 6820
rect 27495 6700 27550 6820
rect 27670 6700 27715 6820
rect 27835 6700 27880 6820
rect 28000 6700 28045 6820
rect 28165 6700 28220 6820
rect 28340 6700 28385 6820
rect 28505 6700 28550 6820
rect 28670 6700 28715 6820
rect 28835 6700 28890 6820
rect 29010 6700 29055 6820
rect 29175 6700 29220 6820
rect 29340 6700 29385 6820
rect 29505 6700 29560 6820
rect 29680 6700 29705 6820
rect 24175 6655 29705 6700
rect 24175 6535 24200 6655
rect 24320 6535 24365 6655
rect 24485 6535 24530 6655
rect 24650 6535 24695 6655
rect 24815 6535 24870 6655
rect 24990 6535 25035 6655
rect 25155 6535 25200 6655
rect 25320 6535 25365 6655
rect 25485 6535 25540 6655
rect 25660 6535 25705 6655
rect 25825 6535 25870 6655
rect 25990 6535 26035 6655
rect 26155 6535 26210 6655
rect 26330 6535 26375 6655
rect 26495 6535 26540 6655
rect 26660 6535 26705 6655
rect 26825 6535 26880 6655
rect 27000 6535 27045 6655
rect 27165 6535 27210 6655
rect 27330 6535 27375 6655
rect 27495 6535 27550 6655
rect 27670 6535 27715 6655
rect 27835 6535 27880 6655
rect 28000 6535 28045 6655
rect 28165 6535 28220 6655
rect 28340 6535 28385 6655
rect 28505 6535 28550 6655
rect 28670 6535 28715 6655
rect 28835 6535 28890 6655
rect 29010 6535 29055 6655
rect 29175 6535 29220 6655
rect 29340 6535 29385 6655
rect 29505 6535 29560 6655
rect 29680 6535 29705 6655
rect 24175 6490 29705 6535
rect 24175 6370 24200 6490
rect 24320 6370 24365 6490
rect 24485 6370 24530 6490
rect 24650 6370 24695 6490
rect 24815 6370 24870 6490
rect 24990 6370 25035 6490
rect 25155 6370 25200 6490
rect 25320 6370 25365 6490
rect 25485 6370 25540 6490
rect 25660 6370 25705 6490
rect 25825 6370 25870 6490
rect 25990 6370 26035 6490
rect 26155 6370 26210 6490
rect 26330 6370 26375 6490
rect 26495 6370 26540 6490
rect 26660 6370 26705 6490
rect 26825 6370 26880 6490
rect 27000 6370 27045 6490
rect 27165 6370 27210 6490
rect 27330 6370 27375 6490
rect 27495 6370 27550 6490
rect 27670 6370 27715 6490
rect 27835 6370 27880 6490
rect 28000 6370 28045 6490
rect 28165 6370 28220 6490
rect 28340 6370 28385 6490
rect 28505 6370 28550 6490
rect 28670 6370 28715 6490
rect 28835 6370 28890 6490
rect 29010 6370 29055 6490
rect 29175 6370 29220 6490
rect 29340 6370 29385 6490
rect 29505 6370 29560 6490
rect 29680 6370 29705 6490
rect 24175 6315 29705 6370
rect 24175 6195 24200 6315
rect 24320 6195 24365 6315
rect 24485 6195 24530 6315
rect 24650 6195 24695 6315
rect 24815 6195 24870 6315
rect 24990 6195 25035 6315
rect 25155 6195 25200 6315
rect 25320 6195 25365 6315
rect 25485 6195 25540 6315
rect 25660 6195 25705 6315
rect 25825 6195 25870 6315
rect 25990 6195 26035 6315
rect 26155 6195 26210 6315
rect 26330 6195 26375 6315
rect 26495 6195 26540 6315
rect 26660 6195 26705 6315
rect 26825 6195 26880 6315
rect 27000 6195 27045 6315
rect 27165 6195 27210 6315
rect 27330 6195 27375 6315
rect 27495 6195 27550 6315
rect 27670 6195 27715 6315
rect 27835 6195 27880 6315
rect 28000 6195 28045 6315
rect 28165 6195 28220 6315
rect 28340 6195 28385 6315
rect 28505 6195 28550 6315
rect 28670 6195 28715 6315
rect 28835 6195 28890 6315
rect 29010 6195 29055 6315
rect 29175 6195 29220 6315
rect 29340 6195 29385 6315
rect 29505 6195 29560 6315
rect 29680 6195 29705 6315
rect 24175 6150 29705 6195
rect 24175 6030 24200 6150
rect 24320 6030 24365 6150
rect 24485 6030 24530 6150
rect 24650 6030 24695 6150
rect 24815 6030 24870 6150
rect 24990 6030 25035 6150
rect 25155 6030 25200 6150
rect 25320 6030 25365 6150
rect 25485 6030 25540 6150
rect 25660 6030 25705 6150
rect 25825 6030 25870 6150
rect 25990 6030 26035 6150
rect 26155 6030 26210 6150
rect 26330 6030 26375 6150
rect 26495 6030 26540 6150
rect 26660 6030 26705 6150
rect 26825 6030 26880 6150
rect 27000 6030 27045 6150
rect 27165 6030 27210 6150
rect 27330 6030 27375 6150
rect 27495 6030 27550 6150
rect 27670 6030 27715 6150
rect 27835 6030 27880 6150
rect 28000 6030 28045 6150
rect 28165 6030 28220 6150
rect 28340 6030 28385 6150
rect 28505 6030 28550 6150
rect 28670 6030 28715 6150
rect 28835 6030 28890 6150
rect 29010 6030 29055 6150
rect 29175 6030 29220 6150
rect 29340 6030 29385 6150
rect 29505 6030 29560 6150
rect 29680 6030 29705 6150
rect 24175 5985 29705 6030
rect 24175 5865 24200 5985
rect 24320 5865 24365 5985
rect 24485 5865 24530 5985
rect 24650 5865 24695 5985
rect 24815 5865 24870 5985
rect 24990 5865 25035 5985
rect 25155 5865 25200 5985
rect 25320 5865 25365 5985
rect 25485 5865 25540 5985
rect 25660 5865 25705 5985
rect 25825 5865 25870 5985
rect 25990 5865 26035 5985
rect 26155 5865 26210 5985
rect 26330 5865 26375 5985
rect 26495 5865 26540 5985
rect 26660 5865 26705 5985
rect 26825 5865 26880 5985
rect 27000 5865 27045 5985
rect 27165 5865 27210 5985
rect 27330 5865 27375 5985
rect 27495 5865 27550 5985
rect 27670 5865 27715 5985
rect 27835 5865 27880 5985
rect 28000 5865 28045 5985
rect 28165 5865 28220 5985
rect 28340 5865 28385 5985
rect 28505 5865 28550 5985
rect 28670 5865 28715 5985
rect 28835 5865 28890 5985
rect 29010 5865 29055 5985
rect 29175 5865 29220 5985
rect 29340 5865 29385 5985
rect 29505 5865 29560 5985
rect 29680 5865 29705 5985
rect 24175 5820 29705 5865
rect 24175 5700 24200 5820
rect 24320 5700 24365 5820
rect 24485 5700 24530 5820
rect 24650 5700 24695 5820
rect 24815 5700 24870 5820
rect 24990 5700 25035 5820
rect 25155 5700 25200 5820
rect 25320 5700 25365 5820
rect 25485 5700 25540 5820
rect 25660 5700 25705 5820
rect 25825 5700 25870 5820
rect 25990 5700 26035 5820
rect 26155 5700 26210 5820
rect 26330 5700 26375 5820
rect 26495 5700 26540 5820
rect 26660 5700 26705 5820
rect 26825 5700 26880 5820
rect 27000 5700 27045 5820
rect 27165 5700 27210 5820
rect 27330 5700 27375 5820
rect 27495 5700 27550 5820
rect 27670 5700 27715 5820
rect 27835 5700 27880 5820
rect 28000 5700 28045 5820
rect 28165 5700 28220 5820
rect 28340 5700 28385 5820
rect 28505 5700 28550 5820
rect 28670 5700 28715 5820
rect 28835 5700 28890 5820
rect 29010 5700 29055 5820
rect 29175 5700 29220 5820
rect 29340 5700 29385 5820
rect 29505 5700 29560 5820
rect 29680 5700 29705 5820
rect 24175 5645 29705 5700
rect 24175 5525 24200 5645
rect 24320 5525 24365 5645
rect 24485 5525 24530 5645
rect 24650 5525 24695 5645
rect 24815 5525 24870 5645
rect 24990 5525 25035 5645
rect 25155 5525 25200 5645
rect 25320 5525 25365 5645
rect 25485 5525 25540 5645
rect 25660 5525 25705 5645
rect 25825 5525 25870 5645
rect 25990 5525 26035 5645
rect 26155 5525 26210 5645
rect 26330 5525 26375 5645
rect 26495 5525 26540 5645
rect 26660 5525 26705 5645
rect 26825 5525 26880 5645
rect 27000 5525 27045 5645
rect 27165 5525 27210 5645
rect 27330 5525 27375 5645
rect 27495 5525 27550 5645
rect 27670 5525 27715 5645
rect 27835 5525 27880 5645
rect 28000 5525 28045 5645
rect 28165 5525 28220 5645
rect 28340 5525 28385 5645
rect 28505 5525 28550 5645
rect 28670 5525 28715 5645
rect 28835 5525 28890 5645
rect 29010 5525 29055 5645
rect 29175 5525 29220 5645
rect 29340 5525 29385 5645
rect 29505 5525 29560 5645
rect 29680 5525 29705 5645
rect 24175 5480 29705 5525
rect 24175 5360 24200 5480
rect 24320 5360 24365 5480
rect 24485 5360 24530 5480
rect 24650 5360 24695 5480
rect 24815 5360 24870 5480
rect 24990 5360 25035 5480
rect 25155 5360 25200 5480
rect 25320 5360 25365 5480
rect 25485 5360 25540 5480
rect 25660 5360 25705 5480
rect 25825 5360 25870 5480
rect 25990 5360 26035 5480
rect 26155 5360 26210 5480
rect 26330 5360 26375 5480
rect 26495 5360 26540 5480
rect 26660 5360 26705 5480
rect 26825 5360 26880 5480
rect 27000 5360 27045 5480
rect 27165 5360 27210 5480
rect 27330 5360 27375 5480
rect 27495 5360 27550 5480
rect 27670 5360 27715 5480
rect 27835 5360 27880 5480
rect 28000 5360 28045 5480
rect 28165 5360 28220 5480
rect 28340 5360 28385 5480
rect 28505 5360 28550 5480
rect 28670 5360 28715 5480
rect 28835 5360 28890 5480
rect 29010 5360 29055 5480
rect 29175 5360 29220 5480
rect 29340 5360 29385 5480
rect 29505 5360 29560 5480
rect 29680 5360 29705 5480
rect 24175 5315 29705 5360
rect 24175 5195 24200 5315
rect 24320 5195 24365 5315
rect 24485 5195 24530 5315
rect 24650 5195 24695 5315
rect 24815 5195 24870 5315
rect 24990 5195 25035 5315
rect 25155 5195 25200 5315
rect 25320 5195 25365 5315
rect 25485 5195 25540 5315
rect 25660 5195 25705 5315
rect 25825 5195 25870 5315
rect 25990 5195 26035 5315
rect 26155 5195 26210 5315
rect 26330 5195 26375 5315
rect 26495 5195 26540 5315
rect 26660 5195 26705 5315
rect 26825 5195 26880 5315
rect 27000 5195 27045 5315
rect 27165 5195 27210 5315
rect 27330 5195 27375 5315
rect 27495 5195 27550 5315
rect 27670 5195 27715 5315
rect 27835 5195 27880 5315
rect 28000 5195 28045 5315
rect 28165 5195 28220 5315
rect 28340 5195 28385 5315
rect 28505 5195 28550 5315
rect 28670 5195 28715 5315
rect 28835 5195 28890 5315
rect 29010 5195 29055 5315
rect 29175 5195 29220 5315
rect 29340 5195 29385 5315
rect 29505 5195 29560 5315
rect 29680 5195 29705 5315
rect 24175 5150 29705 5195
rect 24175 5030 24200 5150
rect 24320 5030 24365 5150
rect 24485 5030 24530 5150
rect 24650 5030 24695 5150
rect 24815 5030 24870 5150
rect 24990 5030 25035 5150
rect 25155 5030 25200 5150
rect 25320 5030 25365 5150
rect 25485 5030 25540 5150
rect 25660 5030 25705 5150
rect 25825 5030 25870 5150
rect 25990 5030 26035 5150
rect 26155 5030 26210 5150
rect 26330 5030 26375 5150
rect 26495 5030 26540 5150
rect 26660 5030 26705 5150
rect 26825 5030 26880 5150
rect 27000 5030 27045 5150
rect 27165 5030 27210 5150
rect 27330 5030 27375 5150
rect 27495 5030 27550 5150
rect 27670 5030 27715 5150
rect 27835 5030 27880 5150
rect 28000 5030 28045 5150
rect 28165 5030 28220 5150
rect 28340 5030 28385 5150
rect 28505 5030 28550 5150
rect 28670 5030 28715 5150
rect 28835 5030 28890 5150
rect 29010 5030 29055 5150
rect 29175 5030 29220 5150
rect 29340 5030 29385 5150
rect 29505 5030 29560 5150
rect 29680 5030 29705 5150
rect 24175 4975 29705 5030
rect 24175 4855 24200 4975
rect 24320 4855 24365 4975
rect 24485 4855 24530 4975
rect 24650 4855 24695 4975
rect 24815 4855 24870 4975
rect 24990 4855 25035 4975
rect 25155 4855 25200 4975
rect 25320 4855 25365 4975
rect 25485 4855 25540 4975
rect 25660 4855 25705 4975
rect 25825 4855 25870 4975
rect 25990 4855 26035 4975
rect 26155 4855 26210 4975
rect 26330 4855 26375 4975
rect 26495 4855 26540 4975
rect 26660 4855 26705 4975
rect 26825 4855 26880 4975
rect 27000 4855 27045 4975
rect 27165 4855 27210 4975
rect 27330 4855 27375 4975
rect 27495 4855 27550 4975
rect 27670 4855 27715 4975
rect 27835 4855 27880 4975
rect 28000 4855 28045 4975
rect 28165 4855 28220 4975
rect 28340 4855 28385 4975
rect 28505 4855 28550 4975
rect 28670 4855 28715 4975
rect 28835 4855 28890 4975
rect 29010 4855 29055 4975
rect 29175 4855 29220 4975
rect 29340 4855 29385 4975
rect 29505 4855 29560 4975
rect 29680 4855 29705 4975
rect 24175 4810 29705 4855
rect 24175 4690 24200 4810
rect 24320 4690 24365 4810
rect 24485 4690 24530 4810
rect 24650 4690 24695 4810
rect 24815 4690 24870 4810
rect 24990 4690 25035 4810
rect 25155 4690 25200 4810
rect 25320 4690 25365 4810
rect 25485 4690 25540 4810
rect 25660 4690 25705 4810
rect 25825 4690 25870 4810
rect 25990 4690 26035 4810
rect 26155 4690 26210 4810
rect 26330 4690 26375 4810
rect 26495 4690 26540 4810
rect 26660 4690 26705 4810
rect 26825 4690 26880 4810
rect 27000 4690 27045 4810
rect 27165 4690 27210 4810
rect 27330 4690 27375 4810
rect 27495 4690 27550 4810
rect 27670 4690 27715 4810
rect 27835 4690 27880 4810
rect 28000 4690 28045 4810
rect 28165 4690 28220 4810
rect 28340 4690 28385 4810
rect 28505 4690 28550 4810
rect 28670 4690 28715 4810
rect 28835 4690 28890 4810
rect 29010 4690 29055 4810
rect 29175 4690 29220 4810
rect 29340 4690 29385 4810
rect 29505 4690 29560 4810
rect 29680 4690 29705 4810
rect 24175 4645 29705 4690
rect 24175 4525 24200 4645
rect 24320 4525 24365 4645
rect 24485 4525 24530 4645
rect 24650 4525 24695 4645
rect 24815 4525 24870 4645
rect 24990 4525 25035 4645
rect 25155 4525 25200 4645
rect 25320 4525 25365 4645
rect 25485 4525 25540 4645
rect 25660 4525 25705 4645
rect 25825 4525 25870 4645
rect 25990 4525 26035 4645
rect 26155 4525 26210 4645
rect 26330 4525 26375 4645
rect 26495 4525 26540 4645
rect 26660 4525 26705 4645
rect 26825 4525 26880 4645
rect 27000 4525 27045 4645
rect 27165 4525 27210 4645
rect 27330 4525 27375 4645
rect 27495 4525 27550 4645
rect 27670 4525 27715 4645
rect 27835 4525 27880 4645
rect 28000 4525 28045 4645
rect 28165 4525 28220 4645
rect 28340 4525 28385 4645
rect 28505 4525 28550 4645
rect 28670 4525 28715 4645
rect 28835 4525 28890 4645
rect 29010 4525 29055 4645
rect 29175 4525 29220 4645
rect 29340 4525 29385 4645
rect 29505 4525 29560 4645
rect 29680 4525 29705 4645
rect 24175 4480 29705 4525
rect 24175 4360 24200 4480
rect 24320 4360 24365 4480
rect 24485 4360 24530 4480
rect 24650 4360 24695 4480
rect 24815 4360 24870 4480
rect 24990 4360 25035 4480
rect 25155 4360 25200 4480
rect 25320 4360 25365 4480
rect 25485 4360 25540 4480
rect 25660 4360 25705 4480
rect 25825 4360 25870 4480
rect 25990 4360 26035 4480
rect 26155 4360 26210 4480
rect 26330 4360 26375 4480
rect 26495 4360 26540 4480
rect 26660 4360 26705 4480
rect 26825 4360 26880 4480
rect 27000 4360 27045 4480
rect 27165 4360 27210 4480
rect 27330 4360 27375 4480
rect 27495 4360 27550 4480
rect 27670 4360 27715 4480
rect 27835 4360 27880 4480
rect 28000 4360 28045 4480
rect 28165 4360 28220 4480
rect 28340 4360 28385 4480
rect 28505 4360 28550 4480
rect 28670 4360 28715 4480
rect 28835 4360 28890 4480
rect 29010 4360 29055 4480
rect 29175 4360 29220 4480
rect 29340 4360 29385 4480
rect 29505 4360 29560 4480
rect 29680 4360 29705 4480
rect 24175 4305 29705 4360
rect 24175 4185 24200 4305
rect 24320 4185 24365 4305
rect 24485 4185 24530 4305
rect 24650 4185 24695 4305
rect 24815 4185 24870 4305
rect 24990 4185 25035 4305
rect 25155 4185 25200 4305
rect 25320 4185 25365 4305
rect 25485 4185 25540 4305
rect 25660 4185 25705 4305
rect 25825 4185 25870 4305
rect 25990 4185 26035 4305
rect 26155 4185 26210 4305
rect 26330 4185 26375 4305
rect 26495 4185 26540 4305
rect 26660 4185 26705 4305
rect 26825 4185 26880 4305
rect 27000 4185 27045 4305
rect 27165 4185 27210 4305
rect 27330 4185 27375 4305
rect 27495 4185 27550 4305
rect 27670 4185 27715 4305
rect 27835 4185 27880 4305
rect 28000 4185 28045 4305
rect 28165 4185 28220 4305
rect 28340 4185 28385 4305
rect 28505 4185 28550 4305
rect 28670 4185 28715 4305
rect 28835 4185 28890 4305
rect 29010 4185 29055 4305
rect 29175 4185 29220 4305
rect 29340 4185 29385 4305
rect 29505 4185 29560 4305
rect 29680 4185 29705 4305
rect 24175 4140 29705 4185
rect 24175 4020 24200 4140
rect 24320 4020 24365 4140
rect 24485 4020 24530 4140
rect 24650 4020 24695 4140
rect 24815 4020 24870 4140
rect 24990 4020 25035 4140
rect 25155 4020 25200 4140
rect 25320 4020 25365 4140
rect 25485 4020 25540 4140
rect 25660 4020 25705 4140
rect 25825 4020 25870 4140
rect 25990 4020 26035 4140
rect 26155 4020 26210 4140
rect 26330 4020 26375 4140
rect 26495 4020 26540 4140
rect 26660 4020 26705 4140
rect 26825 4020 26880 4140
rect 27000 4020 27045 4140
rect 27165 4020 27210 4140
rect 27330 4020 27375 4140
rect 27495 4020 27550 4140
rect 27670 4020 27715 4140
rect 27835 4020 27880 4140
rect 28000 4020 28045 4140
rect 28165 4020 28220 4140
rect 28340 4020 28385 4140
rect 28505 4020 28550 4140
rect 28670 4020 28715 4140
rect 28835 4020 28890 4140
rect 29010 4020 29055 4140
rect 29175 4020 29220 4140
rect 29340 4020 29385 4140
rect 29505 4020 29560 4140
rect 29680 4020 29705 4140
rect 24175 3975 29705 4020
rect 24175 3855 24200 3975
rect 24320 3855 24365 3975
rect 24485 3855 24530 3975
rect 24650 3855 24695 3975
rect 24815 3855 24870 3975
rect 24990 3855 25035 3975
rect 25155 3855 25200 3975
rect 25320 3855 25365 3975
rect 25485 3855 25540 3975
rect 25660 3855 25705 3975
rect 25825 3855 25870 3975
rect 25990 3855 26035 3975
rect 26155 3855 26210 3975
rect 26330 3855 26375 3975
rect 26495 3855 26540 3975
rect 26660 3855 26705 3975
rect 26825 3855 26880 3975
rect 27000 3855 27045 3975
rect 27165 3855 27210 3975
rect 27330 3855 27375 3975
rect 27495 3855 27550 3975
rect 27670 3855 27715 3975
rect 27835 3855 27880 3975
rect 28000 3855 28045 3975
rect 28165 3855 28220 3975
rect 28340 3855 28385 3975
rect 28505 3855 28550 3975
rect 28670 3855 28715 3975
rect 28835 3855 28890 3975
rect 29010 3855 29055 3975
rect 29175 3855 29220 3975
rect 29340 3855 29385 3975
rect 29505 3855 29560 3975
rect 29680 3855 29705 3975
rect 24175 3810 29705 3855
rect 24175 3690 24200 3810
rect 24320 3690 24365 3810
rect 24485 3690 24530 3810
rect 24650 3690 24695 3810
rect 24815 3690 24870 3810
rect 24990 3690 25035 3810
rect 25155 3690 25200 3810
rect 25320 3690 25365 3810
rect 25485 3690 25540 3810
rect 25660 3690 25705 3810
rect 25825 3690 25870 3810
rect 25990 3690 26035 3810
rect 26155 3690 26210 3810
rect 26330 3690 26375 3810
rect 26495 3690 26540 3810
rect 26660 3690 26705 3810
rect 26825 3690 26880 3810
rect 27000 3690 27045 3810
rect 27165 3690 27210 3810
rect 27330 3690 27375 3810
rect 27495 3690 27550 3810
rect 27670 3690 27715 3810
rect 27835 3690 27880 3810
rect 28000 3690 28045 3810
rect 28165 3690 28220 3810
rect 28340 3690 28385 3810
rect 28505 3690 28550 3810
rect 28670 3690 28715 3810
rect 28835 3690 28890 3810
rect 29010 3690 29055 3810
rect 29175 3690 29220 3810
rect 29340 3690 29385 3810
rect 29505 3690 29560 3810
rect 29680 3690 29705 3810
rect 24175 3635 29705 3690
rect 24175 3515 24200 3635
rect 24320 3515 24365 3635
rect 24485 3515 24530 3635
rect 24650 3515 24695 3635
rect 24815 3515 24870 3635
rect 24990 3515 25035 3635
rect 25155 3515 25200 3635
rect 25320 3515 25365 3635
rect 25485 3515 25540 3635
rect 25660 3515 25705 3635
rect 25825 3515 25870 3635
rect 25990 3515 26035 3635
rect 26155 3515 26210 3635
rect 26330 3515 26375 3635
rect 26495 3515 26540 3635
rect 26660 3515 26705 3635
rect 26825 3515 26880 3635
rect 27000 3515 27045 3635
rect 27165 3515 27210 3635
rect 27330 3515 27375 3635
rect 27495 3515 27550 3635
rect 27670 3515 27715 3635
rect 27835 3515 27880 3635
rect 28000 3515 28045 3635
rect 28165 3515 28220 3635
rect 28340 3515 28385 3635
rect 28505 3515 28550 3635
rect 28670 3515 28715 3635
rect 28835 3515 28890 3635
rect 29010 3515 29055 3635
rect 29175 3515 29220 3635
rect 29340 3515 29385 3635
rect 29505 3515 29560 3635
rect 29680 3515 29705 3635
rect 24175 3470 29705 3515
rect 24175 3350 24200 3470
rect 24320 3350 24365 3470
rect 24485 3350 24530 3470
rect 24650 3350 24695 3470
rect 24815 3350 24870 3470
rect 24990 3350 25035 3470
rect 25155 3350 25200 3470
rect 25320 3350 25365 3470
rect 25485 3350 25540 3470
rect 25660 3350 25705 3470
rect 25825 3350 25870 3470
rect 25990 3350 26035 3470
rect 26155 3350 26210 3470
rect 26330 3350 26375 3470
rect 26495 3350 26540 3470
rect 26660 3350 26705 3470
rect 26825 3350 26880 3470
rect 27000 3350 27045 3470
rect 27165 3350 27210 3470
rect 27330 3350 27375 3470
rect 27495 3350 27550 3470
rect 27670 3350 27715 3470
rect 27835 3350 27880 3470
rect 28000 3350 28045 3470
rect 28165 3350 28220 3470
rect 28340 3350 28385 3470
rect 28505 3350 28550 3470
rect 28670 3350 28715 3470
rect 28835 3350 28890 3470
rect 29010 3350 29055 3470
rect 29175 3350 29220 3470
rect 29340 3350 29385 3470
rect 29505 3350 29560 3470
rect 29680 3350 29705 3470
rect 24175 3305 29705 3350
rect 24175 3185 24200 3305
rect 24320 3185 24365 3305
rect 24485 3185 24530 3305
rect 24650 3185 24695 3305
rect 24815 3185 24870 3305
rect 24990 3185 25035 3305
rect 25155 3185 25200 3305
rect 25320 3185 25365 3305
rect 25485 3185 25540 3305
rect 25660 3185 25705 3305
rect 25825 3185 25870 3305
rect 25990 3185 26035 3305
rect 26155 3185 26210 3305
rect 26330 3185 26375 3305
rect 26495 3185 26540 3305
rect 26660 3185 26705 3305
rect 26825 3185 26880 3305
rect 27000 3185 27045 3305
rect 27165 3185 27210 3305
rect 27330 3185 27375 3305
rect 27495 3185 27550 3305
rect 27670 3185 27715 3305
rect 27835 3185 27880 3305
rect 28000 3185 28045 3305
rect 28165 3185 28220 3305
rect 28340 3185 28385 3305
rect 28505 3185 28550 3305
rect 28670 3185 28715 3305
rect 28835 3185 28890 3305
rect 29010 3185 29055 3305
rect 29175 3185 29220 3305
rect 29340 3185 29385 3305
rect 29505 3185 29560 3305
rect 29680 3185 29705 3305
rect 24175 3140 29705 3185
rect 24175 3020 24200 3140
rect 24320 3020 24365 3140
rect 24485 3020 24530 3140
rect 24650 3020 24695 3140
rect 24815 3020 24870 3140
rect 24990 3020 25035 3140
rect 25155 3020 25200 3140
rect 25320 3020 25365 3140
rect 25485 3020 25540 3140
rect 25660 3020 25705 3140
rect 25825 3020 25870 3140
rect 25990 3020 26035 3140
rect 26155 3020 26210 3140
rect 26330 3020 26375 3140
rect 26495 3020 26540 3140
rect 26660 3020 26705 3140
rect 26825 3020 26880 3140
rect 27000 3020 27045 3140
rect 27165 3020 27210 3140
rect 27330 3020 27375 3140
rect 27495 3020 27550 3140
rect 27670 3020 27715 3140
rect 27835 3020 27880 3140
rect 28000 3020 28045 3140
rect 28165 3020 28220 3140
rect 28340 3020 28385 3140
rect 28505 3020 28550 3140
rect 28670 3020 28715 3140
rect 28835 3020 28890 3140
rect 29010 3020 29055 3140
rect 29175 3020 29220 3140
rect 29340 3020 29385 3140
rect 29505 3020 29560 3140
rect 29680 3020 29705 3140
rect 24175 2965 29705 3020
rect 24175 2845 24200 2965
rect 24320 2845 24365 2965
rect 24485 2845 24530 2965
rect 24650 2845 24695 2965
rect 24815 2845 24870 2965
rect 24990 2845 25035 2965
rect 25155 2845 25200 2965
rect 25320 2845 25365 2965
rect 25485 2845 25540 2965
rect 25660 2845 25705 2965
rect 25825 2845 25870 2965
rect 25990 2845 26035 2965
rect 26155 2845 26210 2965
rect 26330 2845 26375 2965
rect 26495 2845 26540 2965
rect 26660 2845 26705 2965
rect 26825 2845 26880 2965
rect 27000 2845 27045 2965
rect 27165 2845 27210 2965
rect 27330 2845 27375 2965
rect 27495 2845 27550 2965
rect 27670 2845 27715 2965
rect 27835 2845 27880 2965
rect 28000 2845 28045 2965
rect 28165 2845 28220 2965
rect 28340 2845 28385 2965
rect 28505 2845 28550 2965
rect 28670 2845 28715 2965
rect 28835 2845 28890 2965
rect 29010 2845 29055 2965
rect 29175 2845 29220 2965
rect 29340 2845 29385 2965
rect 29505 2845 29560 2965
rect 29680 2845 29705 2965
rect 24175 2800 29705 2845
rect 24175 2680 24200 2800
rect 24320 2680 24365 2800
rect 24485 2680 24530 2800
rect 24650 2680 24695 2800
rect 24815 2680 24870 2800
rect 24990 2680 25035 2800
rect 25155 2680 25200 2800
rect 25320 2680 25365 2800
rect 25485 2680 25540 2800
rect 25660 2680 25705 2800
rect 25825 2680 25870 2800
rect 25990 2680 26035 2800
rect 26155 2680 26210 2800
rect 26330 2680 26375 2800
rect 26495 2680 26540 2800
rect 26660 2680 26705 2800
rect 26825 2680 26880 2800
rect 27000 2680 27045 2800
rect 27165 2680 27210 2800
rect 27330 2680 27375 2800
rect 27495 2680 27550 2800
rect 27670 2680 27715 2800
rect 27835 2680 27880 2800
rect 28000 2680 28045 2800
rect 28165 2680 28220 2800
rect 28340 2680 28385 2800
rect 28505 2680 28550 2800
rect 28670 2680 28715 2800
rect 28835 2680 28890 2800
rect 29010 2680 29055 2800
rect 29175 2680 29220 2800
rect 29340 2680 29385 2800
rect 29505 2680 29560 2800
rect 29680 2680 29705 2800
rect 24175 2635 29705 2680
rect 24175 2515 24200 2635
rect 24320 2515 24365 2635
rect 24485 2515 24530 2635
rect 24650 2515 24695 2635
rect 24815 2515 24870 2635
rect 24990 2515 25035 2635
rect 25155 2515 25200 2635
rect 25320 2515 25365 2635
rect 25485 2515 25540 2635
rect 25660 2515 25705 2635
rect 25825 2515 25870 2635
rect 25990 2515 26035 2635
rect 26155 2515 26210 2635
rect 26330 2515 26375 2635
rect 26495 2515 26540 2635
rect 26660 2515 26705 2635
rect 26825 2515 26880 2635
rect 27000 2515 27045 2635
rect 27165 2515 27210 2635
rect 27330 2515 27375 2635
rect 27495 2515 27550 2635
rect 27670 2515 27715 2635
rect 27835 2515 27880 2635
rect 28000 2515 28045 2635
rect 28165 2515 28220 2635
rect 28340 2515 28385 2635
rect 28505 2515 28550 2635
rect 28670 2515 28715 2635
rect 28835 2515 28890 2635
rect 29010 2515 29055 2635
rect 29175 2515 29220 2635
rect 29340 2515 29385 2635
rect 29505 2515 29560 2635
rect 29680 2515 29705 2635
rect 24175 2470 29705 2515
rect 24175 2350 24200 2470
rect 24320 2350 24365 2470
rect 24485 2350 24530 2470
rect 24650 2350 24695 2470
rect 24815 2350 24870 2470
rect 24990 2350 25035 2470
rect 25155 2350 25200 2470
rect 25320 2350 25365 2470
rect 25485 2350 25540 2470
rect 25660 2350 25705 2470
rect 25825 2350 25870 2470
rect 25990 2350 26035 2470
rect 26155 2350 26210 2470
rect 26330 2350 26375 2470
rect 26495 2350 26540 2470
rect 26660 2350 26705 2470
rect 26825 2350 26880 2470
rect 27000 2350 27045 2470
rect 27165 2350 27210 2470
rect 27330 2350 27375 2470
rect 27495 2350 27550 2470
rect 27670 2350 27715 2470
rect 27835 2350 27880 2470
rect 28000 2350 28045 2470
rect 28165 2350 28220 2470
rect 28340 2350 28385 2470
rect 28505 2350 28550 2470
rect 28670 2350 28715 2470
rect 28835 2350 28890 2470
rect 29010 2350 29055 2470
rect 29175 2350 29220 2470
rect 29340 2350 29385 2470
rect 29505 2350 29560 2470
rect 29680 2350 29705 2470
rect 24175 2295 29705 2350
rect 24175 2175 24200 2295
rect 24320 2175 24365 2295
rect 24485 2175 24530 2295
rect 24650 2175 24695 2295
rect 24815 2175 24870 2295
rect 24990 2175 25035 2295
rect 25155 2175 25200 2295
rect 25320 2175 25365 2295
rect 25485 2175 25540 2295
rect 25660 2175 25705 2295
rect 25825 2175 25870 2295
rect 25990 2175 26035 2295
rect 26155 2175 26210 2295
rect 26330 2175 26375 2295
rect 26495 2175 26540 2295
rect 26660 2175 26705 2295
rect 26825 2175 26880 2295
rect 27000 2175 27045 2295
rect 27165 2175 27210 2295
rect 27330 2175 27375 2295
rect 27495 2175 27550 2295
rect 27670 2175 27715 2295
rect 27835 2175 27880 2295
rect 28000 2175 28045 2295
rect 28165 2175 28220 2295
rect 28340 2175 28385 2295
rect 28505 2175 28550 2295
rect 28670 2175 28715 2295
rect 28835 2175 28890 2295
rect 29010 2175 29055 2295
rect 29175 2175 29220 2295
rect 29340 2175 29385 2295
rect 29505 2175 29560 2295
rect 29680 2175 29705 2295
rect 24175 2130 29705 2175
rect 24175 2010 24200 2130
rect 24320 2010 24365 2130
rect 24485 2010 24530 2130
rect 24650 2010 24695 2130
rect 24815 2010 24870 2130
rect 24990 2010 25035 2130
rect 25155 2010 25200 2130
rect 25320 2010 25365 2130
rect 25485 2010 25540 2130
rect 25660 2010 25705 2130
rect 25825 2010 25870 2130
rect 25990 2010 26035 2130
rect 26155 2010 26210 2130
rect 26330 2010 26375 2130
rect 26495 2010 26540 2130
rect 26660 2010 26705 2130
rect 26825 2010 26880 2130
rect 27000 2010 27045 2130
rect 27165 2010 27210 2130
rect 27330 2010 27375 2130
rect 27495 2010 27550 2130
rect 27670 2010 27715 2130
rect 27835 2010 27880 2130
rect 28000 2010 28045 2130
rect 28165 2010 28220 2130
rect 28340 2010 28385 2130
rect 28505 2010 28550 2130
rect 28670 2010 28715 2130
rect 28835 2010 28890 2130
rect 29010 2010 29055 2130
rect 29175 2010 29220 2130
rect 29340 2010 29385 2130
rect 29505 2010 29560 2130
rect 29680 2010 29705 2130
rect 24175 1965 29705 2010
rect 24175 1845 24200 1965
rect 24320 1845 24365 1965
rect 24485 1845 24530 1965
rect 24650 1845 24695 1965
rect 24815 1845 24870 1965
rect 24990 1845 25035 1965
rect 25155 1845 25200 1965
rect 25320 1845 25365 1965
rect 25485 1845 25540 1965
rect 25660 1845 25705 1965
rect 25825 1845 25870 1965
rect 25990 1845 26035 1965
rect 26155 1845 26210 1965
rect 26330 1845 26375 1965
rect 26495 1845 26540 1965
rect 26660 1845 26705 1965
rect 26825 1845 26880 1965
rect 27000 1845 27045 1965
rect 27165 1845 27210 1965
rect 27330 1845 27375 1965
rect 27495 1845 27550 1965
rect 27670 1845 27715 1965
rect 27835 1845 27880 1965
rect 28000 1845 28045 1965
rect 28165 1845 28220 1965
rect 28340 1845 28385 1965
rect 28505 1845 28550 1965
rect 28670 1845 28715 1965
rect 28835 1845 28890 1965
rect 29010 1845 29055 1965
rect 29175 1845 29220 1965
rect 29340 1845 29385 1965
rect 29505 1845 29560 1965
rect 29680 1845 29705 1965
rect 24175 1800 29705 1845
rect 24175 1680 24200 1800
rect 24320 1680 24365 1800
rect 24485 1680 24530 1800
rect 24650 1680 24695 1800
rect 24815 1680 24870 1800
rect 24990 1680 25035 1800
rect 25155 1680 25200 1800
rect 25320 1680 25365 1800
rect 25485 1680 25540 1800
rect 25660 1680 25705 1800
rect 25825 1680 25870 1800
rect 25990 1680 26035 1800
rect 26155 1680 26210 1800
rect 26330 1680 26375 1800
rect 26495 1680 26540 1800
rect 26660 1680 26705 1800
rect 26825 1680 26880 1800
rect 27000 1680 27045 1800
rect 27165 1680 27210 1800
rect 27330 1680 27375 1800
rect 27495 1680 27550 1800
rect 27670 1680 27715 1800
rect 27835 1680 27880 1800
rect 28000 1680 28045 1800
rect 28165 1680 28220 1800
rect 28340 1680 28385 1800
rect 28505 1680 28550 1800
rect 28670 1680 28715 1800
rect 28835 1680 28890 1800
rect 29010 1680 29055 1800
rect 29175 1680 29220 1800
rect 29340 1680 29385 1800
rect 29505 1680 29560 1800
rect 29680 1680 29705 1800
rect 24175 1610 29705 1680
rect 7105 1590 29705 1610
rect 7105 1470 7170 1590
rect 7290 1470 7335 1590
rect 7455 1470 7500 1590
rect 7620 1470 7665 1590
rect 7785 1470 7830 1590
rect 7950 1470 7995 1590
rect 8115 1470 8160 1590
rect 8280 1470 8325 1590
rect 8445 1470 8490 1590
rect 8610 1470 8655 1590
rect 8775 1470 8820 1590
rect 8940 1470 8985 1590
rect 9105 1470 9150 1590
rect 9270 1470 9315 1590
rect 9435 1470 9480 1590
rect 9600 1470 9645 1590
rect 9765 1470 9810 1590
rect 9930 1470 9975 1590
rect 10095 1470 10140 1590
rect 10260 1470 10305 1590
rect 10425 1470 10470 1590
rect 10590 1470 10635 1590
rect 10755 1470 10800 1590
rect 10920 1470 10965 1590
rect 11085 1470 11130 1590
rect 11250 1470 11295 1590
rect 11415 1470 11460 1590
rect 11580 1470 11625 1590
rect 11745 1470 11790 1590
rect 11910 1470 11955 1590
rect 12075 1470 12120 1590
rect 12240 1470 12285 1590
rect 12405 1470 12450 1590
rect 12570 1470 12860 1590
rect 12980 1470 13025 1590
rect 13145 1470 13190 1590
rect 13310 1470 13355 1590
rect 13475 1470 13520 1590
rect 13640 1470 13685 1590
rect 13805 1470 13850 1590
rect 13970 1470 14015 1590
rect 14135 1470 14180 1590
rect 14300 1470 14345 1590
rect 14465 1470 14510 1590
rect 14630 1470 14675 1590
rect 14795 1470 14840 1590
rect 14960 1470 15005 1590
rect 15125 1470 15170 1590
rect 15290 1470 15335 1590
rect 15455 1470 15500 1590
rect 15620 1470 15665 1590
rect 15785 1470 15830 1590
rect 15950 1470 15995 1590
rect 16115 1470 16160 1590
rect 16280 1470 16325 1590
rect 16445 1470 16490 1590
rect 16610 1470 16655 1590
rect 16775 1470 16820 1590
rect 16940 1470 16985 1590
rect 17105 1470 17150 1590
rect 17270 1470 17315 1590
rect 17435 1470 17480 1590
rect 17600 1470 17645 1590
rect 17765 1470 17810 1590
rect 17930 1470 17975 1590
rect 18095 1470 18140 1590
rect 18260 1470 18550 1590
rect 18670 1470 18715 1590
rect 18835 1470 18880 1590
rect 19000 1470 19045 1590
rect 19165 1470 19210 1590
rect 19330 1470 19375 1590
rect 19495 1470 19540 1590
rect 19660 1470 19705 1590
rect 19825 1470 19870 1590
rect 19990 1470 20035 1590
rect 20155 1470 20200 1590
rect 20320 1470 20365 1590
rect 20485 1470 20530 1590
rect 20650 1470 20695 1590
rect 20815 1470 20860 1590
rect 20980 1470 21025 1590
rect 21145 1470 21190 1590
rect 21310 1470 21355 1590
rect 21475 1470 21520 1590
rect 21640 1470 21685 1590
rect 21805 1470 21850 1590
rect 21970 1470 22015 1590
rect 22135 1470 22180 1590
rect 22300 1470 22345 1590
rect 22465 1470 22510 1590
rect 22630 1470 22675 1590
rect 22795 1470 22840 1590
rect 22960 1470 23005 1590
rect 23125 1470 23170 1590
rect 23290 1470 23335 1590
rect 23455 1470 23500 1590
rect 23620 1470 23665 1590
rect 23785 1470 23830 1590
rect 23950 1470 24240 1590
rect 24360 1470 24405 1590
rect 24525 1470 24570 1590
rect 24690 1470 24735 1590
rect 24855 1470 24900 1590
rect 25020 1470 25065 1590
rect 25185 1470 25230 1590
rect 25350 1470 25395 1590
rect 25515 1470 25560 1590
rect 25680 1470 25725 1590
rect 25845 1470 25890 1590
rect 26010 1470 26055 1590
rect 26175 1470 26220 1590
rect 26340 1470 26385 1590
rect 26505 1470 26550 1590
rect 26670 1470 26715 1590
rect 26835 1470 26880 1590
rect 27000 1470 27045 1590
rect 27165 1470 27210 1590
rect 27330 1470 27375 1590
rect 27495 1470 27540 1590
rect 27660 1470 27705 1590
rect 27825 1470 27870 1590
rect 27990 1470 28035 1590
rect 28155 1470 28200 1590
rect 28320 1470 28365 1590
rect 28485 1470 28530 1590
rect 28650 1470 28695 1590
rect 28815 1470 28860 1590
rect 28980 1470 29025 1590
rect 29145 1470 29190 1590
rect 29310 1470 29355 1590
rect 29475 1470 29520 1590
rect 29640 1470 29705 1590
rect 7105 1450 29705 1470
rect 7105 1380 12635 1450
rect 7105 1260 7130 1380
rect 7250 1260 7305 1380
rect 7425 1260 7470 1380
rect 7590 1260 7635 1380
rect 7755 1260 7800 1380
rect 7920 1260 7975 1380
rect 8095 1260 8140 1380
rect 8260 1260 8305 1380
rect 8425 1260 8470 1380
rect 8590 1260 8645 1380
rect 8765 1260 8810 1380
rect 8930 1260 8975 1380
rect 9095 1260 9140 1380
rect 9260 1260 9315 1380
rect 9435 1260 9480 1380
rect 9600 1260 9645 1380
rect 9765 1260 9810 1380
rect 9930 1260 9985 1380
rect 10105 1260 10150 1380
rect 10270 1260 10315 1380
rect 10435 1260 10480 1380
rect 10600 1260 10655 1380
rect 10775 1260 10820 1380
rect 10940 1260 10985 1380
rect 11105 1260 11150 1380
rect 11270 1260 11325 1380
rect 11445 1260 11490 1380
rect 11610 1260 11655 1380
rect 11775 1260 11820 1380
rect 11940 1260 11995 1380
rect 12115 1260 12160 1380
rect 12280 1260 12325 1380
rect 12445 1260 12490 1380
rect 12610 1260 12635 1380
rect 7105 1215 12635 1260
rect 7105 1095 7130 1215
rect 7250 1095 7305 1215
rect 7425 1095 7470 1215
rect 7590 1095 7635 1215
rect 7755 1095 7800 1215
rect 7920 1095 7975 1215
rect 8095 1095 8140 1215
rect 8260 1095 8305 1215
rect 8425 1095 8470 1215
rect 8590 1095 8645 1215
rect 8765 1095 8810 1215
rect 8930 1095 8975 1215
rect 9095 1095 9140 1215
rect 9260 1095 9315 1215
rect 9435 1095 9480 1215
rect 9600 1095 9645 1215
rect 9765 1095 9810 1215
rect 9930 1095 9985 1215
rect 10105 1095 10150 1215
rect 10270 1095 10315 1215
rect 10435 1095 10480 1215
rect 10600 1095 10655 1215
rect 10775 1095 10820 1215
rect 10940 1095 10985 1215
rect 11105 1095 11150 1215
rect 11270 1095 11325 1215
rect 11445 1095 11490 1215
rect 11610 1095 11655 1215
rect 11775 1095 11820 1215
rect 11940 1095 11995 1215
rect 12115 1095 12160 1215
rect 12280 1095 12325 1215
rect 12445 1095 12490 1215
rect 12610 1095 12635 1215
rect 7105 1050 12635 1095
rect 7105 930 7130 1050
rect 7250 930 7305 1050
rect 7425 930 7470 1050
rect 7590 930 7635 1050
rect 7755 930 7800 1050
rect 7920 930 7975 1050
rect 8095 930 8140 1050
rect 8260 930 8305 1050
rect 8425 930 8470 1050
rect 8590 930 8645 1050
rect 8765 930 8810 1050
rect 8930 930 8975 1050
rect 9095 930 9140 1050
rect 9260 930 9315 1050
rect 9435 930 9480 1050
rect 9600 930 9645 1050
rect 9765 930 9810 1050
rect 9930 930 9985 1050
rect 10105 930 10150 1050
rect 10270 930 10315 1050
rect 10435 930 10480 1050
rect 10600 930 10655 1050
rect 10775 930 10820 1050
rect 10940 930 10985 1050
rect 11105 930 11150 1050
rect 11270 930 11325 1050
rect 11445 930 11490 1050
rect 11610 930 11655 1050
rect 11775 930 11820 1050
rect 11940 930 11995 1050
rect 12115 930 12160 1050
rect 12280 930 12325 1050
rect 12445 930 12490 1050
rect 12610 930 12635 1050
rect 7105 885 12635 930
rect 7105 765 7130 885
rect 7250 765 7305 885
rect 7425 765 7470 885
rect 7590 765 7635 885
rect 7755 765 7800 885
rect 7920 765 7975 885
rect 8095 765 8140 885
rect 8260 765 8305 885
rect 8425 765 8470 885
rect 8590 765 8645 885
rect 8765 765 8810 885
rect 8930 765 8975 885
rect 9095 765 9140 885
rect 9260 765 9315 885
rect 9435 765 9480 885
rect 9600 765 9645 885
rect 9765 765 9810 885
rect 9930 765 9985 885
rect 10105 765 10150 885
rect 10270 765 10315 885
rect 10435 765 10480 885
rect 10600 765 10655 885
rect 10775 765 10820 885
rect 10940 765 10985 885
rect 11105 765 11150 885
rect 11270 765 11325 885
rect 11445 765 11490 885
rect 11610 765 11655 885
rect 11775 765 11820 885
rect 11940 765 11995 885
rect 12115 765 12160 885
rect 12280 765 12325 885
rect 12445 765 12490 885
rect 12610 765 12635 885
rect 7105 710 12635 765
rect 7105 590 7130 710
rect 7250 590 7305 710
rect 7425 590 7470 710
rect 7590 590 7635 710
rect 7755 590 7800 710
rect 7920 590 7975 710
rect 8095 590 8140 710
rect 8260 590 8305 710
rect 8425 590 8470 710
rect 8590 590 8645 710
rect 8765 590 8810 710
rect 8930 590 8975 710
rect 9095 590 9140 710
rect 9260 590 9315 710
rect 9435 590 9480 710
rect 9600 590 9645 710
rect 9765 590 9810 710
rect 9930 590 9985 710
rect 10105 590 10150 710
rect 10270 590 10315 710
rect 10435 590 10480 710
rect 10600 590 10655 710
rect 10775 590 10820 710
rect 10940 590 10985 710
rect 11105 590 11150 710
rect 11270 590 11325 710
rect 11445 590 11490 710
rect 11610 590 11655 710
rect 11775 590 11820 710
rect 11940 590 11995 710
rect 12115 590 12160 710
rect 12280 590 12325 710
rect 12445 590 12490 710
rect 12610 590 12635 710
rect 7105 545 12635 590
rect 7105 425 7130 545
rect 7250 425 7305 545
rect 7425 425 7470 545
rect 7590 425 7635 545
rect 7755 425 7800 545
rect 7920 425 7975 545
rect 8095 425 8140 545
rect 8260 425 8305 545
rect 8425 425 8470 545
rect 8590 425 8645 545
rect 8765 425 8810 545
rect 8930 425 8975 545
rect 9095 425 9140 545
rect 9260 425 9315 545
rect 9435 425 9480 545
rect 9600 425 9645 545
rect 9765 425 9810 545
rect 9930 425 9985 545
rect 10105 425 10150 545
rect 10270 425 10315 545
rect 10435 425 10480 545
rect 10600 425 10655 545
rect 10775 425 10820 545
rect 10940 425 10985 545
rect 11105 425 11150 545
rect 11270 425 11325 545
rect 11445 425 11490 545
rect 11610 425 11655 545
rect 11775 425 11820 545
rect 11940 425 11995 545
rect 12115 425 12160 545
rect 12280 425 12325 545
rect 12445 425 12490 545
rect 12610 425 12635 545
rect 7105 380 12635 425
rect 7105 260 7130 380
rect 7250 260 7305 380
rect 7425 260 7470 380
rect 7590 260 7635 380
rect 7755 260 7800 380
rect 7920 260 7975 380
rect 8095 260 8140 380
rect 8260 260 8305 380
rect 8425 260 8470 380
rect 8590 260 8645 380
rect 8765 260 8810 380
rect 8930 260 8975 380
rect 9095 260 9140 380
rect 9260 260 9315 380
rect 9435 260 9480 380
rect 9600 260 9645 380
rect 9765 260 9810 380
rect 9930 260 9985 380
rect 10105 260 10150 380
rect 10270 260 10315 380
rect 10435 260 10480 380
rect 10600 260 10655 380
rect 10775 260 10820 380
rect 10940 260 10985 380
rect 11105 260 11150 380
rect 11270 260 11325 380
rect 11445 260 11490 380
rect 11610 260 11655 380
rect 11775 260 11820 380
rect 11940 260 11995 380
rect 12115 260 12160 380
rect 12280 260 12325 380
rect 12445 260 12490 380
rect 12610 260 12635 380
rect 7105 215 12635 260
rect 7105 95 7130 215
rect 7250 95 7305 215
rect 7425 95 7470 215
rect 7590 95 7635 215
rect 7755 95 7800 215
rect 7920 95 7975 215
rect 8095 95 8140 215
rect 8260 95 8305 215
rect 8425 95 8470 215
rect 8590 95 8645 215
rect 8765 95 8810 215
rect 8930 95 8975 215
rect 9095 95 9140 215
rect 9260 95 9315 215
rect 9435 95 9480 215
rect 9600 95 9645 215
rect 9765 95 9810 215
rect 9930 95 9985 215
rect 10105 95 10150 215
rect 10270 95 10315 215
rect 10435 95 10480 215
rect 10600 95 10655 215
rect 10775 95 10820 215
rect 10940 95 10985 215
rect 11105 95 11150 215
rect 11270 95 11325 215
rect 11445 95 11490 215
rect 11610 95 11655 215
rect 11775 95 11820 215
rect 11940 95 11995 215
rect 12115 95 12160 215
rect 12280 95 12325 215
rect 12445 95 12490 215
rect 12610 95 12635 215
rect 7105 40 12635 95
rect 7105 -80 7130 40
rect 7250 -80 7305 40
rect 7425 -80 7470 40
rect 7590 -80 7635 40
rect 7755 -80 7800 40
rect 7920 -80 7975 40
rect 8095 -80 8140 40
rect 8260 -80 8305 40
rect 8425 -80 8470 40
rect 8590 -80 8645 40
rect 8765 -80 8810 40
rect 8930 -80 8975 40
rect 9095 -80 9140 40
rect 9260 -80 9315 40
rect 9435 -80 9480 40
rect 9600 -80 9645 40
rect 9765 -80 9810 40
rect 9930 -80 9985 40
rect 10105 -80 10150 40
rect 10270 -80 10315 40
rect 10435 -80 10480 40
rect 10600 -80 10655 40
rect 10775 -80 10820 40
rect 10940 -80 10985 40
rect 11105 -80 11150 40
rect 11270 -80 11325 40
rect 11445 -80 11490 40
rect 11610 -80 11655 40
rect 11775 -80 11820 40
rect 11940 -80 11995 40
rect 12115 -80 12160 40
rect 12280 -80 12325 40
rect 12445 -80 12490 40
rect 12610 -80 12635 40
rect 7105 -125 12635 -80
rect 7105 -245 7130 -125
rect 7250 -245 7305 -125
rect 7425 -245 7470 -125
rect 7590 -245 7635 -125
rect 7755 -245 7800 -125
rect 7920 -245 7975 -125
rect 8095 -245 8140 -125
rect 8260 -245 8305 -125
rect 8425 -245 8470 -125
rect 8590 -245 8645 -125
rect 8765 -245 8810 -125
rect 8930 -245 8975 -125
rect 9095 -245 9140 -125
rect 9260 -245 9315 -125
rect 9435 -245 9480 -125
rect 9600 -245 9645 -125
rect 9765 -245 9810 -125
rect 9930 -245 9985 -125
rect 10105 -245 10150 -125
rect 10270 -245 10315 -125
rect 10435 -245 10480 -125
rect 10600 -245 10655 -125
rect 10775 -245 10820 -125
rect 10940 -245 10985 -125
rect 11105 -245 11150 -125
rect 11270 -245 11325 -125
rect 11445 -245 11490 -125
rect 11610 -245 11655 -125
rect 11775 -245 11820 -125
rect 11940 -245 11995 -125
rect 12115 -245 12160 -125
rect 12280 -245 12325 -125
rect 12445 -245 12490 -125
rect 12610 -245 12635 -125
rect 7105 -290 12635 -245
rect 7105 -410 7130 -290
rect 7250 -410 7305 -290
rect 7425 -410 7470 -290
rect 7590 -410 7635 -290
rect 7755 -410 7800 -290
rect 7920 -410 7975 -290
rect 8095 -410 8140 -290
rect 8260 -410 8305 -290
rect 8425 -410 8470 -290
rect 8590 -410 8645 -290
rect 8765 -410 8810 -290
rect 8930 -410 8975 -290
rect 9095 -410 9140 -290
rect 9260 -410 9315 -290
rect 9435 -410 9480 -290
rect 9600 -410 9645 -290
rect 9765 -410 9810 -290
rect 9930 -410 9985 -290
rect 10105 -410 10150 -290
rect 10270 -410 10315 -290
rect 10435 -410 10480 -290
rect 10600 -410 10655 -290
rect 10775 -410 10820 -290
rect 10940 -410 10985 -290
rect 11105 -410 11150 -290
rect 11270 -410 11325 -290
rect 11445 -410 11490 -290
rect 11610 -410 11655 -290
rect 11775 -410 11820 -290
rect 11940 -410 11995 -290
rect 12115 -410 12160 -290
rect 12280 -410 12325 -290
rect 12445 -410 12490 -290
rect 12610 -410 12635 -290
rect 7105 -455 12635 -410
rect 7105 -575 7130 -455
rect 7250 -575 7305 -455
rect 7425 -575 7470 -455
rect 7590 -575 7635 -455
rect 7755 -575 7800 -455
rect 7920 -575 7975 -455
rect 8095 -575 8140 -455
rect 8260 -575 8305 -455
rect 8425 -575 8470 -455
rect 8590 -575 8645 -455
rect 8765 -575 8810 -455
rect 8930 -575 8975 -455
rect 9095 -575 9140 -455
rect 9260 -575 9315 -455
rect 9435 -575 9480 -455
rect 9600 -575 9645 -455
rect 9765 -575 9810 -455
rect 9930 -575 9985 -455
rect 10105 -575 10150 -455
rect 10270 -575 10315 -455
rect 10435 -575 10480 -455
rect 10600 -575 10655 -455
rect 10775 -575 10820 -455
rect 10940 -575 10985 -455
rect 11105 -575 11150 -455
rect 11270 -575 11325 -455
rect 11445 -575 11490 -455
rect 11610 -575 11655 -455
rect 11775 -575 11820 -455
rect 11940 -575 11995 -455
rect 12115 -575 12160 -455
rect 12280 -575 12325 -455
rect 12445 -575 12490 -455
rect 12610 -575 12635 -455
rect 7105 -630 12635 -575
rect 7105 -750 7130 -630
rect 7250 -750 7305 -630
rect 7425 -750 7470 -630
rect 7590 -750 7635 -630
rect 7755 -750 7800 -630
rect 7920 -750 7975 -630
rect 8095 -750 8140 -630
rect 8260 -750 8305 -630
rect 8425 -750 8470 -630
rect 8590 -750 8645 -630
rect 8765 -750 8810 -630
rect 8930 -750 8975 -630
rect 9095 -750 9140 -630
rect 9260 -750 9315 -630
rect 9435 -750 9480 -630
rect 9600 -750 9645 -630
rect 9765 -750 9810 -630
rect 9930 -750 9985 -630
rect 10105 -750 10150 -630
rect 10270 -750 10315 -630
rect 10435 -750 10480 -630
rect 10600 -750 10655 -630
rect 10775 -750 10820 -630
rect 10940 -750 10985 -630
rect 11105 -750 11150 -630
rect 11270 -750 11325 -630
rect 11445 -750 11490 -630
rect 11610 -750 11655 -630
rect 11775 -750 11820 -630
rect 11940 -750 11995 -630
rect 12115 -750 12160 -630
rect 12280 -750 12325 -630
rect 12445 -750 12490 -630
rect 12610 -750 12635 -630
rect 7105 -795 12635 -750
rect 7105 -915 7130 -795
rect 7250 -915 7305 -795
rect 7425 -915 7470 -795
rect 7590 -915 7635 -795
rect 7755 -915 7800 -795
rect 7920 -915 7975 -795
rect 8095 -915 8140 -795
rect 8260 -915 8305 -795
rect 8425 -915 8470 -795
rect 8590 -915 8645 -795
rect 8765 -915 8810 -795
rect 8930 -915 8975 -795
rect 9095 -915 9140 -795
rect 9260 -915 9315 -795
rect 9435 -915 9480 -795
rect 9600 -915 9645 -795
rect 9765 -915 9810 -795
rect 9930 -915 9985 -795
rect 10105 -915 10150 -795
rect 10270 -915 10315 -795
rect 10435 -915 10480 -795
rect 10600 -915 10655 -795
rect 10775 -915 10820 -795
rect 10940 -915 10985 -795
rect 11105 -915 11150 -795
rect 11270 -915 11325 -795
rect 11445 -915 11490 -795
rect 11610 -915 11655 -795
rect 11775 -915 11820 -795
rect 11940 -915 11995 -795
rect 12115 -915 12160 -795
rect 12280 -915 12325 -795
rect 12445 -915 12490 -795
rect 12610 -915 12635 -795
rect 7105 -960 12635 -915
rect 7105 -1080 7130 -960
rect 7250 -1080 7305 -960
rect 7425 -1080 7470 -960
rect 7590 -1080 7635 -960
rect 7755 -1080 7800 -960
rect 7920 -1080 7975 -960
rect 8095 -1080 8140 -960
rect 8260 -1080 8305 -960
rect 8425 -1080 8470 -960
rect 8590 -1080 8645 -960
rect 8765 -1080 8810 -960
rect 8930 -1080 8975 -960
rect 9095 -1080 9140 -960
rect 9260 -1080 9315 -960
rect 9435 -1080 9480 -960
rect 9600 -1080 9645 -960
rect 9765 -1080 9810 -960
rect 9930 -1080 9985 -960
rect 10105 -1080 10150 -960
rect 10270 -1080 10315 -960
rect 10435 -1080 10480 -960
rect 10600 -1080 10655 -960
rect 10775 -1080 10820 -960
rect 10940 -1080 10985 -960
rect 11105 -1080 11150 -960
rect 11270 -1080 11325 -960
rect 11445 -1080 11490 -960
rect 11610 -1080 11655 -960
rect 11775 -1080 11820 -960
rect 11940 -1080 11995 -960
rect 12115 -1080 12160 -960
rect 12280 -1080 12325 -960
rect 12445 -1080 12490 -960
rect 12610 -1080 12635 -960
rect 7105 -1125 12635 -1080
rect 7105 -1245 7130 -1125
rect 7250 -1245 7305 -1125
rect 7425 -1245 7470 -1125
rect 7590 -1245 7635 -1125
rect 7755 -1245 7800 -1125
rect 7920 -1245 7975 -1125
rect 8095 -1245 8140 -1125
rect 8260 -1245 8305 -1125
rect 8425 -1245 8470 -1125
rect 8590 -1245 8645 -1125
rect 8765 -1245 8810 -1125
rect 8930 -1245 8975 -1125
rect 9095 -1245 9140 -1125
rect 9260 -1245 9315 -1125
rect 9435 -1245 9480 -1125
rect 9600 -1245 9645 -1125
rect 9765 -1245 9810 -1125
rect 9930 -1245 9985 -1125
rect 10105 -1245 10150 -1125
rect 10270 -1245 10315 -1125
rect 10435 -1245 10480 -1125
rect 10600 -1245 10655 -1125
rect 10775 -1245 10820 -1125
rect 10940 -1245 10985 -1125
rect 11105 -1245 11150 -1125
rect 11270 -1245 11325 -1125
rect 11445 -1245 11490 -1125
rect 11610 -1245 11655 -1125
rect 11775 -1245 11820 -1125
rect 11940 -1245 11995 -1125
rect 12115 -1245 12160 -1125
rect 12280 -1245 12325 -1125
rect 12445 -1245 12490 -1125
rect 12610 -1245 12635 -1125
rect 7105 -1300 12635 -1245
rect 7105 -1420 7130 -1300
rect 7250 -1420 7305 -1300
rect 7425 -1420 7470 -1300
rect 7590 -1420 7635 -1300
rect 7755 -1420 7800 -1300
rect 7920 -1420 7975 -1300
rect 8095 -1420 8140 -1300
rect 8260 -1420 8305 -1300
rect 8425 -1420 8470 -1300
rect 8590 -1420 8645 -1300
rect 8765 -1420 8810 -1300
rect 8930 -1420 8975 -1300
rect 9095 -1420 9140 -1300
rect 9260 -1420 9315 -1300
rect 9435 -1420 9480 -1300
rect 9600 -1420 9645 -1300
rect 9765 -1420 9810 -1300
rect 9930 -1420 9985 -1300
rect 10105 -1420 10150 -1300
rect 10270 -1420 10315 -1300
rect 10435 -1420 10480 -1300
rect 10600 -1420 10655 -1300
rect 10775 -1420 10820 -1300
rect 10940 -1420 10985 -1300
rect 11105 -1420 11150 -1300
rect 11270 -1420 11325 -1300
rect 11445 -1420 11490 -1300
rect 11610 -1420 11655 -1300
rect 11775 -1420 11820 -1300
rect 11940 -1420 11995 -1300
rect 12115 -1420 12160 -1300
rect 12280 -1420 12325 -1300
rect 12445 -1420 12490 -1300
rect 12610 -1420 12635 -1300
rect 7105 -1465 12635 -1420
rect 7105 -1585 7130 -1465
rect 7250 -1585 7305 -1465
rect 7425 -1585 7470 -1465
rect 7590 -1585 7635 -1465
rect 7755 -1585 7800 -1465
rect 7920 -1585 7975 -1465
rect 8095 -1585 8140 -1465
rect 8260 -1585 8305 -1465
rect 8425 -1585 8470 -1465
rect 8590 -1585 8645 -1465
rect 8765 -1585 8810 -1465
rect 8930 -1585 8975 -1465
rect 9095 -1585 9140 -1465
rect 9260 -1585 9315 -1465
rect 9435 -1585 9480 -1465
rect 9600 -1585 9645 -1465
rect 9765 -1585 9810 -1465
rect 9930 -1585 9985 -1465
rect 10105 -1585 10150 -1465
rect 10270 -1585 10315 -1465
rect 10435 -1585 10480 -1465
rect 10600 -1585 10655 -1465
rect 10775 -1585 10820 -1465
rect 10940 -1585 10985 -1465
rect 11105 -1585 11150 -1465
rect 11270 -1585 11325 -1465
rect 11445 -1585 11490 -1465
rect 11610 -1585 11655 -1465
rect 11775 -1585 11820 -1465
rect 11940 -1585 11995 -1465
rect 12115 -1585 12160 -1465
rect 12280 -1585 12325 -1465
rect 12445 -1585 12490 -1465
rect 12610 -1585 12635 -1465
rect 7105 -1630 12635 -1585
rect 7105 -1750 7130 -1630
rect 7250 -1750 7305 -1630
rect 7425 -1750 7470 -1630
rect 7590 -1750 7635 -1630
rect 7755 -1750 7800 -1630
rect 7920 -1750 7975 -1630
rect 8095 -1750 8140 -1630
rect 8260 -1750 8305 -1630
rect 8425 -1750 8470 -1630
rect 8590 -1750 8645 -1630
rect 8765 -1750 8810 -1630
rect 8930 -1750 8975 -1630
rect 9095 -1750 9140 -1630
rect 9260 -1750 9315 -1630
rect 9435 -1750 9480 -1630
rect 9600 -1750 9645 -1630
rect 9765 -1750 9810 -1630
rect 9930 -1750 9985 -1630
rect 10105 -1750 10150 -1630
rect 10270 -1750 10315 -1630
rect 10435 -1750 10480 -1630
rect 10600 -1750 10655 -1630
rect 10775 -1750 10820 -1630
rect 10940 -1750 10985 -1630
rect 11105 -1750 11150 -1630
rect 11270 -1750 11325 -1630
rect 11445 -1750 11490 -1630
rect 11610 -1750 11655 -1630
rect 11775 -1750 11820 -1630
rect 11940 -1750 11995 -1630
rect 12115 -1750 12160 -1630
rect 12280 -1750 12325 -1630
rect 12445 -1750 12490 -1630
rect 12610 -1750 12635 -1630
rect 7105 -1795 12635 -1750
rect 7105 -1915 7130 -1795
rect 7250 -1915 7305 -1795
rect 7425 -1915 7470 -1795
rect 7590 -1915 7635 -1795
rect 7755 -1915 7800 -1795
rect 7920 -1915 7975 -1795
rect 8095 -1915 8140 -1795
rect 8260 -1915 8305 -1795
rect 8425 -1915 8470 -1795
rect 8590 -1915 8645 -1795
rect 8765 -1915 8810 -1795
rect 8930 -1915 8975 -1795
rect 9095 -1915 9140 -1795
rect 9260 -1915 9315 -1795
rect 9435 -1915 9480 -1795
rect 9600 -1915 9645 -1795
rect 9765 -1915 9810 -1795
rect 9930 -1915 9985 -1795
rect 10105 -1915 10150 -1795
rect 10270 -1915 10315 -1795
rect 10435 -1915 10480 -1795
rect 10600 -1915 10655 -1795
rect 10775 -1915 10820 -1795
rect 10940 -1915 10985 -1795
rect 11105 -1915 11150 -1795
rect 11270 -1915 11325 -1795
rect 11445 -1915 11490 -1795
rect 11610 -1915 11655 -1795
rect 11775 -1915 11820 -1795
rect 11940 -1915 11995 -1795
rect 12115 -1915 12160 -1795
rect 12280 -1915 12325 -1795
rect 12445 -1915 12490 -1795
rect 12610 -1915 12635 -1795
rect 7105 -1970 12635 -1915
rect 7105 -2090 7130 -1970
rect 7250 -2090 7305 -1970
rect 7425 -2090 7470 -1970
rect 7590 -2090 7635 -1970
rect 7755 -2090 7800 -1970
rect 7920 -2090 7975 -1970
rect 8095 -2090 8140 -1970
rect 8260 -2090 8305 -1970
rect 8425 -2090 8470 -1970
rect 8590 -2090 8645 -1970
rect 8765 -2090 8810 -1970
rect 8930 -2090 8975 -1970
rect 9095 -2090 9140 -1970
rect 9260 -2090 9315 -1970
rect 9435 -2090 9480 -1970
rect 9600 -2090 9645 -1970
rect 9765 -2090 9810 -1970
rect 9930 -2090 9985 -1970
rect 10105 -2090 10150 -1970
rect 10270 -2090 10315 -1970
rect 10435 -2090 10480 -1970
rect 10600 -2090 10655 -1970
rect 10775 -2090 10820 -1970
rect 10940 -2090 10985 -1970
rect 11105 -2090 11150 -1970
rect 11270 -2090 11325 -1970
rect 11445 -2090 11490 -1970
rect 11610 -2090 11655 -1970
rect 11775 -2090 11820 -1970
rect 11940 -2090 11995 -1970
rect 12115 -2090 12160 -1970
rect 12280 -2090 12325 -1970
rect 12445 -2090 12490 -1970
rect 12610 -2090 12635 -1970
rect 7105 -2135 12635 -2090
rect 7105 -2255 7130 -2135
rect 7250 -2255 7305 -2135
rect 7425 -2255 7470 -2135
rect 7590 -2255 7635 -2135
rect 7755 -2255 7800 -2135
rect 7920 -2255 7975 -2135
rect 8095 -2255 8140 -2135
rect 8260 -2255 8305 -2135
rect 8425 -2255 8470 -2135
rect 8590 -2255 8645 -2135
rect 8765 -2255 8810 -2135
rect 8930 -2255 8975 -2135
rect 9095 -2255 9140 -2135
rect 9260 -2255 9315 -2135
rect 9435 -2255 9480 -2135
rect 9600 -2255 9645 -2135
rect 9765 -2255 9810 -2135
rect 9930 -2255 9985 -2135
rect 10105 -2255 10150 -2135
rect 10270 -2255 10315 -2135
rect 10435 -2255 10480 -2135
rect 10600 -2255 10655 -2135
rect 10775 -2255 10820 -2135
rect 10940 -2255 10985 -2135
rect 11105 -2255 11150 -2135
rect 11270 -2255 11325 -2135
rect 11445 -2255 11490 -2135
rect 11610 -2255 11655 -2135
rect 11775 -2255 11820 -2135
rect 11940 -2255 11995 -2135
rect 12115 -2255 12160 -2135
rect 12280 -2255 12325 -2135
rect 12445 -2255 12490 -2135
rect 12610 -2255 12635 -2135
rect 7105 -2300 12635 -2255
rect 7105 -2420 7130 -2300
rect 7250 -2420 7305 -2300
rect 7425 -2420 7470 -2300
rect 7590 -2420 7635 -2300
rect 7755 -2420 7800 -2300
rect 7920 -2420 7975 -2300
rect 8095 -2420 8140 -2300
rect 8260 -2420 8305 -2300
rect 8425 -2420 8470 -2300
rect 8590 -2420 8645 -2300
rect 8765 -2420 8810 -2300
rect 8930 -2420 8975 -2300
rect 9095 -2420 9140 -2300
rect 9260 -2420 9315 -2300
rect 9435 -2420 9480 -2300
rect 9600 -2420 9645 -2300
rect 9765 -2420 9810 -2300
rect 9930 -2420 9985 -2300
rect 10105 -2420 10150 -2300
rect 10270 -2420 10315 -2300
rect 10435 -2420 10480 -2300
rect 10600 -2420 10655 -2300
rect 10775 -2420 10820 -2300
rect 10940 -2420 10985 -2300
rect 11105 -2420 11150 -2300
rect 11270 -2420 11325 -2300
rect 11445 -2420 11490 -2300
rect 11610 -2420 11655 -2300
rect 11775 -2420 11820 -2300
rect 11940 -2420 11995 -2300
rect 12115 -2420 12160 -2300
rect 12280 -2420 12325 -2300
rect 12445 -2420 12490 -2300
rect 12610 -2420 12635 -2300
rect 7105 -2465 12635 -2420
rect 7105 -2585 7130 -2465
rect 7250 -2585 7305 -2465
rect 7425 -2585 7470 -2465
rect 7590 -2585 7635 -2465
rect 7755 -2585 7800 -2465
rect 7920 -2585 7975 -2465
rect 8095 -2585 8140 -2465
rect 8260 -2585 8305 -2465
rect 8425 -2585 8470 -2465
rect 8590 -2585 8645 -2465
rect 8765 -2585 8810 -2465
rect 8930 -2585 8975 -2465
rect 9095 -2585 9140 -2465
rect 9260 -2585 9315 -2465
rect 9435 -2585 9480 -2465
rect 9600 -2585 9645 -2465
rect 9765 -2585 9810 -2465
rect 9930 -2585 9985 -2465
rect 10105 -2585 10150 -2465
rect 10270 -2585 10315 -2465
rect 10435 -2585 10480 -2465
rect 10600 -2585 10655 -2465
rect 10775 -2585 10820 -2465
rect 10940 -2585 10985 -2465
rect 11105 -2585 11150 -2465
rect 11270 -2585 11325 -2465
rect 11445 -2585 11490 -2465
rect 11610 -2585 11655 -2465
rect 11775 -2585 11820 -2465
rect 11940 -2585 11995 -2465
rect 12115 -2585 12160 -2465
rect 12280 -2585 12325 -2465
rect 12445 -2585 12490 -2465
rect 12610 -2585 12635 -2465
rect 7105 -2640 12635 -2585
rect 7105 -2760 7130 -2640
rect 7250 -2760 7305 -2640
rect 7425 -2760 7470 -2640
rect 7590 -2760 7635 -2640
rect 7755 -2760 7800 -2640
rect 7920 -2760 7975 -2640
rect 8095 -2760 8140 -2640
rect 8260 -2760 8305 -2640
rect 8425 -2760 8470 -2640
rect 8590 -2760 8645 -2640
rect 8765 -2760 8810 -2640
rect 8930 -2760 8975 -2640
rect 9095 -2760 9140 -2640
rect 9260 -2760 9315 -2640
rect 9435 -2760 9480 -2640
rect 9600 -2760 9645 -2640
rect 9765 -2760 9810 -2640
rect 9930 -2760 9985 -2640
rect 10105 -2760 10150 -2640
rect 10270 -2760 10315 -2640
rect 10435 -2760 10480 -2640
rect 10600 -2760 10655 -2640
rect 10775 -2760 10820 -2640
rect 10940 -2760 10985 -2640
rect 11105 -2760 11150 -2640
rect 11270 -2760 11325 -2640
rect 11445 -2760 11490 -2640
rect 11610 -2760 11655 -2640
rect 11775 -2760 11820 -2640
rect 11940 -2760 11995 -2640
rect 12115 -2760 12160 -2640
rect 12280 -2760 12325 -2640
rect 12445 -2760 12490 -2640
rect 12610 -2760 12635 -2640
rect 7105 -2805 12635 -2760
rect 7105 -2925 7130 -2805
rect 7250 -2925 7305 -2805
rect 7425 -2925 7470 -2805
rect 7590 -2925 7635 -2805
rect 7755 -2925 7800 -2805
rect 7920 -2925 7975 -2805
rect 8095 -2925 8140 -2805
rect 8260 -2925 8305 -2805
rect 8425 -2925 8470 -2805
rect 8590 -2925 8645 -2805
rect 8765 -2925 8810 -2805
rect 8930 -2925 8975 -2805
rect 9095 -2925 9140 -2805
rect 9260 -2925 9315 -2805
rect 9435 -2925 9480 -2805
rect 9600 -2925 9645 -2805
rect 9765 -2925 9810 -2805
rect 9930 -2925 9985 -2805
rect 10105 -2925 10150 -2805
rect 10270 -2925 10315 -2805
rect 10435 -2925 10480 -2805
rect 10600 -2925 10655 -2805
rect 10775 -2925 10820 -2805
rect 10940 -2925 10985 -2805
rect 11105 -2925 11150 -2805
rect 11270 -2925 11325 -2805
rect 11445 -2925 11490 -2805
rect 11610 -2925 11655 -2805
rect 11775 -2925 11820 -2805
rect 11940 -2925 11995 -2805
rect 12115 -2925 12160 -2805
rect 12280 -2925 12325 -2805
rect 12445 -2925 12490 -2805
rect 12610 -2925 12635 -2805
rect 7105 -2970 12635 -2925
rect 7105 -3090 7130 -2970
rect 7250 -3090 7305 -2970
rect 7425 -3090 7470 -2970
rect 7590 -3090 7635 -2970
rect 7755 -3090 7800 -2970
rect 7920 -3090 7975 -2970
rect 8095 -3090 8140 -2970
rect 8260 -3090 8305 -2970
rect 8425 -3090 8470 -2970
rect 8590 -3090 8645 -2970
rect 8765 -3090 8810 -2970
rect 8930 -3090 8975 -2970
rect 9095 -3090 9140 -2970
rect 9260 -3090 9315 -2970
rect 9435 -3090 9480 -2970
rect 9600 -3090 9645 -2970
rect 9765 -3090 9810 -2970
rect 9930 -3090 9985 -2970
rect 10105 -3090 10150 -2970
rect 10270 -3090 10315 -2970
rect 10435 -3090 10480 -2970
rect 10600 -3090 10655 -2970
rect 10775 -3090 10820 -2970
rect 10940 -3090 10985 -2970
rect 11105 -3090 11150 -2970
rect 11270 -3090 11325 -2970
rect 11445 -3090 11490 -2970
rect 11610 -3090 11655 -2970
rect 11775 -3090 11820 -2970
rect 11940 -3090 11995 -2970
rect 12115 -3090 12160 -2970
rect 12280 -3090 12325 -2970
rect 12445 -3090 12490 -2970
rect 12610 -3090 12635 -2970
rect 7105 -3135 12635 -3090
rect 7105 -3255 7130 -3135
rect 7250 -3255 7305 -3135
rect 7425 -3255 7470 -3135
rect 7590 -3255 7635 -3135
rect 7755 -3255 7800 -3135
rect 7920 -3255 7975 -3135
rect 8095 -3255 8140 -3135
rect 8260 -3255 8305 -3135
rect 8425 -3255 8470 -3135
rect 8590 -3255 8645 -3135
rect 8765 -3255 8810 -3135
rect 8930 -3255 8975 -3135
rect 9095 -3255 9140 -3135
rect 9260 -3255 9315 -3135
rect 9435 -3255 9480 -3135
rect 9600 -3255 9645 -3135
rect 9765 -3255 9810 -3135
rect 9930 -3255 9985 -3135
rect 10105 -3255 10150 -3135
rect 10270 -3255 10315 -3135
rect 10435 -3255 10480 -3135
rect 10600 -3255 10655 -3135
rect 10775 -3255 10820 -3135
rect 10940 -3255 10985 -3135
rect 11105 -3255 11150 -3135
rect 11270 -3255 11325 -3135
rect 11445 -3255 11490 -3135
rect 11610 -3255 11655 -3135
rect 11775 -3255 11820 -3135
rect 11940 -3255 11995 -3135
rect 12115 -3255 12160 -3135
rect 12280 -3255 12325 -3135
rect 12445 -3255 12490 -3135
rect 12610 -3255 12635 -3135
rect 7105 -3310 12635 -3255
rect 7105 -3430 7130 -3310
rect 7250 -3430 7305 -3310
rect 7425 -3430 7470 -3310
rect 7590 -3430 7635 -3310
rect 7755 -3430 7800 -3310
rect 7920 -3430 7975 -3310
rect 8095 -3430 8140 -3310
rect 8260 -3430 8305 -3310
rect 8425 -3430 8470 -3310
rect 8590 -3430 8645 -3310
rect 8765 -3430 8810 -3310
rect 8930 -3430 8975 -3310
rect 9095 -3430 9140 -3310
rect 9260 -3430 9315 -3310
rect 9435 -3430 9480 -3310
rect 9600 -3430 9645 -3310
rect 9765 -3430 9810 -3310
rect 9930 -3430 9985 -3310
rect 10105 -3430 10150 -3310
rect 10270 -3430 10315 -3310
rect 10435 -3430 10480 -3310
rect 10600 -3430 10655 -3310
rect 10775 -3430 10820 -3310
rect 10940 -3430 10985 -3310
rect 11105 -3430 11150 -3310
rect 11270 -3430 11325 -3310
rect 11445 -3430 11490 -3310
rect 11610 -3430 11655 -3310
rect 11775 -3430 11820 -3310
rect 11940 -3430 11995 -3310
rect 12115 -3430 12160 -3310
rect 12280 -3430 12325 -3310
rect 12445 -3430 12490 -3310
rect 12610 -3430 12635 -3310
rect 7105 -3475 12635 -3430
rect 7105 -3595 7130 -3475
rect 7250 -3595 7305 -3475
rect 7425 -3595 7470 -3475
rect 7590 -3595 7635 -3475
rect 7755 -3595 7800 -3475
rect 7920 -3595 7975 -3475
rect 8095 -3595 8140 -3475
rect 8260 -3595 8305 -3475
rect 8425 -3595 8470 -3475
rect 8590 -3595 8645 -3475
rect 8765 -3595 8810 -3475
rect 8930 -3595 8975 -3475
rect 9095 -3595 9140 -3475
rect 9260 -3595 9315 -3475
rect 9435 -3595 9480 -3475
rect 9600 -3595 9645 -3475
rect 9765 -3595 9810 -3475
rect 9930 -3595 9985 -3475
rect 10105 -3595 10150 -3475
rect 10270 -3595 10315 -3475
rect 10435 -3595 10480 -3475
rect 10600 -3595 10655 -3475
rect 10775 -3595 10820 -3475
rect 10940 -3595 10985 -3475
rect 11105 -3595 11150 -3475
rect 11270 -3595 11325 -3475
rect 11445 -3595 11490 -3475
rect 11610 -3595 11655 -3475
rect 11775 -3595 11820 -3475
rect 11940 -3595 11995 -3475
rect 12115 -3595 12160 -3475
rect 12280 -3595 12325 -3475
rect 12445 -3595 12490 -3475
rect 12610 -3595 12635 -3475
rect 7105 -3640 12635 -3595
rect 7105 -3760 7130 -3640
rect 7250 -3760 7305 -3640
rect 7425 -3760 7470 -3640
rect 7590 -3760 7635 -3640
rect 7755 -3760 7800 -3640
rect 7920 -3760 7975 -3640
rect 8095 -3760 8140 -3640
rect 8260 -3760 8305 -3640
rect 8425 -3760 8470 -3640
rect 8590 -3760 8645 -3640
rect 8765 -3760 8810 -3640
rect 8930 -3760 8975 -3640
rect 9095 -3760 9140 -3640
rect 9260 -3760 9315 -3640
rect 9435 -3760 9480 -3640
rect 9600 -3760 9645 -3640
rect 9765 -3760 9810 -3640
rect 9930 -3760 9985 -3640
rect 10105 -3760 10150 -3640
rect 10270 -3760 10315 -3640
rect 10435 -3760 10480 -3640
rect 10600 -3760 10655 -3640
rect 10775 -3760 10820 -3640
rect 10940 -3760 10985 -3640
rect 11105 -3760 11150 -3640
rect 11270 -3760 11325 -3640
rect 11445 -3760 11490 -3640
rect 11610 -3760 11655 -3640
rect 11775 -3760 11820 -3640
rect 11940 -3760 11995 -3640
rect 12115 -3760 12160 -3640
rect 12280 -3760 12325 -3640
rect 12445 -3760 12490 -3640
rect 12610 -3760 12635 -3640
rect 7105 -3805 12635 -3760
rect 7105 -3925 7130 -3805
rect 7250 -3925 7305 -3805
rect 7425 -3925 7470 -3805
rect 7590 -3925 7635 -3805
rect 7755 -3925 7800 -3805
rect 7920 -3925 7975 -3805
rect 8095 -3925 8140 -3805
rect 8260 -3925 8305 -3805
rect 8425 -3925 8470 -3805
rect 8590 -3925 8645 -3805
rect 8765 -3925 8810 -3805
rect 8930 -3925 8975 -3805
rect 9095 -3925 9140 -3805
rect 9260 -3925 9315 -3805
rect 9435 -3925 9480 -3805
rect 9600 -3925 9645 -3805
rect 9765 -3925 9810 -3805
rect 9930 -3925 9985 -3805
rect 10105 -3925 10150 -3805
rect 10270 -3925 10315 -3805
rect 10435 -3925 10480 -3805
rect 10600 -3925 10655 -3805
rect 10775 -3925 10820 -3805
rect 10940 -3925 10985 -3805
rect 11105 -3925 11150 -3805
rect 11270 -3925 11325 -3805
rect 11445 -3925 11490 -3805
rect 11610 -3925 11655 -3805
rect 11775 -3925 11820 -3805
rect 11940 -3925 11995 -3805
rect 12115 -3925 12160 -3805
rect 12280 -3925 12325 -3805
rect 12445 -3925 12490 -3805
rect 12610 -3925 12635 -3805
rect 7105 -3980 12635 -3925
rect 7105 -4100 7130 -3980
rect 7250 -4100 7305 -3980
rect 7425 -4100 7470 -3980
rect 7590 -4100 7635 -3980
rect 7755 -4100 7800 -3980
rect 7920 -4100 7975 -3980
rect 8095 -4100 8140 -3980
rect 8260 -4100 8305 -3980
rect 8425 -4100 8470 -3980
rect 8590 -4100 8645 -3980
rect 8765 -4100 8810 -3980
rect 8930 -4100 8975 -3980
rect 9095 -4100 9140 -3980
rect 9260 -4100 9315 -3980
rect 9435 -4100 9480 -3980
rect 9600 -4100 9645 -3980
rect 9765 -4100 9810 -3980
rect 9930 -4100 9985 -3980
rect 10105 -4100 10150 -3980
rect 10270 -4100 10315 -3980
rect 10435 -4100 10480 -3980
rect 10600 -4100 10655 -3980
rect 10775 -4100 10820 -3980
rect 10940 -4100 10985 -3980
rect 11105 -4100 11150 -3980
rect 11270 -4100 11325 -3980
rect 11445 -4100 11490 -3980
rect 11610 -4100 11655 -3980
rect 11775 -4100 11820 -3980
rect 11940 -4100 11995 -3980
rect 12115 -4100 12160 -3980
rect 12280 -4100 12325 -3980
rect 12445 -4100 12490 -3980
rect 12610 -4100 12635 -3980
rect 7105 -4125 12635 -4100
rect 12795 1380 18325 1450
rect 12795 1260 12820 1380
rect 12940 1260 12995 1380
rect 13115 1260 13160 1380
rect 13280 1260 13325 1380
rect 13445 1260 13490 1380
rect 13610 1260 13665 1380
rect 13785 1260 13830 1380
rect 13950 1260 13995 1380
rect 14115 1260 14160 1380
rect 14280 1260 14335 1380
rect 14455 1260 14500 1380
rect 14620 1260 14665 1380
rect 14785 1260 14830 1380
rect 14950 1260 15005 1380
rect 15125 1260 15170 1380
rect 15290 1260 15335 1380
rect 15455 1260 15500 1380
rect 15620 1260 15675 1380
rect 15795 1260 15840 1380
rect 15960 1260 16005 1380
rect 16125 1260 16170 1380
rect 16290 1260 16345 1380
rect 16465 1260 16510 1380
rect 16630 1260 16675 1380
rect 16795 1260 16840 1380
rect 16960 1260 17015 1380
rect 17135 1260 17180 1380
rect 17300 1260 17345 1380
rect 17465 1260 17510 1380
rect 17630 1260 17685 1380
rect 17805 1260 17850 1380
rect 17970 1260 18015 1380
rect 18135 1260 18180 1380
rect 18300 1260 18325 1380
rect 12795 1215 18325 1260
rect 12795 1095 12820 1215
rect 12940 1095 12995 1215
rect 13115 1095 13160 1215
rect 13280 1095 13325 1215
rect 13445 1095 13490 1215
rect 13610 1095 13665 1215
rect 13785 1095 13830 1215
rect 13950 1095 13995 1215
rect 14115 1095 14160 1215
rect 14280 1095 14335 1215
rect 14455 1095 14500 1215
rect 14620 1095 14665 1215
rect 14785 1095 14830 1215
rect 14950 1095 15005 1215
rect 15125 1095 15170 1215
rect 15290 1095 15335 1215
rect 15455 1095 15500 1215
rect 15620 1095 15675 1215
rect 15795 1095 15840 1215
rect 15960 1095 16005 1215
rect 16125 1095 16170 1215
rect 16290 1095 16345 1215
rect 16465 1095 16510 1215
rect 16630 1095 16675 1215
rect 16795 1095 16840 1215
rect 16960 1095 17015 1215
rect 17135 1095 17180 1215
rect 17300 1095 17345 1215
rect 17465 1095 17510 1215
rect 17630 1095 17685 1215
rect 17805 1095 17850 1215
rect 17970 1095 18015 1215
rect 18135 1095 18180 1215
rect 18300 1095 18325 1215
rect 12795 1050 18325 1095
rect 12795 930 12820 1050
rect 12940 930 12995 1050
rect 13115 930 13160 1050
rect 13280 930 13325 1050
rect 13445 930 13490 1050
rect 13610 930 13665 1050
rect 13785 930 13830 1050
rect 13950 930 13995 1050
rect 14115 930 14160 1050
rect 14280 930 14335 1050
rect 14455 930 14500 1050
rect 14620 930 14665 1050
rect 14785 930 14830 1050
rect 14950 930 15005 1050
rect 15125 930 15170 1050
rect 15290 930 15335 1050
rect 15455 930 15500 1050
rect 15620 930 15675 1050
rect 15795 930 15840 1050
rect 15960 930 16005 1050
rect 16125 930 16170 1050
rect 16290 930 16345 1050
rect 16465 930 16510 1050
rect 16630 930 16675 1050
rect 16795 930 16840 1050
rect 16960 930 17015 1050
rect 17135 930 17180 1050
rect 17300 930 17345 1050
rect 17465 930 17510 1050
rect 17630 930 17685 1050
rect 17805 930 17850 1050
rect 17970 930 18015 1050
rect 18135 930 18180 1050
rect 18300 930 18325 1050
rect 12795 885 18325 930
rect 12795 765 12820 885
rect 12940 765 12995 885
rect 13115 765 13160 885
rect 13280 765 13325 885
rect 13445 765 13490 885
rect 13610 765 13665 885
rect 13785 765 13830 885
rect 13950 765 13995 885
rect 14115 765 14160 885
rect 14280 765 14335 885
rect 14455 765 14500 885
rect 14620 765 14665 885
rect 14785 765 14830 885
rect 14950 765 15005 885
rect 15125 765 15170 885
rect 15290 765 15335 885
rect 15455 765 15500 885
rect 15620 765 15675 885
rect 15795 765 15840 885
rect 15960 765 16005 885
rect 16125 765 16170 885
rect 16290 765 16345 885
rect 16465 765 16510 885
rect 16630 765 16675 885
rect 16795 765 16840 885
rect 16960 765 17015 885
rect 17135 765 17180 885
rect 17300 765 17345 885
rect 17465 765 17510 885
rect 17630 765 17685 885
rect 17805 765 17850 885
rect 17970 765 18015 885
rect 18135 765 18180 885
rect 18300 765 18325 885
rect 12795 710 18325 765
rect 12795 590 12820 710
rect 12940 590 12995 710
rect 13115 590 13160 710
rect 13280 590 13325 710
rect 13445 590 13490 710
rect 13610 590 13665 710
rect 13785 590 13830 710
rect 13950 590 13995 710
rect 14115 590 14160 710
rect 14280 590 14335 710
rect 14455 590 14500 710
rect 14620 590 14665 710
rect 14785 590 14830 710
rect 14950 590 15005 710
rect 15125 590 15170 710
rect 15290 590 15335 710
rect 15455 590 15500 710
rect 15620 590 15675 710
rect 15795 590 15840 710
rect 15960 590 16005 710
rect 16125 590 16170 710
rect 16290 590 16345 710
rect 16465 590 16510 710
rect 16630 590 16675 710
rect 16795 590 16840 710
rect 16960 590 17015 710
rect 17135 590 17180 710
rect 17300 590 17345 710
rect 17465 590 17510 710
rect 17630 590 17685 710
rect 17805 590 17850 710
rect 17970 590 18015 710
rect 18135 590 18180 710
rect 18300 590 18325 710
rect 12795 545 18325 590
rect 12795 425 12820 545
rect 12940 425 12995 545
rect 13115 425 13160 545
rect 13280 425 13325 545
rect 13445 425 13490 545
rect 13610 425 13665 545
rect 13785 425 13830 545
rect 13950 425 13995 545
rect 14115 425 14160 545
rect 14280 425 14335 545
rect 14455 425 14500 545
rect 14620 425 14665 545
rect 14785 425 14830 545
rect 14950 425 15005 545
rect 15125 425 15170 545
rect 15290 425 15335 545
rect 15455 425 15500 545
rect 15620 425 15675 545
rect 15795 425 15840 545
rect 15960 425 16005 545
rect 16125 425 16170 545
rect 16290 425 16345 545
rect 16465 425 16510 545
rect 16630 425 16675 545
rect 16795 425 16840 545
rect 16960 425 17015 545
rect 17135 425 17180 545
rect 17300 425 17345 545
rect 17465 425 17510 545
rect 17630 425 17685 545
rect 17805 425 17850 545
rect 17970 425 18015 545
rect 18135 425 18180 545
rect 18300 425 18325 545
rect 12795 380 18325 425
rect 12795 260 12820 380
rect 12940 260 12995 380
rect 13115 260 13160 380
rect 13280 260 13325 380
rect 13445 260 13490 380
rect 13610 260 13665 380
rect 13785 260 13830 380
rect 13950 260 13995 380
rect 14115 260 14160 380
rect 14280 260 14335 380
rect 14455 260 14500 380
rect 14620 260 14665 380
rect 14785 260 14830 380
rect 14950 260 15005 380
rect 15125 260 15170 380
rect 15290 260 15335 380
rect 15455 260 15500 380
rect 15620 260 15675 380
rect 15795 260 15840 380
rect 15960 260 16005 380
rect 16125 260 16170 380
rect 16290 260 16345 380
rect 16465 260 16510 380
rect 16630 260 16675 380
rect 16795 260 16840 380
rect 16960 260 17015 380
rect 17135 260 17180 380
rect 17300 260 17345 380
rect 17465 260 17510 380
rect 17630 260 17685 380
rect 17805 260 17850 380
rect 17970 260 18015 380
rect 18135 260 18180 380
rect 18300 260 18325 380
rect 12795 215 18325 260
rect 12795 95 12820 215
rect 12940 95 12995 215
rect 13115 95 13160 215
rect 13280 95 13325 215
rect 13445 95 13490 215
rect 13610 95 13665 215
rect 13785 95 13830 215
rect 13950 95 13995 215
rect 14115 95 14160 215
rect 14280 95 14335 215
rect 14455 95 14500 215
rect 14620 95 14665 215
rect 14785 95 14830 215
rect 14950 95 15005 215
rect 15125 95 15170 215
rect 15290 95 15335 215
rect 15455 95 15500 215
rect 15620 95 15675 215
rect 15795 95 15840 215
rect 15960 95 16005 215
rect 16125 95 16170 215
rect 16290 95 16345 215
rect 16465 95 16510 215
rect 16630 95 16675 215
rect 16795 95 16840 215
rect 16960 95 17015 215
rect 17135 95 17180 215
rect 17300 95 17345 215
rect 17465 95 17510 215
rect 17630 95 17685 215
rect 17805 95 17850 215
rect 17970 95 18015 215
rect 18135 95 18180 215
rect 18300 95 18325 215
rect 12795 40 18325 95
rect 12795 -80 12820 40
rect 12940 -80 12995 40
rect 13115 -80 13160 40
rect 13280 -80 13325 40
rect 13445 -80 13490 40
rect 13610 -80 13665 40
rect 13785 -80 13830 40
rect 13950 -80 13995 40
rect 14115 -80 14160 40
rect 14280 -80 14335 40
rect 14455 -80 14500 40
rect 14620 -80 14665 40
rect 14785 -80 14830 40
rect 14950 -80 15005 40
rect 15125 -80 15170 40
rect 15290 -80 15335 40
rect 15455 -80 15500 40
rect 15620 -80 15675 40
rect 15795 -80 15840 40
rect 15960 -80 16005 40
rect 16125 -80 16170 40
rect 16290 -80 16345 40
rect 16465 -80 16510 40
rect 16630 -80 16675 40
rect 16795 -80 16840 40
rect 16960 -80 17015 40
rect 17135 -80 17180 40
rect 17300 -80 17345 40
rect 17465 -80 17510 40
rect 17630 -80 17685 40
rect 17805 -80 17850 40
rect 17970 -80 18015 40
rect 18135 -80 18180 40
rect 18300 -80 18325 40
rect 12795 -125 18325 -80
rect 12795 -245 12820 -125
rect 12940 -245 12995 -125
rect 13115 -245 13160 -125
rect 13280 -245 13325 -125
rect 13445 -245 13490 -125
rect 13610 -245 13665 -125
rect 13785 -245 13830 -125
rect 13950 -245 13995 -125
rect 14115 -245 14160 -125
rect 14280 -245 14335 -125
rect 14455 -245 14500 -125
rect 14620 -245 14665 -125
rect 14785 -245 14830 -125
rect 14950 -245 15005 -125
rect 15125 -245 15170 -125
rect 15290 -245 15335 -125
rect 15455 -245 15500 -125
rect 15620 -245 15675 -125
rect 15795 -245 15840 -125
rect 15960 -245 16005 -125
rect 16125 -245 16170 -125
rect 16290 -245 16345 -125
rect 16465 -245 16510 -125
rect 16630 -245 16675 -125
rect 16795 -245 16840 -125
rect 16960 -245 17015 -125
rect 17135 -245 17180 -125
rect 17300 -245 17345 -125
rect 17465 -245 17510 -125
rect 17630 -245 17685 -125
rect 17805 -245 17850 -125
rect 17970 -245 18015 -125
rect 18135 -245 18180 -125
rect 18300 -245 18325 -125
rect 12795 -290 18325 -245
rect 12795 -410 12820 -290
rect 12940 -410 12995 -290
rect 13115 -410 13160 -290
rect 13280 -410 13325 -290
rect 13445 -410 13490 -290
rect 13610 -410 13665 -290
rect 13785 -410 13830 -290
rect 13950 -410 13995 -290
rect 14115 -410 14160 -290
rect 14280 -410 14335 -290
rect 14455 -410 14500 -290
rect 14620 -410 14665 -290
rect 14785 -410 14830 -290
rect 14950 -410 15005 -290
rect 15125 -410 15170 -290
rect 15290 -410 15335 -290
rect 15455 -410 15500 -290
rect 15620 -410 15675 -290
rect 15795 -410 15840 -290
rect 15960 -410 16005 -290
rect 16125 -410 16170 -290
rect 16290 -410 16345 -290
rect 16465 -410 16510 -290
rect 16630 -410 16675 -290
rect 16795 -410 16840 -290
rect 16960 -410 17015 -290
rect 17135 -410 17180 -290
rect 17300 -410 17345 -290
rect 17465 -410 17510 -290
rect 17630 -410 17685 -290
rect 17805 -410 17850 -290
rect 17970 -410 18015 -290
rect 18135 -410 18180 -290
rect 18300 -410 18325 -290
rect 12795 -455 18325 -410
rect 12795 -575 12820 -455
rect 12940 -575 12995 -455
rect 13115 -575 13160 -455
rect 13280 -575 13325 -455
rect 13445 -575 13490 -455
rect 13610 -575 13665 -455
rect 13785 -575 13830 -455
rect 13950 -575 13995 -455
rect 14115 -575 14160 -455
rect 14280 -575 14335 -455
rect 14455 -575 14500 -455
rect 14620 -575 14665 -455
rect 14785 -575 14830 -455
rect 14950 -575 15005 -455
rect 15125 -575 15170 -455
rect 15290 -575 15335 -455
rect 15455 -575 15500 -455
rect 15620 -575 15675 -455
rect 15795 -575 15840 -455
rect 15960 -575 16005 -455
rect 16125 -575 16170 -455
rect 16290 -575 16345 -455
rect 16465 -575 16510 -455
rect 16630 -575 16675 -455
rect 16795 -575 16840 -455
rect 16960 -575 17015 -455
rect 17135 -575 17180 -455
rect 17300 -575 17345 -455
rect 17465 -575 17510 -455
rect 17630 -575 17685 -455
rect 17805 -575 17850 -455
rect 17970 -575 18015 -455
rect 18135 -575 18180 -455
rect 18300 -575 18325 -455
rect 12795 -630 18325 -575
rect 12795 -750 12820 -630
rect 12940 -750 12995 -630
rect 13115 -750 13160 -630
rect 13280 -750 13325 -630
rect 13445 -750 13490 -630
rect 13610 -750 13665 -630
rect 13785 -750 13830 -630
rect 13950 -750 13995 -630
rect 14115 -750 14160 -630
rect 14280 -750 14335 -630
rect 14455 -750 14500 -630
rect 14620 -750 14665 -630
rect 14785 -750 14830 -630
rect 14950 -750 15005 -630
rect 15125 -750 15170 -630
rect 15290 -750 15335 -630
rect 15455 -750 15500 -630
rect 15620 -750 15675 -630
rect 15795 -750 15840 -630
rect 15960 -750 16005 -630
rect 16125 -750 16170 -630
rect 16290 -750 16345 -630
rect 16465 -750 16510 -630
rect 16630 -750 16675 -630
rect 16795 -750 16840 -630
rect 16960 -750 17015 -630
rect 17135 -750 17180 -630
rect 17300 -750 17345 -630
rect 17465 -750 17510 -630
rect 17630 -750 17685 -630
rect 17805 -750 17850 -630
rect 17970 -750 18015 -630
rect 18135 -750 18180 -630
rect 18300 -750 18325 -630
rect 12795 -795 18325 -750
rect 12795 -915 12820 -795
rect 12940 -915 12995 -795
rect 13115 -915 13160 -795
rect 13280 -915 13325 -795
rect 13445 -915 13490 -795
rect 13610 -915 13665 -795
rect 13785 -915 13830 -795
rect 13950 -915 13995 -795
rect 14115 -915 14160 -795
rect 14280 -915 14335 -795
rect 14455 -915 14500 -795
rect 14620 -915 14665 -795
rect 14785 -915 14830 -795
rect 14950 -915 15005 -795
rect 15125 -915 15170 -795
rect 15290 -915 15335 -795
rect 15455 -915 15500 -795
rect 15620 -915 15675 -795
rect 15795 -915 15840 -795
rect 15960 -915 16005 -795
rect 16125 -915 16170 -795
rect 16290 -915 16345 -795
rect 16465 -915 16510 -795
rect 16630 -915 16675 -795
rect 16795 -915 16840 -795
rect 16960 -915 17015 -795
rect 17135 -915 17180 -795
rect 17300 -915 17345 -795
rect 17465 -915 17510 -795
rect 17630 -915 17685 -795
rect 17805 -915 17850 -795
rect 17970 -915 18015 -795
rect 18135 -915 18180 -795
rect 18300 -915 18325 -795
rect 12795 -960 18325 -915
rect 12795 -1080 12820 -960
rect 12940 -1080 12995 -960
rect 13115 -1080 13160 -960
rect 13280 -1080 13325 -960
rect 13445 -1080 13490 -960
rect 13610 -1080 13665 -960
rect 13785 -1080 13830 -960
rect 13950 -1080 13995 -960
rect 14115 -1080 14160 -960
rect 14280 -1080 14335 -960
rect 14455 -1080 14500 -960
rect 14620 -1080 14665 -960
rect 14785 -1080 14830 -960
rect 14950 -1080 15005 -960
rect 15125 -1080 15170 -960
rect 15290 -1080 15335 -960
rect 15455 -1080 15500 -960
rect 15620 -1080 15675 -960
rect 15795 -1080 15840 -960
rect 15960 -1080 16005 -960
rect 16125 -1080 16170 -960
rect 16290 -1080 16345 -960
rect 16465 -1080 16510 -960
rect 16630 -1080 16675 -960
rect 16795 -1080 16840 -960
rect 16960 -1080 17015 -960
rect 17135 -1080 17180 -960
rect 17300 -1080 17345 -960
rect 17465 -1080 17510 -960
rect 17630 -1080 17685 -960
rect 17805 -1080 17850 -960
rect 17970 -1080 18015 -960
rect 18135 -1080 18180 -960
rect 18300 -1080 18325 -960
rect 12795 -1125 18325 -1080
rect 12795 -1245 12820 -1125
rect 12940 -1245 12995 -1125
rect 13115 -1245 13160 -1125
rect 13280 -1245 13325 -1125
rect 13445 -1245 13490 -1125
rect 13610 -1245 13665 -1125
rect 13785 -1245 13830 -1125
rect 13950 -1245 13995 -1125
rect 14115 -1245 14160 -1125
rect 14280 -1245 14335 -1125
rect 14455 -1245 14500 -1125
rect 14620 -1245 14665 -1125
rect 14785 -1245 14830 -1125
rect 14950 -1245 15005 -1125
rect 15125 -1245 15170 -1125
rect 15290 -1245 15335 -1125
rect 15455 -1245 15500 -1125
rect 15620 -1245 15675 -1125
rect 15795 -1245 15840 -1125
rect 15960 -1245 16005 -1125
rect 16125 -1245 16170 -1125
rect 16290 -1245 16345 -1125
rect 16465 -1245 16510 -1125
rect 16630 -1245 16675 -1125
rect 16795 -1245 16840 -1125
rect 16960 -1245 17015 -1125
rect 17135 -1245 17180 -1125
rect 17300 -1245 17345 -1125
rect 17465 -1245 17510 -1125
rect 17630 -1245 17685 -1125
rect 17805 -1245 17850 -1125
rect 17970 -1245 18015 -1125
rect 18135 -1245 18180 -1125
rect 18300 -1245 18325 -1125
rect 12795 -1300 18325 -1245
rect 12795 -1420 12820 -1300
rect 12940 -1420 12995 -1300
rect 13115 -1420 13160 -1300
rect 13280 -1420 13325 -1300
rect 13445 -1420 13490 -1300
rect 13610 -1420 13665 -1300
rect 13785 -1420 13830 -1300
rect 13950 -1420 13995 -1300
rect 14115 -1420 14160 -1300
rect 14280 -1420 14335 -1300
rect 14455 -1420 14500 -1300
rect 14620 -1420 14665 -1300
rect 14785 -1420 14830 -1300
rect 14950 -1420 15005 -1300
rect 15125 -1420 15170 -1300
rect 15290 -1420 15335 -1300
rect 15455 -1420 15500 -1300
rect 15620 -1420 15675 -1300
rect 15795 -1420 15840 -1300
rect 15960 -1420 16005 -1300
rect 16125 -1420 16170 -1300
rect 16290 -1420 16345 -1300
rect 16465 -1420 16510 -1300
rect 16630 -1420 16675 -1300
rect 16795 -1420 16840 -1300
rect 16960 -1420 17015 -1300
rect 17135 -1420 17180 -1300
rect 17300 -1420 17345 -1300
rect 17465 -1420 17510 -1300
rect 17630 -1420 17685 -1300
rect 17805 -1420 17850 -1300
rect 17970 -1420 18015 -1300
rect 18135 -1420 18180 -1300
rect 18300 -1420 18325 -1300
rect 12795 -1465 18325 -1420
rect 12795 -1585 12820 -1465
rect 12940 -1585 12995 -1465
rect 13115 -1585 13160 -1465
rect 13280 -1585 13325 -1465
rect 13445 -1585 13490 -1465
rect 13610 -1585 13665 -1465
rect 13785 -1585 13830 -1465
rect 13950 -1585 13995 -1465
rect 14115 -1585 14160 -1465
rect 14280 -1585 14335 -1465
rect 14455 -1585 14500 -1465
rect 14620 -1585 14665 -1465
rect 14785 -1585 14830 -1465
rect 14950 -1585 15005 -1465
rect 15125 -1585 15170 -1465
rect 15290 -1585 15335 -1465
rect 15455 -1585 15500 -1465
rect 15620 -1585 15675 -1465
rect 15795 -1585 15840 -1465
rect 15960 -1585 16005 -1465
rect 16125 -1585 16170 -1465
rect 16290 -1585 16345 -1465
rect 16465 -1585 16510 -1465
rect 16630 -1585 16675 -1465
rect 16795 -1585 16840 -1465
rect 16960 -1585 17015 -1465
rect 17135 -1585 17180 -1465
rect 17300 -1585 17345 -1465
rect 17465 -1585 17510 -1465
rect 17630 -1585 17685 -1465
rect 17805 -1585 17850 -1465
rect 17970 -1585 18015 -1465
rect 18135 -1585 18180 -1465
rect 18300 -1585 18325 -1465
rect 12795 -1630 18325 -1585
rect 12795 -1750 12820 -1630
rect 12940 -1750 12995 -1630
rect 13115 -1750 13160 -1630
rect 13280 -1750 13325 -1630
rect 13445 -1750 13490 -1630
rect 13610 -1750 13665 -1630
rect 13785 -1750 13830 -1630
rect 13950 -1750 13995 -1630
rect 14115 -1750 14160 -1630
rect 14280 -1750 14335 -1630
rect 14455 -1750 14500 -1630
rect 14620 -1750 14665 -1630
rect 14785 -1750 14830 -1630
rect 14950 -1750 15005 -1630
rect 15125 -1750 15170 -1630
rect 15290 -1750 15335 -1630
rect 15455 -1750 15500 -1630
rect 15620 -1750 15675 -1630
rect 15795 -1750 15840 -1630
rect 15960 -1750 16005 -1630
rect 16125 -1750 16170 -1630
rect 16290 -1750 16345 -1630
rect 16465 -1750 16510 -1630
rect 16630 -1750 16675 -1630
rect 16795 -1750 16840 -1630
rect 16960 -1750 17015 -1630
rect 17135 -1750 17180 -1630
rect 17300 -1750 17345 -1630
rect 17465 -1750 17510 -1630
rect 17630 -1750 17685 -1630
rect 17805 -1750 17850 -1630
rect 17970 -1750 18015 -1630
rect 18135 -1750 18180 -1630
rect 18300 -1750 18325 -1630
rect 12795 -1795 18325 -1750
rect 12795 -1915 12820 -1795
rect 12940 -1915 12995 -1795
rect 13115 -1915 13160 -1795
rect 13280 -1915 13325 -1795
rect 13445 -1915 13490 -1795
rect 13610 -1915 13665 -1795
rect 13785 -1915 13830 -1795
rect 13950 -1915 13995 -1795
rect 14115 -1915 14160 -1795
rect 14280 -1915 14335 -1795
rect 14455 -1915 14500 -1795
rect 14620 -1915 14665 -1795
rect 14785 -1915 14830 -1795
rect 14950 -1915 15005 -1795
rect 15125 -1915 15170 -1795
rect 15290 -1915 15335 -1795
rect 15455 -1915 15500 -1795
rect 15620 -1915 15675 -1795
rect 15795 -1915 15840 -1795
rect 15960 -1915 16005 -1795
rect 16125 -1915 16170 -1795
rect 16290 -1915 16345 -1795
rect 16465 -1915 16510 -1795
rect 16630 -1915 16675 -1795
rect 16795 -1915 16840 -1795
rect 16960 -1915 17015 -1795
rect 17135 -1915 17180 -1795
rect 17300 -1915 17345 -1795
rect 17465 -1915 17510 -1795
rect 17630 -1915 17685 -1795
rect 17805 -1915 17850 -1795
rect 17970 -1915 18015 -1795
rect 18135 -1915 18180 -1795
rect 18300 -1915 18325 -1795
rect 12795 -1970 18325 -1915
rect 12795 -2090 12820 -1970
rect 12940 -2090 12995 -1970
rect 13115 -2090 13160 -1970
rect 13280 -2090 13325 -1970
rect 13445 -2090 13490 -1970
rect 13610 -2090 13665 -1970
rect 13785 -2090 13830 -1970
rect 13950 -2090 13995 -1970
rect 14115 -2090 14160 -1970
rect 14280 -2090 14335 -1970
rect 14455 -2090 14500 -1970
rect 14620 -2090 14665 -1970
rect 14785 -2090 14830 -1970
rect 14950 -2090 15005 -1970
rect 15125 -2090 15170 -1970
rect 15290 -2090 15335 -1970
rect 15455 -2090 15500 -1970
rect 15620 -2090 15675 -1970
rect 15795 -2090 15840 -1970
rect 15960 -2090 16005 -1970
rect 16125 -2090 16170 -1970
rect 16290 -2090 16345 -1970
rect 16465 -2090 16510 -1970
rect 16630 -2090 16675 -1970
rect 16795 -2090 16840 -1970
rect 16960 -2090 17015 -1970
rect 17135 -2090 17180 -1970
rect 17300 -2090 17345 -1970
rect 17465 -2090 17510 -1970
rect 17630 -2090 17685 -1970
rect 17805 -2090 17850 -1970
rect 17970 -2090 18015 -1970
rect 18135 -2090 18180 -1970
rect 18300 -2090 18325 -1970
rect 12795 -2135 18325 -2090
rect 12795 -2255 12820 -2135
rect 12940 -2255 12995 -2135
rect 13115 -2255 13160 -2135
rect 13280 -2255 13325 -2135
rect 13445 -2255 13490 -2135
rect 13610 -2255 13665 -2135
rect 13785 -2255 13830 -2135
rect 13950 -2255 13995 -2135
rect 14115 -2255 14160 -2135
rect 14280 -2255 14335 -2135
rect 14455 -2255 14500 -2135
rect 14620 -2255 14665 -2135
rect 14785 -2255 14830 -2135
rect 14950 -2255 15005 -2135
rect 15125 -2255 15170 -2135
rect 15290 -2255 15335 -2135
rect 15455 -2255 15500 -2135
rect 15620 -2255 15675 -2135
rect 15795 -2255 15840 -2135
rect 15960 -2255 16005 -2135
rect 16125 -2255 16170 -2135
rect 16290 -2255 16345 -2135
rect 16465 -2255 16510 -2135
rect 16630 -2255 16675 -2135
rect 16795 -2255 16840 -2135
rect 16960 -2255 17015 -2135
rect 17135 -2255 17180 -2135
rect 17300 -2255 17345 -2135
rect 17465 -2255 17510 -2135
rect 17630 -2255 17685 -2135
rect 17805 -2255 17850 -2135
rect 17970 -2255 18015 -2135
rect 18135 -2255 18180 -2135
rect 18300 -2255 18325 -2135
rect 12795 -2300 18325 -2255
rect 12795 -2420 12820 -2300
rect 12940 -2420 12995 -2300
rect 13115 -2420 13160 -2300
rect 13280 -2420 13325 -2300
rect 13445 -2420 13490 -2300
rect 13610 -2420 13665 -2300
rect 13785 -2420 13830 -2300
rect 13950 -2420 13995 -2300
rect 14115 -2420 14160 -2300
rect 14280 -2420 14335 -2300
rect 14455 -2420 14500 -2300
rect 14620 -2420 14665 -2300
rect 14785 -2420 14830 -2300
rect 14950 -2420 15005 -2300
rect 15125 -2420 15170 -2300
rect 15290 -2420 15335 -2300
rect 15455 -2420 15500 -2300
rect 15620 -2420 15675 -2300
rect 15795 -2420 15840 -2300
rect 15960 -2420 16005 -2300
rect 16125 -2420 16170 -2300
rect 16290 -2420 16345 -2300
rect 16465 -2420 16510 -2300
rect 16630 -2420 16675 -2300
rect 16795 -2420 16840 -2300
rect 16960 -2420 17015 -2300
rect 17135 -2420 17180 -2300
rect 17300 -2420 17345 -2300
rect 17465 -2420 17510 -2300
rect 17630 -2420 17685 -2300
rect 17805 -2420 17850 -2300
rect 17970 -2420 18015 -2300
rect 18135 -2420 18180 -2300
rect 18300 -2420 18325 -2300
rect 12795 -2465 18325 -2420
rect 12795 -2585 12820 -2465
rect 12940 -2585 12995 -2465
rect 13115 -2585 13160 -2465
rect 13280 -2585 13325 -2465
rect 13445 -2585 13490 -2465
rect 13610 -2585 13665 -2465
rect 13785 -2585 13830 -2465
rect 13950 -2585 13995 -2465
rect 14115 -2585 14160 -2465
rect 14280 -2585 14335 -2465
rect 14455 -2585 14500 -2465
rect 14620 -2585 14665 -2465
rect 14785 -2585 14830 -2465
rect 14950 -2585 15005 -2465
rect 15125 -2585 15170 -2465
rect 15290 -2585 15335 -2465
rect 15455 -2585 15500 -2465
rect 15620 -2585 15675 -2465
rect 15795 -2585 15840 -2465
rect 15960 -2585 16005 -2465
rect 16125 -2585 16170 -2465
rect 16290 -2585 16345 -2465
rect 16465 -2585 16510 -2465
rect 16630 -2585 16675 -2465
rect 16795 -2585 16840 -2465
rect 16960 -2585 17015 -2465
rect 17135 -2585 17180 -2465
rect 17300 -2585 17345 -2465
rect 17465 -2585 17510 -2465
rect 17630 -2585 17685 -2465
rect 17805 -2585 17850 -2465
rect 17970 -2585 18015 -2465
rect 18135 -2585 18180 -2465
rect 18300 -2585 18325 -2465
rect 12795 -2640 18325 -2585
rect 12795 -2760 12820 -2640
rect 12940 -2760 12995 -2640
rect 13115 -2760 13160 -2640
rect 13280 -2760 13325 -2640
rect 13445 -2760 13490 -2640
rect 13610 -2760 13665 -2640
rect 13785 -2760 13830 -2640
rect 13950 -2760 13995 -2640
rect 14115 -2760 14160 -2640
rect 14280 -2760 14335 -2640
rect 14455 -2760 14500 -2640
rect 14620 -2760 14665 -2640
rect 14785 -2760 14830 -2640
rect 14950 -2760 15005 -2640
rect 15125 -2760 15170 -2640
rect 15290 -2760 15335 -2640
rect 15455 -2760 15500 -2640
rect 15620 -2760 15675 -2640
rect 15795 -2760 15840 -2640
rect 15960 -2760 16005 -2640
rect 16125 -2760 16170 -2640
rect 16290 -2760 16345 -2640
rect 16465 -2760 16510 -2640
rect 16630 -2760 16675 -2640
rect 16795 -2760 16840 -2640
rect 16960 -2760 17015 -2640
rect 17135 -2760 17180 -2640
rect 17300 -2760 17345 -2640
rect 17465 -2760 17510 -2640
rect 17630 -2760 17685 -2640
rect 17805 -2760 17850 -2640
rect 17970 -2760 18015 -2640
rect 18135 -2760 18180 -2640
rect 18300 -2760 18325 -2640
rect 12795 -2805 18325 -2760
rect 12795 -2925 12820 -2805
rect 12940 -2925 12995 -2805
rect 13115 -2925 13160 -2805
rect 13280 -2925 13325 -2805
rect 13445 -2925 13490 -2805
rect 13610 -2925 13665 -2805
rect 13785 -2925 13830 -2805
rect 13950 -2925 13995 -2805
rect 14115 -2925 14160 -2805
rect 14280 -2925 14335 -2805
rect 14455 -2925 14500 -2805
rect 14620 -2925 14665 -2805
rect 14785 -2925 14830 -2805
rect 14950 -2925 15005 -2805
rect 15125 -2925 15170 -2805
rect 15290 -2925 15335 -2805
rect 15455 -2925 15500 -2805
rect 15620 -2925 15675 -2805
rect 15795 -2925 15840 -2805
rect 15960 -2925 16005 -2805
rect 16125 -2925 16170 -2805
rect 16290 -2925 16345 -2805
rect 16465 -2925 16510 -2805
rect 16630 -2925 16675 -2805
rect 16795 -2925 16840 -2805
rect 16960 -2925 17015 -2805
rect 17135 -2925 17180 -2805
rect 17300 -2925 17345 -2805
rect 17465 -2925 17510 -2805
rect 17630 -2925 17685 -2805
rect 17805 -2925 17850 -2805
rect 17970 -2925 18015 -2805
rect 18135 -2925 18180 -2805
rect 18300 -2925 18325 -2805
rect 12795 -2970 18325 -2925
rect 12795 -3090 12820 -2970
rect 12940 -3090 12995 -2970
rect 13115 -3090 13160 -2970
rect 13280 -3090 13325 -2970
rect 13445 -3090 13490 -2970
rect 13610 -3090 13665 -2970
rect 13785 -3090 13830 -2970
rect 13950 -3090 13995 -2970
rect 14115 -3090 14160 -2970
rect 14280 -3090 14335 -2970
rect 14455 -3090 14500 -2970
rect 14620 -3090 14665 -2970
rect 14785 -3090 14830 -2970
rect 14950 -3090 15005 -2970
rect 15125 -3090 15170 -2970
rect 15290 -3090 15335 -2970
rect 15455 -3090 15500 -2970
rect 15620 -3090 15675 -2970
rect 15795 -3090 15840 -2970
rect 15960 -3090 16005 -2970
rect 16125 -3090 16170 -2970
rect 16290 -3090 16345 -2970
rect 16465 -3090 16510 -2970
rect 16630 -3090 16675 -2970
rect 16795 -3090 16840 -2970
rect 16960 -3090 17015 -2970
rect 17135 -3090 17180 -2970
rect 17300 -3090 17345 -2970
rect 17465 -3090 17510 -2970
rect 17630 -3090 17685 -2970
rect 17805 -3090 17850 -2970
rect 17970 -3090 18015 -2970
rect 18135 -3090 18180 -2970
rect 18300 -3090 18325 -2970
rect 12795 -3135 18325 -3090
rect 12795 -3255 12820 -3135
rect 12940 -3255 12995 -3135
rect 13115 -3255 13160 -3135
rect 13280 -3255 13325 -3135
rect 13445 -3255 13490 -3135
rect 13610 -3255 13665 -3135
rect 13785 -3255 13830 -3135
rect 13950 -3255 13995 -3135
rect 14115 -3255 14160 -3135
rect 14280 -3255 14335 -3135
rect 14455 -3255 14500 -3135
rect 14620 -3255 14665 -3135
rect 14785 -3255 14830 -3135
rect 14950 -3255 15005 -3135
rect 15125 -3255 15170 -3135
rect 15290 -3255 15335 -3135
rect 15455 -3255 15500 -3135
rect 15620 -3255 15675 -3135
rect 15795 -3255 15840 -3135
rect 15960 -3255 16005 -3135
rect 16125 -3255 16170 -3135
rect 16290 -3255 16345 -3135
rect 16465 -3255 16510 -3135
rect 16630 -3255 16675 -3135
rect 16795 -3255 16840 -3135
rect 16960 -3255 17015 -3135
rect 17135 -3255 17180 -3135
rect 17300 -3255 17345 -3135
rect 17465 -3255 17510 -3135
rect 17630 -3255 17685 -3135
rect 17805 -3255 17850 -3135
rect 17970 -3255 18015 -3135
rect 18135 -3255 18180 -3135
rect 18300 -3255 18325 -3135
rect 12795 -3310 18325 -3255
rect 12795 -3430 12820 -3310
rect 12940 -3430 12995 -3310
rect 13115 -3430 13160 -3310
rect 13280 -3430 13325 -3310
rect 13445 -3430 13490 -3310
rect 13610 -3430 13665 -3310
rect 13785 -3430 13830 -3310
rect 13950 -3430 13995 -3310
rect 14115 -3430 14160 -3310
rect 14280 -3430 14335 -3310
rect 14455 -3430 14500 -3310
rect 14620 -3430 14665 -3310
rect 14785 -3430 14830 -3310
rect 14950 -3430 15005 -3310
rect 15125 -3430 15170 -3310
rect 15290 -3430 15335 -3310
rect 15455 -3430 15500 -3310
rect 15620 -3430 15675 -3310
rect 15795 -3430 15840 -3310
rect 15960 -3430 16005 -3310
rect 16125 -3430 16170 -3310
rect 16290 -3430 16345 -3310
rect 16465 -3430 16510 -3310
rect 16630 -3430 16675 -3310
rect 16795 -3430 16840 -3310
rect 16960 -3430 17015 -3310
rect 17135 -3430 17180 -3310
rect 17300 -3430 17345 -3310
rect 17465 -3430 17510 -3310
rect 17630 -3430 17685 -3310
rect 17805 -3430 17850 -3310
rect 17970 -3430 18015 -3310
rect 18135 -3430 18180 -3310
rect 18300 -3430 18325 -3310
rect 12795 -3475 18325 -3430
rect 12795 -3595 12820 -3475
rect 12940 -3595 12995 -3475
rect 13115 -3595 13160 -3475
rect 13280 -3595 13325 -3475
rect 13445 -3595 13490 -3475
rect 13610 -3595 13665 -3475
rect 13785 -3595 13830 -3475
rect 13950 -3595 13995 -3475
rect 14115 -3595 14160 -3475
rect 14280 -3595 14335 -3475
rect 14455 -3595 14500 -3475
rect 14620 -3595 14665 -3475
rect 14785 -3595 14830 -3475
rect 14950 -3595 15005 -3475
rect 15125 -3595 15170 -3475
rect 15290 -3595 15335 -3475
rect 15455 -3595 15500 -3475
rect 15620 -3595 15675 -3475
rect 15795 -3595 15840 -3475
rect 15960 -3595 16005 -3475
rect 16125 -3595 16170 -3475
rect 16290 -3595 16345 -3475
rect 16465 -3595 16510 -3475
rect 16630 -3595 16675 -3475
rect 16795 -3595 16840 -3475
rect 16960 -3595 17015 -3475
rect 17135 -3595 17180 -3475
rect 17300 -3595 17345 -3475
rect 17465 -3595 17510 -3475
rect 17630 -3595 17685 -3475
rect 17805 -3595 17850 -3475
rect 17970 -3595 18015 -3475
rect 18135 -3595 18180 -3475
rect 18300 -3595 18325 -3475
rect 12795 -3640 18325 -3595
rect 12795 -3760 12820 -3640
rect 12940 -3760 12995 -3640
rect 13115 -3760 13160 -3640
rect 13280 -3760 13325 -3640
rect 13445 -3760 13490 -3640
rect 13610 -3760 13665 -3640
rect 13785 -3760 13830 -3640
rect 13950 -3760 13995 -3640
rect 14115 -3760 14160 -3640
rect 14280 -3760 14335 -3640
rect 14455 -3760 14500 -3640
rect 14620 -3760 14665 -3640
rect 14785 -3760 14830 -3640
rect 14950 -3760 15005 -3640
rect 15125 -3760 15170 -3640
rect 15290 -3760 15335 -3640
rect 15455 -3760 15500 -3640
rect 15620 -3760 15675 -3640
rect 15795 -3760 15840 -3640
rect 15960 -3760 16005 -3640
rect 16125 -3760 16170 -3640
rect 16290 -3760 16345 -3640
rect 16465 -3760 16510 -3640
rect 16630 -3760 16675 -3640
rect 16795 -3760 16840 -3640
rect 16960 -3760 17015 -3640
rect 17135 -3760 17180 -3640
rect 17300 -3760 17345 -3640
rect 17465 -3760 17510 -3640
rect 17630 -3760 17685 -3640
rect 17805 -3760 17850 -3640
rect 17970 -3760 18015 -3640
rect 18135 -3760 18180 -3640
rect 18300 -3760 18325 -3640
rect 12795 -3805 18325 -3760
rect 12795 -3925 12820 -3805
rect 12940 -3925 12995 -3805
rect 13115 -3925 13160 -3805
rect 13280 -3925 13325 -3805
rect 13445 -3925 13490 -3805
rect 13610 -3925 13665 -3805
rect 13785 -3925 13830 -3805
rect 13950 -3925 13995 -3805
rect 14115 -3925 14160 -3805
rect 14280 -3925 14335 -3805
rect 14455 -3925 14500 -3805
rect 14620 -3925 14665 -3805
rect 14785 -3925 14830 -3805
rect 14950 -3925 15005 -3805
rect 15125 -3925 15170 -3805
rect 15290 -3925 15335 -3805
rect 15455 -3925 15500 -3805
rect 15620 -3925 15675 -3805
rect 15795 -3925 15840 -3805
rect 15960 -3925 16005 -3805
rect 16125 -3925 16170 -3805
rect 16290 -3925 16345 -3805
rect 16465 -3925 16510 -3805
rect 16630 -3925 16675 -3805
rect 16795 -3925 16840 -3805
rect 16960 -3925 17015 -3805
rect 17135 -3925 17180 -3805
rect 17300 -3925 17345 -3805
rect 17465 -3925 17510 -3805
rect 17630 -3925 17685 -3805
rect 17805 -3925 17850 -3805
rect 17970 -3925 18015 -3805
rect 18135 -3925 18180 -3805
rect 18300 -3925 18325 -3805
rect 12795 -3980 18325 -3925
rect 12795 -4100 12820 -3980
rect 12940 -4100 12995 -3980
rect 13115 -4100 13160 -3980
rect 13280 -4100 13325 -3980
rect 13445 -4100 13490 -3980
rect 13610 -4100 13665 -3980
rect 13785 -4100 13830 -3980
rect 13950 -4100 13995 -3980
rect 14115 -4100 14160 -3980
rect 14280 -4100 14335 -3980
rect 14455 -4100 14500 -3980
rect 14620 -4100 14665 -3980
rect 14785 -4100 14830 -3980
rect 14950 -4100 15005 -3980
rect 15125 -4100 15170 -3980
rect 15290 -4100 15335 -3980
rect 15455 -4100 15500 -3980
rect 15620 -4100 15675 -3980
rect 15795 -4100 15840 -3980
rect 15960 -4100 16005 -3980
rect 16125 -4100 16170 -3980
rect 16290 -4100 16345 -3980
rect 16465 -4100 16510 -3980
rect 16630 -4100 16675 -3980
rect 16795 -4100 16840 -3980
rect 16960 -4100 17015 -3980
rect 17135 -4100 17180 -3980
rect 17300 -4100 17345 -3980
rect 17465 -4100 17510 -3980
rect 17630 -4100 17685 -3980
rect 17805 -4100 17850 -3980
rect 17970 -4100 18015 -3980
rect 18135 -4100 18180 -3980
rect 18300 -4100 18325 -3980
rect 12795 -4125 18325 -4100
rect 18485 1380 24015 1450
rect 18485 1260 18510 1380
rect 18630 1260 18685 1380
rect 18805 1260 18850 1380
rect 18970 1260 19015 1380
rect 19135 1260 19180 1380
rect 19300 1260 19355 1380
rect 19475 1260 19520 1380
rect 19640 1260 19685 1380
rect 19805 1260 19850 1380
rect 19970 1260 20025 1380
rect 20145 1260 20190 1380
rect 20310 1260 20355 1380
rect 20475 1260 20520 1380
rect 20640 1260 20695 1380
rect 20815 1260 20860 1380
rect 20980 1260 21025 1380
rect 21145 1260 21190 1380
rect 21310 1260 21365 1380
rect 21485 1260 21530 1380
rect 21650 1260 21695 1380
rect 21815 1260 21860 1380
rect 21980 1260 22035 1380
rect 22155 1260 22200 1380
rect 22320 1260 22365 1380
rect 22485 1260 22530 1380
rect 22650 1260 22705 1380
rect 22825 1260 22870 1380
rect 22990 1260 23035 1380
rect 23155 1260 23200 1380
rect 23320 1260 23375 1380
rect 23495 1260 23540 1380
rect 23660 1260 23705 1380
rect 23825 1260 23870 1380
rect 23990 1260 24015 1380
rect 18485 1215 24015 1260
rect 18485 1095 18510 1215
rect 18630 1095 18685 1215
rect 18805 1095 18850 1215
rect 18970 1095 19015 1215
rect 19135 1095 19180 1215
rect 19300 1095 19355 1215
rect 19475 1095 19520 1215
rect 19640 1095 19685 1215
rect 19805 1095 19850 1215
rect 19970 1095 20025 1215
rect 20145 1095 20190 1215
rect 20310 1095 20355 1215
rect 20475 1095 20520 1215
rect 20640 1095 20695 1215
rect 20815 1095 20860 1215
rect 20980 1095 21025 1215
rect 21145 1095 21190 1215
rect 21310 1095 21365 1215
rect 21485 1095 21530 1215
rect 21650 1095 21695 1215
rect 21815 1095 21860 1215
rect 21980 1095 22035 1215
rect 22155 1095 22200 1215
rect 22320 1095 22365 1215
rect 22485 1095 22530 1215
rect 22650 1095 22705 1215
rect 22825 1095 22870 1215
rect 22990 1095 23035 1215
rect 23155 1095 23200 1215
rect 23320 1095 23375 1215
rect 23495 1095 23540 1215
rect 23660 1095 23705 1215
rect 23825 1095 23870 1215
rect 23990 1095 24015 1215
rect 18485 1050 24015 1095
rect 18485 930 18510 1050
rect 18630 930 18685 1050
rect 18805 930 18850 1050
rect 18970 930 19015 1050
rect 19135 930 19180 1050
rect 19300 930 19355 1050
rect 19475 930 19520 1050
rect 19640 930 19685 1050
rect 19805 930 19850 1050
rect 19970 930 20025 1050
rect 20145 930 20190 1050
rect 20310 930 20355 1050
rect 20475 930 20520 1050
rect 20640 930 20695 1050
rect 20815 930 20860 1050
rect 20980 930 21025 1050
rect 21145 930 21190 1050
rect 21310 930 21365 1050
rect 21485 930 21530 1050
rect 21650 930 21695 1050
rect 21815 930 21860 1050
rect 21980 930 22035 1050
rect 22155 930 22200 1050
rect 22320 930 22365 1050
rect 22485 930 22530 1050
rect 22650 930 22705 1050
rect 22825 930 22870 1050
rect 22990 930 23035 1050
rect 23155 930 23200 1050
rect 23320 930 23375 1050
rect 23495 930 23540 1050
rect 23660 930 23705 1050
rect 23825 930 23870 1050
rect 23990 930 24015 1050
rect 18485 885 24015 930
rect 18485 765 18510 885
rect 18630 765 18685 885
rect 18805 765 18850 885
rect 18970 765 19015 885
rect 19135 765 19180 885
rect 19300 765 19355 885
rect 19475 765 19520 885
rect 19640 765 19685 885
rect 19805 765 19850 885
rect 19970 765 20025 885
rect 20145 765 20190 885
rect 20310 765 20355 885
rect 20475 765 20520 885
rect 20640 765 20695 885
rect 20815 765 20860 885
rect 20980 765 21025 885
rect 21145 765 21190 885
rect 21310 765 21365 885
rect 21485 765 21530 885
rect 21650 765 21695 885
rect 21815 765 21860 885
rect 21980 765 22035 885
rect 22155 765 22200 885
rect 22320 765 22365 885
rect 22485 765 22530 885
rect 22650 765 22705 885
rect 22825 765 22870 885
rect 22990 765 23035 885
rect 23155 765 23200 885
rect 23320 765 23375 885
rect 23495 765 23540 885
rect 23660 765 23705 885
rect 23825 765 23870 885
rect 23990 765 24015 885
rect 18485 710 24015 765
rect 18485 590 18510 710
rect 18630 590 18685 710
rect 18805 590 18850 710
rect 18970 590 19015 710
rect 19135 590 19180 710
rect 19300 590 19355 710
rect 19475 590 19520 710
rect 19640 590 19685 710
rect 19805 590 19850 710
rect 19970 590 20025 710
rect 20145 590 20190 710
rect 20310 590 20355 710
rect 20475 590 20520 710
rect 20640 590 20695 710
rect 20815 590 20860 710
rect 20980 590 21025 710
rect 21145 590 21190 710
rect 21310 590 21365 710
rect 21485 590 21530 710
rect 21650 590 21695 710
rect 21815 590 21860 710
rect 21980 590 22035 710
rect 22155 590 22200 710
rect 22320 590 22365 710
rect 22485 590 22530 710
rect 22650 590 22705 710
rect 22825 590 22870 710
rect 22990 590 23035 710
rect 23155 590 23200 710
rect 23320 590 23375 710
rect 23495 590 23540 710
rect 23660 590 23705 710
rect 23825 590 23870 710
rect 23990 590 24015 710
rect 18485 545 24015 590
rect 18485 425 18510 545
rect 18630 425 18685 545
rect 18805 425 18850 545
rect 18970 425 19015 545
rect 19135 425 19180 545
rect 19300 425 19355 545
rect 19475 425 19520 545
rect 19640 425 19685 545
rect 19805 425 19850 545
rect 19970 425 20025 545
rect 20145 425 20190 545
rect 20310 425 20355 545
rect 20475 425 20520 545
rect 20640 425 20695 545
rect 20815 425 20860 545
rect 20980 425 21025 545
rect 21145 425 21190 545
rect 21310 425 21365 545
rect 21485 425 21530 545
rect 21650 425 21695 545
rect 21815 425 21860 545
rect 21980 425 22035 545
rect 22155 425 22200 545
rect 22320 425 22365 545
rect 22485 425 22530 545
rect 22650 425 22705 545
rect 22825 425 22870 545
rect 22990 425 23035 545
rect 23155 425 23200 545
rect 23320 425 23375 545
rect 23495 425 23540 545
rect 23660 425 23705 545
rect 23825 425 23870 545
rect 23990 425 24015 545
rect 18485 380 24015 425
rect 18485 260 18510 380
rect 18630 260 18685 380
rect 18805 260 18850 380
rect 18970 260 19015 380
rect 19135 260 19180 380
rect 19300 260 19355 380
rect 19475 260 19520 380
rect 19640 260 19685 380
rect 19805 260 19850 380
rect 19970 260 20025 380
rect 20145 260 20190 380
rect 20310 260 20355 380
rect 20475 260 20520 380
rect 20640 260 20695 380
rect 20815 260 20860 380
rect 20980 260 21025 380
rect 21145 260 21190 380
rect 21310 260 21365 380
rect 21485 260 21530 380
rect 21650 260 21695 380
rect 21815 260 21860 380
rect 21980 260 22035 380
rect 22155 260 22200 380
rect 22320 260 22365 380
rect 22485 260 22530 380
rect 22650 260 22705 380
rect 22825 260 22870 380
rect 22990 260 23035 380
rect 23155 260 23200 380
rect 23320 260 23375 380
rect 23495 260 23540 380
rect 23660 260 23705 380
rect 23825 260 23870 380
rect 23990 260 24015 380
rect 18485 215 24015 260
rect 18485 95 18510 215
rect 18630 95 18685 215
rect 18805 95 18850 215
rect 18970 95 19015 215
rect 19135 95 19180 215
rect 19300 95 19355 215
rect 19475 95 19520 215
rect 19640 95 19685 215
rect 19805 95 19850 215
rect 19970 95 20025 215
rect 20145 95 20190 215
rect 20310 95 20355 215
rect 20475 95 20520 215
rect 20640 95 20695 215
rect 20815 95 20860 215
rect 20980 95 21025 215
rect 21145 95 21190 215
rect 21310 95 21365 215
rect 21485 95 21530 215
rect 21650 95 21695 215
rect 21815 95 21860 215
rect 21980 95 22035 215
rect 22155 95 22200 215
rect 22320 95 22365 215
rect 22485 95 22530 215
rect 22650 95 22705 215
rect 22825 95 22870 215
rect 22990 95 23035 215
rect 23155 95 23200 215
rect 23320 95 23375 215
rect 23495 95 23540 215
rect 23660 95 23705 215
rect 23825 95 23870 215
rect 23990 95 24015 215
rect 18485 40 24015 95
rect 18485 -80 18510 40
rect 18630 -80 18685 40
rect 18805 -80 18850 40
rect 18970 -80 19015 40
rect 19135 -80 19180 40
rect 19300 -80 19355 40
rect 19475 -80 19520 40
rect 19640 -80 19685 40
rect 19805 -80 19850 40
rect 19970 -80 20025 40
rect 20145 -80 20190 40
rect 20310 -80 20355 40
rect 20475 -80 20520 40
rect 20640 -80 20695 40
rect 20815 -80 20860 40
rect 20980 -80 21025 40
rect 21145 -80 21190 40
rect 21310 -80 21365 40
rect 21485 -80 21530 40
rect 21650 -80 21695 40
rect 21815 -80 21860 40
rect 21980 -80 22035 40
rect 22155 -80 22200 40
rect 22320 -80 22365 40
rect 22485 -80 22530 40
rect 22650 -80 22705 40
rect 22825 -80 22870 40
rect 22990 -80 23035 40
rect 23155 -80 23200 40
rect 23320 -80 23375 40
rect 23495 -80 23540 40
rect 23660 -80 23705 40
rect 23825 -80 23870 40
rect 23990 -80 24015 40
rect 18485 -125 24015 -80
rect 18485 -245 18510 -125
rect 18630 -245 18685 -125
rect 18805 -245 18850 -125
rect 18970 -245 19015 -125
rect 19135 -245 19180 -125
rect 19300 -245 19355 -125
rect 19475 -245 19520 -125
rect 19640 -245 19685 -125
rect 19805 -245 19850 -125
rect 19970 -245 20025 -125
rect 20145 -245 20190 -125
rect 20310 -245 20355 -125
rect 20475 -245 20520 -125
rect 20640 -245 20695 -125
rect 20815 -245 20860 -125
rect 20980 -245 21025 -125
rect 21145 -245 21190 -125
rect 21310 -245 21365 -125
rect 21485 -245 21530 -125
rect 21650 -245 21695 -125
rect 21815 -245 21860 -125
rect 21980 -245 22035 -125
rect 22155 -245 22200 -125
rect 22320 -245 22365 -125
rect 22485 -245 22530 -125
rect 22650 -245 22705 -125
rect 22825 -245 22870 -125
rect 22990 -245 23035 -125
rect 23155 -245 23200 -125
rect 23320 -245 23375 -125
rect 23495 -245 23540 -125
rect 23660 -245 23705 -125
rect 23825 -245 23870 -125
rect 23990 -245 24015 -125
rect 18485 -290 24015 -245
rect 18485 -410 18510 -290
rect 18630 -410 18685 -290
rect 18805 -410 18850 -290
rect 18970 -410 19015 -290
rect 19135 -410 19180 -290
rect 19300 -410 19355 -290
rect 19475 -410 19520 -290
rect 19640 -410 19685 -290
rect 19805 -410 19850 -290
rect 19970 -410 20025 -290
rect 20145 -410 20190 -290
rect 20310 -410 20355 -290
rect 20475 -410 20520 -290
rect 20640 -410 20695 -290
rect 20815 -410 20860 -290
rect 20980 -410 21025 -290
rect 21145 -410 21190 -290
rect 21310 -410 21365 -290
rect 21485 -410 21530 -290
rect 21650 -410 21695 -290
rect 21815 -410 21860 -290
rect 21980 -410 22035 -290
rect 22155 -410 22200 -290
rect 22320 -410 22365 -290
rect 22485 -410 22530 -290
rect 22650 -410 22705 -290
rect 22825 -410 22870 -290
rect 22990 -410 23035 -290
rect 23155 -410 23200 -290
rect 23320 -410 23375 -290
rect 23495 -410 23540 -290
rect 23660 -410 23705 -290
rect 23825 -410 23870 -290
rect 23990 -410 24015 -290
rect 18485 -455 24015 -410
rect 18485 -575 18510 -455
rect 18630 -575 18685 -455
rect 18805 -575 18850 -455
rect 18970 -575 19015 -455
rect 19135 -575 19180 -455
rect 19300 -575 19355 -455
rect 19475 -575 19520 -455
rect 19640 -575 19685 -455
rect 19805 -575 19850 -455
rect 19970 -575 20025 -455
rect 20145 -575 20190 -455
rect 20310 -575 20355 -455
rect 20475 -575 20520 -455
rect 20640 -575 20695 -455
rect 20815 -575 20860 -455
rect 20980 -575 21025 -455
rect 21145 -575 21190 -455
rect 21310 -575 21365 -455
rect 21485 -575 21530 -455
rect 21650 -575 21695 -455
rect 21815 -575 21860 -455
rect 21980 -575 22035 -455
rect 22155 -575 22200 -455
rect 22320 -575 22365 -455
rect 22485 -575 22530 -455
rect 22650 -575 22705 -455
rect 22825 -575 22870 -455
rect 22990 -575 23035 -455
rect 23155 -575 23200 -455
rect 23320 -575 23375 -455
rect 23495 -575 23540 -455
rect 23660 -575 23705 -455
rect 23825 -575 23870 -455
rect 23990 -575 24015 -455
rect 18485 -630 24015 -575
rect 18485 -750 18510 -630
rect 18630 -750 18685 -630
rect 18805 -750 18850 -630
rect 18970 -750 19015 -630
rect 19135 -750 19180 -630
rect 19300 -750 19355 -630
rect 19475 -750 19520 -630
rect 19640 -750 19685 -630
rect 19805 -750 19850 -630
rect 19970 -750 20025 -630
rect 20145 -750 20190 -630
rect 20310 -750 20355 -630
rect 20475 -750 20520 -630
rect 20640 -750 20695 -630
rect 20815 -750 20860 -630
rect 20980 -750 21025 -630
rect 21145 -750 21190 -630
rect 21310 -750 21365 -630
rect 21485 -750 21530 -630
rect 21650 -750 21695 -630
rect 21815 -750 21860 -630
rect 21980 -750 22035 -630
rect 22155 -750 22200 -630
rect 22320 -750 22365 -630
rect 22485 -750 22530 -630
rect 22650 -750 22705 -630
rect 22825 -750 22870 -630
rect 22990 -750 23035 -630
rect 23155 -750 23200 -630
rect 23320 -750 23375 -630
rect 23495 -750 23540 -630
rect 23660 -750 23705 -630
rect 23825 -750 23870 -630
rect 23990 -750 24015 -630
rect 18485 -795 24015 -750
rect 18485 -915 18510 -795
rect 18630 -915 18685 -795
rect 18805 -915 18850 -795
rect 18970 -915 19015 -795
rect 19135 -915 19180 -795
rect 19300 -915 19355 -795
rect 19475 -915 19520 -795
rect 19640 -915 19685 -795
rect 19805 -915 19850 -795
rect 19970 -915 20025 -795
rect 20145 -915 20190 -795
rect 20310 -915 20355 -795
rect 20475 -915 20520 -795
rect 20640 -915 20695 -795
rect 20815 -915 20860 -795
rect 20980 -915 21025 -795
rect 21145 -915 21190 -795
rect 21310 -915 21365 -795
rect 21485 -915 21530 -795
rect 21650 -915 21695 -795
rect 21815 -915 21860 -795
rect 21980 -915 22035 -795
rect 22155 -915 22200 -795
rect 22320 -915 22365 -795
rect 22485 -915 22530 -795
rect 22650 -915 22705 -795
rect 22825 -915 22870 -795
rect 22990 -915 23035 -795
rect 23155 -915 23200 -795
rect 23320 -915 23375 -795
rect 23495 -915 23540 -795
rect 23660 -915 23705 -795
rect 23825 -915 23870 -795
rect 23990 -915 24015 -795
rect 18485 -960 24015 -915
rect 18485 -1080 18510 -960
rect 18630 -1080 18685 -960
rect 18805 -1080 18850 -960
rect 18970 -1080 19015 -960
rect 19135 -1080 19180 -960
rect 19300 -1080 19355 -960
rect 19475 -1080 19520 -960
rect 19640 -1080 19685 -960
rect 19805 -1080 19850 -960
rect 19970 -1080 20025 -960
rect 20145 -1080 20190 -960
rect 20310 -1080 20355 -960
rect 20475 -1080 20520 -960
rect 20640 -1080 20695 -960
rect 20815 -1080 20860 -960
rect 20980 -1080 21025 -960
rect 21145 -1080 21190 -960
rect 21310 -1080 21365 -960
rect 21485 -1080 21530 -960
rect 21650 -1080 21695 -960
rect 21815 -1080 21860 -960
rect 21980 -1080 22035 -960
rect 22155 -1080 22200 -960
rect 22320 -1080 22365 -960
rect 22485 -1080 22530 -960
rect 22650 -1080 22705 -960
rect 22825 -1080 22870 -960
rect 22990 -1080 23035 -960
rect 23155 -1080 23200 -960
rect 23320 -1080 23375 -960
rect 23495 -1080 23540 -960
rect 23660 -1080 23705 -960
rect 23825 -1080 23870 -960
rect 23990 -1080 24015 -960
rect 18485 -1125 24015 -1080
rect 18485 -1245 18510 -1125
rect 18630 -1245 18685 -1125
rect 18805 -1245 18850 -1125
rect 18970 -1245 19015 -1125
rect 19135 -1245 19180 -1125
rect 19300 -1245 19355 -1125
rect 19475 -1245 19520 -1125
rect 19640 -1245 19685 -1125
rect 19805 -1245 19850 -1125
rect 19970 -1245 20025 -1125
rect 20145 -1245 20190 -1125
rect 20310 -1245 20355 -1125
rect 20475 -1245 20520 -1125
rect 20640 -1245 20695 -1125
rect 20815 -1245 20860 -1125
rect 20980 -1245 21025 -1125
rect 21145 -1245 21190 -1125
rect 21310 -1245 21365 -1125
rect 21485 -1245 21530 -1125
rect 21650 -1245 21695 -1125
rect 21815 -1245 21860 -1125
rect 21980 -1245 22035 -1125
rect 22155 -1245 22200 -1125
rect 22320 -1245 22365 -1125
rect 22485 -1245 22530 -1125
rect 22650 -1245 22705 -1125
rect 22825 -1245 22870 -1125
rect 22990 -1245 23035 -1125
rect 23155 -1245 23200 -1125
rect 23320 -1245 23375 -1125
rect 23495 -1245 23540 -1125
rect 23660 -1245 23705 -1125
rect 23825 -1245 23870 -1125
rect 23990 -1245 24015 -1125
rect 18485 -1300 24015 -1245
rect 18485 -1420 18510 -1300
rect 18630 -1420 18685 -1300
rect 18805 -1420 18850 -1300
rect 18970 -1420 19015 -1300
rect 19135 -1420 19180 -1300
rect 19300 -1420 19355 -1300
rect 19475 -1420 19520 -1300
rect 19640 -1420 19685 -1300
rect 19805 -1420 19850 -1300
rect 19970 -1420 20025 -1300
rect 20145 -1420 20190 -1300
rect 20310 -1420 20355 -1300
rect 20475 -1420 20520 -1300
rect 20640 -1420 20695 -1300
rect 20815 -1420 20860 -1300
rect 20980 -1420 21025 -1300
rect 21145 -1420 21190 -1300
rect 21310 -1420 21365 -1300
rect 21485 -1420 21530 -1300
rect 21650 -1420 21695 -1300
rect 21815 -1420 21860 -1300
rect 21980 -1420 22035 -1300
rect 22155 -1420 22200 -1300
rect 22320 -1420 22365 -1300
rect 22485 -1420 22530 -1300
rect 22650 -1420 22705 -1300
rect 22825 -1420 22870 -1300
rect 22990 -1420 23035 -1300
rect 23155 -1420 23200 -1300
rect 23320 -1420 23375 -1300
rect 23495 -1420 23540 -1300
rect 23660 -1420 23705 -1300
rect 23825 -1420 23870 -1300
rect 23990 -1420 24015 -1300
rect 18485 -1465 24015 -1420
rect 18485 -1585 18510 -1465
rect 18630 -1585 18685 -1465
rect 18805 -1585 18850 -1465
rect 18970 -1585 19015 -1465
rect 19135 -1585 19180 -1465
rect 19300 -1585 19355 -1465
rect 19475 -1585 19520 -1465
rect 19640 -1585 19685 -1465
rect 19805 -1585 19850 -1465
rect 19970 -1585 20025 -1465
rect 20145 -1585 20190 -1465
rect 20310 -1585 20355 -1465
rect 20475 -1585 20520 -1465
rect 20640 -1585 20695 -1465
rect 20815 -1585 20860 -1465
rect 20980 -1585 21025 -1465
rect 21145 -1585 21190 -1465
rect 21310 -1585 21365 -1465
rect 21485 -1585 21530 -1465
rect 21650 -1585 21695 -1465
rect 21815 -1585 21860 -1465
rect 21980 -1585 22035 -1465
rect 22155 -1585 22200 -1465
rect 22320 -1585 22365 -1465
rect 22485 -1585 22530 -1465
rect 22650 -1585 22705 -1465
rect 22825 -1585 22870 -1465
rect 22990 -1585 23035 -1465
rect 23155 -1585 23200 -1465
rect 23320 -1585 23375 -1465
rect 23495 -1585 23540 -1465
rect 23660 -1585 23705 -1465
rect 23825 -1585 23870 -1465
rect 23990 -1585 24015 -1465
rect 18485 -1630 24015 -1585
rect 18485 -1750 18510 -1630
rect 18630 -1750 18685 -1630
rect 18805 -1750 18850 -1630
rect 18970 -1750 19015 -1630
rect 19135 -1750 19180 -1630
rect 19300 -1750 19355 -1630
rect 19475 -1750 19520 -1630
rect 19640 -1750 19685 -1630
rect 19805 -1750 19850 -1630
rect 19970 -1750 20025 -1630
rect 20145 -1750 20190 -1630
rect 20310 -1750 20355 -1630
rect 20475 -1750 20520 -1630
rect 20640 -1750 20695 -1630
rect 20815 -1750 20860 -1630
rect 20980 -1750 21025 -1630
rect 21145 -1750 21190 -1630
rect 21310 -1750 21365 -1630
rect 21485 -1750 21530 -1630
rect 21650 -1750 21695 -1630
rect 21815 -1750 21860 -1630
rect 21980 -1750 22035 -1630
rect 22155 -1750 22200 -1630
rect 22320 -1750 22365 -1630
rect 22485 -1750 22530 -1630
rect 22650 -1750 22705 -1630
rect 22825 -1750 22870 -1630
rect 22990 -1750 23035 -1630
rect 23155 -1750 23200 -1630
rect 23320 -1750 23375 -1630
rect 23495 -1750 23540 -1630
rect 23660 -1750 23705 -1630
rect 23825 -1750 23870 -1630
rect 23990 -1750 24015 -1630
rect 18485 -1795 24015 -1750
rect 18485 -1915 18510 -1795
rect 18630 -1915 18685 -1795
rect 18805 -1915 18850 -1795
rect 18970 -1915 19015 -1795
rect 19135 -1915 19180 -1795
rect 19300 -1915 19355 -1795
rect 19475 -1915 19520 -1795
rect 19640 -1915 19685 -1795
rect 19805 -1915 19850 -1795
rect 19970 -1915 20025 -1795
rect 20145 -1915 20190 -1795
rect 20310 -1915 20355 -1795
rect 20475 -1915 20520 -1795
rect 20640 -1915 20695 -1795
rect 20815 -1915 20860 -1795
rect 20980 -1915 21025 -1795
rect 21145 -1915 21190 -1795
rect 21310 -1915 21365 -1795
rect 21485 -1915 21530 -1795
rect 21650 -1915 21695 -1795
rect 21815 -1915 21860 -1795
rect 21980 -1915 22035 -1795
rect 22155 -1915 22200 -1795
rect 22320 -1915 22365 -1795
rect 22485 -1915 22530 -1795
rect 22650 -1915 22705 -1795
rect 22825 -1915 22870 -1795
rect 22990 -1915 23035 -1795
rect 23155 -1915 23200 -1795
rect 23320 -1915 23375 -1795
rect 23495 -1915 23540 -1795
rect 23660 -1915 23705 -1795
rect 23825 -1915 23870 -1795
rect 23990 -1915 24015 -1795
rect 18485 -1970 24015 -1915
rect 18485 -2090 18510 -1970
rect 18630 -2090 18685 -1970
rect 18805 -2090 18850 -1970
rect 18970 -2090 19015 -1970
rect 19135 -2090 19180 -1970
rect 19300 -2090 19355 -1970
rect 19475 -2090 19520 -1970
rect 19640 -2090 19685 -1970
rect 19805 -2090 19850 -1970
rect 19970 -2090 20025 -1970
rect 20145 -2090 20190 -1970
rect 20310 -2090 20355 -1970
rect 20475 -2090 20520 -1970
rect 20640 -2090 20695 -1970
rect 20815 -2090 20860 -1970
rect 20980 -2090 21025 -1970
rect 21145 -2090 21190 -1970
rect 21310 -2090 21365 -1970
rect 21485 -2090 21530 -1970
rect 21650 -2090 21695 -1970
rect 21815 -2090 21860 -1970
rect 21980 -2090 22035 -1970
rect 22155 -2090 22200 -1970
rect 22320 -2090 22365 -1970
rect 22485 -2090 22530 -1970
rect 22650 -2090 22705 -1970
rect 22825 -2090 22870 -1970
rect 22990 -2090 23035 -1970
rect 23155 -2090 23200 -1970
rect 23320 -2090 23375 -1970
rect 23495 -2090 23540 -1970
rect 23660 -2090 23705 -1970
rect 23825 -2090 23870 -1970
rect 23990 -2090 24015 -1970
rect 18485 -2135 24015 -2090
rect 18485 -2255 18510 -2135
rect 18630 -2255 18685 -2135
rect 18805 -2255 18850 -2135
rect 18970 -2255 19015 -2135
rect 19135 -2255 19180 -2135
rect 19300 -2255 19355 -2135
rect 19475 -2255 19520 -2135
rect 19640 -2255 19685 -2135
rect 19805 -2255 19850 -2135
rect 19970 -2255 20025 -2135
rect 20145 -2255 20190 -2135
rect 20310 -2255 20355 -2135
rect 20475 -2255 20520 -2135
rect 20640 -2255 20695 -2135
rect 20815 -2255 20860 -2135
rect 20980 -2255 21025 -2135
rect 21145 -2255 21190 -2135
rect 21310 -2255 21365 -2135
rect 21485 -2255 21530 -2135
rect 21650 -2255 21695 -2135
rect 21815 -2255 21860 -2135
rect 21980 -2255 22035 -2135
rect 22155 -2255 22200 -2135
rect 22320 -2255 22365 -2135
rect 22485 -2255 22530 -2135
rect 22650 -2255 22705 -2135
rect 22825 -2255 22870 -2135
rect 22990 -2255 23035 -2135
rect 23155 -2255 23200 -2135
rect 23320 -2255 23375 -2135
rect 23495 -2255 23540 -2135
rect 23660 -2255 23705 -2135
rect 23825 -2255 23870 -2135
rect 23990 -2255 24015 -2135
rect 18485 -2300 24015 -2255
rect 18485 -2420 18510 -2300
rect 18630 -2420 18685 -2300
rect 18805 -2420 18850 -2300
rect 18970 -2420 19015 -2300
rect 19135 -2420 19180 -2300
rect 19300 -2420 19355 -2300
rect 19475 -2420 19520 -2300
rect 19640 -2420 19685 -2300
rect 19805 -2420 19850 -2300
rect 19970 -2420 20025 -2300
rect 20145 -2420 20190 -2300
rect 20310 -2420 20355 -2300
rect 20475 -2420 20520 -2300
rect 20640 -2420 20695 -2300
rect 20815 -2420 20860 -2300
rect 20980 -2420 21025 -2300
rect 21145 -2420 21190 -2300
rect 21310 -2420 21365 -2300
rect 21485 -2420 21530 -2300
rect 21650 -2420 21695 -2300
rect 21815 -2420 21860 -2300
rect 21980 -2420 22035 -2300
rect 22155 -2420 22200 -2300
rect 22320 -2420 22365 -2300
rect 22485 -2420 22530 -2300
rect 22650 -2420 22705 -2300
rect 22825 -2420 22870 -2300
rect 22990 -2420 23035 -2300
rect 23155 -2420 23200 -2300
rect 23320 -2420 23375 -2300
rect 23495 -2420 23540 -2300
rect 23660 -2420 23705 -2300
rect 23825 -2420 23870 -2300
rect 23990 -2420 24015 -2300
rect 18485 -2465 24015 -2420
rect 18485 -2585 18510 -2465
rect 18630 -2585 18685 -2465
rect 18805 -2585 18850 -2465
rect 18970 -2585 19015 -2465
rect 19135 -2585 19180 -2465
rect 19300 -2585 19355 -2465
rect 19475 -2585 19520 -2465
rect 19640 -2585 19685 -2465
rect 19805 -2585 19850 -2465
rect 19970 -2585 20025 -2465
rect 20145 -2585 20190 -2465
rect 20310 -2585 20355 -2465
rect 20475 -2585 20520 -2465
rect 20640 -2585 20695 -2465
rect 20815 -2585 20860 -2465
rect 20980 -2585 21025 -2465
rect 21145 -2585 21190 -2465
rect 21310 -2585 21365 -2465
rect 21485 -2585 21530 -2465
rect 21650 -2585 21695 -2465
rect 21815 -2585 21860 -2465
rect 21980 -2585 22035 -2465
rect 22155 -2585 22200 -2465
rect 22320 -2585 22365 -2465
rect 22485 -2585 22530 -2465
rect 22650 -2585 22705 -2465
rect 22825 -2585 22870 -2465
rect 22990 -2585 23035 -2465
rect 23155 -2585 23200 -2465
rect 23320 -2585 23375 -2465
rect 23495 -2585 23540 -2465
rect 23660 -2585 23705 -2465
rect 23825 -2585 23870 -2465
rect 23990 -2585 24015 -2465
rect 18485 -2640 24015 -2585
rect 18485 -2760 18510 -2640
rect 18630 -2760 18685 -2640
rect 18805 -2760 18850 -2640
rect 18970 -2760 19015 -2640
rect 19135 -2760 19180 -2640
rect 19300 -2760 19355 -2640
rect 19475 -2760 19520 -2640
rect 19640 -2760 19685 -2640
rect 19805 -2760 19850 -2640
rect 19970 -2760 20025 -2640
rect 20145 -2760 20190 -2640
rect 20310 -2760 20355 -2640
rect 20475 -2760 20520 -2640
rect 20640 -2760 20695 -2640
rect 20815 -2760 20860 -2640
rect 20980 -2760 21025 -2640
rect 21145 -2760 21190 -2640
rect 21310 -2760 21365 -2640
rect 21485 -2760 21530 -2640
rect 21650 -2760 21695 -2640
rect 21815 -2760 21860 -2640
rect 21980 -2760 22035 -2640
rect 22155 -2760 22200 -2640
rect 22320 -2760 22365 -2640
rect 22485 -2760 22530 -2640
rect 22650 -2760 22705 -2640
rect 22825 -2760 22870 -2640
rect 22990 -2760 23035 -2640
rect 23155 -2760 23200 -2640
rect 23320 -2760 23375 -2640
rect 23495 -2760 23540 -2640
rect 23660 -2760 23705 -2640
rect 23825 -2760 23870 -2640
rect 23990 -2760 24015 -2640
rect 18485 -2805 24015 -2760
rect 18485 -2925 18510 -2805
rect 18630 -2925 18685 -2805
rect 18805 -2925 18850 -2805
rect 18970 -2925 19015 -2805
rect 19135 -2925 19180 -2805
rect 19300 -2925 19355 -2805
rect 19475 -2925 19520 -2805
rect 19640 -2925 19685 -2805
rect 19805 -2925 19850 -2805
rect 19970 -2925 20025 -2805
rect 20145 -2925 20190 -2805
rect 20310 -2925 20355 -2805
rect 20475 -2925 20520 -2805
rect 20640 -2925 20695 -2805
rect 20815 -2925 20860 -2805
rect 20980 -2925 21025 -2805
rect 21145 -2925 21190 -2805
rect 21310 -2925 21365 -2805
rect 21485 -2925 21530 -2805
rect 21650 -2925 21695 -2805
rect 21815 -2925 21860 -2805
rect 21980 -2925 22035 -2805
rect 22155 -2925 22200 -2805
rect 22320 -2925 22365 -2805
rect 22485 -2925 22530 -2805
rect 22650 -2925 22705 -2805
rect 22825 -2925 22870 -2805
rect 22990 -2925 23035 -2805
rect 23155 -2925 23200 -2805
rect 23320 -2925 23375 -2805
rect 23495 -2925 23540 -2805
rect 23660 -2925 23705 -2805
rect 23825 -2925 23870 -2805
rect 23990 -2925 24015 -2805
rect 18485 -2970 24015 -2925
rect 18485 -3090 18510 -2970
rect 18630 -3090 18685 -2970
rect 18805 -3090 18850 -2970
rect 18970 -3090 19015 -2970
rect 19135 -3090 19180 -2970
rect 19300 -3090 19355 -2970
rect 19475 -3090 19520 -2970
rect 19640 -3090 19685 -2970
rect 19805 -3090 19850 -2970
rect 19970 -3090 20025 -2970
rect 20145 -3090 20190 -2970
rect 20310 -3090 20355 -2970
rect 20475 -3090 20520 -2970
rect 20640 -3090 20695 -2970
rect 20815 -3090 20860 -2970
rect 20980 -3090 21025 -2970
rect 21145 -3090 21190 -2970
rect 21310 -3090 21365 -2970
rect 21485 -3090 21530 -2970
rect 21650 -3090 21695 -2970
rect 21815 -3090 21860 -2970
rect 21980 -3090 22035 -2970
rect 22155 -3090 22200 -2970
rect 22320 -3090 22365 -2970
rect 22485 -3090 22530 -2970
rect 22650 -3090 22705 -2970
rect 22825 -3090 22870 -2970
rect 22990 -3090 23035 -2970
rect 23155 -3090 23200 -2970
rect 23320 -3090 23375 -2970
rect 23495 -3090 23540 -2970
rect 23660 -3090 23705 -2970
rect 23825 -3090 23870 -2970
rect 23990 -3090 24015 -2970
rect 18485 -3135 24015 -3090
rect 18485 -3255 18510 -3135
rect 18630 -3255 18685 -3135
rect 18805 -3255 18850 -3135
rect 18970 -3255 19015 -3135
rect 19135 -3255 19180 -3135
rect 19300 -3255 19355 -3135
rect 19475 -3255 19520 -3135
rect 19640 -3255 19685 -3135
rect 19805 -3255 19850 -3135
rect 19970 -3255 20025 -3135
rect 20145 -3255 20190 -3135
rect 20310 -3255 20355 -3135
rect 20475 -3255 20520 -3135
rect 20640 -3255 20695 -3135
rect 20815 -3255 20860 -3135
rect 20980 -3255 21025 -3135
rect 21145 -3255 21190 -3135
rect 21310 -3255 21365 -3135
rect 21485 -3255 21530 -3135
rect 21650 -3255 21695 -3135
rect 21815 -3255 21860 -3135
rect 21980 -3255 22035 -3135
rect 22155 -3255 22200 -3135
rect 22320 -3255 22365 -3135
rect 22485 -3255 22530 -3135
rect 22650 -3255 22705 -3135
rect 22825 -3255 22870 -3135
rect 22990 -3255 23035 -3135
rect 23155 -3255 23200 -3135
rect 23320 -3255 23375 -3135
rect 23495 -3255 23540 -3135
rect 23660 -3255 23705 -3135
rect 23825 -3255 23870 -3135
rect 23990 -3255 24015 -3135
rect 18485 -3310 24015 -3255
rect 18485 -3430 18510 -3310
rect 18630 -3430 18685 -3310
rect 18805 -3430 18850 -3310
rect 18970 -3430 19015 -3310
rect 19135 -3430 19180 -3310
rect 19300 -3430 19355 -3310
rect 19475 -3430 19520 -3310
rect 19640 -3430 19685 -3310
rect 19805 -3430 19850 -3310
rect 19970 -3430 20025 -3310
rect 20145 -3430 20190 -3310
rect 20310 -3430 20355 -3310
rect 20475 -3430 20520 -3310
rect 20640 -3430 20695 -3310
rect 20815 -3430 20860 -3310
rect 20980 -3430 21025 -3310
rect 21145 -3430 21190 -3310
rect 21310 -3430 21365 -3310
rect 21485 -3430 21530 -3310
rect 21650 -3430 21695 -3310
rect 21815 -3430 21860 -3310
rect 21980 -3430 22035 -3310
rect 22155 -3430 22200 -3310
rect 22320 -3430 22365 -3310
rect 22485 -3430 22530 -3310
rect 22650 -3430 22705 -3310
rect 22825 -3430 22870 -3310
rect 22990 -3430 23035 -3310
rect 23155 -3430 23200 -3310
rect 23320 -3430 23375 -3310
rect 23495 -3430 23540 -3310
rect 23660 -3430 23705 -3310
rect 23825 -3430 23870 -3310
rect 23990 -3430 24015 -3310
rect 18485 -3475 24015 -3430
rect 18485 -3595 18510 -3475
rect 18630 -3595 18685 -3475
rect 18805 -3595 18850 -3475
rect 18970 -3595 19015 -3475
rect 19135 -3595 19180 -3475
rect 19300 -3595 19355 -3475
rect 19475 -3595 19520 -3475
rect 19640 -3595 19685 -3475
rect 19805 -3595 19850 -3475
rect 19970 -3595 20025 -3475
rect 20145 -3595 20190 -3475
rect 20310 -3595 20355 -3475
rect 20475 -3595 20520 -3475
rect 20640 -3595 20695 -3475
rect 20815 -3595 20860 -3475
rect 20980 -3595 21025 -3475
rect 21145 -3595 21190 -3475
rect 21310 -3595 21365 -3475
rect 21485 -3595 21530 -3475
rect 21650 -3595 21695 -3475
rect 21815 -3595 21860 -3475
rect 21980 -3595 22035 -3475
rect 22155 -3595 22200 -3475
rect 22320 -3595 22365 -3475
rect 22485 -3595 22530 -3475
rect 22650 -3595 22705 -3475
rect 22825 -3595 22870 -3475
rect 22990 -3595 23035 -3475
rect 23155 -3595 23200 -3475
rect 23320 -3595 23375 -3475
rect 23495 -3595 23540 -3475
rect 23660 -3595 23705 -3475
rect 23825 -3595 23870 -3475
rect 23990 -3595 24015 -3475
rect 18485 -3640 24015 -3595
rect 18485 -3760 18510 -3640
rect 18630 -3760 18685 -3640
rect 18805 -3760 18850 -3640
rect 18970 -3760 19015 -3640
rect 19135 -3760 19180 -3640
rect 19300 -3760 19355 -3640
rect 19475 -3760 19520 -3640
rect 19640 -3760 19685 -3640
rect 19805 -3760 19850 -3640
rect 19970 -3760 20025 -3640
rect 20145 -3760 20190 -3640
rect 20310 -3760 20355 -3640
rect 20475 -3760 20520 -3640
rect 20640 -3760 20695 -3640
rect 20815 -3760 20860 -3640
rect 20980 -3760 21025 -3640
rect 21145 -3760 21190 -3640
rect 21310 -3760 21365 -3640
rect 21485 -3760 21530 -3640
rect 21650 -3760 21695 -3640
rect 21815 -3760 21860 -3640
rect 21980 -3760 22035 -3640
rect 22155 -3760 22200 -3640
rect 22320 -3760 22365 -3640
rect 22485 -3760 22530 -3640
rect 22650 -3760 22705 -3640
rect 22825 -3760 22870 -3640
rect 22990 -3760 23035 -3640
rect 23155 -3760 23200 -3640
rect 23320 -3760 23375 -3640
rect 23495 -3760 23540 -3640
rect 23660 -3760 23705 -3640
rect 23825 -3760 23870 -3640
rect 23990 -3760 24015 -3640
rect 18485 -3805 24015 -3760
rect 18485 -3925 18510 -3805
rect 18630 -3925 18685 -3805
rect 18805 -3925 18850 -3805
rect 18970 -3925 19015 -3805
rect 19135 -3925 19180 -3805
rect 19300 -3925 19355 -3805
rect 19475 -3925 19520 -3805
rect 19640 -3925 19685 -3805
rect 19805 -3925 19850 -3805
rect 19970 -3925 20025 -3805
rect 20145 -3925 20190 -3805
rect 20310 -3925 20355 -3805
rect 20475 -3925 20520 -3805
rect 20640 -3925 20695 -3805
rect 20815 -3925 20860 -3805
rect 20980 -3925 21025 -3805
rect 21145 -3925 21190 -3805
rect 21310 -3925 21365 -3805
rect 21485 -3925 21530 -3805
rect 21650 -3925 21695 -3805
rect 21815 -3925 21860 -3805
rect 21980 -3925 22035 -3805
rect 22155 -3925 22200 -3805
rect 22320 -3925 22365 -3805
rect 22485 -3925 22530 -3805
rect 22650 -3925 22705 -3805
rect 22825 -3925 22870 -3805
rect 22990 -3925 23035 -3805
rect 23155 -3925 23200 -3805
rect 23320 -3925 23375 -3805
rect 23495 -3925 23540 -3805
rect 23660 -3925 23705 -3805
rect 23825 -3925 23870 -3805
rect 23990 -3925 24015 -3805
rect 18485 -3980 24015 -3925
rect 18485 -4100 18510 -3980
rect 18630 -4100 18685 -3980
rect 18805 -4100 18850 -3980
rect 18970 -4100 19015 -3980
rect 19135 -4100 19180 -3980
rect 19300 -4100 19355 -3980
rect 19475 -4100 19520 -3980
rect 19640 -4100 19685 -3980
rect 19805 -4100 19850 -3980
rect 19970 -4100 20025 -3980
rect 20145 -4100 20190 -3980
rect 20310 -4100 20355 -3980
rect 20475 -4100 20520 -3980
rect 20640 -4100 20695 -3980
rect 20815 -4100 20860 -3980
rect 20980 -4100 21025 -3980
rect 21145 -4100 21190 -3980
rect 21310 -4100 21365 -3980
rect 21485 -4100 21530 -3980
rect 21650 -4100 21695 -3980
rect 21815 -4100 21860 -3980
rect 21980 -4100 22035 -3980
rect 22155 -4100 22200 -3980
rect 22320 -4100 22365 -3980
rect 22485 -4100 22530 -3980
rect 22650 -4100 22705 -3980
rect 22825 -4100 22870 -3980
rect 22990 -4100 23035 -3980
rect 23155 -4100 23200 -3980
rect 23320 -4100 23375 -3980
rect 23495 -4100 23540 -3980
rect 23660 -4100 23705 -3980
rect 23825 -4100 23870 -3980
rect 23990 -4100 24015 -3980
rect 18485 -4125 24015 -4100
rect 24175 1380 29705 1450
rect 24175 1260 24200 1380
rect 24320 1260 24375 1380
rect 24495 1260 24540 1380
rect 24660 1260 24705 1380
rect 24825 1260 24870 1380
rect 24990 1260 25045 1380
rect 25165 1260 25210 1380
rect 25330 1260 25375 1380
rect 25495 1260 25540 1380
rect 25660 1260 25715 1380
rect 25835 1260 25880 1380
rect 26000 1260 26045 1380
rect 26165 1260 26210 1380
rect 26330 1260 26385 1380
rect 26505 1260 26550 1380
rect 26670 1260 26715 1380
rect 26835 1260 26880 1380
rect 27000 1260 27055 1380
rect 27175 1260 27220 1380
rect 27340 1260 27385 1380
rect 27505 1260 27550 1380
rect 27670 1260 27725 1380
rect 27845 1260 27890 1380
rect 28010 1260 28055 1380
rect 28175 1260 28220 1380
rect 28340 1260 28395 1380
rect 28515 1260 28560 1380
rect 28680 1260 28725 1380
rect 28845 1260 28890 1380
rect 29010 1260 29065 1380
rect 29185 1260 29230 1380
rect 29350 1260 29395 1380
rect 29515 1260 29560 1380
rect 29680 1260 29705 1380
rect 24175 1215 29705 1260
rect 24175 1095 24200 1215
rect 24320 1095 24375 1215
rect 24495 1095 24540 1215
rect 24660 1095 24705 1215
rect 24825 1095 24870 1215
rect 24990 1095 25045 1215
rect 25165 1095 25210 1215
rect 25330 1095 25375 1215
rect 25495 1095 25540 1215
rect 25660 1095 25715 1215
rect 25835 1095 25880 1215
rect 26000 1095 26045 1215
rect 26165 1095 26210 1215
rect 26330 1095 26385 1215
rect 26505 1095 26550 1215
rect 26670 1095 26715 1215
rect 26835 1095 26880 1215
rect 27000 1095 27055 1215
rect 27175 1095 27220 1215
rect 27340 1095 27385 1215
rect 27505 1095 27550 1215
rect 27670 1095 27725 1215
rect 27845 1095 27890 1215
rect 28010 1095 28055 1215
rect 28175 1095 28220 1215
rect 28340 1095 28395 1215
rect 28515 1095 28560 1215
rect 28680 1095 28725 1215
rect 28845 1095 28890 1215
rect 29010 1095 29065 1215
rect 29185 1095 29230 1215
rect 29350 1095 29395 1215
rect 29515 1095 29560 1215
rect 29680 1095 29705 1215
rect 24175 1050 29705 1095
rect 24175 930 24200 1050
rect 24320 930 24375 1050
rect 24495 930 24540 1050
rect 24660 930 24705 1050
rect 24825 930 24870 1050
rect 24990 930 25045 1050
rect 25165 930 25210 1050
rect 25330 930 25375 1050
rect 25495 930 25540 1050
rect 25660 930 25715 1050
rect 25835 930 25880 1050
rect 26000 930 26045 1050
rect 26165 930 26210 1050
rect 26330 930 26385 1050
rect 26505 930 26550 1050
rect 26670 930 26715 1050
rect 26835 930 26880 1050
rect 27000 930 27055 1050
rect 27175 930 27220 1050
rect 27340 930 27385 1050
rect 27505 930 27550 1050
rect 27670 930 27725 1050
rect 27845 930 27890 1050
rect 28010 930 28055 1050
rect 28175 930 28220 1050
rect 28340 930 28395 1050
rect 28515 930 28560 1050
rect 28680 930 28725 1050
rect 28845 930 28890 1050
rect 29010 930 29065 1050
rect 29185 930 29230 1050
rect 29350 930 29395 1050
rect 29515 930 29560 1050
rect 29680 930 29705 1050
rect 24175 885 29705 930
rect 24175 765 24200 885
rect 24320 765 24375 885
rect 24495 765 24540 885
rect 24660 765 24705 885
rect 24825 765 24870 885
rect 24990 765 25045 885
rect 25165 765 25210 885
rect 25330 765 25375 885
rect 25495 765 25540 885
rect 25660 765 25715 885
rect 25835 765 25880 885
rect 26000 765 26045 885
rect 26165 765 26210 885
rect 26330 765 26385 885
rect 26505 765 26550 885
rect 26670 765 26715 885
rect 26835 765 26880 885
rect 27000 765 27055 885
rect 27175 765 27220 885
rect 27340 765 27385 885
rect 27505 765 27550 885
rect 27670 765 27725 885
rect 27845 765 27890 885
rect 28010 765 28055 885
rect 28175 765 28220 885
rect 28340 765 28395 885
rect 28515 765 28560 885
rect 28680 765 28725 885
rect 28845 765 28890 885
rect 29010 765 29065 885
rect 29185 765 29230 885
rect 29350 765 29395 885
rect 29515 765 29560 885
rect 29680 765 29705 885
rect 24175 710 29705 765
rect 24175 590 24200 710
rect 24320 590 24375 710
rect 24495 590 24540 710
rect 24660 590 24705 710
rect 24825 590 24870 710
rect 24990 590 25045 710
rect 25165 590 25210 710
rect 25330 590 25375 710
rect 25495 590 25540 710
rect 25660 590 25715 710
rect 25835 590 25880 710
rect 26000 590 26045 710
rect 26165 590 26210 710
rect 26330 590 26385 710
rect 26505 590 26550 710
rect 26670 590 26715 710
rect 26835 590 26880 710
rect 27000 590 27055 710
rect 27175 590 27220 710
rect 27340 590 27385 710
rect 27505 590 27550 710
rect 27670 590 27725 710
rect 27845 590 27890 710
rect 28010 590 28055 710
rect 28175 590 28220 710
rect 28340 590 28395 710
rect 28515 590 28560 710
rect 28680 590 28725 710
rect 28845 590 28890 710
rect 29010 590 29065 710
rect 29185 590 29230 710
rect 29350 590 29395 710
rect 29515 590 29560 710
rect 29680 590 29705 710
rect 24175 545 29705 590
rect 24175 425 24200 545
rect 24320 425 24375 545
rect 24495 425 24540 545
rect 24660 425 24705 545
rect 24825 425 24870 545
rect 24990 425 25045 545
rect 25165 425 25210 545
rect 25330 425 25375 545
rect 25495 425 25540 545
rect 25660 425 25715 545
rect 25835 425 25880 545
rect 26000 425 26045 545
rect 26165 425 26210 545
rect 26330 425 26385 545
rect 26505 425 26550 545
rect 26670 425 26715 545
rect 26835 425 26880 545
rect 27000 425 27055 545
rect 27175 425 27220 545
rect 27340 425 27385 545
rect 27505 425 27550 545
rect 27670 425 27725 545
rect 27845 425 27890 545
rect 28010 425 28055 545
rect 28175 425 28220 545
rect 28340 425 28395 545
rect 28515 425 28560 545
rect 28680 425 28725 545
rect 28845 425 28890 545
rect 29010 425 29065 545
rect 29185 425 29230 545
rect 29350 425 29395 545
rect 29515 425 29560 545
rect 29680 425 29705 545
rect 24175 380 29705 425
rect 24175 260 24200 380
rect 24320 260 24375 380
rect 24495 260 24540 380
rect 24660 260 24705 380
rect 24825 260 24870 380
rect 24990 260 25045 380
rect 25165 260 25210 380
rect 25330 260 25375 380
rect 25495 260 25540 380
rect 25660 260 25715 380
rect 25835 260 25880 380
rect 26000 260 26045 380
rect 26165 260 26210 380
rect 26330 260 26385 380
rect 26505 260 26550 380
rect 26670 260 26715 380
rect 26835 260 26880 380
rect 27000 260 27055 380
rect 27175 260 27220 380
rect 27340 260 27385 380
rect 27505 260 27550 380
rect 27670 260 27725 380
rect 27845 260 27890 380
rect 28010 260 28055 380
rect 28175 260 28220 380
rect 28340 260 28395 380
rect 28515 260 28560 380
rect 28680 260 28725 380
rect 28845 260 28890 380
rect 29010 260 29065 380
rect 29185 260 29230 380
rect 29350 260 29395 380
rect 29515 260 29560 380
rect 29680 260 29705 380
rect 24175 215 29705 260
rect 24175 95 24200 215
rect 24320 95 24375 215
rect 24495 95 24540 215
rect 24660 95 24705 215
rect 24825 95 24870 215
rect 24990 95 25045 215
rect 25165 95 25210 215
rect 25330 95 25375 215
rect 25495 95 25540 215
rect 25660 95 25715 215
rect 25835 95 25880 215
rect 26000 95 26045 215
rect 26165 95 26210 215
rect 26330 95 26385 215
rect 26505 95 26550 215
rect 26670 95 26715 215
rect 26835 95 26880 215
rect 27000 95 27055 215
rect 27175 95 27220 215
rect 27340 95 27385 215
rect 27505 95 27550 215
rect 27670 95 27725 215
rect 27845 95 27890 215
rect 28010 95 28055 215
rect 28175 95 28220 215
rect 28340 95 28395 215
rect 28515 95 28560 215
rect 28680 95 28725 215
rect 28845 95 28890 215
rect 29010 95 29065 215
rect 29185 95 29230 215
rect 29350 95 29395 215
rect 29515 95 29560 215
rect 29680 95 29705 215
rect 24175 40 29705 95
rect 24175 -80 24200 40
rect 24320 -80 24375 40
rect 24495 -80 24540 40
rect 24660 -80 24705 40
rect 24825 -80 24870 40
rect 24990 -80 25045 40
rect 25165 -80 25210 40
rect 25330 -80 25375 40
rect 25495 -80 25540 40
rect 25660 -80 25715 40
rect 25835 -80 25880 40
rect 26000 -80 26045 40
rect 26165 -80 26210 40
rect 26330 -80 26385 40
rect 26505 -80 26550 40
rect 26670 -80 26715 40
rect 26835 -80 26880 40
rect 27000 -80 27055 40
rect 27175 -80 27220 40
rect 27340 -80 27385 40
rect 27505 -80 27550 40
rect 27670 -80 27725 40
rect 27845 -80 27890 40
rect 28010 -80 28055 40
rect 28175 -80 28220 40
rect 28340 -80 28395 40
rect 28515 -80 28560 40
rect 28680 -80 28725 40
rect 28845 -80 28890 40
rect 29010 -80 29065 40
rect 29185 -80 29230 40
rect 29350 -80 29395 40
rect 29515 -80 29560 40
rect 29680 -80 29705 40
rect 24175 -125 29705 -80
rect 24175 -245 24200 -125
rect 24320 -245 24375 -125
rect 24495 -245 24540 -125
rect 24660 -245 24705 -125
rect 24825 -245 24870 -125
rect 24990 -245 25045 -125
rect 25165 -245 25210 -125
rect 25330 -245 25375 -125
rect 25495 -245 25540 -125
rect 25660 -245 25715 -125
rect 25835 -245 25880 -125
rect 26000 -245 26045 -125
rect 26165 -245 26210 -125
rect 26330 -245 26385 -125
rect 26505 -245 26550 -125
rect 26670 -245 26715 -125
rect 26835 -245 26880 -125
rect 27000 -245 27055 -125
rect 27175 -245 27220 -125
rect 27340 -245 27385 -125
rect 27505 -245 27550 -125
rect 27670 -245 27725 -125
rect 27845 -245 27890 -125
rect 28010 -245 28055 -125
rect 28175 -245 28220 -125
rect 28340 -245 28395 -125
rect 28515 -245 28560 -125
rect 28680 -245 28725 -125
rect 28845 -245 28890 -125
rect 29010 -245 29065 -125
rect 29185 -245 29230 -125
rect 29350 -245 29395 -125
rect 29515 -245 29560 -125
rect 29680 -245 29705 -125
rect 24175 -290 29705 -245
rect 24175 -410 24200 -290
rect 24320 -410 24375 -290
rect 24495 -410 24540 -290
rect 24660 -410 24705 -290
rect 24825 -410 24870 -290
rect 24990 -410 25045 -290
rect 25165 -410 25210 -290
rect 25330 -410 25375 -290
rect 25495 -410 25540 -290
rect 25660 -410 25715 -290
rect 25835 -410 25880 -290
rect 26000 -410 26045 -290
rect 26165 -410 26210 -290
rect 26330 -410 26385 -290
rect 26505 -410 26550 -290
rect 26670 -410 26715 -290
rect 26835 -410 26880 -290
rect 27000 -410 27055 -290
rect 27175 -410 27220 -290
rect 27340 -410 27385 -290
rect 27505 -410 27550 -290
rect 27670 -410 27725 -290
rect 27845 -410 27890 -290
rect 28010 -410 28055 -290
rect 28175 -410 28220 -290
rect 28340 -410 28395 -290
rect 28515 -410 28560 -290
rect 28680 -410 28725 -290
rect 28845 -410 28890 -290
rect 29010 -410 29065 -290
rect 29185 -410 29230 -290
rect 29350 -410 29395 -290
rect 29515 -410 29560 -290
rect 29680 -410 29705 -290
rect 24175 -455 29705 -410
rect 24175 -575 24200 -455
rect 24320 -575 24375 -455
rect 24495 -575 24540 -455
rect 24660 -575 24705 -455
rect 24825 -575 24870 -455
rect 24990 -575 25045 -455
rect 25165 -575 25210 -455
rect 25330 -575 25375 -455
rect 25495 -575 25540 -455
rect 25660 -575 25715 -455
rect 25835 -575 25880 -455
rect 26000 -575 26045 -455
rect 26165 -575 26210 -455
rect 26330 -575 26385 -455
rect 26505 -575 26550 -455
rect 26670 -575 26715 -455
rect 26835 -575 26880 -455
rect 27000 -575 27055 -455
rect 27175 -575 27220 -455
rect 27340 -575 27385 -455
rect 27505 -575 27550 -455
rect 27670 -575 27725 -455
rect 27845 -575 27890 -455
rect 28010 -575 28055 -455
rect 28175 -575 28220 -455
rect 28340 -575 28395 -455
rect 28515 -575 28560 -455
rect 28680 -575 28725 -455
rect 28845 -575 28890 -455
rect 29010 -575 29065 -455
rect 29185 -575 29230 -455
rect 29350 -575 29395 -455
rect 29515 -575 29560 -455
rect 29680 -575 29705 -455
rect 24175 -630 29705 -575
rect 24175 -750 24200 -630
rect 24320 -750 24375 -630
rect 24495 -750 24540 -630
rect 24660 -750 24705 -630
rect 24825 -750 24870 -630
rect 24990 -750 25045 -630
rect 25165 -750 25210 -630
rect 25330 -750 25375 -630
rect 25495 -750 25540 -630
rect 25660 -750 25715 -630
rect 25835 -750 25880 -630
rect 26000 -750 26045 -630
rect 26165 -750 26210 -630
rect 26330 -750 26385 -630
rect 26505 -750 26550 -630
rect 26670 -750 26715 -630
rect 26835 -750 26880 -630
rect 27000 -750 27055 -630
rect 27175 -750 27220 -630
rect 27340 -750 27385 -630
rect 27505 -750 27550 -630
rect 27670 -750 27725 -630
rect 27845 -750 27890 -630
rect 28010 -750 28055 -630
rect 28175 -750 28220 -630
rect 28340 -750 28395 -630
rect 28515 -750 28560 -630
rect 28680 -750 28725 -630
rect 28845 -750 28890 -630
rect 29010 -750 29065 -630
rect 29185 -750 29230 -630
rect 29350 -750 29395 -630
rect 29515 -750 29560 -630
rect 29680 -750 29705 -630
rect 24175 -795 29705 -750
rect 24175 -915 24200 -795
rect 24320 -915 24375 -795
rect 24495 -915 24540 -795
rect 24660 -915 24705 -795
rect 24825 -915 24870 -795
rect 24990 -915 25045 -795
rect 25165 -915 25210 -795
rect 25330 -915 25375 -795
rect 25495 -915 25540 -795
rect 25660 -915 25715 -795
rect 25835 -915 25880 -795
rect 26000 -915 26045 -795
rect 26165 -915 26210 -795
rect 26330 -915 26385 -795
rect 26505 -915 26550 -795
rect 26670 -915 26715 -795
rect 26835 -915 26880 -795
rect 27000 -915 27055 -795
rect 27175 -915 27220 -795
rect 27340 -915 27385 -795
rect 27505 -915 27550 -795
rect 27670 -915 27725 -795
rect 27845 -915 27890 -795
rect 28010 -915 28055 -795
rect 28175 -915 28220 -795
rect 28340 -915 28395 -795
rect 28515 -915 28560 -795
rect 28680 -915 28725 -795
rect 28845 -915 28890 -795
rect 29010 -915 29065 -795
rect 29185 -915 29230 -795
rect 29350 -915 29395 -795
rect 29515 -915 29560 -795
rect 29680 -915 29705 -795
rect 24175 -960 29705 -915
rect 24175 -1080 24200 -960
rect 24320 -1080 24375 -960
rect 24495 -1080 24540 -960
rect 24660 -1080 24705 -960
rect 24825 -1080 24870 -960
rect 24990 -1080 25045 -960
rect 25165 -1080 25210 -960
rect 25330 -1080 25375 -960
rect 25495 -1080 25540 -960
rect 25660 -1080 25715 -960
rect 25835 -1080 25880 -960
rect 26000 -1080 26045 -960
rect 26165 -1080 26210 -960
rect 26330 -1080 26385 -960
rect 26505 -1080 26550 -960
rect 26670 -1080 26715 -960
rect 26835 -1080 26880 -960
rect 27000 -1080 27055 -960
rect 27175 -1080 27220 -960
rect 27340 -1080 27385 -960
rect 27505 -1080 27550 -960
rect 27670 -1080 27725 -960
rect 27845 -1080 27890 -960
rect 28010 -1080 28055 -960
rect 28175 -1080 28220 -960
rect 28340 -1080 28395 -960
rect 28515 -1080 28560 -960
rect 28680 -1080 28725 -960
rect 28845 -1080 28890 -960
rect 29010 -1080 29065 -960
rect 29185 -1080 29230 -960
rect 29350 -1080 29395 -960
rect 29515 -1080 29560 -960
rect 29680 -1080 29705 -960
rect 24175 -1125 29705 -1080
rect 24175 -1245 24200 -1125
rect 24320 -1245 24375 -1125
rect 24495 -1245 24540 -1125
rect 24660 -1245 24705 -1125
rect 24825 -1245 24870 -1125
rect 24990 -1245 25045 -1125
rect 25165 -1245 25210 -1125
rect 25330 -1245 25375 -1125
rect 25495 -1245 25540 -1125
rect 25660 -1245 25715 -1125
rect 25835 -1245 25880 -1125
rect 26000 -1245 26045 -1125
rect 26165 -1245 26210 -1125
rect 26330 -1245 26385 -1125
rect 26505 -1245 26550 -1125
rect 26670 -1245 26715 -1125
rect 26835 -1245 26880 -1125
rect 27000 -1245 27055 -1125
rect 27175 -1245 27220 -1125
rect 27340 -1245 27385 -1125
rect 27505 -1245 27550 -1125
rect 27670 -1245 27725 -1125
rect 27845 -1245 27890 -1125
rect 28010 -1245 28055 -1125
rect 28175 -1245 28220 -1125
rect 28340 -1245 28395 -1125
rect 28515 -1245 28560 -1125
rect 28680 -1245 28725 -1125
rect 28845 -1245 28890 -1125
rect 29010 -1245 29065 -1125
rect 29185 -1245 29230 -1125
rect 29350 -1245 29395 -1125
rect 29515 -1245 29560 -1125
rect 29680 -1245 29705 -1125
rect 24175 -1300 29705 -1245
rect 24175 -1420 24200 -1300
rect 24320 -1420 24375 -1300
rect 24495 -1420 24540 -1300
rect 24660 -1420 24705 -1300
rect 24825 -1420 24870 -1300
rect 24990 -1420 25045 -1300
rect 25165 -1420 25210 -1300
rect 25330 -1420 25375 -1300
rect 25495 -1420 25540 -1300
rect 25660 -1420 25715 -1300
rect 25835 -1420 25880 -1300
rect 26000 -1420 26045 -1300
rect 26165 -1420 26210 -1300
rect 26330 -1420 26385 -1300
rect 26505 -1420 26550 -1300
rect 26670 -1420 26715 -1300
rect 26835 -1420 26880 -1300
rect 27000 -1420 27055 -1300
rect 27175 -1420 27220 -1300
rect 27340 -1420 27385 -1300
rect 27505 -1420 27550 -1300
rect 27670 -1420 27725 -1300
rect 27845 -1420 27890 -1300
rect 28010 -1420 28055 -1300
rect 28175 -1420 28220 -1300
rect 28340 -1420 28395 -1300
rect 28515 -1420 28560 -1300
rect 28680 -1420 28725 -1300
rect 28845 -1420 28890 -1300
rect 29010 -1420 29065 -1300
rect 29185 -1420 29230 -1300
rect 29350 -1420 29395 -1300
rect 29515 -1420 29560 -1300
rect 29680 -1420 29705 -1300
rect 24175 -1465 29705 -1420
rect 24175 -1585 24200 -1465
rect 24320 -1585 24375 -1465
rect 24495 -1585 24540 -1465
rect 24660 -1585 24705 -1465
rect 24825 -1585 24870 -1465
rect 24990 -1585 25045 -1465
rect 25165 -1585 25210 -1465
rect 25330 -1585 25375 -1465
rect 25495 -1585 25540 -1465
rect 25660 -1585 25715 -1465
rect 25835 -1585 25880 -1465
rect 26000 -1585 26045 -1465
rect 26165 -1585 26210 -1465
rect 26330 -1585 26385 -1465
rect 26505 -1585 26550 -1465
rect 26670 -1585 26715 -1465
rect 26835 -1585 26880 -1465
rect 27000 -1585 27055 -1465
rect 27175 -1585 27220 -1465
rect 27340 -1585 27385 -1465
rect 27505 -1585 27550 -1465
rect 27670 -1585 27725 -1465
rect 27845 -1585 27890 -1465
rect 28010 -1585 28055 -1465
rect 28175 -1585 28220 -1465
rect 28340 -1585 28395 -1465
rect 28515 -1585 28560 -1465
rect 28680 -1585 28725 -1465
rect 28845 -1585 28890 -1465
rect 29010 -1585 29065 -1465
rect 29185 -1585 29230 -1465
rect 29350 -1585 29395 -1465
rect 29515 -1585 29560 -1465
rect 29680 -1585 29705 -1465
rect 24175 -1630 29705 -1585
rect 24175 -1750 24200 -1630
rect 24320 -1750 24375 -1630
rect 24495 -1750 24540 -1630
rect 24660 -1750 24705 -1630
rect 24825 -1750 24870 -1630
rect 24990 -1750 25045 -1630
rect 25165 -1750 25210 -1630
rect 25330 -1750 25375 -1630
rect 25495 -1750 25540 -1630
rect 25660 -1750 25715 -1630
rect 25835 -1750 25880 -1630
rect 26000 -1750 26045 -1630
rect 26165 -1750 26210 -1630
rect 26330 -1750 26385 -1630
rect 26505 -1750 26550 -1630
rect 26670 -1750 26715 -1630
rect 26835 -1750 26880 -1630
rect 27000 -1750 27055 -1630
rect 27175 -1750 27220 -1630
rect 27340 -1750 27385 -1630
rect 27505 -1750 27550 -1630
rect 27670 -1750 27725 -1630
rect 27845 -1750 27890 -1630
rect 28010 -1750 28055 -1630
rect 28175 -1750 28220 -1630
rect 28340 -1750 28395 -1630
rect 28515 -1750 28560 -1630
rect 28680 -1750 28725 -1630
rect 28845 -1750 28890 -1630
rect 29010 -1750 29065 -1630
rect 29185 -1750 29230 -1630
rect 29350 -1750 29395 -1630
rect 29515 -1750 29560 -1630
rect 29680 -1750 29705 -1630
rect 24175 -1795 29705 -1750
rect 24175 -1915 24200 -1795
rect 24320 -1915 24375 -1795
rect 24495 -1915 24540 -1795
rect 24660 -1915 24705 -1795
rect 24825 -1915 24870 -1795
rect 24990 -1915 25045 -1795
rect 25165 -1915 25210 -1795
rect 25330 -1915 25375 -1795
rect 25495 -1915 25540 -1795
rect 25660 -1915 25715 -1795
rect 25835 -1915 25880 -1795
rect 26000 -1915 26045 -1795
rect 26165 -1915 26210 -1795
rect 26330 -1915 26385 -1795
rect 26505 -1915 26550 -1795
rect 26670 -1915 26715 -1795
rect 26835 -1915 26880 -1795
rect 27000 -1915 27055 -1795
rect 27175 -1915 27220 -1795
rect 27340 -1915 27385 -1795
rect 27505 -1915 27550 -1795
rect 27670 -1915 27725 -1795
rect 27845 -1915 27890 -1795
rect 28010 -1915 28055 -1795
rect 28175 -1915 28220 -1795
rect 28340 -1915 28395 -1795
rect 28515 -1915 28560 -1795
rect 28680 -1915 28725 -1795
rect 28845 -1915 28890 -1795
rect 29010 -1915 29065 -1795
rect 29185 -1915 29230 -1795
rect 29350 -1915 29395 -1795
rect 29515 -1915 29560 -1795
rect 29680 -1915 29705 -1795
rect 24175 -1970 29705 -1915
rect 24175 -2090 24200 -1970
rect 24320 -2090 24375 -1970
rect 24495 -2090 24540 -1970
rect 24660 -2090 24705 -1970
rect 24825 -2090 24870 -1970
rect 24990 -2090 25045 -1970
rect 25165 -2090 25210 -1970
rect 25330 -2090 25375 -1970
rect 25495 -2090 25540 -1970
rect 25660 -2090 25715 -1970
rect 25835 -2090 25880 -1970
rect 26000 -2090 26045 -1970
rect 26165 -2090 26210 -1970
rect 26330 -2090 26385 -1970
rect 26505 -2090 26550 -1970
rect 26670 -2090 26715 -1970
rect 26835 -2090 26880 -1970
rect 27000 -2090 27055 -1970
rect 27175 -2090 27220 -1970
rect 27340 -2090 27385 -1970
rect 27505 -2090 27550 -1970
rect 27670 -2090 27725 -1970
rect 27845 -2090 27890 -1970
rect 28010 -2090 28055 -1970
rect 28175 -2090 28220 -1970
rect 28340 -2090 28395 -1970
rect 28515 -2090 28560 -1970
rect 28680 -2090 28725 -1970
rect 28845 -2090 28890 -1970
rect 29010 -2090 29065 -1970
rect 29185 -2090 29230 -1970
rect 29350 -2090 29395 -1970
rect 29515 -2090 29560 -1970
rect 29680 -2090 29705 -1970
rect 24175 -2135 29705 -2090
rect 24175 -2255 24200 -2135
rect 24320 -2255 24375 -2135
rect 24495 -2255 24540 -2135
rect 24660 -2255 24705 -2135
rect 24825 -2255 24870 -2135
rect 24990 -2255 25045 -2135
rect 25165 -2255 25210 -2135
rect 25330 -2255 25375 -2135
rect 25495 -2255 25540 -2135
rect 25660 -2255 25715 -2135
rect 25835 -2255 25880 -2135
rect 26000 -2255 26045 -2135
rect 26165 -2255 26210 -2135
rect 26330 -2255 26385 -2135
rect 26505 -2255 26550 -2135
rect 26670 -2255 26715 -2135
rect 26835 -2255 26880 -2135
rect 27000 -2255 27055 -2135
rect 27175 -2255 27220 -2135
rect 27340 -2255 27385 -2135
rect 27505 -2255 27550 -2135
rect 27670 -2255 27725 -2135
rect 27845 -2255 27890 -2135
rect 28010 -2255 28055 -2135
rect 28175 -2255 28220 -2135
rect 28340 -2255 28395 -2135
rect 28515 -2255 28560 -2135
rect 28680 -2255 28725 -2135
rect 28845 -2255 28890 -2135
rect 29010 -2255 29065 -2135
rect 29185 -2255 29230 -2135
rect 29350 -2255 29395 -2135
rect 29515 -2255 29560 -2135
rect 29680 -2255 29705 -2135
rect 24175 -2300 29705 -2255
rect 24175 -2420 24200 -2300
rect 24320 -2420 24375 -2300
rect 24495 -2420 24540 -2300
rect 24660 -2420 24705 -2300
rect 24825 -2420 24870 -2300
rect 24990 -2420 25045 -2300
rect 25165 -2420 25210 -2300
rect 25330 -2420 25375 -2300
rect 25495 -2420 25540 -2300
rect 25660 -2420 25715 -2300
rect 25835 -2420 25880 -2300
rect 26000 -2420 26045 -2300
rect 26165 -2420 26210 -2300
rect 26330 -2420 26385 -2300
rect 26505 -2420 26550 -2300
rect 26670 -2420 26715 -2300
rect 26835 -2420 26880 -2300
rect 27000 -2420 27055 -2300
rect 27175 -2420 27220 -2300
rect 27340 -2420 27385 -2300
rect 27505 -2420 27550 -2300
rect 27670 -2420 27725 -2300
rect 27845 -2420 27890 -2300
rect 28010 -2420 28055 -2300
rect 28175 -2420 28220 -2300
rect 28340 -2420 28395 -2300
rect 28515 -2420 28560 -2300
rect 28680 -2420 28725 -2300
rect 28845 -2420 28890 -2300
rect 29010 -2420 29065 -2300
rect 29185 -2420 29230 -2300
rect 29350 -2420 29395 -2300
rect 29515 -2420 29560 -2300
rect 29680 -2420 29705 -2300
rect 24175 -2465 29705 -2420
rect 24175 -2585 24200 -2465
rect 24320 -2585 24375 -2465
rect 24495 -2585 24540 -2465
rect 24660 -2585 24705 -2465
rect 24825 -2585 24870 -2465
rect 24990 -2585 25045 -2465
rect 25165 -2585 25210 -2465
rect 25330 -2585 25375 -2465
rect 25495 -2585 25540 -2465
rect 25660 -2585 25715 -2465
rect 25835 -2585 25880 -2465
rect 26000 -2585 26045 -2465
rect 26165 -2585 26210 -2465
rect 26330 -2585 26385 -2465
rect 26505 -2585 26550 -2465
rect 26670 -2585 26715 -2465
rect 26835 -2585 26880 -2465
rect 27000 -2585 27055 -2465
rect 27175 -2585 27220 -2465
rect 27340 -2585 27385 -2465
rect 27505 -2585 27550 -2465
rect 27670 -2585 27725 -2465
rect 27845 -2585 27890 -2465
rect 28010 -2585 28055 -2465
rect 28175 -2585 28220 -2465
rect 28340 -2585 28395 -2465
rect 28515 -2585 28560 -2465
rect 28680 -2585 28725 -2465
rect 28845 -2585 28890 -2465
rect 29010 -2585 29065 -2465
rect 29185 -2585 29230 -2465
rect 29350 -2585 29395 -2465
rect 29515 -2585 29560 -2465
rect 29680 -2585 29705 -2465
rect 24175 -2640 29705 -2585
rect 24175 -2760 24200 -2640
rect 24320 -2760 24375 -2640
rect 24495 -2760 24540 -2640
rect 24660 -2760 24705 -2640
rect 24825 -2760 24870 -2640
rect 24990 -2760 25045 -2640
rect 25165 -2760 25210 -2640
rect 25330 -2760 25375 -2640
rect 25495 -2760 25540 -2640
rect 25660 -2760 25715 -2640
rect 25835 -2760 25880 -2640
rect 26000 -2760 26045 -2640
rect 26165 -2760 26210 -2640
rect 26330 -2760 26385 -2640
rect 26505 -2760 26550 -2640
rect 26670 -2760 26715 -2640
rect 26835 -2760 26880 -2640
rect 27000 -2760 27055 -2640
rect 27175 -2760 27220 -2640
rect 27340 -2760 27385 -2640
rect 27505 -2760 27550 -2640
rect 27670 -2760 27725 -2640
rect 27845 -2760 27890 -2640
rect 28010 -2760 28055 -2640
rect 28175 -2760 28220 -2640
rect 28340 -2760 28395 -2640
rect 28515 -2760 28560 -2640
rect 28680 -2760 28725 -2640
rect 28845 -2760 28890 -2640
rect 29010 -2760 29065 -2640
rect 29185 -2760 29230 -2640
rect 29350 -2760 29395 -2640
rect 29515 -2760 29560 -2640
rect 29680 -2760 29705 -2640
rect 24175 -2805 29705 -2760
rect 24175 -2925 24200 -2805
rect 24320 -2925 24375 -2805
rect 24495 -2925 24540 -2805
rect 24660 -2925 24705 -2805
rect 24825 -2925 24870 -2805
rect 24990 -2925 25045 -2805
rect 25165 -2925 25210 -2805
rect 25330 -2925 25375 -2805
rect 25495 -2925 25540 -2805
rect 25660 -2925 25715 -2805
rect 25835 -2925 25880 -2805
rect 26000 -2925 26045 -2805
rect 26165 -2925 26210 -2805
rect 26330 -2925 26385 -2805
rect 26505 -2925 26550 -2805
rect 26670 -2925 26715 -2805
rect 26835 -2925 26880 -2805
rect 27000 -2925 27055 -2805
rect 27175 -2925 27220 -2805
rect 27340 -2925 27385 -2805
rect 27505 -2925 27550 -2805
rect 27670 -2925 27725 -2805
rect 27845 -2925 27890 -2805
rect 28010 -2925 28055 -2805
rect 28175 -2925 28220 -2805
rect 28340 -2925 28395 -2805
rect 28515 -2925 28560 -2805
rect 28680 -2925 28725 -2805
rect 28845 -2925 28890 -2805
rect 29010 -2925 29065 -2805
rect 29185 -2925 29230 -2805
rect 29350 -2925 29395 -2805
rect 29515 -2925 29560 -2805
rect 29680 -2925 29705 -2805
rect 24175 -2970 29705 -2925
rect 24175 -3090 24200 -2970
rect 24320 -3090 24375 -2970
rect 24495 -3090 24540 -2970
rect 24660 -3090 24705 -2970
rect 24825 -3090 24870 -2970
rect 24990 -3090 25045 -2970
rect 25165 -3090 25210 -2970
rect 25330 -3090 25375 -2970
rect 25495 -3090 25540 -2970
rect 25660 -3090 25715 -2970
rect 25835 -3090 25880 -2970
rect 26000 -3090 26045 -2970
rect 26165 -3090 26210 -2970
rect 26330 -3090 26385 -2970
rect 26505 -3090 26550 -2970
rect 26670 -3090 26715 -2970
rect 26835 -3090 26880 -2970
rect 27000 -3090 27055 -2970
rect 27175 -3090 27220 -2970
rect 27340 -3090 27385 -2970
rect 27505 -3090 27550 -2970
rect 27670 -3090 27725 -2970
rect 27845 -3090 27890 -2970
rect 28010 -3090 28055 -2970
rect 28175 -3090 28220 -2970
rect 28340 -3090 28395 -2970
rect 28515 -3090 28560 -2970
rect 28680 -3090 28725 -2970
rect 28845 -3090 28890 -2970
rect 29010 -3090 29065 -2970
rect 29185 -3090 29230 -2970
rect 29350 -3090 29395 -2970
rect 29515 -3090 29560 -2970
rect 29680 -3090 29705 -2970
rect 24175 -3135 29705 -3090
rect 24175 -3255 24200 -3135
rect 24320 -3255 24375 -3135
rect 24495 -3255 24540 -3135
rect 24660 -3255 24705 -3135
rect 24825 -3255 24870 -3135
rect 24990 -3255 25045 -3135
rect 25165 -3255 25210 -3135
rect 25330 -3255 25375 -3135
rect 25495 -3255 25540 -3135
rect 25660 -3255 25715 -3135
rect 25835 -3255 25880 -3135
rect 26000 -3255 26045 -3135
rect 26165 -3255 26210 -3135
rect 26330 -3255 26385 -3135
rect 26505 -3255 26550 -3135
rect 26670 -3255 26715 -3135
rect 26835 -3255 26880 -3135
rect 27000 -3255 27055 -3135
rect 27175 -3255 27220 -3135
rect 27340 -3255 27385 -3135
rect 27505 -3255 27550 -3135
rect 27670 -3255 27725 -3135
rect 27845 -3255 27890 -3135
rect 28010 -3255 28055 -3135
rect 28175 -3255 28220 -3135
rect 28340 -3255 28395 -3135
rect 28515 -3255 28560 -3135
rect 28680 -3255 28725 -3135
rect 28845 -3255 28890 -3135
rect 29010 -3255 29065 -3135
rect 29185 -3255 29230 -3135
rect 29350 -3255 29395 -3135
rect 29515 -3255 29560 -3135
rect 29680 -3255 29705 -3135
rect 24175 -3310 29705 -3255
rect 24175 -3430 24200 -3310
rect 24320 -3430 24375 -3310
rect 24495 -3430 24540 -3310
rect 24660 -3430 24705 -3310
rect 24825 -3430 24870 -3310
rect 24990 -3430 25045 -3310
rect 25165 -3430 25210 -3310
rect 25330 -3430 25375 -3310
rect 25495 -3430 25540 -3310
rect 25660 -3430 25715 -3310
rect 25835 -3430 25880 -3310
rect 26000 -3430 26045 -3310
rect 26165 -3430 26210 -3310
rect 26330 -3430 26385 -3310
rect 26505 -3430 26550 -3310
rect 26670 -3430 26715 -3310
rect 26835 -3430 26880 -3310
rect 27000 -3430 27055 -3310
rect 27175 -3430 27220 -3310
rect 27340 -3430 27385 -3310
rect 27505 -3430 27550 -3310
rect 27670 -3430 27725 -3310
rect 27845 -3430 27890 -3310
rect 28010 -3430 28055 -3310
rect 28175 -3430 28220 -3310
rect 28340 -3430 28395 -3310
rect 28515 -3430 28560 -3310
rect 28680 -3430 28725 -3310
rect 28845 -3430 28890 -3310
rect 29010 -3430 29065 -3310
rect 29185 -3430 29230 -3310
rect 29350 -3430 29395 -3310
rect 29515 -3430 29560 -3310
rect 29680 -3430 29705 -3310
rect 24175 -3475 29705 -3430
rect 24175 -3595 24200 -3475
rect 24320 -3595 24375 -3475
rect 24495 -3595 24540 -3475
rect 24660 -3595 24705 -3475
rect 24825 -3595 24870 -3475
rect 24990 -3595 25045 -3475
rect 25165 -3595 25210 -3475
rect 25330 -3595 25375 -3475
rect 25495 -3595 25540 -3475
rect 25660 -3595 25715 -3475
rect 25835 -3595 25880 -3475
rect 26000 -3595 26045 -3475
rect 26165 -3595 26210 -3475
rect 26330 -3595 26385 -3475
rect 26505 -3595 26550 -3475
rect 26670 -3595 26715 -3475
rect 26835 -3595 26880 -3475
rect 27000 -3595 27055 -3475
rect 27175 -3595 27220 -3475
rect 27340 -3595 27385 -3475
rect 27505 -3595 27550 -3475
rect 27670 -3595 27725 -3475
rect 27845 -3595 27890 -3475
rect 28010 -3595 28055 -3475
rect 28175 -3595 28220 -3475
rect 28340 -3595 28395 -3475
rect 28515 -3595 28560 -3475
rect 28680 -3595 28725 -3475
rect 28845 -3595 28890 -3475
rect 29010 -3595 29065 -3475
rect 29185 -3595 29230 -3475
rect 29350 -3595 29395 -3475
rect 29515 -3595 29560 -3475
rect 29680 -3595 29705 -3475
rect 24175 -3640 29705 -3595
rect 24175 -3760 24200 -3640
rect 24320 -3760 24375 -3640
rect 24495 -3760 24540 -3640
rect 24660 -3760 24705 -3640
rect 24825 -3760 24870 -3640
rect 24990 -3760 25045 -3640
rect 25165 -3760 25210 -3640
rect 25330 -3760 25375 -3640
rect 25495 -3760 25540 -3640
rect 25660 -3760 25715 -3640
rect 25835 -3760 25880 -3640
rect 26000 -3760 26045 -3640
rect 26165 -3760 26210 -3640
rect 26330 -3760 26385 -3640
rect 26505 -3760 26550 -3640
rect 26670 -3760 26715 -3640
rect 26835 -3760 26880 -3640
rect 27000 -3760 27055 -3640
rect 27175 -3760 27220 -3640
rect 27340 -3760 27385 -3640
rect 27505 -3760 27550 -3640
rect 27670 -3760 27725 -3640
rect 27845 -3760 27890 -3640
rect 28010 -3760 28055 -3640
rect 28175 -3760 28220 -3640
rect 28340 -3760 28395 -3640
rect 28515 -3760 28560 -3640
rect 28680 -3760 28725 -3640
rect 28845 -3760 28890 -3640
rect 29010 -3760 29065 -3640
rect 29185 -3760 29230 -3640
rect 29350 -3760 29395 -3640
rect 29515 -3760 29560 -3640
rect 29680 -3760 29705 -3640
rect 24175 -3805 29705 -3760
rect 24175 -3925 24200 -3805
rect 24320 -3925 24375 -3805
rect 24495 -3925 24540 -3805
rect 24660 -3925 24705 -3805
rect 24825 -3925 24870 -3805
rect 24990 -3925 25045 -3805
rect 25165 -3925 25210 -3805
rect 25330 -3925 25375 -3805
rect 25495 -3925 25540 -3805
rect 25660 -3925 25715 -3805
rect 25835 -3925 25880 -3805
rect 26000 -3925 26045 -3805
rect 26165 -3925 26210 -3805
rect 26330 -3925 26385 -3805
rect 26505 -3925 26550 -3805
rect 26670 -3925 26715 -3805
rect 26835 -3925 26880 -3805
rect 27000 -3925 27055 -3805
rect 27175 -3925 27220 -3805
rect 27340 -3925 27385 -3805
rect 27505 -3925 27550 -3805
rect 27670 -3925 27725 -3805
rect 27845 -3925 27890 -3805
rect 28010 -3925 28055 -3805
rect 28175 -3925 28220 -3805
rect 28340 -3925 28395 -3805
rect 28515 -3925 28560 -3805
rect 28680 -3925 28725 -3805
rect 28845 -3925 28890 -3805
rect 29010 -3925 29065 -3805
rect 29185 -3925 29230 -3805
rect 29350 -3925 29395 -3805
rect 29515 -3925 29560 -3805
rect 29680 -3925 29705 -3805
rect 24175 -3980 29705 -3925
rect 24175 -4100 24200 -3980
rect 24320 -4100 24375 -3980
rect 24495 -4100 24540 -3980
rect 24660 -4100 24705 -3980
rect 24825 -4100 24870 -3980
rect 24990 -4100 25045 -3980
rect 25165 -4100 25210 -3980
rect 25330 -4100 25375 -3980
rect 25495 -4100 25540 -3980
rect 25660 -4100 25715 -3980
rect 25835 -4100 25880 -3980
rect 26000 -4100 26045 -3980
rect 26165 -4100 26210 -3980
rect 26330 -4100 26385 -3980
rect 26505 -4100 26550 -3980
rect 26670 -4100 26715 -3980
rect 26835 -4100 26880 -3980
rect 27000 -4100 27055 -3980
rect 27175 -4100 27220 -3980
rect 27340 -4100 27385 -3980
rect 27505 -4100 27550 -3980
rect 27670 -4100 27725 -3980
rect 27845 -4100 27890 -3980
rect 28010 -4100 28055 -3980
rect 28175 -4100 28220 -3980
rect 28340 -4100 28395 -3980
rect 28515 -4100 28560 -3980
rect 28680 -4100 28725 -3980
rect 28845 -4100 28890 -3980
rect 29010 -4100 29065 -3980
rect 29185 -4100 29230 -3980
rect 29350 -4100 29395 -3980
rect 29515 -4100 29560 -3980
rect 29680 -4100 29705 -3980
rect 24175 -4125 29705 -4100
rect 7105 -4310 12635 -4285
rect 7105 -4430 7130 -4310
rect 7250 -4430 7295 -4310
rect 7415 -4430 7460 -4310
rect 7580 -4430 7625 -4310
rect 7745 -4430 7800 -4310
rect 7920 -4430 7965 -4310
rect 8085 -4430 8130 -4310
rect 8250 -4430 8295 -4310
rect 8415 -4430 8470 -4310
rect 8590 -4430 8635 -4310
rect 8755 -4430 8800 -4310
rect 8920 -4430 8965 -4310
rect 9085 -4430 9140 -4310
rect 9260 -4430 9305 -4310
rect 9425 -4430 9470 -4310
rect 9590 -4430 9635 -4310
rect 9755 -4430 9810 -4310
rect 9930 -4430 9975 -4310
rect 10095 -4430 10140 -4310
rect 10260 -4430 10305 -4310
rect 10425 -4430 10480 -4310
rect 10600 -4430 10645 -4310
rect 10765 -4430 10810 -4310
rect 10930 -4430 10975 -4310
rect 11095 -4430 11150 -4310
rect 11270 -4430 11315 -4310
rect 11435 -4430 11480 -4310
rect 11600 -4430 11645 -4310
rect 11765 -4430 11820 -4310
rect 11940 -4430 11985 -4310
rect 12105 -4430 12150 -4310
rect 12270 -4430 12315 -4310
rect 12435 -4430 12490 -4310
rect 12610 -4430 12635 -4310
rect 7105 -4485 12635 -4430
rect 7105 -4605 7130 -4485
rect 7250 -4605 7295 -4485
rect 7415 -4605 7460 -4485
rect 7580 -4605 7625 -4485
rect 7745 -4605 7800 -4485
rect 7920 -4605 7965 -4485
rect 8085 -4605 8130 -4485
rect 8250 -4605 8295 -4485
rect 8415 -4605 8470 -4485
rect 8590 -4605 8635 -4485
rect 8755 -4605 8800 -4485
rect 8920 -4605 8965 -4485
rect 9085 -4605 9140 -4485
rect 9260 -4605 9305 -4485
rect 9425 -4605 9470 -4485
rect 9590 -4605 9635 -4485
rect 9755 -4605 9810 -4485
rect 9930 -4605 9975 -4485
rect 10095 -4605 10140 -4485
rect 10260 -4605 10305 -4485
rect 10425 -4605 10480 -4485
rect 10600 -4605 10645 -4485
rect 10765 -4605 10810 -4485
rect 10930 -4605 10975 -4485
rect 11095 -4605 11150 -4485
rect 11270 -4605 11315 -4485
rect 11435 -4605 11480 -4485
rect 11600 -4605 11645 -4485
rect 11765 -4605 11820 -4485
rect 11940 -4605 11985 -4485
rect 12105 -4605 12150 -4485
rect 12270 -4605 12315 -4485
rect 12435 -4605 12490 -4485
rect 12610 -4605 12635 -4485
rect 7105 -4650 12635 -4605
rect 7105 -4770 7130 -4650
rect 7250 -4770 7295 -4650
rect 7415 -4770 7460 -4650
rect 7580 -4770 7625 -4650
rect 7745 -4770 7800 -4650
rect 7920 -4770 7965 -4650
rect 8085 -4770 8130 -4650
rect 8250 -4770 8295 -4650
rect 8415 -4770 8470 -4650
rect 8590 -4770 8635 -4650
rect 8755 -4770 8800 -4650
rect 8920 -4770 8965 -4650
rect 9085 -4770 9140 -4650
rect 9260 -4770 9305 -4650
rect 9425 -4770 9470 -4650
rect 9590 -4770 9635 -4650
rect 9755 -4770 9810 -4650
rect 9930 -4770 9975 -4650
rect 10095 -4770 10140 -4650
rect 10260 -4770 10305 -4650
rect 10425 -4770 10480 -4650
rect 10600 -4770 10645 -4650
rect 10765 -4770 10810 -4650
rect 10930 -4770 10975 -4650
rect 11095 -4770 11150 -4650
rect 11270 -4770 11315 -4650
rect 11435 -4770 11480 -4650
rect 11600 -4770 11645 -4650
rect 11765 -4770 11820 -4650
rect 11940 -4770 11985 -4650
rect 12105 -4770 12150 -4650
rect 12270 -4770 12315 -4650
rect 12435 -4770 12490 -4650
rect 12610 -4770 12635 -4650
rect 7105 -4815 12635 -4770
rect 7105 -4935 7130 -4815
rect 7250 -4935 7295 -4815
rect 7415 -4935 7460 -4815
rect 7580 -4935 7625 -4815
rect 7745 -4935 7800 -4815
rect 7920 -4935 7965 -4815
rect 8085 -4935 8130 -4815
rect 8250 -4935 8295 -4815
rect 8415 -4935 8470 -4815
rect 8590 -4935 8635 -4815
rect 8755 -4935 8800 -4815
rect 8920 -4935 8965 -4815
rect 9085 -4935 9140 -4815
rect 9260 -4935 9305 -4815
rect 9425 -4935 9470 -4815
rect 9590 -4935 9635 -4815
rect 9755 -4935 9810 -4815
rect 9930 -4935 9975 -4815
rect 10095 -4935 10140 -4815
rect 10260 -4935 10305 -4815
rect 10425 -4935 10480 -4815
rect 10600 -4935 10645 -4815
rect 10765 -4935 10810 -4815
rect 10930 -4935 10975 -4815
rect 11095 -4935 11150 -4815
rect 11270 -4935 11315 -4815
rect 11435 -4935 11480 -4815
rect 11600 -4935 11645 -4815
rect 11765 -4935 11820 -4815
rect 11940 -4935 11985 -4815
rect 12105 -4935 12150 -4815
rect 12270 -4935 12315 -4815
rect 12435 -4935 12490 -4815
rect 12610 -4935 12635 -4815
rect 7105 -4980 12635 -4935
rect 7105 -5100 7130 -4980
rect 7250 -5100 7295 -4980
rect 7415 -5100 7460 -4980
rect 7580 -5100 7625 -4980
rect 7745 -5100 7800 -4980
rect 7920 -5100 7965 -4980
rect 8085 -5100 8130 -4980
rect 8250 -5100 8295 -4980
rect 8415 -5100 8470 -4980
rect 8590 -5100 8635 -4980
rect 8755 -5100 8800 -4980
rect 8920 -5100 8965 -4980
rect 9085 -5100 9140 -4980
rect 9260 -5100 9305 -4980
rect 9425 -5100 9470 -4980
rect 9590 -5100 9635 -4980
rect 9755 -5100 9810 -4980
rect 9930 -5100 9975 -4980
rect 10095 -5100 10140 -4980
rect 10260 -5100 10305 -4980
rect 10425 -5100 10480 -4980
rect 10600 -5100 10645 -4980
rect 10765 -5100 10810 -4980
rect 10930 -5100 10975 -4980
rect 11095 -5100 11150 -4980
rect 11270 -5100 11315 -4980
rect 11435 -5100 11480 -4980
rect 11600 -5100 11645 -4980
rect 11765 -5100 11820 -4980
rect 11940 -5100 11985 -4980
rect 12105 -5100 12150 -4980
rect 12270 -5100 12315 -4980
rect 12435 -5100 12490 -4980
rect 12610 -5100 12635 -4980
rect 7105 -5155 12635 -5100
rect 7105 -5275 7130 -5155
rect 7250 -5275 7295 -5155
rect 7415 -5275 7460 -5155
rect 7580 -5275 7625 -5155
rect 7745 -5275 7800 -5155
rect 7920 -5275 7965 -5155
rect 8085 -5275 8130 -5155
rect 8250 -5275 8295 -5155
rect 8415 -5275 8470 -5155
rect 8590 -5275 8635 -5155
rect 8755 -5275 8800 -5155
rect 8920 -5275 8965 -5155
rect 9085 -5275 9140 -5155
rect 9260 -5275 9305 -5155
rect 9425 -5275 9470 -5155
rect 9590 -5275 9635 -5155
rect 9755 -5275 9810 -5155
rect 9930 -5275 9975 -5155
rect 10095 -5275 10140 -5155
rect 10260 -5275 10305 -5155
rect 10425 -5275 10480 -5155
rect 10600 -5275 10645 -5155
rect 10765 -5275 10810 -5155
rect 10930 -5275 10975 -5155
rect 11095 -5275 11150 -5155
rect 11270 -5275 11315 -5155
rect 11435 -5275 11480 -5155
rect 11600 -5275 11645 -5155
rect 11765 -5275 11820 -5155
rect 11940 -5275 11985 -5155
rect 12105 -5275 12150 -5155
rect 12270 -5275 12315 -5155
rect 12435 -5275 12490 -5155
rect 12610 -5275 12635 -5155
rect 7105 -5320 12635 -5275
rect 7105 -5440 7130 -5320
rect 7250 -5440 7295 -5320
rect 7415 -5440 7460 -5320
rect 7580 -5440 7625 -5320
rect 7745 -5440 7800 -5320
rect 7920 -5440 7965 -5320
rect 8085 -5440 8130 -5320
rect 8250 -5440 8295 -5320
rect 8415 -5440 8470 -5320
rect 8590 -5440 8635 -5320
rect 8755 -5440 8800 -5320
rect 8920 -5440 8965 -5320
rect 9085 -5440 9140 -5320
rect 9260 -5440 9305 -5320
rect 9425 -5440 9470 -5320
rect 9590 -5440 9635 -5320
rect 9755 -5440 9810 -5320
rect 9930 -5440 9975 -5320
rect 10095 -5440 10140 -5320
rect 10260 -5440 10305 -5320
rect 10425 -5440 10480 -5320
rect 10600 -5440 10645 -5320
rect 10765 -5440 10810 -5320
rect 10930 -5440 10975 -5320
rect 11095 -5440 11150 -5320
rect 11270 -5440 11315 -5320
rect 11435 -5440 11480 -5320
rect 11600 -5440 11645 -5320
rect 11765 -5440 11820 -5320
rect 11940 -5440 11985 -5320
rect 12105 -5440 12150 -5320
rect 12270 -5440 12315 -5320
rect 12435 -5440 12490 -5320
rect 12610 -5440 12635 -5320
rect 7105 -5485 12635 -5440
rect 7105 -5605 7130 -5485
rect 7250 -5605 7295 -5485
rect 7415 -5605 7460 -5485
rect 7580 -5605 7625 -5485
rect 7745 -5605 7800 -5485
rect 7920 -5605 7965 -5485
rect 8085 -5605 8130 -5485
rect 8250 -5605 8295 -5485
rect 8415 -5605 8470 -5485
rect 8590 -5605 8635 -5485
rect 8755 -5605 8800 -5485
rect 8920 -5605 8965 -5485
rect 9085 -5605 9140 -5485
rect 9260 -5605 9305 -5485
rect 9425 -5605 9470 -5485
rect 9590 -5605 9635 -5485
rect 9755 -5605 9810 -5485
rect 9930 -5605 9975 -5485
rect 10095 -5605 10140 -5485
rect 10260 -5605 10305 -5485
rect 10425 -5605 10480 -5485
rect 10600 -5605 10645 -5485
rect 10765 -5605 10810 -5485
rect 10930 -5605 10975 -5485
rect 11095 -5605 11150 -5485
rect 11270 -5605 11315 -5485
rect 11435 -5605 11480 -5485
rect 11600 -5605 11645 -5485
rect 11765 -5605 11820 -5485
rect 11940 -5605 11985 -5485
rect 12105 -5605 12150 -5485
rect 12270 -5605 12315 -5485
rect 12435 -5605 12490 -5485
rect 12610 -5605 12635 -5485
rect 7105 -5650 12635 -5605
rect 7105 -5770 7130 -5650
rect 7250 -5770 7295 -5650
rect 7415 -5770 7460 -5650
rect 7580 -5770 7625 -5650
rect 7745 -5770 7800 -5650
rect 7920 -5770 7965 -5650
rect 8085 -5770 8130 -5650
rect 8250 -5770 8295 -5650
rect 8415 -5770 8470 -5650
rect 8590 -5770 8635 -5650
rect 8755 -5770 8800 -5650
rect 8920 -5770 8965 -5650
rect 9085 -5770 9140 -5650
rect 9260 -5770 9305 -5650
rect 9425 -5770 9470 -5650
rect 9590 -5770 9635 -5650
rect 9755 -5770 9810 -5650
rect 9930 -5770 9975 -5650
rect 10095 -5770 10140 -5650
rect 10260 -5770 10305 -5650
rect 10425 -5770 10480 -5650
rect 10600 -5770 10645 -5650
rect 10765 -5770 10810 -5650
rect 10930 -5770 10975 -5650
rect 11095 -5770 11150 -5650
rect 11270 -5770 11315 -5650
rect 11435 -5770 11480 -5650
rect 11600 -5770 11645 -5650
rect 11765 -5770 11820 -5650
rect 11940 -5770 11985 -5650
rect 12105 -5770 12150 -5650
rect 12270 -5770 12315 -5650
rect 12435 -5770 12490 -5650
rect 12610 -5770 12635 -5650
rect 7105 -5825 12635 -5770
rect 7105 -5945 7130 -5825
rect 7250 -5945 7295 -5825
rect 7415 -5945 7460 -5825
rect 7580 -5945 7625 -5825
rect 7745 -5945 7800 -5825
rect 7920 -5945 7965 -5825
rect 8085 -5945 8130 -5825
rect 8250 -5945 8295 -5825
rect 8415 -5945 8470 -5825
rect 8590 -5945 8635 -5825
rect 8755 -5945 8800 -5825
rect 8920 -5945 8965 -5825
rect 9085 -5945 9140 -5825
rect 9260 -5945 9305 -5825
rect 9425 -5945 9470 -5825
rect 9590 -5945 9635 -5825
rect 9755 -5945 9810 -5825
rect 9930 -5945 9975 -5825
rect 10095 -5945 10140 -5825
rect 10260 -5945 10305 -5825
rect 10425 -5945 10480 -5825
rect 10600 -5945 10645 -5825
rect 10765 -5945 10810 -5825
rect 10930 -5945 10975 -5825
rect 11095 -5945 11150 -5825
rect 11270 -5945 11315 -5825
rect 11435 -5945 11480 -5825
rect 11600 -5945 11645 -5825
rect 11765 -5945 11820 -5825
rect 11940 -5945 11985 -5825
rect 12105 -5945 12150 -5825
rect 12270 -5945 12315 -5825
rect 12435 -5945 12490 -5825
rect 12610 -5945 12635 -5825
rect 7105 -5990 12635 -5945
rect 7105 -6110 7130 -5990
rect 7250 -6110 7295 -5990
rect 7415 -6110 7460 -5990
rect 7580 -6110 7625 -5990
rect 7745 -6110 7800 -5990
rect 7920 -6110 7965 -5990
rect 8085 -6110 8130 -5990
rect 8250 -6110 8295 -5990
rect 8415 -6110 8470 -5990
rect 8590 -6110 8635 -5990
rect 8755 -6110 8800 -5990
rect 8920 -6110 8965 -5990
rect 9085 -6110 9140 -5990
rect 9260 -6110 9305 -5990
rect 9425 -6110 9470 -5990
rect 9590 -6110 9635 -5990
rect 9755 -6110 9810 -5990
rect 9930 -6110 9975 -5990
rect 10095 -6110 10140 -5990
rect 10260 -6110 10305 -5990
rect 10425 -6110 10480 -5990
rect 10600 -6110 10645 -5990
rect 10765 -6110 10810 -5990
rect 10930 -6110 10975 -5990
rect 11095 -6110 11150 -5990
rect 11270 -6110 11315 -5990
rect 11435 -6110 11480 -5990
rect 11600 -6110 11645 -5990
rect 11765 -6110 11820 -5990
rect 11940 -6110 11985 -5990
rect 12105 -6110 12150 -5990
rect 12270 -6110 12315 -5990
rect 12435 -6110 12490 -5990
rect 12610 -6110 12635 -5990
rect 7105 -6155 12635 -6110
rect 7105 -6275 7130 -6155
rect 7250 -6275 7295 -6155
rect 7415 -6275 7460 -6155
rect 7580 -6275 7625 -6155
rect 7745 -6275 7800 -6155
rect 7920 -6275 7965 -6155
rect 8085 -6275 8130 -6155
rect 8250 -6275 8295 -6155
rect 8415 -6275 8470 -6155
rect 8590 -6275 8635 -6155
rect 8755 -6275 8800 -6155
rect 8920 -6275 8965 -6155
rect 9085 -6275 9140 -6155
rect 9260 -6275 9305 -6155
rect 9425 -6275 9470 -6155
rect 9590 -6275 9635 -6155
rect 9755 -6275 9810 -6155
rect 9930 -6275 9975 -6155
rect 10095 -6275 10140 -6155
rect 10260 -6275 10305 -6155
rect 10425 -6275 10480 -6155
rect 10600 -6275 10645 -6155
rect 10765 -6275 10810 -6155
rect 10930 -6275 10975 -6155
rect 11095 -6275 11150 -6155
rect 11270 -6275 11315 -6155
rect 11435 -6275 11480 -6155
rect 11600 -6275 11645 -6155
rect 11765 -6275 11820 -6155
rect 11940 -6275 11985 -6155
rect 12105 -6275 12150 -6155
rect 12270 -6275 12315 -6155
rect 12435 -6275 12490 -6155
rect 12610 -6275 12635 -6155
rect 7105 -6320 12635 -6275
rect 7105 -6440 7130 -6320
rect 7250 -6440 7295 -6320
rect 7415 -6440 7460 -6320
rect 7580 -6440 7625 -6320
rect 7745 -6440 7800 -6320
rect 7920 -6440 7965 -6320
rect 8085 -6440 8130 -6320
rect 8250 -6440 8295 -6320
rect 8415 -6440 8470 -6320
rect 8590 -6440 8635 -6320
rect 8755 -6440 8800 -6320
rect 8920 -6440 8965 -6320
rect 9085 -6440 9140 -6320
rect 9260 -6440 9305 -6320
rect 9425 -6440 9470 -6320
rect 9590 -6440 9635 -6320
rect 9755 -6440 9810 -6320
rect 9930 -6440 9975 -6320
rect 10095 -6440 10140 -6320
rect 10260 -6440 10305 -6320
rect 10425 -6440 10480 -6320
rect 10600 -6440 10645 -6320
rect 10765 -6440 10810 -6320
rect 10930 -6440 10975 -6320
rect 11095 -6440 11150 -6320
rect 11270 -6440 11315 -6320
rect 11435 -6440 11480 -6320
rect 11600 -6440 11645 -6320
rect 11765 -6440 11820 -6320
rect 11940 -6440 11985 -6320
rect 12105 -6440 12150 -6320
rect 12270 -6440 12315 -6320
rect 12435 -6440 12490 -6320
rect 12610 -6440 12635 -6320
rect 7105 -6495 12635 -6440
rect 7105 -6615 7130 -6495
rect 7250 -6615 7295 -6495
rect 7415 -6615 7460 -6495
rect 7580 -6615 7625 -6495
rect 7745 -6615 7800 -6495
rect 7920 -6615 7965 -6495
rect 8085 -6615 8130 -6495
rect 8250 -6615 8295 -6495
rect 8415 -6615 8470 -6495
rect 8590 -6615 8635 -6495
rect 8755 -6615 8800 -6495
rect 8920 -6615 8965 -6495
rect 9085 -6615 9140 -6495
rect 9260 -6615 9305 -6495
rect 9425 -6615 9470 -6495
rect 9590 -6615 9635 -6495
rect 9755 -6615 9810 -6495
rect 9930 -6615 9975 -6495
rect 10095 -6615 10140 -6495
rect 10260 -6615 10305 -6495
rect 10425 -6615 10480 -6495
rect 10600 -6615 10645 -6495
rect 10765 -6615 10810 -6495
rect 10930 -6615 10975 -6495
rect 11095 -6615 11150 -6495
rect 11270 -6615 11315 -6495
rect 11435 -6615 11480 -6495
rect 11600 -6615 11645 -6495
rect 11765 -6615 11820 -6495
rect 11940 -6615 11985 -6495
rect 12105 -6615 12150 -6495
rect 12270 -6615 12315 -6495
rect 12435 -6615 12490 -6495
rect 12610 -6615 12635 -6495
rect 7105 -6660 12635 -6615
rect 7105 -6780 7130 -6660
rect 7250 -6780 7295 -6660
rect 7415 -6780 7460 -6660
rect 7580 -6780 7625 -6660
rect 7745 -6780 7800 -6660
rect 7920 -6780 7965 -6660
rect 8085 -6780 8130 -6660
rect 8250 -6780 8295 -6660
rect 8415 -6780 8470 -6660
rect 8590 -6780 8635 -6660
rect 8755 -6780 8800 -6660
rect 8920 -6780 8965 -6660
rect 9085 -6780 9140 -6660
rect 9260 -6780 9305 -6660
rect 9425 -6780 9470 -6660
rect 9590 -6780 9635 -6660
rect 9755 -6780 9810 -6660
rect 9930 -6780 9975 -6660
rect 10095 -6780 10140 -6660
rect 10260 -6780 10305 -6660
rect 10425 -6780 10480 -6660
rect 10600 -6780 10645 -6660
rect 10765 -6780 10810 -6660
rect 10930 -6780 10975 -6660
rect 11095 -6780 11150 -6660
rect 11270 -6780 11315 -6660
rect 11435 -6780 11480 -6660
rect 11600 -6780 11645 -6660
rect 11765 -6780 11820 -6660
rect 11940 -6780 11985 -6660
rect 12105 -6780 12150 -6660
rect 12270 -6780 12315 -6660
rect 12435 -6780 12490 -6660
rect 12610 -6780 12635 -6660
rect 7105 -6825 12635 -6780
rect 7105 -6945 7130 -6825
rect 7250 -6945 7295 -6825
rect 7415 -6945 7460 -6825
rect 7580 -6945 7625 -6825
rect 7745 -6945 7800 -6825
rect 7920 -6945 7965 -6825
rect 8085 -6945 8130 -6825
rect 8250 -6945 8295 -6825
rect 8415 -6945 8470 -6825
rect 8590 -6945 8635 -6825
rect 8755 -6945 8800 -6825
rect 8920 -6945 8965 -6825
rect 9085 -6945 9140 -6825
rect 9260 -6945 9305 -6825
rect 9425 -6945 9470 -6825
rect 9590 -6945 9635 -6825
rect 9755 -6945 9810 -6825
rect 9930 -6945 9975 -6825
rect 10095 -6945 10140 -6825
rect 10260 -6945 10305 -6825
rect 10425 -6945 10480 -6825
rect 10600 -6945 10645 -6825
rect 10765 -6945 10810 -6825
rect 10930 -6945 10975 -6825
rect 11095 -6945 11150 -6825
rect 11270 -6945 11315 -6825
rect 11435 -6945 11480 -6825
rect 11600 -6945 11645 -6825
rect 11765 -6945 11820 -6825
rect 11940 -6945 11985 -6825
rect 12105 -6945 12150 -6825
rect 12270 -6945 12315 -6825
rect 12435 -6945 12490 -6825
rect 12610 -6945 12635 -6825
rect 7105 -6990 12635 -6945
rect 7105 -7110 7130 -6990
rect 7250 -7110 7295 -6990
rect 7415 -7110 7460 -6990
rect 7580 -7110 7625 -6990
rect 7745 -7110 7800 -6990
rect 7920 -7110 7965 -6990
rect 8085 -7110 8130 -6990
rect 8250 -7110 8295 -6990
rect 8415 -7110 8470 -6990
rect 8590 -7110 8635 -6990
rect 8755 -7110 8800 -6990
rect 8920 -7110 8965 -6990
rect 9085 -7110 9140 -6990
rect 9260 -7110 9305 -6990
rect 9425 -7110 9470 -6990
rect 9590 -7110 9635 -6990
rect 9755 -7110 9810 -6990
rect 9930 -7110 9975 -6990
rect 10095 -7110 10140 -6990
rect 10260 -7110 10305 -6990
rect 10425 -7110 10480 -6990
rect 10600 -7110 10645 -6990
rect 10765 -7110 10810 -6990
rect 10930 -7110 10975 -6990
rect 11095 -7110 11150 -6990
rect 11270 -7110 11315 -6990
rect 11435 -7110 11480 -6990
rect 11600 -7110 11645 -6990
rect 11765 -7110 11820 -6990
rect 11940 -7110 11985 -6990
rect 12105 -7110 12150 -6990
rect 12270 -7110 12315 -6990
rect 12435 -7110 12490 -6990
rect 12610 -7110 12635 -6990
rect 7105 -7165 12635 -7110
rect 7105 -7285 7130 -7165
rect 7250 -7285 7295 -7165
rect 7415 -7285 7460 -7165
rect 7580 -7285 7625 -7165
rect 7745 -7285 7800 -7165
rect 7920 -7285 7965 -7165
rect 8085 -7285 8130 -7165
rect 8250 -7285 8295 -7165
rect 8415 -7285 8470 -7165
rect 8590 -7285 8635 -7165
rect 8755 -7285 8800 -7165
rect 8920 -7285 8965 -7165
rect 9085 -7285 9140 -7165
rect 9260 -7285 9305 -7165
rect 9425 -7285 9470 -7165
rect 9590 -7285 9635 -7165
rect 9755 -7285 9810 -7165
rect 9930 -7285 9975 -7165
rect 10095 -7285 10140 -7165
rect 10260 -7285 10305 -7165
rect 10425 -7285 10480 -7165
rect 10600 -7285 10645 -7165
rect 10765 -7285 10810 -7165
rect 10930 -7285 10975 -7165
rect 11095 -7285 11150 -7165
rect 11270 -7285 11315 -7165
rect 11435 -7285 11480 -7165
rect 11600 -7285 11645 -7165
rect 11765 -7285 11820 -7165
rect 11940 -7285 11985 -7165
rect 12105 -7285 12150 -7165
rect 12270 -7285 12315 -7165
rect 12435 -7285 12490 -7165
rect 12610 -7285 12635 -7165
rect 7105 -7330 12635 -7285
rect 7105 -7450 7130 -7330
rect 7250 -7450 7295 -7330
rect 7415 -7450 7460 -7330
rect 7580 -7450 7625 -7330
rect 7745 -7450 7800 -7330
rect 7920 -7450 7965 -7330
rect 8085 -7450 8130 -7330
rect 8250 -7450 8295 -7330
rect 8415 -7450 8470 -7330
rect 8590 -7450 8635 -7330
rect 8755 -7450 8800 -7330
rect 8920 -7450 8965 -7330
rect 9085 -7450 9140 -7330
rect 9260 -7450 9305 -7330
rect 9425 -7450 9470 -7330
rect 9590 -7450 9635 -7330
rect 9755 -7450 9810 -7330
rect 9930 -7450 9975 -7330
rect 10095 -7450 10140 -7330
rect 10260 -7450 10305 -7330
rect 10425 -7450 10480 -7330
rect 10600 -7450 10645 -7330
rect 10765 -7450 10810 -7330
rect 10930 -7450 10975 -7330
rect 11095 -7450 11150 -7330
rect 11270 -7450 11315 -7330
rect 11435 -7450 11480 -7330
rect 11600 -7450 11645 -7330
rect 11765 -7450 11820 -7330
rect 11940 -7450 11985 -7330
rect 12105 -7450 12150 -7330
rect 12270 -7450 12315 -7330
rect 12435 -7450 12490 -7330
rect 12610 -7450 12635 -7330
rect 7105 -7495 12635 -7450
rect 7105 -7615 7130 -7495
rect 7250 -7615 7295 -7495
rect 7415 -7615 7460 -7495
rect 7580 -7615 7625 -7495
rect 7745 -7615 7800 -7495
rect 7920 -7615 7965 -7495
rect 8085 -7615 8130 -7495
rect 8250 -7615 8295 -7495
rect 8415 -7615 8470 -7495
rect 8590 -7615 8635 -7495
rect 8755 -7615 8800 -7495
rect 8920 -7615 8965 -7495
rect 9085 -7615 9140 -7495
rect 9260 -7615 9305 -7495
rect 9425 -7615 9470 -7495
rect 9590 -7615 9635 -7495
rect 9755 -7615 9810 -7495
rect 9930 -7615 9975 -7495
rect 10095 -7615 10140 -7495
rect 10260 -7615 10305 -7495
rect 10425 -7615 10480 -7495
rect 10600 -7615 10645 -7495
rect 10765 -7615 10810 -7495
rect 10930 -7615 10975 -7495
rect 11095 -7615 11150 -7495
rect 11270 -7615 11315 -7495
rect 11435 -7615 11480 -7495
rect 11600 -7615 11645 -7495
rect 11765 -7615 11820 -7495
rect 11940 -7615 11985 -7495
rect 12105 -7615 12150 -7495
rect 12270 -7615 12315 -7495
rect 12435 -7615 12490 -7495
rect 12610 -7615 12635 -7495
rect 7105 -7660 12635 -7615
rect 7105 -7780 7130 -7660
rect 7250 -7780 7295 -7660
rect 7415 -7780 7460 -7660
rect 7580 -7780 7625 -7660
rect 7745 -7780 7800 -7660
rect 7920 -7780 7965 -7660
rect 8085 -7780 8130 -7660
rect 8250 -7780 8295 -7660
rect 8415 -7780 8470 -7660
rect 8590 -7780 8635 -7660
rect 8755 -7780 8800 -7660
rect 8920 -7780 8965 -7660
rect 9085 -7780 9140 -7660
rect 9260 -7780 9305 -7660
rect 9425 -7780 9470 -7660
rect 9590 -7780 9635 -7660
rect 9755 -7780 9810 -7660
rect 9930 -7780 9975 -7660
rect 10095 -7780 10140 -7660
rect 10260 -7780 10305 -7660
rect 10425 -7780 10480 -7660
rect 10600 -7780 10645 -7660
rect 10765 -7780 10810 -7660
rect 10930 -7780 10975 -7660
rect 11095 -7780 11150 -7660
rect 11270 -7780 11315 -7660
rect 11435 -7780 11480 -7660
rect 11600 -7780 11645 -7660
rect 11765 -7780 11820 -7660
rect 11940 -7780 11985 -7660
rect 12105 -7780 12150 -7660
rect 12270 -7780 12315 -7660
rect 12435 -7780 12490 -7660
rect 12610 -7780 12635 -7660
rect 7105 -7835 12635 -7780
rect 7105 -7955 7130 -7835
rect 7250 -7955 7295 -7835
rect 7415 -7955 7460 -7835
rect 7580 -7955 7625 -7835
rect 7745 -7955 7800 -7835
rect 7920 -7955 7965 -7835
rect 8085 -7955 8130 -7835
rect 8250 -7955 8295 -7835
rect 8415 -7955 8470 -7835
rect 8590 -7955 8635 -7835
rect 8755 -7955 8800 -7835
rect 8920 -7955 8965 -7835
rect 9085 -7955 9140 -7835
rect 9260 -7955 9305 -7835
rect 9425 -7955 9470 -7835
rect 9590 -7955 9635 -7835
rect 9755 -7955 9810 -7835
rect 9930 -7955 9975 -7835
rect 10095 -7955 10140 -7835
rect 10260 -7955 10305 -7835
rect 10425 -7955 10480 -7835
rect 10600 -7955 10645 -7835
rect 10765 -7955 10810 -7835
rect 10930 -7955 10975 -7835
rect 11095 -7955 11150 -7835
rect 11270 -7955 11315 -7835
rect 11435 -7955 11480 -7835
rect 11600 -7955 11645 -7835
rect 11765 -7955 11820 -7835
rect 11940 -7955 11985 -7835
rect 12105 -7955 12150 -7835
rect 12270 -7955 12315 -7835
rect 12435 -7955 12490 -7835
rect 12610 -7955 12635 -7835
rect 7105 -8000 12635 -7955
rect 7105 -8120 7130 -8000
rect 7250 -8120 7295 -8000
rect 7415 -8120 7460 -8000
rect 7580 -8120 7625 -8000
rect 7745 -8120 7800 -8000
rect 7920 -8120 7965 -8000
rect 8085 -8120 8130 -8000
rect 8250 -8120 8295 -8000
rect 8415 -8120 8470 -8000
rect 8590 -8120 8635 -8000
rect 8755 -8120 8800 -8000
rect 8920 -8120 8965 -8000
rect 9085 -8120 9140 -8000
rect 9260 -8120 9305 -8000
rect 9425 -8120 9470 -8000
rect 9590 -8120 9635 -8000
rect 9755 -8120 9810 -8000
rect 9930 -8120 9975 -8000
rect 10095 -8120 10140 -8000
rect 10260 -8120 10305 -8000
rect 10425 -8120 10480 -8000
rect 10600 -8120 10645 -8000
rect 10765 -8120 10810 -8000
rect 10930 -8120 10975 -8000
rect 11095 -8120 11150 -8000
rect 11270 -8120 11315 -8000
rect 11435 -8120 11480 -8000
rect 11600 -8120 11645 -8000
rect 11765 -8120 11820 -8000
rect 11940 -8120 11985 -8000
rect 12105 -8120 12150 -8000
rect 12270 -8120 12315 -8000
rect 12435 -8120 12490 -8000
rect 12610 -8120 12635 -8000
rect 7105 -8165 12635 -8120
rect 7105 -8285 7130 -8165
rect 7250 -8285 7295 -8165
rect 7415 -8285 7460 -8165
rect 7580 -8285 7625 -8165
rect 7745 -8285 7800 -8165
rect 7920 -8285 7965 -8165
rect 8085 -8285 8130 -8165
rect 8250 -8285 8295 -8165
rect 8415 -8285 8470 -8165
rect 8590 -8285 8635 -8165
rect 8755 -8285 8800 -8165
rect 8920 -8285 8965 -8165
rect 9085 -8285 9140 -8165
rect 9260 -8285 9305 -8165
rect 9425 -8285 9470 -8165
rect 9590 -8285 9635 -8165
rect 9755 -8285 9810 -8165
rect 9930 -8285 9975 -8165
rect 10095 -8285 10140 -8165
rect 10260 -8285 10305 -8165
rect 10425 -8285 10480 -8165
rect 10600 -8285 10645 -8165
rect 10765 -8285 10810 -8165
rect 10930 -8285 10975 -8165
rect 11095 -8285 11150 -8165
rect 11270 -8285 11315 -8165
rect 11435 -8285 11480 -8165
rect 11600 -8285 11645 -8165
rect 11765 -8285 11820 -8165
rect 11940 -8285 11985 -8165
rect 12105 -8285 12150 -8165
rect 12270 -8285 12315 -8165
rect 12435 -8285 12490 -8165
rect 12610 -8285 12635 -8165
rect 7105 -8330 12635 -8285
rect 7105 -8450 7130 -8330
rect 7250 -8450 7295 -8330
rect 7415 -8450 7460 -8330
rect 7580 -8450 7625 -8330
rect 7745 -8450 7800 -8330
rect 7920 -8450 7965 -8330
rect 8085 -8450 8130 -8330
rect 8250 -8450 8295 -8330
rect 8415 -8450 8470 -8330
rect 8590 -8450 8635 -8330
rect 8755 -8450 8800 -8330
rect 8920 -8450 8965 -8330
rect 9085 -8450 9140 -8330
rect 9260 -8450 9305 -8330
rect 9425 -8450 9470 -8330
rect 9590 -8450 9635 -8330
rect 9755 -8450 9810 -8330
rect 9930 -8450 9975 -8330
rect 10095 -8450 10140 -8330
rect 10260 -8450 10305 -8330
rect 10425 -8450 10480 -8330
rect 10600 -8450 10645 -8330
rect 10765 -8450 10810 -8330
rect 10930 -8450 10975 -8330
rect 11095 -8450 11150 -8330
rect 11270 -8450 11315 -8330
rect 11435 -8450 11480 -8330
rect 11600 -8450 11645 -8330
rect 11765 -8450 11820 -8330
rect 11940 -8450 11985 -8330
rect 12105 -8450 12150 -8330
rect 12270 -8450 12315 -8330
rect 12435 -8450 12490 -8330
rect 12610 -8450 12635 -8330
rect 7105 -8505 12635 -8450
rect 7105 -8625 7130 -8505
rect 7250 -8625 7295 -8505
rect 7415 -8625 7460 -8505
rect 7580 -8625 7625 -8505
rect 7745 -8625 7800 -8505
rect 7920 -8625 7965 -8505
rect 8085 -8625 8130 -8505
rect 8250 -8625 8295 -8505
rect 8415 -8625 8470 -8505
rect 8590 -8625 8635 -8505
rect 8755 -8625 8800 -8505
rect 8920 -8625 8965 -8505
rect 9085 -8625 9140 -8505
rect 9260 -8625 9305 -8505
rect 9425 -8625 9470 -8505
rect 9590 -8625 9635 -8505
rect 9755 -8625 9810 -8505
rect 9930 -8625 9975 -8505
rect 10095 -8625 10140 -8505
rect 10260 -8625 10305 -8505
rect 10425 -8625 10480 -8505
rect 10600 -8625 10645 -8505
rect 10765 -8625 10810 -8505
rect 10930 -8625 10975 -8505
rect 11095 -8625 11150 -8505
rect 11270 -8625 11315 -8505
rect 11435 -8625 11480 -8505
rect 11600 -8625 11645 -8505
rect 11765 -8625 11820 -8505
rect 11940 -8625 11985 -8505
rect 12105 -8625 12150 -8505
rect 12270 -8625 12315 -8505
rect 12435 -8625 12490 -8505
rect 12610 -8625 12635 -8505
rect 7105 -8670 12635 -8625
rect 7105 -8790 7130 -8670
rect 7250 -8790 7295 -8670
rect 7415 -8790 7460 -8670
rect 7580 -8790 7625 -8670
rect 7745 -8790 7800 -8670
rect 7920 -8790 7965 -8670
rect 8085 -8790 8130 -8670
rect 8250 -8790 8295 -8670
rect 8415 -8790 8470 -8670
rect 8590 -8790 8635 -8670
rect 8755 -8790 8800 -8670
rect 8920 -8790 8965 -8670
rect 9085 -8790 9140 -8670
rect 9260 -8790 9305 -8670
rect 9425 -8790 9470 -8670
rect 9590 -8790 9635 -8670
rect 9755 -8790 9810 -8670
rect 9930 -8790 9975 -8670
rect 10095 -8790 10140 -8670
rect 10260 -8790 10305 -8670
rect 10425 -8790 10480 -8670
rect 10600 -8790 10645 -8670
rect 10765 -8790 10810 -8670
rect 10930 -8790 10975 -8670
rect 11095 -8790 11150 -8670
rect 11270 -8790 11315 -8670
rect 11435 -8790 11480 -8670
rect 11600 -8790 11645 -8670
rect 11765 -8790 11820 -8670
rect 11940 -8790 11985 -8670
rect 12105 -8790 12150 -8670
rect 12270 -8790 12315 -8670
rect 12435 -8790 12490 -8670
rect 12610 -8790 12635 -8670
rect 7105 -8835 12635 -8790
rect 7105 -8955 7130 -8835
rect 7250 -8955 7295 -8835
rect 7415 -8955 7460 -8835
rect 7580 -8955 7625 -8835
rect 7745 -8955 7800 -8835
rect 7920 -8955 7965 -8835
rect 8085 -8955 8130 -8835
rect 8250 -8955 8295 -8835
rect 8415 -8955 8470 -8835
rect 8590 -8955 8635 -8835
rect 8755 -8955 8800 -8835
rect 8920 -8955 8965 -8835
rect 9085 -8955 9140 -8835
rect 9260 -8955 9305 -8835
rect 9425 -8955 9470 -8835
rect 9590 -8955 9635 -8835
rect 9755 -8955 9810 -8835
rect 9930 -8955 9975 -8835
rect 10095 -8955 10140 -8835
rect 10260 -8955 10305 -8835
rect 10425 -8955 10480 -8835
rect 10600 -8955 10645 -8835
rect 10765 -8955 10810 -8835
rect 10930 -8955 10975 -8835
rect 11095 -8955 11150 -8835
rect 11270 -8955 11315 -8835
rect 11435 -8955 11480 -8835
rect 11600 -8955 11645 -8835
rect 11765 -8955 11820 -8835
rect 11940 -8955 11985 -8835
rect 12105 -8955 12150 -8835
rect 12270 -8955 12315 -8835
rect 12435 -8955 12490 -8835
rect 12610 -8955 12635 -8835
rect 7105 -9000 12635 -8955
rect 7105 -9120 7130 -9000
rect 7250 -9120 7295 -9000
rect 7415 -9120 7460 -9000
rect 7580 -9120 7625 -9000
rect 7745 -9120 7800 -9000
rect 7920 -9120 7965 -9000
rect 8085 -9120 8130 -9000
rect 8250 -9120 8295 -9000
rect 8415 -9120 8470 -9000
rect 8590 -9120 8635 -9000
rect 8755 -9120 8800 -9000
rect 8920 -9120 8965 -9000
rect 9085 -9120 9140 -9000
rect 9260 -9120 9305 -9000
rect 9425 -9120 9470 -9000
rect 9590 -9120 9635 -9000
rect 9755 -9120 9810 -9000
rect 9930 -9120 9975 -9000
rect 10095 -9120 10140 -9000
rect 10260 -9120 10305 -9000
rect 10425 -9120 10480 -9000
rect 10600 -9120 10645 -9000
rect 10765 -9120 10810 -9000
rect 10930 -9120 10975 -9000
rect 11095 -9120 11150 -9000
rect 11270 -9120 11315 -9000
rect 11435 -9120 11480 -9000
rect 11600 -9120 11645 -9000
rect 11765 -9120 11820 -9000
rect 11940 -9120 11985 -9000
rect 12105 -9120 12150 -9000
rect 12270 -9120 12315 -9000
rect 12435 -9120 12490 -9000
rect 12610 -9120 12635 -9000
rect 7105 -9175 12635 -9120
rect 7105 -9295 7130 -9175
rect 7250 -9295 7295 -9175
rect 7415 -9295 7460 -9175
rect 7580 -9295 7625 -9175
rect 7745 -9295 7800 -9175
rect 7920 -9295 7965 -9175
rect 8085 -9295 8130 -9175
rect 8250 -9295 8295 -9175
rect 8415 -9295 8470 -9175
rect 8590 -9295 8635 -9175
rect 8755 -9295 8800 -9175
rect 8920 -9295 8965 -9175
rect 9085 -9295 9140 -9175
rect 9260 -9295 9305 -9175
rect 9425 -9295 9470 -9175
rect 9590 -9295 9635 -9175
rect 9755 -9295 9810 -9175
rect 9930 -9295 9975 -9175
rect 10095 -9295 10140 -9175
rect 10260 -9295 10305 -9175
rect 10425 -9295 10480 -9175
rect 10600 -9295 10645 -9175
rect 10765 -9295 10810 -9175
rect 10930 -9295 10975 -9175
rect 11095 -9295 11150 -9175
rect 11270 -9295 11315 -9175
rect 11435 -9295 11480 -9175
rect 11600 -9295 11645 -9175
rect 11765 -9295 11820 -9175
rect 11940 -9295 11985 -9175
rect 12105 -9295 12150 -9175
rect 12270 -9295 12315 -9175
rect 12435 -9295 12490 -9175
rect 12610 -9295 12635 -9175
rect 7105 -9340 12635 -9295
rect 7105 -9460 7130 -9340
rect 7250 -9460 7295 -9340
rect 7415 -9460 7460 -9340
rect 7580 -9460 7625 -9340
rect 7745 -9460 7800 -9340
rect 7920 -9460 7965 -9340
rect 8085 -9460 8130 -9340
rect 8250 -9460 8295 -9340
rect 8415 -9460 8470 -9340
rect 8590 -9460 8635 -9340
rect 8755 -9460 8800 -9340
rect 8920 -9460 8965 -9340
rect 9085 -9460 9140 -9340
rect 9260 -9460 9305 -9340
rect 9425 -9460 9470 -9340
rect 9590 -9460 9635 -9340
rect 9755 -9460 9810 -9340
rect 9930 -9460 9975 -9340
rect 10095 -9460 10140 -9340
rect 10260 -9460 10305 -9340
rect 10425 -9460 10480 -9340
rect 10600 -9460 10645 -9340
rect 10765 -9460 10810 -9340
rect 10930 -9460 10975 -9340
rect 11095 -9460 11150 -9340
rect 11270 -9460 11315 -9340
rect 11435 -9460 11480 -9340
rect 11600 -9460 11645 -9340
rect 11765 -9460 11820 -9340
rect 11940 -9460 11985 -9340
rect 12105 -9460 12150 -9340
rect 12270 -9460 12315 -9340
rect 12435 -9460 12490 -9340
rect 12610 -9460 12635 -9340
rect 7105 -9505 12635 -9460
rect 7105 -9625 7130 -9505
rect 7250 -9625 7295 -9505
rect 7415 -9625 7460 -9505
rect 7580 -9625 7625 -9505
rect 7745 -9625 7800 -9505
rect 7920 -9625 7965 -9505
rect 8085 -9625 8130 -9505
rect 8250 -9625 8295 -9505
rect 8415 -9625 8470 -9505
rect 8590 -9625 8635 -9505
rect 8755 -9625 8800 -9505
rect 8920 -9625 8965 -9505
rect 9085 -9625 9140 -9505
rect 9260 -9625 9305 -9505
rect 9425 -9625 9470 -9505
rect 9590 -9625 9635 -9505
rect 9755 -9625 9810 -9505
rect 9930 -9625 9975 -9505
rect 10095 -9625 10140 -9505
rect 10260 -9625 10305 -9505
rect 10425 -9625 10480 -9505
rect 10600 -9625 10645 -9505
rect 10765 -9625 10810 -9505
rect 10930 -9625 10975 -9505
rect 11095 -9625 11150 -9505
rect 11270 -9625 11315 -9505
rect 11435 -9625 11480 -9505
rect 11600 -9625 11645 -9505
rect 11765 -9625 11820 -9505
rect 11940 -9625 11985 -9505
rect 12105 -9625 12150 -9505
rect 12270 -9625 12315 -9505
rect 12435 -9625 12490 -9505
rect 12610 -9625 12635 -9505
rect 7105 -9670 12635 -9625
rect 7105 -9790 7130 -9670
rect 7250 -9790 7295 -9670
rect 7415 -9790 7460 -9670
rect 7580 -9790 7625 -9670
rect 7745 -9790 7800 -9670
rect 7920 -9790 7965 -9670
rect 8085 -9790 8130 -9670
rect 8250 -9790 8295 -9670
rect 8415 -9790 8470 -9670
rect 8590 -9790 8635 -9670
rect 8755 -9790 8800 -9670
rect 8920 -9790 8965 -9670
rect 9085 -9790 9140 -9670
rect 9260 -9790 9305 -9670
rect 9425 -9790 9470 -9670
rect 9590 -9790 9635 -9670
rect 9755 -9790 9810 -9670
rect 9930 -9790 9975 -9670
rect 10095 -9790 10140 -9670
rect 10260 -9790 10305 -9670
rect 10425 -9790 10480 -9670
rect 10600 -9790 10645 -9670
rect 10765 -9790 10810 -9670
rect 10930 -9790 10975 -9670
rect 11095 -9790 11150 -9670
rect 11270 -9790 11315 -9670
rect 11435 -9790 11480 -9670
rect 11600 -9790 11645 -9670
rect 11765 -9790 11820 -9670
rect 11940 -9790 11985 -9670
rect 12105 -9790 12150 -9670
rect 12270 -9790 12315 -9670
rect 12435 -9790 12490 -9670
rect 12610 -9790 12635 -9670
rect 7105 -9860 12635 -9790
rect 12795 -4310 18325 -4285
rect 12795 -4430 12820 -4310
rect 12940 -4430 12985 -4310
rect 13105 -4430 13150 -4310
rect 13270 -4430 13315 -4310
rect 13435 -4430 13490 -4310
rect 13610 -4430 13655 -4310
rect 13775 -4430 13820 -4310
rect 13940 -4430 13985 -4310
rect 14105 -4430 14160 -4310
rect 14280 -4430 14325 -4310
rect 14445 -4430 14490 -4310
rect 14610 -4430 14655 -4310
rect 14775 -4430 14830 -4310
rect 14950 -4430 14995 -4310
rect 15115 -4430 15160 -4310
rect 15280 -4430 15325 -4310
rect 15445 -4430 15500 -4310
rect 15620 -4430 15665 -4310
rect 15785 -4430 15830 -4310
rect 15950 -4430 15995 -4310
rect 16115 -4430 16170 -4310
rect 16290 -4430 16335 -4310
rect 16455 -4430 16500 -4310
rect 16620 -4430 16665 -4310
rect 16785 -4430 16840 -4310
rect 16960 -4430 17005 -4310
rect 17125 -4430 17170 -4310
rect 17290 -4430 17335 -4310
rect 17455 -4430 17510 -4310
rect 17630 -4430 17675 -4310
rect 17795 -4430 17840 -4310
rect 17960 -4430 18005 -4310
rect 18125 -4430 18180 -4310
rect 18300 -4430 18325 -4310
rect 12795 -4485 18325 -4430
rect 12795 -4605 12820 -4485
rect 12940 -4605 12985 -4485
rect 13105 -4605 13150 -4485
rect 13270 -4605 13315 -4485
rect 13435 -4605 13490 -4485
rect 13610 -4605 13655 -4485
rect 13775 -4605 13820 -4485
rect 13940 -4605 13985 -4485
rect 14105 -4605 14160 -4485
rect 14280 -4605 14325 -4485
rect 14445 -4605 14490 -4485
rect 14610 -4605 14655 -4485
rect 14775 -4605 14830 -4485
rect 14950 -4605 14995 -4485
rect 15115 -4605 15160 -4485
rect 15280 -4605 15325 -4485
rect 15445 -4605 15500 -4485
rect 15620 -4605 15665 -4485
rect 15785 -4605 15830 -4485
rect 15950 -4605 15995 -4485
rect 16115 -4605 16170 -4485
rect 16290 -4605 16335 -4485
rect 16455 -4605 16500 -4485
rect 16620 -4605 16665 -4485
rect 16785 -4605 16840 -4485
rect 16960 -4605 17005 -4485
rect 17125 -4605 17170 -4485
rect 17290 -4605 17335 -4485
rect 17455 -4605 17510 -4485
rect 17630 -4605 17675 -4485
rect 17795 -4605 17840 -4485
rect 17960 -4605 18005 -4485
rect 18125 -4605 18180 -4485
rect 18300 -4605 18325 -4485
rect 12795 -4650 18325 -4605
rect 12795 -4770 12820 -4650
rect 12940 -4770 12985 -4650
rect 13105 -4770 13150 -4650
rect 13270 -4770 13315 -4650
rect 13435 -4770 13490 -4650
rect 13610 -4770 13655 -4650
rect 13775 -4770 13820 -4650
rect 13940 -4770 13985 -4650
rect 14105 -4770 14160 -4650
rect 14280 -4770 14325 -4650
rect 14445 -4770 14490 -4650
rect 14610 -4770 14655 -4650
rect 14775 -4770 14830 -4650
rect 14950 -4770 14995 -4650
rect 15115 -4770 15160 -4650
rect 15280 -4770 15325 -4650
rect 15445 -4770 15500 -4650
rect 15620 -4770 15665 -4650
rect 15785 -4770 15830 -4650
rect 15950 -4770 15995 -4650
rect 16115 -4770 16170 -4650
rect 16290 -4770 16335 -4650
rect 16455 -4770 16500 -4650
rect 16620 -4770 16665 -4650
rect 16785 -4770 16840 -4650
rect 16960 -4770 17005 -4650
rect 17125 -4770 17170 -4650
rect 17290 -4770 17335 -4650
rect 17455 -4770 17510 -4650
rect 17630 -4770 17675 -4650
rect 17795 -4770 17840 -4650
rect 17960 -4770 18005 -4650
rect 18125 -4770 18180 -4650
rect 18300 -4770 18325 -4650
rect 12795 -4815 18325 -4770
rect 12795 -4935 12820 -4815
rect 12940 -4935 12985 -4815
rect 13105 -4935 13150 -4815
rect 13270 -4935 13315 -4815
rect 13435 -4935 13490 -4815
rect 13610 -4935 13655 -4815
rect 13775 -4935 13820 -4815
rect 13940 -4935 13985 -4815
rect 14105 -4935 14160 -4815
rect 14280 -4935 14325 -4815
rect 14445 -4935 14490 -4815
rect 14610 -4935 14655 -4815
rect 14775 -4935 14830 -4815
rect 14950 -4935 14995 -4815
rect 15115 -4935 15160 -4815
rect 15280 -4935 15325 -4815
rect 15445 -4935 15500 -4815
rect 15620 -4935 15665 -4815
rect 15785 -4935 15830 -4815
rect 15950 -4935 15995 -4815
rect 16115 -4935 16170 -4815
rect 16290 -4935 16335 -4815
rect 16455 -4935 16500 -4815
rect 16620 -4935 16665 -4815
rect 16785 -4935 16840 -4815
rect 16960 -4935 17005 -4815
rect 17125 -4935 17170 -4815
rect 17290 -4935 17335 -4815
rect 17455 -4935 17510 -4815
rect 17630 -4935 17675 -4815
rect 17795 -4935 17840 -4815
rect 17960 -4935 18005 -4815
rect 18125 -4935 18180 -4815
rect 18300 -4935 18325 -4815
rect 12795 -4980 18325 -4935
rect 12795 -5100 12820 -4980
rect 12940 -5100 12985 -4980
rect 13105 -5100 13150 -4980
rect 13270 -5100 13315 -4980
rect 13435 -5100 13490 -4980
rect 13610 -5100 13655 -4980
rect 13775 -5100 13820 -4980
rect 13940 -5100 13985 -4980
rect 14105 -5100 14160 -4980
rect 14280 -5100 14325 -4980
rect 14445 -5100 14490 -4980
rect 14610 -5100 14655 -4980
rect 14775 -5100 14830 -4980
rect 14950 -5100 14995 -4980
rect 15115 -5100 15160 -4980
rect 15280 -5100 15325 -4980
rect 15445 -5100 15500 -4980
rect 15620 -5100 15665 -4980
rect 15785 -5100 15830 -4980
rect 15950 -5100 15995 -4980
rect 16115 -5100 16170 -4980
rect 16290 -5100 16335 -4980
rect 16455 -5100 16500 -4980
rect 16620 -5100 16665 -4980
rect 16785 -5100 16840 -4980
rect 16960 -5100 17005 -4980
rect 17125 -5100 17170 -4980
rect 17290 -5100 17335 -4980
rect 17455 -5100 17510 -4980
rect 17630 -5100 17675 -4980
rect 17795 -5100 17840 -4980
rect 17960 -5100 18005 -4980
rect 18125 -5100 18180 -4980
rect 18300 -5100 18325 -4980
rect 12795 -5155 18325 -5100
rect 12795 -5275 12820 -5155
rect 12940 -5275 12985 -5155
rect 13105 -5275 13150 -5155
rect 13270 -5275 13315 -5155
rect 13435 -5275 13490 -5155
rect 13610 -5275 13655 -5155
rect 13775 -5275 13820 -5155
rect 13940 -5275 13985 -5155
rect 14105 -5275 14160 -5155
rect 14280 -5275 14325 -5155
rect 14445 -5275 14490 -5155
rect 14610 -5275 14655 -5155
rect 14775 -5275 14830 -5155
rect 14950 -5275 14995 -5155
rect 15115 -5275 15160 -5155
rect 15280 -5275 15325 -5155
rect 15445 -5275 15500 -5155
rect 15620 -5275 15665 -5155
rect 15785 -5275 15830 -5155
rect 15950 -5275 15995 -5155
rect 16115 -5275 16170 -5155
rect 16290 -5275 16335 -5155
rect 16455 -5275 16500 -5155
rect 16620 -5275 16665 -5155
rect 16785 -5275 16840 -5155
rect 16960 -5275 17005 -5155
rect 17125 -5275 17170 -5155
rect 17290 -5275 17335 -5155
rect 17455 -5275 17510 -5155
rect 17630 -5275 17675 -5155
rect 17795 -5275 17840 -5155
rect 17960 -5275 18005 -5155
rect 18125 -5275 18180 -5155
rect 18300 -5275 18325 -5155
rect 12795 -5320 18325 -5275
rect 12795 -5440 12820 -5320
rect 12940 -5440 12985 -5320
rect 13105 -5440 13150 -5320
rect 13270 -5440 13315 -5320
rect 13435 -5440 13490 -5320
rect 13610 -5440 13655 -5320
rect 13775 -5440 13820 -5320
rect 13940 -5440 13985 -5320
rect 14105 -5440 14160 -5320
rect 14280 -5440 14325 -5320
rect 14445 -5440 14490 -5320
rect 14610 -5440 14655 -5320
rect 14775 -5440 14830 -5320
rect 14950 -5440 14995 -5320
rect 15115 -5440 15160 -5320
rect 15280 -5440 15325 -5320
rect 15445 -5440 15500 -5320
rect 15620 -5440 15665 -5320
rect 15785 -5440 15830 -5320
rect 15950 -5440 15995 -5320
rect 16115 -5440 16170 -5320
rect 16290 -5440 16335 -5320
rect 16455 -5440 16500 -5320
rect 16620 -5440 16665 -5320
rect 16785 -5440 16840 -5320
rect 16960 -5440 17005 -5320
rect 17125 -5440 17170 -5320
rect 17290 -5440 17335 -5320
rect 17455 -5440 17510 -5320
rect 17630 -5440 17675 -5320
rect 17795 -5440 17840 -5320
rect 17960 -5440 18005 -5320
rect 18125 -5440 18180 -5320
rect 18300 -5440 18325 -5320
rect 12795 -5485 18325 -5440
rect 12795 -5605 12820 -5485
rect 12940 -5605 12985 -5485
rect 13105 -5605 13150 -5485
rect 13270 -5605 13315 -5485
rect 13435 -5605 13490 -5485
rect 13610 -5605 13655 -5485
rect 13775 -5605 13820 -5485
rect 13940 -5605 13985 -5485
rect 14105 -5605 14160 -5485
rect 14280 -5605 14325 -5485
rect 14445 -5605 14490 -5485
rect 14610 -5605 14655 -5485
rect 14775 -5605 14830 -5485
rect 14950 -5605 14995 -5485
rect 15115 -5605 15160 -5485
rect 15280 -5605 15325 -5485
rect 15445 -5605 15500 -5485
rect 15620 -5605 15665 -5485
rect 15785 -5605 15830 -5485
rect 15950 -5605 15995 -5485
rect 16115 -5605 16170 -5485
rect 16290 -5605 16335 -5485
rect 16455 -5605 16500 -5485
rect 16620 -5605 16665 -5485
rect 16785 -5605 16840 -5485
rect 16960 -5605 17005 -5485
rect 17125 -5605 17170 -5485
rect 17290 -5605 17335 -5485
rect 17455 -5605 17510 -5485
rect 17630 -5605 17675 -5485
rect 17795 -5605 17840 -5485
rect 17960 -5605 18005 -5485
rect 18125 -5605 18180 -5485
rect 18300 -5605 18325 -5485
rect 12795 -5650 18325 -5605
rect 12795 -5770 12820 -5650
rect 12940 -5770 12985 -5650
rect 13105 -5770 13150 -5650
rect 13270 -5770 13315 -5650
rect 13435 -5770 13490 -5650
rect 13610 -5770 13655 -5650
rect 13775 -5770 13820 -5650
rect 13940 -5770 13985 -5650
rect 14105 -5770 14160 -5650
rect 14280 -5770 14325 -5650
rect 14445 -5770 14490 -5650
rect 14610 -5770 14655 -5650
rect 14775 -5770 14830 -5650
rect 14950 -5770 14995 -5650
rect 15115 -5770 15160 -5650
rect 15280 -5770 15325 -5650
rect 15445 -5770 15500 -5650
rect 15620 -5770 15665 -5650
rect 15785 -5770 15830 -5650
rect 15950 -5770 15995 -5650
rect 16115 -5770 16170 -5650
rect 16290 -5770 16335 -5650
rect 16455 -5770 16500 -5650
rect 16620 -5770 16665 -5650
rect 16785 -5770 16840 -5650
rect 16960 -5770 17005 -5650
rect 17125 -5770 17170 -5650
rect 17290 -5770 17335 -5650
rect 17455 -5770 17510 -5650
rect 17630 -5770 17675 -5650
rect 17795 -5770 17840 -5650
rect 17960 -5770 18005 -5650
rect 18125 -5770 18180 -5650
rect 18300 -5770 18325 -5650
rect 12795 -5825 18325 -5770
rect 12795 -5945 12820 -5825
rect 12940 -5945 12985 -5825
rect 13105 -5945 13150 -5825
rect 13270 -5945 13315 -5825
rect 13435 -5945 13490 -5825
rect 13610 -5945 13655 -5825
rect 13775 -5945 13820 -5825
rect 13940 -5945 13985 -5825
rect 14105 -5945 14160 -5825
rect 14280 -5945 14325 -5825
rect 14445 -5945 14490 -5825
rect 14610 -5945 14655 -5825
rect 14775 -5945 14830 -5825
rect 14950 -5945 14995 -5825
rect 15115 -5945 15160 -5825
rect 15280 -5945 15325 -5825
rect 15445 -5945 15500 -5825
rect 15620 -5945 15665 -5825
rect 15785 -5945 15830 -5825
rect 15950 -5945 15995 -5825
rect 16115 -5945 16170 -5825
rect 16290 -5945 16335 -5825
rect 16455 -5945 16500 -5825
rect 16620 -5945 16665 -5825
rect 16785 -5945 16840 -5825
rect 16960 -5945 17005 -5825
rect 17125 -5945 17170 -5825
rect 17290 -5945 17335 -5825
rect 17455 -5945 17510 -5825
rect 17630 -5945 17675 -5825
rect 17795 -5945 17840 -5825
rect 17960 -5945 18005 -5825
rect 18125 -5945 18180 -5825
rect 18300 -5945 18325 -5825
rect 12795 -5990 18325 -5945
rect 12795 -6110 12820 -5990
rect 12940 -6110 12985 -5990
rect 13105 -6110 13150 -5990
rect 13270 -6110 13315 -5990
rect 13435 -6110 13490 -5990
rect 13610 -6110 13655 -5990
rect 13775 -6110 13820 -5990
rect 13940 -6110 13985 -5990
rect 14105 -6110 14160 -5990
rect 14280 -6110 14325 -5990
rect 14445 -6110 14490 -5990
rect 14610 -6110 14655 -5990
rect 14775 -6110 14830 -5990
rect 14950 -6110 14995 -5990
rect 15115 -6110 15160 -5990
rect 15280 -6110 15325 -5990
rect 15445 -6110 15500 -5990
rect 15620 -6110 15665 -5990
rect 15785 -6110 15830 -5990
rect 15950 -6110 15995 -5990
rect 16115 -6110 16170 -5990
rect 16290 -6110 16335 -5990
rect 16455 -6110 16500 -5990
rect 16620 -6110 16665 -5990
rect 16785 -6110 16840 -5990
rect 16960 -6110 17005 -5990
rect 17125 -6110 17170 -5990
rect 17290 -6110 17335 -5990
rect 17455 -6110 17510 -5990
rect 17630 -6110 17675 -5990
rect 17795 -6110 17840 -5990
rect 17960 -6110 18005 -5990
rect 18125 -6110 18180 -5990
rect 18300 -6110 18325 -5990
rect 12795 -6155 18325 -6110
rect 12795 -6275 12820 -6155
rect 12940 -6275 12985 -6155
rect 13105 -6275 13150 -6155
rect 13270 -6275 13315 -6155
rect 13435 -6275 13490 -6155
rect 13610 -6275 13655 -6155
rect 13775 -6275 13820 -6155
rect 13940 -6275 13985 -6155
rect 14105 -6275 14160 -6155
rect 14280 -6275 14325 -6155
rect 14445 -6275 14490 -6155
rect 14610 -6275 14655 -6155
rect 14775 -6275 14830 -6155
rect 14950 -6275 14995 -6155
rect 15115 -6275 15160 -6155
rect 15280 -6275 15325 -6155
rect 15445 -6275 15500 -6155
rect 15620 -6275 15665 -6155
rect 15785 -6275 15830 -6155
rect 15950 -6275 15995 -6155
rect 16115 -6275 16170 -6155
rect 16290 -6275 16335 -6155
rect 16455 -6275 16500 -6155
rect 16620 -6275 16665 -6155
rect 16785 -6275 16840 -6155
rect 16960 -6275 17005 -6155
rect 17125 -6275 17170 -6155
rect 17290 -6275 17335 -6155
rect 17455 -6275 17510 -6155
rect 17630 -6275 17675 -6155
rect 17795 -6275 17840 -6155
rect 17960 -6275 18005 -6155
rect 18125 -6275 18180 -6155
rect 18300 -6275 18325 -6155
rect 12795 -6320 18325 -6275
rect 12795 -6440 12820 -6320
rect 12940 -6440 12985 -6320
rect 13105 -6440 13150 -6320
rect 13270 -6440 13315 -6320
rect 13435 -6440 13490 -6320
rect 13610 -6440 13655 -6320
rect 13775 -6440 13820 -6320
rect 13940 -6440 13985 -6320
rect 14105 -6440 14160 -6320
rect 14280 -6440 14325 -6320
rect 14445 -6440 14490 -6320
rect 14610 -6440 14655 -6320
rect 14775 -6440 14830 -6320
rect 14950 -6440 14995 -6320
rect 15115 -6440 15160 -6320
rect 15280 -6440 15325 -6320
rect 15445 -6440 15500 -6320
rect 15620 -6440 15665 -6320
rect 15785 -6440 15830 -6320
rect 15950 -6440 15995 -6320
rect 16115 -6440 16170 -6320
rect 16290 -6440 16335 -6320
rect 16455 -6440 16500 -6320
rect 16620 -6440 16665 -6320
rect 16785 -6440 16840 -6320
rect 16960 -6440 17005 -6320
rect 17125 -6440 17170 -6320
rect 17290 -6440 17335 -6320
rect 17455 -6440 17510 -6320
rect 17630 -6440 17675 -6320
rect 17795 -6440 17840 -6320
rect 17960 -6440 18005 -6320
rect 18125 -6440 18180 -6320
rect 18300 -6440 18325 -6320
rect 12795 -6495 18325 -6440
rect 12795 -6615 12820 -6495
rect 12940 -6615 12985 -6495
rect 13105 -6615 13150 -6495
rect 13270 -6615 13315 -6495
rect 13435 -6615 13490 -6495
rect 13610 -6615 13655 -6495
rect 13775 -6615 13820 -6495
rect 13940 -6615 13985 -6495
rect 14105 -6615 14160 -6495
rect 14280 -6615 14325 -6495
rect 14445 -6615 14490 -6495
rect 14610 -6615 14655 -6495
rect 14775 -6615 14830 -6495
rect 14950 -6615 14995 -6495
rect 15115 -6615 15160 -6495
rect 15280 -6615 15325 -6495
rect 15445 -6615 15500 -6495
rect 15620 -6615 15665 -6495
rect 15785 -6615 15830 -6495
rect 15950 -6615 15995 -6495
rect 16115 -6615 16170 -6495
rect 16290 -6615 16335 -6495
rect 16455 -6615 16500 -6495
rect 16620 -6615 16665 -6495
rect 16785 -6615 16840 -6495
rect 16960 -6615 17005 -6495
rect 17125 -6615 17170 -6495
rect 17290 -6615 17335 -6495
rect 17455 -6615 17510 -6495
rect 17630 -6615 17675 -6495
rect 17795 -6615 17840 -6495
rect 17960 -6615 18005 -6495
rect 18125 -6615 18180 -6495
rect 18300 -6615 18325 -6495
rect 12795 -6660 18325 -6615
rect 12795 -6780 12820 -6660
rect 12940 -6780 12985 -6660
rect 13105 -6780 13150 -6660
rect 13270 -6780 13315 -6660
rect 13435 -6780 13490 -6660
rect 13610 -6780 13655 -6660
rect 13775 -6780 13820 -6660
rect 13940 -6780 13985 -6660
rect 14105 -6780 14160 -6660
rect 14280 -6780 14325 -6660
rect 14445 -6780 14490 -6660
rect 14610 -6780 14655 -6660
rect 14775 -6780 14830 -6660
rect 14950 -6780 14995 -6660
rect 15115 -6780 15160 -6660
rect 15280 -6780 15325 -6660
rect 15445 -6780 15500 -6660
rect 15620 -6780 15665 -6660
rect 15785 -6780 15830 -6660
rect 15950 -6780 15995 -6660
rect 16115 -6780 16170 -6660
rect 16290 -6780 16335 -6660
rect 16455 -6780 16500 -6660
rect 16620 -6780 16665 -6660
rect 16785 -6780 16840 -6660
rect 16960 -6780 17005 -6660
rect 17125 -6780 17170 -6660
rect 17290 -6780 17335 -6660
rect 17455 -6780 17510 -6660
rect 17630 -6780 17675 -6660
rect 17795 -6780 17840 -6660
rect 17960 -6780 18005 -6660
rect 18125 -6780 18180 -6660
rect 18300 -6780 18325 -6660
rect 12795 -6825 18325 -6780
rect 12795 -6945 12820 -6825
rect 12940 -6945 12985 -6825
rect 13105 -6945 13150 -6825
rect 13270 -6945 13315 -6825
rect 13435 -6945 13490 -6825
rect 13610 -6945 13655 -6825
rect 13775 -6945 13820 -6825
rect 13940 -6945 13985 -6825
rect 14105 -6945 14160 -6825
rect 14280 -6945 14325 -6825
rect 14445 -6945 14490 -6825
rect 14610 -6945 14655 -6825
rect 14775 -6945 14830 -6825
rect 14950 -6945 14995 -6825
rect 15115 -6945 15160 -6825
rect 15280 -6945 15325 -6825
rect 15445 -6945 15500 -6825
rect 15620 -6945 15665 -6825
rect 15785 -6945 15830 -6825
rect 15950 -6945 15995 -6825
rect 16115 -6945 16170 -6825
rect 16290 -6945 16335 -6825
rect 16455 -6945 16500 -6825
rect 16620 -6945 16665 -6825
rect 16785 -6945 16840 -6825
rect 16960 -6945 17005 -6825
rect 17125 -6945 17170 -6825
rect 17290 -6945 17335 -6825
rect 17455 -6945 17510 -6825
rect 17630 -6945 17675 -6825
rect 17795 -6945 17840 -6825
rect 17960 -6945 18005 -6825
rect 18125 -6945 18180 -6825
rect 18300 -6945 18325 -6825
rect 12795 -6990 18325 -6945
rect 12795 -7110 12820 -6990
rect 12940 -7110 12985 -6990
rect 13105 -7110 13150 -6990
rect 13270 -7110 13315 -6990
rect 13435 -7110 13490 -6990
rect 13610 -7110 13655 -6990
rect 13775 -7110 13820 -6990
rect 13940 -7110 13985 -6990
rect 14105 -7110 14160 -6990
rect 14280 -7110 14325 -6990
rect 14445 -7110 14490 -6990
rect 14610 -7110 14655 -6990
rect 14775 -7110 14830 -6990
rect 14950 -7110 14995 -6990
rect 15115 -7110 15160 -6990
rect 15280 -7110 15325 -6990
rect 15445 -7110 15500 -6990
rect 15620 -7110 15665 -6990
rect 15785 -7110 15830 -6990
rect 15950 -7110 15995 -6990
rect 16115 -7110 16170 -6990
rect 16290 -7110 16335 -6990
rect 16455 -7110 16500 -6990
rect 16620 -7110 16665 -6990
rect 16785 -7110 16840 -6990
rect 16960 -7110 17005 -6990
rect 17125 -7110 17170 -6990
rect 17290 -7110 17335 -6990
rect 17455 -7110 17510 -6990
rect 17630 -7110 17675 -6990
rect 17795 -7110 17840 -6990
rect 17960 -7110 18005 -6990
rect 18125 -7110 18180 -6990
rect 18300 -7110 18325 -6990
rect 12795 -7165 18325 -7110
rect 12795 -7285 12820 -7165
rect 12940 -7285 12985 -7165
rect 13105 -7285 13150 -7165
rect 13270 -7285 13315 -7165
rect 13435 -7285 13490 -7165
rect 13610 -7285 13655 -7165
rect 13775 -7285 13820 -7165
rect 13940 -7285 13985 -7165
rect 14105 -7285 14160 -7165
rect 14280 -7285 14325 -7165
rect 14445 -7285 14490 -7165
rect 14610 -7285 14655 -7165
rect 14775 -7285 14830 -7165
rect 14950 -7285 14995 -7165
rect 15115 -7285 15160 -7165
rect 15280 -7285 15325 -7165
rect 15445 -7285 15500 -7165
rect 15620 -7285 15665 -7165
rect 15785 -7285 15830 -7165
rect 15950 -7285 15995 -7165
rect 16115 -7285 16170 -7165
rect 16290 -7285 16335 -7165
rect 16455 -7285 16500 -7165
rect 16620 -7285 16665 -7165
rect 16785 -7285 16840 -7165
rect 16960 -7285 17005 -7165
rect 17125 -7285 17170 -7165
rect 17290 -7285 17335 -7165
rect 17455 -7285 17510 -7165
rect 17630 -7285 17675 -7165
rect 17795 -7285 17840 -7165
rect 17960 -7285 18005 -7165
rect 18125 -7285 18180 -7165
rect 18300 -7285 18325 -7165
rect 12795 -7330 18325 -7285
rect 12795 -7450 12820 -7330
rect 12940 -7450 12985 -7330
rect 13105 -7450 13150 -7330
rect 13270 -7450 13315 -7330
rect 13435 -7450 13490 -7330
rect 13610 -7450 13655 -7330
rect 13775 -7450 13820 -7330
rect 13940 -7450 13985 -7330
rect 14105 -7450 14160 -7330
rect 14280 -7450 14325 -7330
rect 14445 -7450 14490 -7330
rect 14610 -7450 14655 -7330
rect 14775 -7450 14830 -7330
rect 14950 -7450 14995 -7330
rect 15115 -7450 15160 -7330
rect 15280 -7450 15325 -7330
rect 15445 -7450 15500 -7330
rect 15620 -7450 15665 -7330
rect 15785 -7450 15830 -7330
rect 15950 -7450 15995 -7330
rect 16115 -7450 16170 -7330
rect 16290 -7450 16335 -7330
rect 16455 -7450 16500 -7330
rect 16620 -7450 16665 -7330
rect 16785 -7450 16840 -7330
rect 16960 -7450 17005 -7330
rect 17125 -7450 17170 -7330
rect 17290 -7450 17335 -7330
rect 17455 -7450 17510 -7330
rect 17630 -7450 17675 -7330
rect 17795 -7450 17840 -7330
rect 17960 -7450 18005 -7330
rect 18125 -7450 18180 -7330
rect 18300 -7450 18325 -7330
rect 12795 -7495 18325 -7450
rect 12795 -7615 12820 -7495
rect 12940 -7615 12985 -7495
rect 13105 -7615 13150 -7495
rect 13270 -7615 13315 -7495
rect 13435 -7615 13490 -7495
rect 13610 -7615 13655 -7495
rect 13775 -7615 13820 -7495
rect 13940 -7615 13985 -7495
rect 14105 -7615 14160 -7495
rect 14280 -7615 14325 -7495
rect 14445 -7615 14490 -7495
rect 14610 -7615 14655 -7495
rect 14775 -7615 14830 -7495
rect 14950 -7615 14995 -7495
rect 15115 -7615 15160 -7495
rect 15280 -7615 15325 -7495
rect 15445 -7615 15500 -7495
rect 15620 -7615 15665 -7495
rect 15785 -7615 15830 -7495
rect 15950 -7615 15995 -7495
rect 16115 -7615 16170 -7495
rect 16290 -7615 16335 -7495
rect 16455 -7615 16500 -7495
rect 16620 -7615 16665 -7495
rect 16785 -7615 16840 -7495
rect 16960 -7615 17005 -7495
rect 17125 -7615 17170 -7495
rect 17290 -7615 17335 -7495
rect 17455 -7615 17510 -7495
rect 17630 -7615 17675 -7495
rect 17795 -7615 17840 -7495
rect 17960 -7615 18005 -7495
rect 18125 -7615 18180 -7495
rect 18300 -7615 18325 -7495
rect 12795 -7660 18325 -7615
rect 12795 -7780 12820 -7660
rect 12940 -7780 12985 -7660
rect 13105 -7780 13150 -7660
rect 13270 -7780 13315 -7660
rect 13435 -7780 13490 -7660
rect 13610 -7780 13655 -7660
rect 13775 -7780 13820 -7660
rect 13940 -7780 13985 -7660
rect 14105 -7780 14160 -7660
rect 14280 -7780 14325 -7660
rect 14445 -7780 14490 -7660
rect 14610 -7780 14655 -7660
rect 14775 -7780 14830 -7660
rect 14950 -7780 14995 -7660
rect 15115 -7780 15160 -7660
rect 15280 -7780 15325 -7660
rect 15445 -7780 15500 -7660
rect 15620 -7780 15665 -7660
rect 15785 -7780 15830 -7660
rect 15950 -7780 15995 -7660
rect 16115 -7780 16170 -7660
rect 16290 -7780 16335 -7660
rect 16455 -7780 16500 -7660
rect 16620 -7780 16665 -7660
rect 16785 -7780 16840 -7660
rect 16960 -7780 17005 -7660
rect 17125 -7780 17170 -7660
rect 17290 -7780 17335 -7660
rect 17455 -7780 17510 -7660
rect 17630 -7780 17675 -7660
rect 17795 -7780 17840 -7660
rect 17960 -7780 18005 -7660
rect 18125 -7780 18180 -7660
rect 18300 -7780 18325 -7660
rect 12795 -7835 18325 -7780
rect 12795 -7955 12820 -7835
rect 12940 -7955 12985 -7835
rect 13105 -7955 13150 -7835
rect 13270 -7955 13315 -7835
rect 13435 -7955 13490 -7835
rect 13610 -7955 13655 -7835
rect 13775 -7955 13820 -7835
rect 13940 -7955 13985 -7835
rect 14105 -7955 14160 -7835
rect 14280 -7955 14325 -7835
rect 14445 -7955 14490 -7835
rect 14610 -7955 14655 -7835
rect 14775 -7955 14830 -7835
rect 14950 -7955 14995 -7835
rect 15115 -7955 15160 -7835
rect 15280 -7955 15325 -7835
rect 15445 -7955 15500 -7835
rect 15620 -7955 15665 -7835
rect 15785 -7955 15830 -7835
rect 15950 -7955 15995 -7835
rect 16115 -7955 16170 -7835
rect 16290 -7955 16335 -7835
rect 16455 -7955 16500 -7835
rect 16620 -7955 16665 -7835
rect 16785 -7955 16840 -7835
rect 16960 -7955 17005 -7835
rect 17125 -7955 17170 -7835
rect 17290 -7955 17335 -7835
rect 17455 -7955 17510 -7835
rect 17630 -7955 17675 -7835
rect 17795 -7955 17840 -7835
rect 17960 -7955 18005 -7835
rect 18125 -7955 18180 -7835
rect 18300 -7955 18325 -7835
rect 12795 -8000 18325 -7955
rect 12795 -8120 12820 -8000
rect 12940 -8120 12985 -8000
rect 13105 -8120 13150 -8000
rect 13270 -8120 13315 -8000
rect 13435 -8120 13490 -8000
rect 13610 -8120 13655 -8000
rect 13775 -8120 13820 -8000
rect 13940 -8120 13985 -8000
rect 14105 -8120 14160 -8000
rect 14280 -8120 14325 -8000
rect 14445 -8120 14490 -8000
rect 14610 -8120 14655 -8000
rect 14775 -8120 14830 -8000
rect 14950 -8120 14995 -8000
rect 15115 -8120 15160 -8000
rect 15280 -8120 15325 -8000
rect 15445 -8120 15500 -8000
rect 15620 -8120 15665 -8000
rect 15785 -8120 15830 -8000
rect 15950 -8120 15995 -8000
rect 16115 -8120 16170 -8000
rect 16290 -8120 16335 -8000
rect 16455 -8120 16500 -8000
rect 16620 -8120 16665 -8000
rect 16785 -8120 16840 -8000
rect 16960 -8120 17005 -8000
rect 17125 -8120 17170 -8000
rect 17290 -8120 17335 -8000
rect 17455 -8120 17510 -8000
rect 17630 -8120 17675 -8000
rect 17795 -8120 17840 -8000
rect 17960 -8120 18005 -8000
rect 18125 -8120 18180 -8000
rect 18300 -8120 18325 -8000
rect 12795 -8165 18325 -8120
rect 12795 -8285 12820 -8165
rect 12940 -8285 12985 -8165
rect 13105 -8285 13150 -8165
rect 13270 -8285 13315 -8165
rect 13435 -8285 13490 -8165
rect 13610 -8285 13655 -8165
rect 13775 -8285 13820 -8165
rect 13940 -8285 13985 -8165
rect 14105 -8285 14160 -8165
rect 14280 -8285 14325 -8165
rect 14445 -8285 14490 -8165
rect 14610 -8285 14655 -8165
rect 14775 -8285 14830 -8165
rect 14950 -8285 14995 -8165
rect 15115 -8285 15160 -8165
rect 15280 -8285 15325 -8165
rect 15445 -8285 15500 -8165
rect 15620 -8285 15665 -8165
rect 15785 -8285 15830 -8165
rect 15950 -8285 15995 -8165
rect 16115 -8285 16170 -8165
rect 16290 -8285 16335 -8165
rect 16455 -8285 16500 -8165
rect 16620 -8285 16665 -8165
rect 16785 -8285 16840 -8165
rect 16960 -8285 17005 -8165
rect 17125 -8285 17170 -8165
rect 17290 -8285 17335 -8165
rect 17455 -8285 17510 -8165
rect 17630 -8285 17675 -8165
rect 17795 -8285 17840 -8165
rect 17960 -8285 18005 -8165
rect 18125 -8285 18180 -8165
rect 18300 -8285 18325 -8165
rect 12795 -8330 18325 -8285
rect 12795 -8450 12820 -8330
rect 12940 -8450 12985 -8330
rect 13105 -8450 13150 -8330
rect 13270 -8450 13315 -8330
rect 13435 -8450 13490 -8330
rect 13610 -8450 13655 -8330
rect 13775 -8450 13820 -8330
rect 13940 -8450 13985 -8330
rect 14105 -8450 14160 -8330
rect 14280 -8450 14325 -8330
rect 14445 -8450 14490 -8330
rect 14610 -8450 14655 -8330
rect 14775 -8450 14830 -8330
rect 14950 -8450 14995 -8330
rect 15115 -8450 15160 -8330
rect 15280 -8450 15325 -8330
rect 15445 -8450 15500 -8330
rect 15620 -8450 15665 -8330
rect 15785 -8450 15830 -8330
rect 15950 -8450 15995 -8330
rect 16115 -8450 16170 -8330
rect 16290 -8450 16335 -8330
rect 16455 -8450 16500 -8330
rect 16620 -8450 16665 -8330
rect 16785 -8450 16840 -8330
rect 16960 -8450 17005 -8330
rect 17125 -8450 17170 -8330
rect 17290 -8450 17335 -8330
rect 17455 -8450 17510 -8330
rect 17630 -8450 17675 -8330
rect 17795 -8450 17840 -8330
rect 17960 -8450 18005 -8330
rect 18125 -8450 18180 -8330
rect 18300 -8450 18325 -8330
rect 12795 -8505 18325 -8450
rect 12795 -8625 12820 -8505
rect 12940 -8625 12985 -8505
rect 13105 -8625 13150 -8505
rect 13270 -8625 13315 -8505
rect 13435 -8625 13490 -8505
rect 13610 -8625 13655 -8505
rect 13775 -8625 13820 -8505
rect 13940 -8625 13985 -8505
rect 14105 -8625 14160 -8505
rect 14280 -8625 14325 -8505
rect 14445 -8625 14490 -8505
rect 14610 -8625 14655 -8505
rect 14775 -8625 14830 -8505
rect 14950 -8625 14995 -8505
rect 15115 -8625 15160 -8505
rect 15280 -8625 15325 -8505
rect 15445 -8625 15500 -8505
rect 15620 -8625 15665 -8505
rect 15785 -8625 15830 -8505
rect 15950 -8625 15995 -8505
rect 16115 -8625 16170 -8505
rect 16290 -8625 16335 -8505
rect 16455 -8625 16500 -8505
rect 16620 -8625 16665 -8505
rect 16785 -8625 16840 -8505
rect 16960 -8625 17005 -8505
rect 17125 -8625 17170 -8505
rect 17290 -8625 17335 -8505
rect 17455 -8625 17510 -8505
rect 17630 -8625 17675 -8505
rect 17795 -8625 17840 -8505
rect 17960 -8625 18005 -8505
rect 18125 -8625 18180 -8505
rect 18300 -8625 18325 -8505
rect 12795 -8670 18325 -8625
rect 12795 -8790 12820 -8670
rect 12940 -8790 12985 -8670
rect 13105 -8790 13150 -8670
rect 13270 -8790 13315 -8670
rect 13435 -8790 13490 -8670
rect 13610 -8790 13655 -8670
rect 13775 -8790 13820 -8670
rect 13940 -8790 13985 -8670
rect 14105 -8790 14160 -8670
rect 14280 -8790 14325 -8670
rect 14445 -8790 14490 -8670
rect 14610 -8790 14655 -8670
rect 14775 -8790 14830 -8670
rect 14950 -8790 14995 -8670
rect 15115 -8790 15160 -8670
rect 15280 -8790 15325 -8670
rect 15445 -8790 15500 -8670
rect 15620 -8790 15665 -8670
rect 15785 -8790 15830 -8670
rect 15950 -8790 15995 -8670
rect 16115 -8790 16170 -8670
rect 16290 -8790 16335 -8670
rect 16455 -8790 16500 -8670
rect 16620 -8790 16665 -8670
rect 16785 -8790 16840 -8670
rect 16960 -8790 17005 -8670
rect 17125 -8790 17170 -8670
rect 17290 -8790 17335 -8670
rect 17455 -8790 17510 -8670
rect 17630 -8790 17675 -8670
rect 17795 -8790 17840 -8670
rect 17960 -8790 18005 -8670
rect 18125 -8790 18180 -8670
rect 18300 -8790 18325 -8670
rect 12795 -8835 18325 -8790
rect 12795 -8955 12820 -8835
rect 12940 -8955 12985 -8835
rect 13105 -8955 13150 -8835
rect 13270 -8955 13315 -8835
rect 13435 -8955 13490 -8835
rect 13610 -8955 13655 -8835
rect 13775 -8955 13820 -8835
rect 13940 -8955 13985 -8835
rect 14105 -8955 14160 -8835
rect 14280 -8955 14325 -8835
rect 14445 -8955 14490 -8835
rect 14610 -8955 14655 -8835
rect 14775 -8955 14830 -8835
rect 14950 -8955 14995 -8835
rect 15115 -8955 15160 -8835
rect 15280 -8955 15325 -8835
rect 15445 -8955 15500 -8835
rect 15620 -8955 15665 -8835
rect 15785 -8955 15830 -8835
rect 15950 -8955 15995 -8835
rect 16115 -8955 16170 -8835
rect 16290 -8955 16335 -8835
rect 16455 -8955 16500 -8835
rect 16620 -8955 16665 -8835
rect 16785 -8955 16840 -8835
rect 16960 -8955 17005 -8835
rect 17125 -8955 17170 -8835
rect 17290 -8955 17335 -8835
rect 17455 -8955 17510 -8835
rect 17630 -8955 17675 -8835
rect 17795 -8955 17840 -8835
rect 17960 -8955 18005 -8835
rect 18125 -8955 18180 -8835
rect 18300 -8955 18325 -8835
rect 12795 -9000 18325 -8955
rect 12795 -9120 12820 -9000
rect 12940 -9120 12985 -9000
rect 13105 -9120 13150 -9000
rect 13270 -9120 13315 -9000
rect 13435 -9120 13490 -9000
rect 13610 -9120 13655 -9000
rect 13775 -9120 13820 -9000
rect 13940 -9120 13985 -9000
rect 14105 -9120 14160 -9000
rect 14280 -9120 14325 -9000
rect 14445 -9120 14490 -9000
rect 14610 -9120 14655 -9000
rect 14775 -9120 14830 -9000
rect 14950 -9120 14995 -9000
rect 15115 -9120 15160 -9000
rect 15280 -9120 15325 -9000
rect 15445 -9120 15500 -9000
rect 15620 -9120 15665 -9000
rect 15785 -9120 15830 -9000
rect 15950 -9120 15995 -9000
rect 16115 -9120 16170 -9000
rect 16290 -9120 16335 -9000
rect 16455 -9120 16500 -9000
rect 16620 -9120 16665 -9000
rect 16785 -9120 16840 -9000
rect 16960 -9120 17005 -9000
rect 17125 -9120 17170 -9000
rect 17290 -9120 17335 -9000
rect 17455 -9120 17510 -9000
rect 17630 -9120 17675 -9000
rect 17795 -9120 17840 -9000
rect 17960 -9120 18005 -9000
rect 18125 -9120 18180 -9000
rect 18300 -9120 18325 -9000
rect 12795 -9175 18325 -9120
rect 12795 -9295 12820 -9175
rect 12940 -9295 12985 -9175
rect 13105 -9295 13150 -9175
rect 13270 -9295 13315 -9175
rect 13435 -9295 13490 -9175
rect 13610 -9295 13655 -9175
rect 13775 -9295 13820 -9175
rect 13940 -9295 13985 -9175
rect 14105 -9295 14160 -9175
rect 14280 -9295 14325 -9175
rect 14445 -9295 14490 -9175
rect 14610 -9295 14655 -9175
rect 14775 -9295 14830 -9175
rect 14950 -9295 14995 -9175
rect 15115 -9295 15160 -9175
rect 15280 -9295 15325 -9175
rect 15445 -9295 15500 -9175
rect 15620 -9295 15665 -9175
rect 15785 -9295 15830 -9175
rect 15950 -9295 15995 -9175
rect 16115 -9295 16170 -9175
rect 16290 -9295 16335 -9175
rect 16455 -9295 16500 -9175
rect 16620 -9295 16665 -9175
rect 16785 -9295 16840 -9175
rect 16960 -9295 17005 -9175
rect 17125 -9295 17170 -9175
rect 17290 -9295 17335 -9175
rect 17455 -9295 17510 -9175
rect 17630 -9295 17675 -9175
rect 17795 -9295 17840 -9175
rect 17960 -9295 18005 -9175
rect 18125 -9295 18180 -9175
rect 18300 -9295 18325 -9175
rect 12795 -9340 18325 -9295
rect 12795 -9460 12820 -9340
rect 12940 -9460 12985 -9340
rect 13105 -9460 13150 -9340
rect 13270 -9460 13315 -9340
rect 13435 -9460 13490 -9340
rect 13610 -9460 13655 -9340
rect 13775 -9460 13820 -9340
rect 13940 -9460 13985 -9340
rect 14105 -9460 14160 -9340
rect 14280 -9460 14325 -9340
rect 14445 -9460 14490 -9340
rect 14610 -9460 14655 -9340
rect 14775 -9460 14830 -9340
rect 14950 -9460 14995 -9340
rect 15115 -9460 15160 -9340
rect 15280 -9460 15325 -9340
rect 15445 -9460 15500 -9340
rect 15620 -9460 15665 -9340
rect 15785 -9460 15830 -9340
rect 15950 -9460 15995 -9340
rect 16115 -9460 16170 -9340
rect 16290 -9460 16335 -9340
rect 16455 -9460 16500 -9340
rect 16620 -9460 16665 -9340
rect 16785 -9460 16840 -9340
rect 16960 -9460 17005 -9340
rect 17125 -9460 17170 -9340
rect 17290 -9460 17335 -9340
rect 17455 -9460 17510 -9340
rect 17630 -9460 17675 -9340
rect 17795 -9460 17840 -9340
rect 17960 -9460 18005 -9340
rect 18125 -9460 18180 -9340
rect 18300 -9460 18325 -9340
rect 12795 -9505 18325 -9460
rect 12795 -9625 12820 -9505
rect 12940 -9625 12985 -9505
rect 13105 -9625 13150 -9505
rect 13270 -9625 13315 -9505
rect 13435 -9625 13490 -9505
rect 13610 -9625 13655 -9505
rect 13775 -9625 13820 -9505
rect 13940 -9625 13985 -9505
rect 14105 -9625 14160 -9505
rect 14280 -9625 14325 -9505
rect 14445 -9625 14490 -9505
rect 14610 -9625 14655 -9505
rect 14775 -9625 14830 -9505
rect 14950 -9625 14995 -9505
rect 15115 -9625 15160 -9505
rect 15280 -9625 15325 -9505
rect 15445 -9625 15500 -9505
rect 15620 -9625 15665 -9505
rect 15785 -9625 15830 -9505
rect 15950 -9625 15995 -9505
rect 16115 -9625 16170 -9505
rect 16290 -9625 16335 -9505
rect 16455 -9625 16500 -9505
rect 16620 -9625 16665 -9505
rect 16785 -9625 16840 -9505
rect 16960 -9625 17005 -9505
rect 17125 -9625 17170 -9505
rect 17290 -9625 17335 -9505
rect 17455 -9625 17510 -9505
rect 17630 -9625 17675 -9505
rect 17795 -9625 17840 -9505
rect 17960 -9625 18005 -9505
rect 18125 -9625 18180 -9505
rect 18300 -9625 18325 -9505
rect 12795 -9670 18325 -9625
rect 12795 -9790 12820 -9670
rect 12940 -9790 12985 -9670
rect 13105 -9790 13150 -9670
rect 13270 -9790 13315 -9670
rect 13435 -9790 13490 -9670
rect 13610 -9790 13655 -9670
rect 13775 -9790 13820 -9670
rect 13940 -9790 13985 -9670
rect 14105 -9790 14160 -9670
rect 14280 -9790 14325 -9670
rect 14445 -9790 14490 -9670
rect 14610 -9790 14655 -9670
rect 14775 -9790 14830 -9670
rect 14950 -9790 14995 -9670
rect 15115 -9790 15160 -9670
rect 15280 -9790 15325 -9670
rect 15445 -9790 15500 -9670
rect 15620 -9790 15665 -9670
rect 15785 -9790 15830 -9670
rect 15950 -9790 15995 -9670
rect 16115 -9790 16170 -9670
rect 16290 -9790 16335 -9670
rect 16455 -9790 16500 -9670
rect 16620 -9790 16665 -9670
rect 16785 -9790 16840 -9670
rect 16960 -9790 17005 -9670
rect 17125 -9790 17170 -9670
rect 17290 -9790 17335 -9670
rect 17455 -9790 17510 -9670
rect 17630 -9790 17675 -9670
rect 17795 -9790 17840 -9670
rect 17960 -9790 18005 -9670
rect 18125 -9790 18180 -9670
rect 18300 -9790 18325 -9670
rect 12795 -9860 18325 -9790
rect 18485 -4310 24015 -4285
rect 18485 -4430 18510 -4310
rect 18630 -4430 18675 -4310
rect 18795 -4430 18840 -4310
rect 18960 -4430 19005 -4310
rect 19125 -4430 19180 -4310
rect 19300 -4430 19345 -4310
rect 19465 -4430 19510 -4310
rect 19630 -4430 19675 -4310
rect 19795 -4430 19850 -4310
rect 19970 -4430 20015 -4310
rect 20135 -4430 20180 -4310
rect 20300 -4430 20345 -4310
rect 20465 -4430 20520 -4310
rect 20640 -4430 20685 -4310
rect 20805 -4430 20850 -4310
rect 20970 -4430 21015 -4310
rect 21135 -4430 21190 -4310
rect 21310 -4430 21355 -4310
rect 21475 -4430 21520 -4310
rect 21640 -4430 21685 -4310
rect 21805 -4430 21860 -4310
rect 21980 -4430 22025 -4310
rect 22145 -4430 22190 -4310
rect 22310 -4430 22355 -4310
rect 22475 -4430 22530 -4310
rect 22650 -4430 22695 -4310
rect 22815 -4430 22860 -4310
rect 22980 -4430 23025 -4310
rect 23145 -4430 23200 -4310
rect 23320 -4430 23365 -4310
rect 23485 -4430 23530 -4310
rect 23650 -4430 23695 -4310
rect 23815 -4430 23870 -4310
rect 23990 -4430 24015 -4310
rect 18485 -4485 24015 -4430
rect 18485 -4605 18510 -4485
rect 18630 -4605 18675 -4485
rect 18795 -4605 18840 -4485
rect 18960 -4605 19005 -4485
rect 19125 -4605 19180 -4485
rect 19300 -4605 19345 -4485
rect 19465 -4605 19510 -4485
rect 19630 -4605 19675 -4485
rect 19795 -4605 19850 -4485
rect 19970 -4605 20015 -4485
rect 20135 -4605 20180 -4485
rect 20300 -4605 20345 -4485
rect 20465 -4605 20520 -4485
rect 20640 -4605 20685 -4485
rect 20805 -4605 20850 -4485
rect 20970 -4605 21015 -4485
rect 21135 -4605 21190 -4485
rect 21310 -4605 21355 -4485
rect 21475 -4605 21520 -4485
rect 21640 -4605 21685 -4485
rect 21805 -4605 21860 -4485
rect 21980 -4605 22025 -4485
rect 22145 -4605 22190 -4485
rect 22310 -4605 22355 -4485
rect 22475 -4605 22530 -4485
rect 22650 -4605 22695 -4485
rect 22815 -4605 22860 -4485
rect 22980 -4605 23025 -4485
rect 23145 -4605 23200 -4485
rect 23320 -4605 23365 -4485
rect 23485 -4605 23530 -4485
rect 23650 -4605 23695 -4485
rect 23815 -4605 23870 -4485
rect 23990 -4605 24015 -4485
rect 18485 -4650 24015 -4605
rect 18485 -4770 18510 -4650
rect 18630 -4770 18675 -4650
rect 18795 -4770 18840 -4650
rect 18960 -4770 19005 -4650
rect 19125 -4770 19180 -4650
rect 19300 -4770 19345 -4650
rect 19465 -4770 19510 -4650
rect 19630 -4770 19675 -4650
rect 19795 -4770 19850 -4650
rect 19970 -4770 20015 -4650
rect 20135 -4770 20180 -4650
rect 20300 -4770 20345 -4650
rect 20465 -4770 20520 -4650
rect 20640 -4770 20685 -4650
rect 20805 -4770 20850 -4650
rect 20970 -4770 21015 -4650
rect 21135 -4770 21190 -4650
rect 21310 -4770 21355 -4650
rect 21475 -4770 21520 -4650
rect 21640 -4770 21685 -4650
rect 21805 -4770 21860 -4650
rect 21980 -4770 22025 -4650
rect 22145 -4770 22190 -4650
rect 22310 -4770 22355 -4650
rect 22475 -4770 22530 -4650
rect 22650 -4770 22695 -4650
rect 22815 -4770 22860 -4650
rect 22980 -4770 23025 -4650
rect 23145 -4770 23200 -4650
rect 23320 -4770 23365 -4650
rect 23485 -4770 23530 -4650
rect 23650 -4770 23695 -4650
rect 23815 -4770 23870 -4650
rect 23990 -4770 24015 -4650
rect 18485 -4815 24015 -4770
rect 18485 -4935 18510 -4815
rect 18630 -4935 18675 -4815
rect 18795 -4935 18840 -4815
rect 18960 -4935 19005 -4815
rect 19125 -4935 19180 -4815
rect 19300 -4935 19345 -4815
rect 19465 -4935 19510 -4815
rect 19630 -4935 19675 -4815
rect 19795 -4935 19850 -4815
rect 19970 -4935 20015 -4815
rect 20135 -4935 20180 -4815
rect 20300 -4935 20345 -4815
rect 20465 -4935 20520 -4815
rect 20640 -4935 20685 -4815
rect 20805 -4935 20850 -4815
rect 20970 -4935 21015 -4815
rect 21135 -4935 21190 -4815
rect 21310 -4935 21355 -4815
rect 21475 -4935 21520 -4815
rect 21640 -4935 21685 -4815
rect 21805 -4935 21860 -4815
rect 21980 -4935 22025 -4815
rect 22145 -4935 22190 -4815
rect 22310 -4935 22355 -4815
rect 22475 -4935 22530 -4815
rect 22650 -4935 22695 -4815
rect 22815 -4935 22860 -4815
rect 22980 -4935 23025 -4815
rect 23145 -4935 23200 -4815
rect 23320 -4935 23365 -4815
rect 23485 -4935 23530 -4815
rect 23650 -4935 23695 -4815
rect 23815 -4935 23870 -4815
rect 23990 -4935 24015 -4815
rect 18485 -4980 24015 -4935
rect 18485 -5100 18510 -4980
rect 18630 -5100 18675 -4980
rect 18795 -5100 18840 -4980
rect 18960 -5100 19005 -4980
rect 19125 -5100 19180 -4980
rect 19300 -5100 19345 -4980
rect 19465 -5100 19510 -4980
rect 19630 -5100 19675 -4980
rect 19795 -5100 19850 -4980
rect 19970 -5100 20015 -4980
rect 20135 -5100 20180 -4980
rect 20300 -5100 20345 -4980
rect 20465 -5100 20520 -4980
rect 20640 -5100 20685 -4980
rect 20805 -5100 20850 -4980
rect 20970 -5100 21015 -4980
rect 21135 -5100 21190 -4980
rect 21310 -5100 21355 -4980
rect 21475 -5100 21520 -4980
rect 21640 -5100 21685 -4980
rect 21805 -5100 21860 -4980
rect 21980 -5100 22025 -4980
rect 22145 -5100 22190 -4980
rect 22310 -5100 22355 -4980
rect 22475 -5100 22530 -4980
rect 22650 -5100 22695 -4980
rect 22815 -5100 22860 -4980
rect 22980 -5100 23025 -4980
rect 23145 -5100 23200 -4980
rect 23320 -5100 23365 -4980
rect 23485 -5100 23530 -4980
rect 23650 -5100 23695 -4980
rect 23815 -5100 23870 -4980
rect 23990 -5100 24015 -4980
rect 18485 -5155 24015 -5100
rect 18485 -5275 18510 -5155
rect 18630 -5275 18675 -5155
rect 18795 -5275 18840 -5155
rect 18960 -5275 19005 -5155
rect 19125 -5275 19180 -5155
rect 19300 -5275 19345 -5155
rect 19465 -5275 19510 -5155
rect 19630 -5275 19675 -5155
rect 19795 -5275 19850 -5155
rect 19970 -5275 20015 -5155
rect 20135 -5275 20180 -5155
rect 20300 -5275 20345 -5155
rect 20465 -5275 20520 -5155
rect 20640 -5275 20685 -5155
rect 20805 -5275 20850 -5155
rect 20970 -5275 21015 -5155
rect 21135 -5275 21190 -5155
rect 21310 -5275 21355 -5155
rect 21475 -5275 21520 -5155
rect 21640 -5275 21685 -5155
rect 21805 -5275 21860 -5155
rect 21980 -5275 22025 -5155
rect 22145 -5275 22190 -5155
rect 22310 -5275 22355 -5155
rect 22475 -5275 22530 -5155
rect 22650 -5275 22695 -5155
rect 22815 -5275 22860 -5155
rect 22980 -5275 23025 -5155
rect 23145 -5275 23200 -5155
rect 23320 -5275 23365 -5155
rect 23485 -5275 23530 -5155
rect 23650 -5275 23695 -5155
rect 23815 -5275 23870 -5155
rect 23990 -5275 24015 -5155
rect 18485 -5320 24015 -5275
rect 18485 -5440 18510 -5320
rect 18630 -5440 18675 -5320
rect 18795 -5440 18840 -5320
rect 18960 -5440 19005 -5320
rect 19125 -5440 19180 -5320
rect 19300 -5440 19345 -5320
rect 19465 -5440 19510 -5320
rect 19630 -5440 19675 -5320
rect 19795 -5440 19850 -5320
rect 19970 -5440 20015 -5320
rect 20135 -5440 20180 -5320
rect 20300 -5440 20345 -5320
rect 20465 -5440 20520 -5320
rect 20640 -5440 20685 -5320
rect 20805 -5440 20850 -5320
rect 20970 -5440 21015 -5320
rect 21135 -5440 21190 -5320
rect 21310 -5440 21355 -5320
rect 21475 -5440 21520 -5320
rect 21640 -5440 21685 -5320
rect 21805 -5440 21860 -5320
rect 21980 -5440 22025 -5320
rect 22145 -5440 22190 -5320
rect 22310 -5440 22355 -5320
rect 22475 -5440 22530 -5320
rect 22650 -5440 22695 -5320
rect 22815 -5440 22860 -5320
rect 22980 -5440 23025 -5320
rect 23145 -5440 23200 -5320
rect 23320 -5440 23365 -5320
rect 23485 -5440 23530 -5320
rect 23650 -5440 23695 -5320
rect 23815 -5440 23870 -5320
rect 23990 -5440 24015 -5320
rect 18485 -5485 24015 -5440
rect 18485 -5605 18510 -5485
rect 18630 -5605 18675 -5485
rect 18795 -5605 18840 -5485
rect 18960 -5605 19005 -5485
rect 19125 -5605 19180 -5485
rect 19300 -5605 19345 -5485
rect 19465 -5605 19510 -5485
rect 19630 -5605 19675 -5485
rect 19795 -5605 19850 -5485
rect 19970 -5605 20015 -5485
rect 20135 -5605 20180 -5485
rect 20300 -5605 20345 -5485
rect 20465 -5605 20520 -5485
rect 20640 -5605 20685 -5485
rect 20805 -5605 20850 -5485
rect 20970 -5605 21015 -5485
rect 21135 -5605 21190 -5485
rect 21310 -5605 21355 -5485
rect 21475 -5605 21520 -5485
rect 21640 -5605 21685 -5485
rect 21805 -5605 21860 -5485
rect 21980 -5605 22025 -5485
rect 22145 -5605 22190 -5485
rect 22310 -5605 22355 -5485
rect 22475 -5605 22530 -5485
rect 22650 -5605 22695 -5485
rect 22815 -5605 22860 -5485
rect 22980 -5605 23025 -5485
rect 23145 -5605 23200 -5485
rect 23320 -5605 23365 -5485
rect 23485 -5605 23530 -5485
rect 23650 -5605 23695 -5485
rect 23815 -5605 23870 -5485
rect 23990 -5605 24015 -5485
rect 18485 -5650 24015 -5605
rect 18485 -5770 18510 -5650
rect 18630 -5770 18675 -5650
rect 18795 -5770 18840 -5650
rect 18960 -5770 19005 -5650
rect 19125 -5770 19180 -5650
rect 19300 -5770 19345 -5650
rect 19465 -5770 19510 -5650
rect 19630 -5770 19675 -5650
rect 19795 -5770 19850 -5650
rect 19970 -5770 20015 -5650
rect 20135 -5770 20180 -5650
rect 20300 -5770 20345 -5650
rect 20465 -5770 20520 -5650
rect 20640 -5770 20685 -5650
rect 20805 -5770 20850 -5650
rect 20970 -5770 21015 -5650
rect 21135 -5770 21190 -5650
rect 21310 -5770 21355 -5650
rect 21475 -5770 21520 -5650
rect 21640 -5770 21685 -5650
rect 21805 -5770 21860 -5650
rect 21980 -5770 22025 -5650
rect 22145 -5770 22190 -5650
rect 22310 -5770 22355 -5650
rect 22475 -5770 22530 -5650
rect 22650 -5770 22695 -5650
rect 22815 -5770 22860 -5650
rect 22980 -5770 23025 -5650
rect 23145 -5770 23200 -5650
rect 23320 -5770 23365 -5650
rect 23485 -5770 23530 -5650
rect 23650 -5770 23695 -5650
rect 23815 -5770 23870 -5650
rect 23990 -5770 24015 -5650
rect 18485 -5825 24015 -5770
rect 18485 -5945 18510 -5825
rect 18630 -5945 18675 -5825
rect 18795 -5945 18840 -5825
rect 18960 -5945 19005 -5825
rect 19125 -5945 19180 -5825
rect 19300 -5945 19345 -5825
rect 19465 -5945 19510 -5825
rect 19630 -5945 19675 -5825
rect 19795 -5945 19850 -5825
rect 19970 -5945 20015 -5825
rect 20135 -5945 20180 -5825
rect 20300 -5945 20345 -5825
rect 20465 -5945 20520 -5825
rect 20640 -5945 20685 -5825
rect 20805 -5945 20850 -5825
rect 20970 -5945 21015 -5825
rect 21135 -5945 21190 -5825
rect 21310 -5945 21355 -5825
rect 21475 -5945 21520 -5825
rect 21640 -5945 21685 -5825
rect 21805 -5945 21860 -5825
rect 21980 -5945 22025 -5825
rect 22145 -5945 22190 -5825
rect 22310 -5945 22355 -5825
rect 22475 -5945 22530 -5825
rect 22650 -5945 22695 -5825
rect 22815 -5945 22860 -5825
rect 22980 -5945 23025 -5825
rect 23145 -5945 23200 -5825
rect 23320 -5945 23365 -5825
rect 23485 -5945 23530 -5825
rect 23650 -5945 23695 -5825
rect 23815 -5945 23870 -5825
rect 23990 -5945 24015 -5825
rect 18485 -5990 24015 -5945
rect 18485 -6110 18510 -5990
rect 18630 -6110 18675 -5990
rect 18795 -6110 18840 -5990
rect 18960 -6110 19005 -5990
rect 19125 -6110 19180 -5990
rect 19300 -6110 19345 -5990
rect 19465 -6110 19510 -5990
rect 19630 -6110 19675 -5990
rect 19795 -6110 19850 -5990
rect 19970 -6110 20015 -5990
rect 20135 -6110 20180 -5990
rect 20300 -6110 20345 -5990
rect 20465 -6110 20520 -5990
rect 20640 -6110 20685 -5990
rect 20805 -6110 20850 -5990
rect 20970 -6110 21015 -5990
rect 21135 -6110 21190 -5990
rect 21310 -6110 21355 -5990
rect 21475 -6110 21520 -5990
rect 21640 -6110 21685 -5990
rect 21805 -6110 21860 -5990
rect 21980 -6110 22025 -5990
rect 22145 -6110 22190 -5990
rect 22310 -6110 22355 -5990
rect 22475 -6110 22530 -5990
rect 22650 -6110 22695 -5990
rect 22815 -6110 22860 -5990
rect 22980 -6110 23025 -5990
rect 23145 -6110 23200 -5990
rect 23320 -6110 23365 -5990
rect 23485 -6110 23530 -5990
rect 23650 -6110 23695 -5990
rect 23815 -6110 23870 -5990
rect 23990 -6110 24015 -5990
rect 18485 -6155 24015 -6110
rect 18485 -6275 18510 -6155
rect 18630 -6275 18675 -6155
rect 18795 -6275 18840 -6155
rect 18960 -6275 19005 -6155
rect 19125 -6275 19180 -6155
rect 19300 -6275 19345 -6155
rect 19465 -6275 19510 -6155
rect 19630 -6275 19675 -6155
rect 19795 -6275 19850 -6155
rect 19970 -6275 20015 -6155
rect 20135 -6275 20180 -6155
rect 20300 -6275 20345 -6155
rect 20465 -6275 20520 -6155
rect 20640 -6275 20685 -6155
rect 20805 -6275 20850 -6155
rect 20970 -6275 21015 -6155
rect 21135 -6275 21190 -6155
rect 21310 -6275 21355 -6155
rect 21475 -6275 21520 -6155
rect 21640 -6275 21685 -6155
rect 21805 -6275 21860 -6155
rect 21980 -6275 22025 -6155
rect 22145 -6275 22190 -6155
rect 22310 -6275 22355 -6155
rect 22475 -6275 22530 -6155
rect 22650 -6275 22695 -6155
rect 22815 -6275 22860 -6155
rect 22980 -6275 23025 -6155
rect 23145 -6275 23200 -6155
rect 23320 -6275 23365 -6155
rect 23485 -6275 23530 -6155
rect 23650 -6275 23695 -6155
rect 23815 -6275 23870 -6155
rect 23990 -6275 24015 -6155
rect 18485 -6320 24015 -6275
rect 18485 -6440 18510 -6320
rect 18630 -6440 18675 -6320
rect 18795 -6440 18840 -6320
rect 18960 -6440 19005 -6320
rect 19125 -6440 19180 -6320
rect 19300 -6440 19345 -6320
rect 19465 -6440 19510 -6320
rect 19630 -6440 19675 -6320
rect 19795 -6440 19850 -6320
rect 19970 -6440 20015 -6320
rect 20135 -6440 20180 -6320
rect 20300 -6440 20345 -6320
rect 20465 -6440 20520 -6320
rect 20640 -6440 20685 -6320
rect 20805 -6440 20850 -6320
rect 20970 -6440 21015 -6320
rect 21135 -6440 21190 -6320
rect 21310 -6440 21355 -6320
rect 21475 -6440 21520 -6320
rect 21640 -6440 21685 -6320
rect 21805 -6440 21860 -6320
rect 21980 -6440 22025 -6320
rect 22145 -6440 22190 -6320
rect 22310 -6440 22355 -6320
rect 22475 -6440 22530 -6320
rect 22650 -6440 22695 -6320
rect 22815 -6440 22860 -6320
rect 22980 -6440 23025 -6320
rect 23145 -6440 23200 -6320
rect 23320 -6440 23365 -6320
rect 23485 -6440 23530 -6320
rect 23650 -6440 23695 -6320
rect 23815 -6440 23870 -6320
rect 23990 -6440 24015 -6320
rect 18485 -6495 24015 -6440
rect 18485 -6615 18510 -6495
rect 18630 -6615 18675 -6495
rect 18795 -6615 18840 -6495
rect 18960 -6615 19005 -6495
rect 19125 -6615 19180 -6495
rect 19300 -6615 19345 -6495
rect 19465 -6615 19510 -6495
rect 19630 -6615 19675 -6495
rect 19795 -6615 19850 -6495
rect 19970 -6615 20015 -6495
rect 20135 -6615 20180 -6495
rect 20300 -6615 20345 -6495
rect 20465 -6615 20520 -6495
rect 20640 -6615 20685 -6495
rect 20805 -6615 20850 -6495
rect 20970 -6615 21015 -6495
rect 21135 -6615 21190 -6495
rect 21310 -6615 21355 -6495
rect 21475 -6615 21520 -6495
rect 21640 -6615 21685 -6495
rect 21805 -6615 21860 -6495
rect 21980 -6615 22025 -6495
rect 22145 -6615 22190 -6495
rect 22310 -6615 22355 -6495
rect 22475 -6615 22530 -6495
rect 22650 -6615 22695 -6495
rect 22815 -6615 22860 -6495
rect 22980 -6615 23025 -6495
rect 23145 -6615 23200 -6495
rect 23320 -6615 23365 -6495
rect 23485 -6615 23530 -6495
rect 23650 -6615 23695 -6495
rect 23815 -6615 23870 -6495
rect 23990 -6615 24015 -6495
rect 18485 -6660 24015 -6615
rect 18485 -6780 18510 -6660
rect 18630 -6780 18675 -6660
rect 18795 -6780 18840 -6660
rect 18960 -6780 19005 -6660
rect 19125 -6780 19180 -6660
rect 19300 -6780 19345 -6660
rect 19465 -6780 19510 -6660
rect 19630 -6780 19675 -6660
rect 19795 -6780 19850 -6660
rect 19970 -6780 20015 -6660
rect 20135 -6780 20180 -6660
rect 20300 -6780 20345 -6660
rect 20465 -6780 20520 -6660
rect 20640 -6780 20685 -6660
rect 20805 -6780 20850 -6660
rect 20970 -6780 21015 -6660
rect 21135 -6780 21190 -6660
rect 21310 -6780 21355 -6660
rect 21475 -6780 21520 -6660
rect 21640 -6780 21685 -6660
rect 21805 -6780 21860 -6660
rect 21980 -6780 22025 -6660
rect 22145 -6780 22190 -6660
rect 22310 -6780 22355 -6660
rect 22475 -6780 22530 -6660
rect 22650 -6780 22695 -6660
rect 22815 -6780 22860 -6660
rect 22980 -6780 23025 -6660
rect 23145 -6780 23200 -6660
rect 23320 -6780 23365 -6660
rect 23485 -6780 23530 -6660
rect 23650 -6780 23695 -6660
rect 23815 -6780 23870 -6660
rect 23990 -6780 24015 -6660
rect 18485 -6825 24015 -6780
rect 18485 -6945 18510 -6825
rect 18630 -6945 18675 -6825
rect 18795 -6945 18840 -6825
rect 18960 -6945 19005 -6825
rect 19125 -6945 19180 -6825
rect 19300 -6945 19345 -6825
rect 19465 -6945 19510 -6825
rect 19630 -6945 19675 -6825
rect 19795 -6945 19850 -6825
rect 19970 -6945 20015 -6825
rect 20135 -6945 20180 -6825
rect 20300 -6945 20345 -6825
rect 20465 -6945 20520 -6825
rect 20640 -6945 20685 -6825
rect 20805 -6945 20850 -6825
rect 20970 -6945 21015 -6825
rect 21135 -6945 21190 -6825
rect 21310 -6945 21355 -6825
rect 21475 -6945 21520 -6825
rect 21640 -6945 21685 -6825
rect 21805 -6945 21860 -6825
rect 21980 -6945 22025 -6825
rect 22145 -6945 22190 -6825
rect 22310 -6945 22355 -6825
rect 22475 -6945 22530 -6825
rect 22650 -6945 22695 -6825
rect 22815 -6945 22860 -6825
rect 22980 -6945 23025 -6825
rect 23145 -6945 23200 -6825
rect 23320 -6945 23365 -6825
rect 23485 -6945 23530 -6825
rect 23650 -6945 23695 -6825
rect 23815 -6945 23870 -6825
rect 23990 -6945 24015 -6825
rect 18485 -6990 24015 -6945
rect 18485 -7110 18510 -6990
rect 18630 -7110 18675 -6990
rect 18795 -7110 18840 -6990
rect 18960 -7110 19005 -6990
rect 19125 -7110 19180 -6990
rect 19300 -7110 19345 -6990
rect 19465 -7110 19510 -6990
rect 19630 -7110 19675 -6990
rect 19795 -7110 19850 -6990
rect 19970 -7110 20015 -6990
rect 20135 -7110 20180 -6990
rect 20300 -7110 20345 -6990
rect 20465 -7110 20520 -6990
rect 20640 -7110 20685 -6990
rect 20805 -7110 20850 -6990
rect 20970 -7110 21015 -6990
rect 21135 -7110 21190 -6990
rect 21310 -7110 21355 -6990
rect 21475 -7110 21520 -6990
rect 21640 -7110 21685 -6990
rect 21805 -7110 21860 -6990
rect 21980 -7110 22025 -6990
rect 22145 -7110 22190 -6990
rect 22310 -7110 22355 -6990
rect 22475 -7110 22530 -6990
rect 22650 -7110 22695 -6990
rect 22815 -7110 22860 -6990
rect 22980 -7110 23025 -6990
rect 23145 -7110 23200 -6990
rect 23320 -7110 23365 -6990
rect 23485 -7110 23530 -6990
rect 23650 -7110 23695 -6990
rect 23815 -7110 23870 -6990
rect 23990 -7110 24015 -6990
rect 18485 -7165 24015 -7110
rect 18485 -7285 18510 -7165
rect 18630 -7285 18675 -7165
rect 18795 -7285 18840 -7165
rect 18960 -7285 19005 -7165
rect 19125 -7285 19180 -7165
rect 19300 -7285 19345 -7165
rect 19465 -7285 19510 -7165
rect 19630 -7285 19675 -7165
rect 19795 -7285 19850 -7165
rect 19970 -7285 20015 -7165
rect 20135 -7285 20180 -7165
rect 20300 -7285 20345 -7165
rect 20465 -7285 20520 -7165
rect 20640 -7285 20685 -7165
rect 20805 -7285 20850 -7165
rect 20970 -7285 21015 -7165
rect 21135 -7285 21190 -7165
rect 21310 -7285 21355 -7165
rect 21475 -7285 21520 -7165
rect 21640 -7285 21685 -7165
rect 21805 -7285 21860 -7165
rect 21980 -7285 22025 -7165
rect 22145 -7285 22190 -7165
rect 22310 -7285 22355 -7165
rect 22475 -7285 22530 -7165
rect 22650 -7285 22695 -7165
rect 22815 -7285 22860 -7165
rect 22980 -7285 23025 -7165
rect 23145 -7285 23200 -7165
rect 23320 -7285 23365 -7165
rect 23485 -7285 23530 -7165
rect 23650 -7285 23695 -7165
rect 23815 -7285 23870 -7165
rect 23990 -7285 24015 -7165
rect 18485 -7330 24015 -7285
rect 18485 -7450 18510 -7330
rect 18630 -7450 18675 -7330
rect 18795 -7450 18840 -7330
rect 18960 -7450 19005 -7330
rect 19125 -7450 19180 -7330
rect 19300 -7450 19345 -7330
rect 19465 -7450 19510 -7330
rect 19630 -7450 19675 -7330
rect 19795 -7450 19850 -7330
rect 19970 -7450 20015 -7330
rect 20135 -7450 20180 -7330
rect 20300 -7450 20345 -7330
rect 20465 -7450 20520 -7330
rect 20640 -7450 20685 -7330
rect 20805 -7450 20850 -7330
rect 20970 -7450 21015 -7330
rect 21135 -7450 21190 -7330
rect 21310 -7450 21355 -7330
rect 21475 -7450 21520 -7330
rect 21640 -7450 21685 -7330
rect 21805 -7450 21860 -7330
rect 21980 -7450 22025 -7330
rect 22145 -7450 22190 -7330
rect 22310 -7450 22355 -7330
rect 22475 -7450 22530 -7330
rect 22650 -7450 22695 -7330
rect 22815 -7450 22860 -7330
rect 22980 -7450 23025 -7330
rect 23145 -7450 23200 -7330
rect 23320 -7450 23365 -7330
rect 23485 -7450 23530 -7330
rect 23650 -7450 23695 -7330
rect 23815 -7450 23870 -7330
rect 23990 -7450 24015 -7330
rect 18485 -7495 24015 -7450
rect 18485 -7615 18510 -7495
rect 18630 -7615 18675 -7495
rect 18795 -7615 18840 -7495
rect 18960 -7615 19005 -7495
rect 19125 -7615 19180 -7495
rect 19300 -7615 19345 -7495
rect 19465 -7615 19510 -7495
rect 19630 -7615 19675 -7495
rect 19795 -7615 19850 -7495
rect 19970 -7615 20015 -7495
rect 20135 -7615 20180 -7495
rect 20300 -7615 20345 -7495
rect 20465 -7615 20520 -7495
rect 20640 -7615 20685 -7495
rect 20805 -7615 20850 -7495
rect 20970 -7615 21015 -7495
rect 21135 -7615 21190 -7495
rect 21310 -7615 21355 -7495
rect 21475 -7615 21520 -7495
rect 21640 -7615 21685 -7495
rect 21805 -7615 21860 -7495
rect 21980 -7615 22025 -7495
rect 22145 -7615 22190 -7495
rect 22310 -7615 22355 -7495
rect 22475 -7615 22530 -7495
rect 22650 -7615 22695 -7495
rect 22815 -7615 22860 -7495
rect 22980 -7615 23025 -7495
rect 23145 -7615 23200 -7495
rect 23320 -7615 23365 -7495
rect 23485 -7615 23530 -7495
rect 23650 -7615 23695 -7495
rect 23815 -7615 23870 -7495
rect 23990 -7615 24015 -7495
rect 18485 -7660 24015 -7615
rect 18485 -7780 18510 -7660
rect 18630 -7780 18675 -7660
rect 18795 -7780 18840 -7660
rect 18960 -7780 19005 -7660
rect 19125 -7780 19180 -7660
rect 19300 -7780 19345 -7660
rect 19465 -7780 19510 -7660
rect 19630 -7780 19675 -7660
rect 19795 -7780 19850 -7660
rect 19970 -7780 20015 -7660
rect 20135 -7780 20180 -7660
rect 20300 -7780 20345 -7660
rect 20465 -7780 20520 -7660
rect 20640 -7780 20685 -7660
rect 20805 -7780 20850 -7660
rect 20970 -7780 21015 -7660
rect 21135 -7780 21190 -7660
rect 21310 -7780 21355 -7660
rect 21475 -7780 21520 -7660
rect 21640 -7780 21685 -7660
rect 21805 -7780 21860 -7660
rect 21980 -7780 22025 -7660
rect 22145 -7780 22190 -7660
rect 22310 -7780 22355 -7660
rect 22475 -7780 22530 -7660
rect 22650 -7780 22695 -7660
rect 22815 -7780 22860 -7660
rect 22980 -7780 23025 -7660
rect 23145 -7780 23200 -7660
rect 23320 -7780 23365 -7660
rect 23485 -7780 23530 -7660
rect 23650 -7780 23695 -7660
rect 23815 -7780 23870 -7660
rect 23990 -7780 24015 -7660
rect 18485 -7835 24015 -7780
rect 18485 -7955 18510 -7835
rect 18630 -7955 18675 -7835
rect 18795 -7955 18840 -7835
rect 18960 -7955 19005 -7835
rect 19125 -7955 19180 -7835
rect 19300 -7955 19345 -7835
rect 19465 -7955 19510 -7835
rect 19630 -7955 19675 -7835
rect 19795 -7955 19850 -7835
rect 19970 -7955 20015 -7835
rect 20135 -7955 20180 -7835
rect 20300 -7955 20345 -7835
rect 20465 -7955 20520 -7835
rect 20640 -7955 20685 -7835
rect 20805 -7955 20850 -7835
rect 20970 -7955 21015 -7835
rect 21135 -7955 21190 -7835
rect 21310 -7955 21355 -7835
rect 21475 -7955 21520 -7835
rect 21640 -7955 21685 -7835
rect 21805 -7955 21860 -7835
rect 21980 -7955 22025 -7835
rect 22145 -7955 22190 -7835
rect 22310 -7955 22355 -7835
rect 22475 -7955 22530 -7835
rect 22650 -7955 22695 -7835
rect 22815 -7955 22860 -7835
rect 22980 -7955 23025 -7835
rect 23145 -7955 23200 -7835
rect 23320 -7955 23365 -7835
rect 23485 -7955 23530 -7835
rect 23650 -7955 23695 -7835
rect 23815 -7955 23870 -7835
rect 23990 -7955 24015 -7835
rect 18485 -8000 24015 -7955
rect 18485 -8120 18510 -8000
rect 18630 -8120 18675 -8000
rect 18795 -8120 18840 -8000
rect 18960 -8120 19005 -8000
rect 19125 -8120 19180 -8000
rect 19300 -8120 19345 -8000
rect 19465 -8120 19510 -8000
rect 19630 -8120 19675 -8000
rect 19795 -8120 19850 -8000
rect 19970 -8120 20015 -8000
rect 20135 -8120 20180 -8000
rect 20300 -8120 20345 -8000
rect 20465 -8120 20520 -8000
rect 20640 -8120 20685 -8000
rect 20805 -8120 20850 -8000
rect 20970 -8120 21015 -8000
rect 21135 -8120 21190 -8000
rect 21310 -8120 21355 -8000
rect 21475 -8120 21520 -8000
rect 21640 -8120 21685 -8000
rect 21805 -8120 21860 -8000
rect 21980 -8120 22025 -8000
rect 22145 -8120 22190 -8000
rect 22310 -8120 22355 -8000
rect 22475 -8120 22530 -8000
rect 22650 -8120 22695 -8000
rect 22815 -8120 22860 -8000
rect 22980 -8120 23025 -8000
rect 23145 -8120 23200 -8000
rect 23320 -8120 23365 -8000
rect 23485 -8120 23530 -8000
rect 23650 -8120 23695 -8000
rect 23815 -8120 23870 -8000
rect 23990 -8120 24015 -8000
rect 18485 -8165 24015 -8120
rect 18485 -8285 18510 -8165
rect 18630 -8285 18675 -8165
rect 18795 -8285 18840 -8165
rect 18960 -8285 19005 -8165
rect 19125 -8285 19180 -8165
rect 19300 -8285 19345 -8165
rect 19465 -8285 19510 -8165
rect 19630 -8285 19675 -8165
rect 19795 -8285 19850 -8165
rect 19970 -8285 20015 -8165
rect 20135 -8285 20180 -8165
rect 20300 -8285 20345 -8165
rect 20465 -8285 20520 -8165
rect 20640 -8285 20685 -8165
rect 20805 -8285 20850 -8165
rect 20970 -8285 21015 -8165
rect 21135 -8285 21190 -8165
rect 21310 -8285 21355 -8165
rect 21475 -8285 21520 -8165
rect 21640 -8285 21685 -8165
rect 21805 -8285 21860 -8165
rect 21980 -8285 22025 -8165
rect 22145 -8285 22190 -8165
rect 22310 -8285 22355 -8165
rect 22475 -8285 22530 -8165
rect 22650 -8285 22695 -8165
rect 22815 -8285 22860 -8165
rect 22980 -8285 23025 -8165
rect 23145 -8285 23200 -8165
rect 23320 -8285 23365 -8165
rect 23485 -8285 23530 -8165
rect 23650 -8285 23695 -8165
rect 23815 -8285 23870 -8165
rect 23990 -8285 24015 -8165
rect 18485 -8330 24015 -8285
rect 18485 -8450 18510 -8330
rect 18630 -8450 18675 -8330
rect 18795 -8450 18840 -8330
rect 18960 -8450 19005 -8330
rect 19125 -8450 19180 -8330
rect 19300 -8450 19345 -8330
rect 19465 -8450 19510 -8330
rect 19630 -8450 19675 -8330
rect 19795 -8450 19850 -8330
rect 19970 -8450 20015 -8330
rect 20135 -8450 20180 -8330
rect 20300 -8450 20345 -8330
rect 20465 -8450 20520 -8330
rect 20640 -8450 20685 -8330
rect 20805 -8450 20850 -8330
rect 20970 -8450 21015 -8330
rect 21135 -8450 21190 -8330
rect 21310 -8450 21355 -8330
rect 21475 -8450 21520 -8330
rect 21640 -8450 21685 -8330
rect 21805 -8450 21860 -8330
rect 21980 -8450 22025 -8330
rect 22145 -8450 22190 -8330
rect 22310 -8450 22355 -8330
rect 22475 -8450 22530 -8330
rect 22650 -8450 22695 -8330
rect 22815 -8450 22860 -8330
rect 22980 -8450 23025 -8330
rect 23145 -8450 23200 -8330
rect 23320 -8450 23365 -8330
rect 23485 -8450 23530 -8330
rect 23650 -8450 23695 -8330
rect 23815 -8450 23870 -8330
rect 23990 -8450 24015 -8330
rect 18485 -8505 24015 -8450
rect 18485 -8625 18510 -8505
rect 18630 -8625 18675 -8505
rect 18795 -8625 18840 -8505
rect 18960 -8625 19005 -8505
rect 19125 -8625 19180 -8505
rect 19300 -8625 19345 -8505
rect 19465 -8625 19510 -8505
rect 19630 -8625 19675 -8505
rect 19795 -8625 19850 -8505
rect 19970 -8625 20015 -8505
rect 20135 -8625 20180 -8505
rect 20300 -8625 20345 -8505
rect 20465 -8625 20520 -8505
rect 20640 -8625 20685 -8505
rect 20805 -8625 20850 -8505
rect 20970 -8625 21015 -8505
rect 21135 -8625 21190 -8505
rect 21310 -8625 21355 -8505
rect 21475 -8625 21520 -8505
rect 21640 -8625 21685 -8505
rect 21805 -8625 21860 -8505
rect 21980 -8625 22025 -8505
rect 22145 -8625 22190 -8505
rect 22310 -8625 22355 -8505
rect 22475 -8625 22530 -8505
rect 22650 -8625 22695 -8505
rect 22815 -8625 22860 -8505
rect 22980 -8625 23025 -8505
rect 23145 -8625 23200 -8505
rect 23320 -8625 23365 -8505
rect 23485 -8625 23530 -8505
rect 23650 -8625 23695 -8505
rect 23815 -8625 23870 -8505
rect 23990 -8625 24015 -8505
rect 18485 -8670 24015 -8625
rect 18485 -8790 18510 -8670
rect 18630 -8790 18675 -8670
rect 18795 -8790 18840 -8670
rect 18960 -8790 19005 -8670
rect 19125 -8790 19180 -8670
rect 19300 -8790 19345 -8670
rect 19465 -8790 19510 -8670
rect 19630 -8790 19675 -8670
rect 19795 -8790 19850 -8670
rect 19970 -8790 20015 -8670
rect 20135 -8790 20180 -8670
rect 20300 -8790 20345 -8670
rect 20465 -8790 20520 -8670
rect 20640 -8790 20685 -8670
rect 20805 -8790 20850 -8670
rect 20970 -8790 21015 -8670
rect 21135 -8790 21190 -8670
rect 21310 -8790 21355 -8670
rect 21475 -8790 21520 -8670
rect 21640 -8790 21685 -8670
rect 21805 -8790 21860 -8670
rect 21980 -8790 22025 -8670
rect 22145 -8790 22190 -8670
rect 22310 -8790 22355 -8670
rect 22475 -8790 22530 -8670
rect 22650 -8790 22695 -8670
rect 22815 -8790 22860 -8670
rect 22980 -8790 23025 -8670
rect 23145 -8790 23200 -8670
rect 23320 -8790 23365 -8670
rect 23485 -8790 23530 -8670
rect 23650 -8790 23695 -8670
rect 23815 -8790 23870 -8670
rect 23990 -8790 24015 -8670
rect 18485 -8835 24015 -8790
rect 18485 -8955 18510 -8835
rect 18630 -8955 18675 -8835
rect 18795 -8955 18840 -8835
rect 18960 -8955 19005 -8835
rect 19125 -8955 19180 -8835
rect 19300 -8955 19345 -8835
rect 19465 -8955 19510 -8835
rect 19630 -8955 19675 -8835
rect 19795 -8955 19850 -8835
rect 19970 -8955 20015 -8835
rect 20135 -8955 20180 -8835
rect 20300 -8955 20345 -8835
rect 20465 -8955 20520 -8835
rect 20640 -8955 20685 -8835
rect 20805 -8955 20850 -8835
rect 20970 -8955 21015 -8835
rect 21135 -8955 21190 -8835
rect 21310 -8955 21355 -8835
rect 21475 -8955 21520 -8835
rect 21640 -8955 21685 -8835
rect 21805 -8955 21860 -8835
rect 21980 -8955 22025 -8835
rect 22145 -8955 22190 -8835
rect 22310 -8955 22355 -8835
rect 22475 -8955 22530 -8835
rect 22650 -8955 22695 -8835
rect 22815 -8955 22860 -8835
rect 22980 -8955 23025 -8835
rect 23145 -8955 23200 -8835
rect 23320 -8955 23365 -8835
rect 23485 -8955 23530 -8835
rect 23650 -8955 23695 -8835
rect 23815 -8955 23870 -8835
rect 23990 -8955 24015 -8835
rect 18485 -9000 24015 -8955
rect 18485 -9120 18510 -9000
rect 18630 -9120 18675 -9000
rect 18795 -9120 18840 -9000
rect 18960 -9120 19005 -9000
rect 19125 -9120 19180 -9000
rect 19300 -9120 19345 -9000
rect 19465 -9120 19510 -9000
rect 19630 -9120 19675 -9000
rect 19795 -9120 19850 -9000
rect 19970 -9120 20015 -9000
rect 20135 -9120 20180 -9000
rect 20300 -9120 20345 -9000
rect 20465 -9120 20520 -9000
rect 20640 -9120 20685 -9000
rect 20805 -9120 20850 -9000
rect 20970 -9120 21015 -9000
rect 21135 -9120 21190 -9000
rect 21310 -9120 21355 -9000
rect 21475 -9120 21520 -9000
rect 21640 -9120 21685 -9000
rect 21805 -9120 21860 -9000
rect 21980 -9120 22025 -9000
rect 22145 -9120 22190 -9000
rect 22310 -9120 22355 -9000
rect 22475 -9120 22530 -9000
rect 22650 -9120 22695 -9000
rect 22815 -9120 22860 -9000
rect 22980 -9120 23025 -9000
rect 23145 -9120 23200 -9000
rect 23320 -9120 23365 -9000
rect 23485 -9120 23530 -9000
rect 23650 -9120 23695 -9000
rect 23815 -9120 23870 -9000
rect 23990 -9120 24015 -9000
rect 18485 -9175 24015 -9120
rect 18485 -9295 18510 -9175
rect 18630 -9295 18675 -9175
rect 18795 -9295 18840 -9175
rect 18960 -9295 19005 -9175
rect 19125 -9295 19180 -9175
rect 19300 -9295 19345 -9175
rect 19465 -9295 19510 -9175
rect 19630 -9295 19675 -9175
rect 19795 -9295 19850 -9175
rect 19970 -9295 20015 -9175
rect 20135 -9295 20180 -9175
rect 20300 -9295 20345 -9175
rect 20465 -9295 20520 -9175
rect 20640 -9295 20685 -9175
rect 20805 -9295 20850 -9175
rect 20970 -9295 21015 -9175
rect 21135 -9295 21190 -9175
rect 21310 -9295 21355 -9175
rect 21475 -9295 21520 -9175
rect 21640 -9295 21685 -9175
rect 21805 -9295 21860 -9175
rect 21980 -9295 22025 -9175
rect 22145 -9295 22190 -9175
rect 22310 -9295 22355 -9175
rect 22475 -9295 22530 -9175
rect 22650 -9295 22695 -9175
rect 22815 -9295 22860 -9175
rect 22980 -9295 23025 -9175
rect 23145 -9295 23200 -9175
rect 23320 -9295 23365 -9175
rect 23485 -9295 23530 -9175
rect 23650 -9295 23695 -9175
rect 23815 -9295 23870 -9175
rect 23990 -9295 24015 -9175
rect 18485 -9340 24015 -9295
rect 18485 -9460 18510 -9340
rect 18630 -9460 18675 -9340
rect 18795 -9460 18840 -9340
rect 18960 -9460 19005 -9340
rect 19125 -9460 19180 -9340
rect 19300 -9460 19345 -9340
rect 19465 -9460 19510 -9340
rect 19630 -9460 19675 -9340
rect 19795 -9460 19850 -9340
rect 19970 -9460 20015 -9340
rect 20135 -9460 20180 -9340
rect 20300 -9460 20345 -9340
rect 20465 -9460 20520 -9340
rect 20640 -9460 20685 -9340
rect 20805 -9460 20850 -9340
rect 20970 -9460 21015 -9340
rect 21135 -9460 21190 -9340
rect 21310 -9460 21355 -9340
rect 21475 -9460 21520 -9340
rect 21640 -9460 21685 -9340
rect 21805 -9460 21860 -9340
rect 21980 -9460 22025 -9340
rect 22145 -9460 22190 -9340
rect 22310 -9460 22355 -9340
rect 22475 -9460 22530 -9340
rect 22650 -9460 22695 -9340
rect 22815 -9460 22860 -9340
rect 22980 -9460 23025 -9340
rect 23145 -9460 23200 -9340
rect 23320 -9460 23365 -9340
rect 23485 -9460 23530 -9340
rect 23650 -9460 23695 -9340
rect 23815 -9460 23870 -9340
rect 23990 -9460 24015 -9340
rect 18485 -9505 24015 -9460
rect 18485 -9625 18510 -9505
rect 18630 -9625 18675 -9505
rect 18795 -9625 18840 -9505
rect 18960 -9625 19005 -9505
rect 19125 -9625 19180 -9505
rect 19300 -9625 19345 -9505
rect 19465 -9625 19510 -9505
rect 19630 -9625 19675 -9505
rect 19795 -9625 19850 -9505
rect 19970 -9625 20015 -9505
rect 20135 -9625 20180 -9505
rect 20300 -9625 20345 -9505
rect 20465 -9625 20520 -9505
rect 20640 -9625 20685 -9505
rect 20805 -9625 20850 -9505
rect 20970 -9625 21015 -9505
rect 21135 -9625 21190 -9505
rect 21310 -9625 21355 -9505
rect 21475 -9625 21520 -9505
rect 21640 -9625 21685 -9505
rect 21805 -9625 21860 -9505
rect 21980 -9625 22025 -9505
rect 22145 -9625 22190 -9505
rect 22310 -9625 22355 -9505
rect 22475 -9625 22530 -9505
rect 22650 -9625 22695 -9505
rect 22815 -9625 22860 -9505
rect 22980 -9625 23025 -9505
rect 23145 -9625 23200 -9505
rect 23320 -9625 23365 -9505
rect 23485 -9625 23530 -9505
rect 23650 -9625 23695 -9505
rect 23815 -9625 23870 -9505
rect 23990 -9625 24015 -9505
rect 18485 -9670 24015 -9625
rect 18485 -9790 18510 -9670
rect 18630 -9790 18675 -9670
rect 18795 -9790 18840 -9670
rect 18960 -9790 19005 -9670
rect 19125 -9790 19180 -9670
rect 19300 -9790 19345 -9670
rect 19465 -9790 19510 -9670
rect 19630 -9790 19675 -9670
rect 19795 -9790 19850 -9670
rect 19970 -9790 20015 -9670
rect 20135 -9790 20180 -9670
rect 20300 -9790 20345 -9670
rect 20465 -9790 20520 -9670
rect 20640 -9790 20685 -9670
rect 20805 -9790 20850 -9670
rect 20970 -9790 21015 -9670
rect 21135 -9790 21190 -9670
rect 21310 -9790 21355 -9670
rect 21475 -9790 21520 -9670
rect 21640 -9790 21685 -9670
rect 21805 -9790 21860 -9670
rect 21980 -9790 22025 -9670
rect 22145 -9790 22190 -9670
rect 22310 -9790 22355 -9670
rect 22475 -9790 22530 -9670
rect 22650 -9790 22695 -9670
rect 22815 -9790 22860 -9670
rect 22980 -9790 23025 -9670
rect 23145 -9790 23200 -9670
rect 23320 -9790 23365 -9670
rect 23485 -9790 23530 -9670
rect 23650 -9790 23695 -9670
rect 23815 -9790 23870 -9670
rect 23990 -9790 24015 -9670
rect 18485 -9860 24015 -9790
rect 24175 -4310 29705 -4285
rect 24175 -4430 24200 -4310
rect 24320 -4430 24365 -4310
rect 24485 -4430 24530 -4310
rect 24650 -4430 24695 -4310
rect 24815 -4430 24870 -4310
rect 24990 -4430 25035 -4310
rect 25155 -4430 25200 -4310
rect 25320 -4430 25365 -4310
rect 25485 -4430 25540 -4310
rect 25660 -4430 25705 -4310
rect 25825 -4430 25870 -4310
rect 25990 -4430 26035 -4310
rect 26155 -4430 26210 -4310
rect 26330 -4430 26375 -4310
rect 26495 -4430 26540 -4310
rect 26660 -4430 26705 -4310
rect 26825 -4430 26880 -4310
rect 27000 -4430 27045 -4310
rect 27165 -4430 27210 -4310
rect 27330 -4430 27375 -4310
rect 27495 -4430 27550 -4310
rect 27670 -4430 27715 -4310
rect 27835 -4430 27880 -4310
rect 28000 -4430 28045 -4310
rect 28165 -4430 28220 -4310
rect 28340 -4430 28385 -4310
rect 28505 -4430 28550 -4310
rect 28670 -4430 28715 -4310
rect 28835 -4430 28890 -4310
rect 29010 -4430 29055 -4310
rect 29175 -4430 29220 -4310
rect 29340 -4430 29385 -4310
rect 29505 -4430 29560 -4310
rect 29680 -4430 29705 -4310
rect 24175 -4485 29705 -4430
rect 24175 -4605 24200 -4485
rect 24320 -4605 24365 -4485
rect 24485 -4605 24530 -4485
rect 24650 -4605 24695 -4485
rect 24815 -4605 24870 -4485
rect 24990 -4605 25035 -4485
rect 25155 -4605 25200 -4485
rect 25320 -4605 25365 -4485
rect 25485 -4605 25540 -4485
rect 25660 -4605 25705 -4485
rect 25825 -4605 25870 -4485
rect 25990 -4605 26035 -4485
rect 26155 -4605 26210 -4485
rect 26330 -4605 26375 -4485
rect 26495 -4605 26540 -4485
rect 26660 -4605 26705 -4485
rect 26825 -4605 26880 -4485
rect 27000 -4605 27045 -4485
rect 27165 -4605 27210 -4485
rect 27330 -4605 27375 -4485
rect 27495 -4605 27550 -4485
rect 27670 -4605 27715 -4485
rect 27835 -4605 27880 -4485
rect 28000 -4605 28045 -4485
rect 28165 -4605 28220 -4485
rect 28340 -4605 28385 -4485
rect 28505 -4605 28550 -4485
rect 28670 -4605 28715 -4485
rect 28835 -4605 28890 -4485
rect 29010 -4605 29055 -4485
rect 29175 -4605 29220 -4485
rect 29340 -4605 29385 -4485
rect 29505 -4605 29560 -4485
rect 29680 -4605 29705 -4485
rect 24175 -4650 29705 -4605
rect 24175 -4770 24200 -4650
rect 24320 -4770 24365 -4650
rect 24485 -4770 24530 -4650
rect 24650 -4770 24695 -4650
rect 24815 -4770 24870 -4650
rect 24990 -4770 25035 -4650
rect 25155 -4770 25200 -4650
rect 25320 -4770 25365 -4650
rect 25485 -4770 25540 -4650
rect 25660 -4770 25705 -4650
rect 25825 -4770 25870 -4650
rect 25990 -4770 26035 -4650
rect 26155 -4770 26210 -4650
rect 26330 -4770 26375 -4650
rect 26495 -4770 26540 -4650
rect 26660 -4770 26705 -4650
rect 26825 -4770 26880 -4650
rect 27000 -4770 27045 -4650
rect 27165 -4770 27210 -4650
rect 27330 -4770 27375 -4650
rect 27495 -4770 27550 -4650
rect 27670 -4770 27715 -4650
rect 27835 -4770 27880 -4650
rect 28000 -4770 28045 -4650
rect 28165 -4770 28220 -4650
rect 28340 -4770 28385 -4650
rect 28505 -4770 28550 -4650
rect 28670 -4770 28715 -4650
rect 28835 -4770 28890 -4650
rect 29010 -4770 29055 -4650
rect 29175 -4770 29220 -4650
rect 29340 -4770 29385 -4650
rect 29505 -4770 29560 -4650
rect 29680 -4770 29705 -4650
rect 24175 -4815 29705 -4770
rect 24175 -4935 24200 -4815
rect 24320 -4935 24365 -4815
rect 24485 -4935 24530 -4815
rect 24650 -4935 24695 -4815
rect 24815 -4935 24870 -4815
rect 24990 -4935 25035 -4815
rect 25155 -4935 25200 -4815
rect 25320 -4935 25365 -4815
rect 25485 -4935 25540 -4815
rect 25660 -4935 25705 -4815
rect 25825 -4935 25870 -4815
rect 25990 -4935 26035 -4815
rect 26155 -4935 26210 -4815
rect 26330 -4935 26375 -4815
rect 26495 -4935 26540 -4815
rect 26660 -4935 26705 -4815
rect 26825 -4935 26880 -4815
rect 27000 -4935 27045 -4815
rect 27165 -4935 27210 -4815
rect 27330 -4935 27375 -4815
rect 27495 -4935 27550 -4815
rect 27670 -4935 27715 -4815
rect 27835 -4935 27880 -4815
rect 28000 -4935 28045 -4815
rect 28165 -4935 28220 -4815
rect 28340 -4935 28385 -4815
rect 28505 -4935 28550 -4815
rect 28670 -4935 28715 -4815
rect 28835 -4935 28890 -4815
rect 29010 -4935 29055 -4815
rect 29175 -4935 29220 -4815
rect 29340 -4935 29385 -4815
rect 29505 -4935 29560 -4815
rect 29680 -4935 29705 -4815
rect 24175 -4980 29705 -4935
rect 24175 -5100 24200 -4980
rect 24320 -5100 24365 -4980
rect 24485 -5100 24530 -4980
rect 24650 -5100 24695 -4980
rect 24815 -5100 24870 -4980
rect 24990 -5100 25035 -4980
rect 25155 -5100 25200 -4980
rect 25320 -5100 25365 -4980
rect 25485 -5100 25540 -4980
rect 25660 -5100 25705 -4980
rect 25825 -5100 25870 -4980
rect 25990 -5100 26035 -4980
rect 26155 -5100 26210 -4980
rect 26330 -5100 26375 -4980
rect 26495 -5100 26540 -4980
rect 26660 -5100 26705 -4980
rect 26825 -5100 26880 -4980
rect 27000 -5100 27045 -4980
rect 27165 -5100 27210 -4980
rect 27330 -5100 27375 -4980
rect 27495 -5100 27550 -4980
rect 27670 -5100 27715 -4980
rect 27835 -5100 27880 -4980
rect 28000 -5100 28045 -4980
rect 28165 -5100 28220 -4980
rect 28340 -5100 28385 -4980
rect 28505 -5100 28550 -4980
rect 28670 -5100 28715 -4980
rect 28835 -5100 28890 -4980
rect 29010 -5100 29055 -4980
rect 29175 -5100 29220 -4980
rect 29340 -5100 29385 -4980
rect 29505 -5100 29560 -4980
rect 29680 -5100 29705 -4980
rect 24175 -5155 29705 -5100
rect 24175 -5275 24200 -5155
rect 24320 -5275 24365 -5155
rect 24485 -5275 24530 -5155
rect 24650 -5275 24695 -5155
rect 24815 -5275 24870 -5155
rect 24990 -5275 25035 -5155
rect 25155 -5275 25200 -5155
rect 25320 -5275 25365 -5155
rect 25485 -5275 25540 -5155
rect 25660 -5275 25705 -5155
rect 25825 -5275 25870 -5155
rect 25990 -5275 26035 -5155
rect 26155 -5275 26210 -5155
rect 26330 -5275 26375 -5155
rect 26495 -5275 26540 -5155
rect 26660 -5275 26705 -5155
rect 26825 -5275 26880 -5155
rect 27000 -5275 27045 -5155
rect 27165 -5275 27210 -5155
rect 27330 -5275 27375 -5155
rect 27495 -5275 27550 -5155
rect 27670 -5275 27715 -5155
rect 27835 -5275 27880 -5155
rect 28000 -5275 28045 -5155
rect 28165 -5275 28220 -5155
rect 28340 -5275 28385 -5155
rect 28505 -5275 28550 -5155
rect 28670 -5275 28715 -5155
rect 28835 -5275 28890 -5155
rect 29010 -5275 29055 -5155
rect 29175 -5275 29220 -5155
rect 29340 -5275 29385 -5155
rect 29505 -5275 29560 -5155
rect 29680 -5275 29705 -5155
rect 24175 -5320 29705 -5275
rect 24175 -5440 24200 -5320
rect 24320 -5440 24365 -5320
rect 24485 -5440 24530 -5320
rect 24650 -5440 24695 -5320
rect 24815 -5440 24870 -5320
rect 24990 -5440 25035 -5320
rect 25155 -5440 25200 -5320
rect 25320 -5440 25365 -5320
rect 25485 -5440 25540 -5320
rect 25660 -5440 25705 -5320
rect 25825 -5440 25870 -5320
rect 25990 -5440 26035 -5320
rect 26155 -5440 26210 -5320
rect 26330 -5440 26375 -5320
rect 26495 -5440 26540 -5320
rect 26660 -5440 26705 -5320
rect 26825 -5440 26880 -5320
rect 27000 -5440 27045 -5320
rect 27165 -5440 27210 -5320
rect 27330 -5440 27375 -5320
rect 27495 -5440 27550 -5320
rect 27670 -5440 27715 -5320
rect 27835 -5440 27880 -5320
rect 28000 -5440 28045 -5320
rect 28165 -5440 28220 -5320
rect 28340 -5440 28385 -5320
rect 28505 -5440 28550 -5320
rect 28670 -5440 28715 -5320
rect 28835 -5440 28890 -5320
rect 29010 -5440 29055 -5320
rect 29175 -5440 29220 -5320
rect 29340 -5440 29385 -5320
rect 29505 -5440 29560 -5320
rect 29680 -5440 29705 -5320
rect 24175 -5485 29705 -5440
rect 24175 -5605 24200 -5485
rect 24320 -5605 24365 -5485
rect 24485 -5605 24530 -5485
rect 24650 -5605 24695 -5485
rect 24815 -5605 24870 -5485
rect 24990 -5605 25035 -5485
rect 25155 -5605 25200 -5485
rect 25320 -5605 25365 -5485
rect 25485 -5605 25540 -5485
rect 25660 -5605 25705 -5485
rect 25825 -5605 25870 -5485
rect 25990 -5605 26035 -5485
rect 26155 -5605 26210 -5485
rect 26330 -5605 26375 -5485
rect 26495 -5605 26540 -5485
rect 26660 -5605 26705 -5485
rect 26825 -5605 26880 -5485
rect 27000 -5605 27045 -5485
rect 27165 -5605 27210 -5485
rect 27330 -5605 27375 -5485
rect 27495 -5605 27550 -5485
rect 27670 -5605 27715 -5485
rect 27835 -5605 27880 -5485
rect 28000 -5605 28045 -5485
rect 28165 -5605 28220 -5485
rect 28340 -5605 28385 -5485
rect 28505 -5605 28550 -5485
rect 28670 -5605 28715 -5485
rect 28835 -5605 28890 -5485
rect 29010 -5605 29055 -5485
rect 29175 -5605 29220 -5485
rect 29340 -5605 29385 -5485
rect 29505 -5605 29560 -5485
rect 29680 -5605 29705 -5485
rect 24175 -5650 29705 -5605
rect 24175 -5770 24200 -5650
rect 24320 -5770 24365 -5650
rect 24485 -5770 24530 -5650
rect 24650 -5770 24695 -5650
rect 24815 -5770 24870 -5650
rect 24990 -5770 25035 -5650
rect 25155 -5770 25200 -5650
rect 25320 -5770 25365 -5650
rect 25485 -5770 25540 -5650
rect 25660 -5770 25705 -5650
rect 25825 -5770 25870 -5650
rect 25990 -5770 26035 -5650
rect 26155 -5770 26210 -5650
rect 26330 -5770 26375 -5650
rect 26495 -5770 26540 -5650
rect 26660 -5770 26705 -5650
rect 26825 -5770 26880 -5650
rect 27000 -5770 27045 -5650
rect 27165 -5770 27210 -5650
rect 27330 -5770 27375 -5650
rect 27495 -5770 27550 -5650
rect 27670 -5770 27715 -5650
rect 27835 -5770 27880 -5650
rect 28000 -5770 28045 -5650
rect 28165 -5770 28220 -5650
rect 28340 -5770 28385 -5650
rect 28505 -5770 28550 -5650
rect 28670 -5770 28715 -5650
rect 28835 -5770 28890 -5650
rect 29010 -5770 29055 -5650
rect 29175 -5770 29220 -5650
rect 29340 -5770 29385 -5650
rect 29505 -5770 29560 -5650
rect 29680 -5770 29705 -5650
rect 24175 -5825 29705 -5770
rect 24175 -5945 24200 -5825
rect 24320 -5945 24365 -5825
rect 24485 -5945 24530 -5825
rect 24650 -5945 24695 -5825
rect 24815 -5945 24870 -5825
rect 24990 -5945 25035 -5825
rect 25155 -5945 25200 -5825
rect 25320 -5945 25365 -5825
rect 25485 -5945 25540 -5825
rect 25660 -5945 25705 -5825
rect 25825 -5945 25870 -5825
rect 25990 -5945 26035 -5825
rect 26155 -5945 26210 -5825
rect 26330 -5945 26375 -5825
rect 26495 -5945 26540 -5825
rect 26660 -5945 26705 -5825
rect 26825 -5945 26880 -5825
rect 27000 -5945 27045 -5825
rect 27165 -5945 27210 -5825
rect 27330 -5945 27375 -5825
rect 27495 -5945 27550 -5825
rect 27670 -5945 27715 -5825
rect 27835 -5945 27880 -5825
rect 28000 -5945 28045 -5825
rect 28165 -5945 28220 -5825
rect 28340 -5945 28385 -5825
rect 28505 -5945 28550 -5825
rect 28670 -5945 28715 -5825
rect 28835 -5945 28890 -5825
rect 29010 -5945 29055 -5825
rect 29175 -5945 29220 -5825
rect 29340 -5945 29385 -5825
rect 29505 -5945 29560 -5825
rect 29680 -5945 29705 -5825
rect 24175 -5990 29705 -5945
rect 24175 -6110 24200 -5990
rect 24320 -6110 24365 -5990
rect 24485 -6110 24530 -5990
rect 24650 -6110 24695 -5990
rect 24815 -6110 24870 -5990
rect 24990 -6110 25035 -5990
rect 25155 -6110 25200 -5990
rect 25320 -6110 25365 -5990
rect 25485 -6110 25540 -5990
rect 25660 -6110 25705 -5990
rect 25825 -6110 25870 -5990
rect 25990 -6110 26035 -5990
rect 26155 -6110 26210 -5990
rect 26330 -6110 26375 -5990
rect 26495 -6110 26540 -5990
rect 26660 -6110 26705 -5990
rect 26825 -6110 26880 -5990
rect 27000 -6110 27045 -5990
rect 27165 -6110 27210 -5990
rect 27330 -6110 27375 -5990
rect 27495 -6110 27550 -5990
rect 27670 -6110 27715 -5990
rect 27835 -6110 27880 -5990
rect 28000 -6110 28045 -5990
rect 28165 -6110 28220 -5990
rect 28340 -6110 28385 -5990
rect 28505 -6110 28550 -5990
rect 28670 -6110 28715 -5990
rect 28835 -6110 28890 -5990
rect 29010 -6110 29055 -5990
rect 29175 -6110 29220 -5990
rect 29340 -6110 29385 -5990
rect 29505 -6110 29560 -5990
rect 29680 -6110 29705 -5990
rect 24175 -6155 29705 -6110
rect 24175 -6275 24200 -6155
rect 24320 -6275 24365 -6155
rect 24485 -6275 24530 -6155
rect 24650 -6275 24695 -6155
rect 24815 -6275 24870 -6155
rect 24990 -6275 25035 -6155
rect 25155 -6275 25200 -6155
rect 25320 -6275 25365 -6155
rect 25485 -6275 25540 -6155
rect 25660 -6275 25705 -6155
rect 25825 -6275 25870 -6155
rect 25990 -6275 26035 -6155
rect 26155 -6275 26210 -6155
rect 26330 -6275 26375 -6155
rect 26495 -6275 26540 -6155
rect 26660 -6275 26705 -6155
rect 26825 -6275 26880 -6155
rect 27000 -6275 27045 -6155
rect 27165 -6275 27210 -6155
rect 27330 -6275 27375 -6155
rect 27495 -6275 27550 -6155
rect 27670 -6275 27715 -6155
rect 27835 -6275 27880 -6155
rect 28000 -6275 28045 -6155
rect 28165 -6275 28220 -6155
rect 28340 -6275 28385 -6155
rect 28505 -6275 28550 -6155
rect 28670 -6275 28715 -6155
rect 28835 -6275 28890 -6155
rect 29010 -6275 29055 -6155
rect 29175 -6275 29220 -6155
rect 29340 -6275 29385 -6155
rect 29505 -6275 29560 -6155
rect 29680 -6275 29705 -6155
rect 24175 -6320 29705 -6275
rect 24175 -6440 24200 -6320
rect 24320 -6440 24365 -6320
rect 24485 -6440 24530 -6320
rect 24650 -6440 24695 -6320
rect 24815 -6440 24870 -6320
rect 24990 -6440 25035 -6320
rect 25155 -6440 25200 -6320
rect 25320 -6440 25365 -6320
rect 25485 -6440 25540 -6320
rect 25660 -6440 25705 -6320
rect 25825 -6440 25870 -6320
rect 25990 -6440 26035 -6320
rect 26155 -6440 26210 -6320
rect 26330 -6440 26375 -6320
rect 26495 -6440 26540 -6320
rect 26660 -6440 26705 -6320
rect 26825 -6440 26880 -6320
rect 27000 -6440 27045 -6320
rect 27165 -6440 27210 -6320
rect 27330 -6440 27375 -6320
rect 27495 -6440 27550 -6320
rect 27670 -6440 27715 -6320
rect 27835 -6440 27880 -6320
rect 28000 -6440 28045 -6320
rect 28165 -6440 28220 -6320
rect 28340 -6440 28385 -6320
rect 28505 -6440 28550 -6320
rect 28670 -6440 28715 -6320
rect 28835 -6440 28890 -6320
rect 29010 -6440 29055 -6320
rect 29175 -6440 29220 -6320
rect 29340 -6440 29385 -6320
rect 29505 -6440 29560 -6320
rect 29680 -6440 29705 -6320
rect 24175 -6495 29705 -6440
rect 24175 -6615 24200 -6495
rect 24320 -6615 24365 -6495
rect 24485 -6615 24530 -6495
rect 24650 -6615 24695 -6495
rect 24815 -6615 24870 -6495
rect 24990 -6615 25035 -6495
rect 25155 -6615 25200 -6495
rect 25320 -6615 25365 -6495
rect 25485 -6615 25540 -6495
rect 25660 -6615 25705 -6495
rect 25825 -6615 25870 -6495
rect 25990 -6615 26035 -6495
rect 26155 -6615 26210 -6495
rect 26330 -6615 26375 -6495
rect 26495 -6615 26540 -6495
rect 26660 -6615 26705 -6495
rect 26825 -6615 26880 -6495
rect 27000 -6615 27045 -6495
rect 27165 -6615 27210 -6495
rect 27330 -6615 27375 -6495
rect 27495 -6615 27550 -6495
rect 27670 -6615 27715 -6495
rect 27835 -6615 27880 -6495
rect 28000 -6615 28045 -6495
rect 28165 -6615 28220 -6495
rect 28340 -6615 28385 -6495
rect 28505 -6615 28550 -6495
rect 28670 -6615 28715 -6495
rect 28835 -6615 28890 -6495
rect 29010 -6615 29055 -6495
rect 29175 -6615 29220 -6495
rect 29340 -6615 29385 -6495
rect 29505 -6615 29560 -6495
rect 29680 -6615 29705 -6495
rect 24175 -6660 29705 -6615
rect 24175 -6780 24200 -6660
rect 24320 -6780 24365 -6660
rect 24485 -6780 24530 -6660
rect 24650 -6780 24695 -6660
rect 24815 -6780 24870 -6660
rect 24990 -6780 25035 -6660
rect 25155 -6780 25200 -6660
rect 25320 -6780 25365 -6660
rect 25485 -6780 25540 -6660
rect 25660 -6780 25705 -6660
rect 25825 -6780 25870 -6660
rect 25990 -6780 26035 -6660
rect 26155 -6780 26210 -6660
rect 26330 -6780 26375 -6660
rect 26495 -6780 26540 -6660
rect 26660 -6780 26705 -6660
rect 26825 -6780 26880 -6660
rect 27000 -6780 27045 -6660
rect 27165 -6780 27210 -6660
rect 27330 -6780 27375 -6660
rect 27495 -6780 27550 -6660
rect 27670 -6780 27715 -6660
rect 27835 -6780 27880 -6660
rect 28000 -6780 28045 -6660
rect 28165 -6780 28220 -6660
rect 28340 -6780 28385 -6660
rect 28505 -6780 28550 -6660
rect 28670 -6780 28715 -6660
rect 28835 -6780 28890 -6660
rect 29010 -6780 29055 -6660
rect 29175 -6780 29220 -6660
rect 29340 -6780 29385 -6660
rect 29505 -6780 29560 -6660
rect 29680 -6780 29705 -6660
rect 24175 -6825 29705 -6780
rect 24175 -6945 24200 -6825
rect 24320 -6945 24365 -6825
rect 24485 -6945 24530 -6825
rect 24650 -6945 24695 -6825
rect 24815 -6945 24870 -6825
rect 24990 -6945 25035 -6825
rect 25155 -6945 25200 -6825
rect 25320 -6945 25365 -6825
rect 25485 -6945 25540 -6825
rect 25660 -6945 25705 -6825
rect 25825 -6945 25870 -6825
rect 25990 -6945 26035 -6825
rect 26155 -6945 26210 -6825
rect 26330 -6945 26375 -6825
rect 26495 -6945 26540 -6825
rect 26660 -6945 26705 -6825
rect 26825 -6945 26880 -6825
rect 27000 -6945 27045 -6825
rect 27165 -6945 27210 -6825
rect 27330 -6945 27375 -6825
rect 27495 -6945 27550 -6825
rect 27670 -6945 27715 -6825
rect 27835 -6945 27880 -6825
rect 28000 -6945 28045 -6825
rect 28165 -6945 28220 -6825
rect 28340 -6945 28385 -6825
rect 28505 -6945 28550 -6825
rect 28670 -6945 28715 -6825
rect 28835 -6945 28890 -6825
rect 29010 -6945 29055 -6825
rect 29175 -6945 29220 -6825
rect 29340 -6945 29385 -6825
rect 29505 -6945 29560 -6825
rect 29680 -6945 29705 -6825
rect 24175 -6990 29705 -6945
rect 24175 -7110 24200 -6990
rect 24320 -7110 24365 -6990
rect 24485 -7110 24530 -6990
rect 24650 -7110 24695 -6990
rect 24815 -7110 24870 -6990
rect 24990 -7110 25035 -6990
rect 25155 -7110 25200 -6990
rect 25320 -7110 25365 -6990
rect 25485 -7110 25540 -6990
rect 25660 -7110 25705 -6990
rect 25825 -7110 25870 -6990
rect 25990 -7110 26035 -6990
rect 26155 -7110 26210 -6990
rect 26330 -7110 26375 -6990
rect 26495 -7110 26540 -6990
rect 26660 -7110 26705 -6990
rect 26825 -7110 26880 -6990
rect 27000 -7110 27045 -6990
rect 27165 -7110 27210 -6990
rect 27330 -7110 27375 -6990
rect 27495 -7110 27550 -6990
rect 27670 -7110 27715 -6990
rect 27835 -7110 27880 -6990
rect 28000 -7110 28045 -6990
rect 28165 -7110 28220 -6990
rect 28340 -7110 28385 -6990
rect 28505 -7110 28550 -6990
rect 28670 -7110 28715 -6990
rect 28835 -7110 28890 -6990
rect 29010 -7110 29055 -6990
rect 29175 -7110 29220 -6990
rect 29340 -7110 29385 -6990
rect 29505 -7110 29560 -6990
rect 29680 -7110 29705 -6990
rect 24175 -7165 29705 -7110
rect 24175 -7285 24200 -7165
rect 24320 -7285 24365 -7165
rect 24485 -7285 24530 -7165
rect 24650 -7285 24695 -7165
rect 24815 -7285 24870 -7165
rect 24990 -7285 25035 -7165
rect 25155 -7285 25200 -7165
rect 25320 -7285 25365 -7165
rect 25485 -7285 25540 -7165
rect 25660 -7285 25705 -7165
rect 25825 -7285 25870 -7165
rect 25990 -7285 26035 -7165
rect 26155 -7285 26210 -7165
rect 26330 -7285 26375 -7165
rect 26495 -7285 26540 -7165
rect 26660 -7285 26705 -7165
rect 26825 -7285 26880 -7165
rect 27000 -7285 27045 -7165
rect 27165 -7285 27210 -7165
rect 27330 -7285 27375 -7165
rect 27495 -7285 27550 -7165
rect 27670 -7285 27715 -7165
rect 27835 -7285 27880 -7165
rect 28000 -7285 28045 -7165
rect 28165 -7285 28220 -7165
rect 28340 -7285 28385 -7165
rect 28505 -7285 28550 -7165
rect 28670 -7285 28715 -7165
rect 28835 -7285 28890 -7165
rect 29010 -7285 29055 -7165
rect 29175 -7285 29220 -7165
rect 29340 -7285 29385 -7165
rect 29505 -7285 29560 -7165
rect 29680 -7285 29705 -7165
rect 24175 -7330 29705 -7285
rect 24175 -7450 24200 -7330
rect 24320 -7450 24365 -7330
rect 24485 -7450 24530 -7330
rect 24650 -7450 24695 -7330
rect 24815 -7450 24870 -7330
rect 24990 -7450 25035 -7330
rect 25155 -7450 25200 -7330
rect 25320 -7450 25365 -7330
rect 25485 -7450 25540 -7330
rect 25660 -7450 25705 -7330
rect 25825 -7450 25870 -7330
rect 25990 -7450 26035 -7330
rect 26155 -7450 26210 -7330
rect 26330 -7450 26375 -7330
rect 26495 -7450 26540 -7330
rect 26660 -7450 26705 -7330
rect 26825 -7450 26880 -7330
rect 27000 -7450 27045 -7330
rect 27165 -7450 27210 -7330
rect 27330 -7450 27375 -7330
rect 27495 -7450 27550 -7330
rect 27670 -7450 27715 -7330
rect 27835 -7450 27880 -7330
rect 28000 -7450 28045 -7330
rect 28165 -7450 28220 -7330
rect 28340 -7450 28385 -7330
rect 28505 -7450 28550 -7330
rect 28670 -7450 28715 -7330
rect 28835 -7450 28890 -7330
rect 29010 -7450 29055 -7330
rect 29175 -7450 29220 -7330
rect 29340 -7450 29385 -7330
rect 29505 -7450 29560 -7330
rect 29680 -7450 29705 -7330
rect 24175 -7495 29705 -7450
rect 24175 -7615 24200 -7495
rect 24320 -7615 24365 -7495
rect 24485 -7615 24530 -7495
rect 24650 -7615 24695 -7495
rect 24815 -7615 24870 -7495
rect 24990 -7615 25035 -7495
rect 25155 -7615 25200 -7495
rect 25320 -7615 25365 -7495
rect 25485 -7615 25540 -7495
rect 25660 -7615 25705 -7495
rect 25825 -7615 25870 -7495
rect 25990 -7615 26035 -7495
rect 26155 -7615 26210 -7495
rect 26330 -7615 26375 -7495
rect 26495 -7615 26540 -7495
rect 26660 -7615 26705 -7495
rect 26825 -7615 26880 -7495
rect 27000 -7615 27045 -7495
rect 27165 -7615 27210 -7495
rect 27330 -7615 27375 -7495
rect 27495 -7615 27550 -7495
rect 27670 -7615 27715 -7495
rect 27835 -7615 27880 -7495
rect 28000 -7615 28045 -7495
rect 28165 -7615 28220 -7495
rect 28340 -7615 28385 -7495
rect 28505 -7615 28550 -7495
rect 28670 -7615 28715 -7495
rect 28835 -7615 28890 -7495
rect 29010 -7615 29055 -7495
rect 29175 -7615 29220 -7495
rect 29340 -7615 29385 -7495
rect 29505 -7615 29560 -7495
rect 29680 -7615 29705 -7495
rect 24175 -7660 29705 -7615
rect 24175 -7780 24200 -7660
rect 24320 -7780 24365 -7660
rect 24485 -7780 24530 -7660
rect 24650 -7780 24695 -7660
rect 24815 -7780 24870 -7660
rect 24990 -7780 25035 -7660
rect 25155 -7780 25200 -7660
rect 25320 -7780 25365 -7660
rect 25485 -7780 25540 -7660
rect 25660 -7780 25705 -7660
rect 25825 -7780 25870 -7660
rect 25990 -7780 26035 -7660
rect 26155 -7780 26210 -7660
rect 26330 -7780 26375 -7660
rect 26495 -7780 26540 -7660
rect 26660 -7780 26705 -7660
rect 26825 -7780 26880 -7660
rect 27000 -7780 27045 -7660
rect 27165 -7780 27210 -7660
rect 27330 -7780 27375 -7660
rect 27495 -7780 27550 -7660
rect 27670 -7780 27715 -7660
rect 27835 -7780 27880 -7660
rect 28000 -7780 28045 -7660
rect 28165 -7780 28220 -7660
rect 28340 -7780 28385 -7660
rect 28505 -7780 28550 -7660
rect 28670 -7780 28715 -7660
rect 28835 -7780 28890 -7660
rect 29010 -7780 29055 -7660
rect 29175 -7780 29220 -7660
rect 29340 -7780 29385 -7660
rect 29505 -7780 29560 -7660
rect 29680 -7780 29705 -7660
rect 24175 -7835 29705 -7780
rect 24175 -7955 24200 -7835
rect 24320 -7955 24365 -7835
rect 24485 -7955 24530 -7835
rect 24650 -7955 24695 -7835
rect 24815 -7955 24870 -7835
rect 24990 -7955 25035 -7835
rect 25155 -7955 25200 -7835
rect 25320 -7955 25365 -7835
rect 25485 -7955 25540 -7835
rect 25660 -7955 25705 -7835
rect 25825 -7955 25870 -7835
rect 25990 -7955 26035 -7835
rect 26155 -7955 26210 -7835
rect 26330 -7955 26375 -7835
rect 26495 -7955 26540 -7835
rect 26660 -7955 26705 -7835
rect 26825 -7955 26880 -7835
rect 27000 -7955 27045 -7835
rect 27165 -7955 27210 -7835
rect 27330 -7955 27375 -7835
rect 27495 -7955 27550 -7835
rect 27670 -7955 27715 -7835
rect 27835 -7955 27880 -7835
rect 28000 -7955 28045 -7835
rect 28165 -7955 28220 -7835
rect 28340 -7955 28385 -7835
rect 28505 -7955 28550 -7835
rect 28670 -7955 28715 -7835
rect 28835 -7955 28890 -7835
rect 29010 -7955 29055 -7835
rect 29175 -7955 29220 -7835
rect 29340 -7955 29385 -7835
rect 29505 -7955 29560 -7835
rect 29680 -7955 29705 -7835
rect 24175 -8000 29705 -7955
rect 24175 -8120 24200 -8000
rect 24320 -8120 24365 -8000
rect 24485 -8120 24530 -8000
rect 24650 -8120 24695 -8000
rect 24815 -8120 24870 -8000
rect 24990 -8120 25035 -8000
rect 25155 -8120 25200 -8000
rect 25320 -8120 25365 -8000
rect 25485 -8120 25540 -8000
rect 25660 -8120 25705 -8000
rect 25825 -8120 25870 -8000
rect 25990 -8120 26035 -8000
rect 26155 -8120 26210 -8000
rect 26330 -8120 26375 -8000
rect 26495 -8120 26540 -8000
rect 26660 -8120 26705 -8000
rect 26825 -8120 26880 -8000
rect 27000 -8120 27045 -8000
rect 27165 -8120 27210 -8000
rect 27330 -8120 27375 -8000
rect 27495 -8120 27550 -8000
rect 27670 -8120 27715 -8000
rect 27835 -8120 27880 -8000
rect 28000 -8120 28045 -8000
rect 28165 -8120 28220 -8000
rect 28340 -8120 28385 -8000
rect 28505 -8120 28550 -8000
rect 28670 -8120 28715 -8000
rect 28835 -8120 28890 -8000
rect 29010 -8120 29055 -8000
rect 29175 -8120 29220 -8000
rect 29340 -8120 29385 -8000
rect 29505 -8120 29560 -8000
rect 29680 -8120 29705 -8000
rect 24175 -8165 29705 -8120
rect 24175 -8285 24200 -8165
rect 24320 -8285 24365 -8165
rect 24485 -8285 24530 -8165
rect 24650 -8285 24695 -8165
rect 24815 -8285 24870 -8165
rect 24990 -8285 25035 -8165
rect 25155 -8285 25200 -8165
rect 25320 -8285 25365 -8165
rect 25485 -8285 25540 -8165
rect 25660 -8285 25705 -8165
rect 25825 -8285 25870 -8165
rect 25990 -8285 26035 -8165
rect 26155 -8285 26210 -8165
rect 26330 -8285 26375 -8165
rect 26495 -8285 26540 -8165
rect 26660 -8285 26705 -8165
rect 26825 -8285 26880 -8165
rect 27000 -8285 27045 -8165
rect 27165 -8285 27210 -8165
rect 27330 -8285 27375 -8165
rect 27495 -8285 27550 -8165
rect 27670 -8285 27715 -8165
rect 27835 -8285 27880 -8165
rect 28000 -8285 28045 -8165
rect 28165 -8285 28220 -8165
rect 28340 -8285 28385 -8165
rect 28505 -8285 28550 -8165
rect 28670 -8285 28715 -8165
rect 28835 -8285 28890 -8165
rect 29010 -8285 29055 -8165
rect 29175 -8285 29220 -8165
rect 29340 -8285 29385 -8165
rect 29505 -8285 29560 -8165
rect 29680 -8285 29705 -8165
rect 24175 -8330 29705 -8285
rect 24175 -8450 24200 -8330
rect 24320 -8450 24365 -8330
rect 24485 -8450 24530 -8330
rect 24650 -8450 24695 -8330
rect 24815 -8450 24870 -8330
rect 24990 -8450 25035 -8330
rect 25155 -8450 25200 -8330
rect 25320 -8450 25365 -8330
rect 25485 -8450 25540 -8330
rect 25660 -8450 25705 -8330
rect 25825 -8450 25870 -8330
rect 25990 -8450 26035 -8330
rect 26155 -8450 26210 -8330
rect 26330 -8450 26375 -8330
rect 26495 -8450 26540 -8330
rect 26660 -8450 26705 -8330
rect 26825 -8450 26880 -8330
rect 27000 -8450 27045 -8330
rect 27165 -8450 27210 -8330
rect 27330 -8450 27375 -8330
rect 27495 -8450 27550 -8330
rect 27670 -8450 27715 -8330
rect 27835 -8450 27880 -8330
rect 28000 -8450 28045 -8330
rect 28165 -8450 28220 -8330
rect 28340 -8450 28385 -8330
rect 28505 -8450 28550 -8330
rect 28670 -8450 28715 -8330
rect 28835 -8450 28890 -8330
rect 29010 -8450 29055 -8330
rect 29175 -8450 29220 -8330
rect 29340 -8450 29385 -8330
rect 29505 -8450 29560 -8330
rect 29680 -8450 29705 -8330
rect 24175 -8505 29705 -8450
rect 24175 -8625 24200 -8505
rect 24320 -8625 24365 -8505
rect 24485 -8625 24530 -8505
rect 24650 -8625 24695 -8505
rect 24815 -8625 24870 -8505
rect 24990 -8625 25035 -8505
rect 25155 -8625 25200 -8505
rect 25320 -8625 25365 -8505
rect 25485 -8625 25540 -8505
rect 25660 -8625 25705 -8505
rect 25825 -8625 25870 -8505
rect 25990 -8625 26035 -8505
rect 26155 -8625 26210 -8505
rect 26330 -8625 26375 -8505
rect 26495 -8625 26540 -8505
rect 26660 -8625 26705 -8505
rect 26825 -8625 26880 -8505
rect 27000 -8625 27045 -8505
rect 27165 -8625 27210 -8505
rect 27330 -8625 27375 -8505
rect 27495 -8625 27550 -8505
rect 27670 -8625 27715 -8505
rect 27835 -8625 27880 -8505
rect 28000 -8625 28045 -8505
rect 28165 -8625 28220 -8505
rect 28340 -8625 28385 -8505
rect 28505 -8625 28550 -8505
rect 28670 -8625 28715 -8505
rect 28835 -8625 28890 -8505
rect 29010 -8625 29055 -8505
rect 29175 -8625 29220 -8505
rect 29340 -8625 29385 -8505
rect 29505 -8625 29560 -8505
rect 29680 -8625 29705 -8505
rect 24175 -8670 29705 -8625
rect 24175 -8790 24200 -8670
rect 24320 -8790 24365 -8670
rect 24485 -8790 24530 -8670
rect 24650 -8790 24695 -8670
rect 24815 -8790 24870 -8670
rect 24990 -8790 25035 -8670
rect 25155 -8790 25200 -8670
rect 25320 -8790 25365 -8670
rect 25485 -8790 25540 -8670
rect 25660 -8790 25705 -8670
rect 25825 -8790 25870 -8670
rect 25990 -8790 26035 -8670
rect 26155 -8790 26210 -8670
rect 26330 -8790 26375 -8670
rect 26495 -8790 26540 -8670
rect 26660 -8790 26705 -8670
rect 26825 -8790 26880 -8670
rect 27000 -8790 27045 -8670
rect 27165 -8790 27210 -8670
rect 27330 -8790 27375 -8670
rect 27495 -8790 27550 -8670
rect 27670 -8790 27715 -8670
rect 27835 -8790 27880 -8670
rect 28000 -8790 28045 -8670
rect 28165 -8790 28220 -8670
rect 28340 -8790 28385 -8670
rect 28505 -8790 28550 -8670
rect 28670 -8790 28715 -8670
rect 28835 -8790 28890 -8670
rect 29010 -8790 29055 -8670
rect 29175 -8790 29220 -8670
rect 29340 -8790 29385 -8670
rect 29505 -8790 29560 -8670
rect 29680 -8790 29705 -8670
rect 24175 -8835 29705 -8790
rect 24175 -8955 24200 -8835
rect 24320 -8955 24365 -8835
rect 24485 -8955 24530 -8835
rect 24650 -8955 24695 -8835
rect 24815 -8955 24870 -8835
rect 24990 -8955 25035 -8835
rect 25155 -8955 25200 -8835
rect 25320 -8955 25365 -8835
rect 25485 -8955 25540 -8835
rect 25660 -8955 25705 -8835
rect 25825 -8955 25870 -8835
rect 25990 -8955 26035 -8835
rect 26155 -8955 26210 -8835
rect 26330 -8955 26375 -8835
rect 26495 -8955 26540 -8835
rect 26660 -8955 26705 -8835
rect 26825 -8955 26880 -8835
rect 27000 -8955 27045 -8835
rect 27165 -8955 27210 -8835
rect 27330 -8955 27375 -8835
rect 27495 -8955 27550 -8835
rect 27670 -8955 27715 -8835
rect 27835 -8955 27880 -8835
rect 28000 -8955 28045 -8835
rect 28165 -8955 28220 -8835
rect 28340 -8955 28385 -8835
rect 28505 -8955 28550 -8835
rect 28670 -8955 28715 -8835
rect 28835 -8955 28890 -8835
rect 29010 -8955 29055 -8835
rect 29175 -8955 29220 -8835
rect 29340 -8955 29385 -8835
rect 29505 -8955 29560 -8835
rect 29680 -8955 29705 -8835
rect 24175 -9000 29705 -8955
rect 24175 -9120 24200 -9000
rect 24320 -9120 24365 -9000
rect 24485 -9120 24530 -9000
rect 24650 -9120 24695 -9000
rect 24815 -9120 24870 -9000
rect 24990 -9120 25035 -9000
rect 25155 -9120 25200 -9000
rect 25320 -9120 25365 -9000
rect 25485 -9120 25540 -9000
rect 25660 -9120 25705 -9000
rect 25825 -9120 25870 -9000
rect 25990 -9120 26035 -9000
rect 26155 -9120 26210 -9000
rect 26330 -9120 26375 -9000
rect 26495 -9120 26540 -9000
rect 26660 -9120 26705 -9000
rect 26825 -9120 26880 -9000
rect 27000 -9120 27045 -9000
rect 27165 -9120 27210 -9000
rect 27330 -9120 27375 -9000
rect 27495 -9120 27550 -9000
rect 27670 -9120 27715 -9000
rect 27835 -9120 27880 -9000
rect 28000 -9120 28045 -9000
rect 28165 -9120 28220 -9000
rect 28340 -9120 28385 -9000
rect 28505 -9120 28550 -9000
rect 28670 -9120 28715 -9000
rect 28835 -9120 28890 -9000
rect 29010 -9120 29055 -9000
rect 29175 -9120 29220 -9000
rect 29340 -9120 29385 -9000
rect 29505 -9120 29560 -9000
rect 29680 -9120 29705 -9000
rect 24175 -9175 29705 -9120
rect 24175 -9295 24200 -9175
rect 24320 -9295 24365 -9175
rect 24485 -9295 24530 -9175
rect 24650 -9295 24695 -9175
rect 24815 -9295 24870 -9175
rect 24990 -9295 25035 -9175
rect 25155 -9295 25200 -9175
rect 25320 -9295 25365 -9175
rect 25485 -9295 25540 -9175
rect 25660 -9295 25705 -9175
rect 25825 -9295 25870 -9175
rect 25990 -9295 26035 -9175
rect 26155 -9295 26210 -9175
rect 26330 -9295 26375 -9175
rect 26495 -9295 26540 -9175
rect 26660 -9295 26705 -9175
rect 26825 -9295 26880 -9175
rect 27000 -9295 27045 -9175
rect 27165 -9295 27210 -9175
rect 27330 -9295 27375 -9175
rect 27495 -9295 27550 -9175
rect 27670 -9295 27715 -9175
rect 27835 -9295 27880 -9175
rect 28000 -9295 28045 -9175
rect 28165 -9295 28220 -9175
rect 28340 -9295 28385 -9175
rect 28505 -9295 28550 -9175
rect 28670 -9295 28715 -9175
rect 28835 -9295 28890 -9175
rect 29010 -9295 29055 -9175
rect 29175 -9295 29220 -9175
rect 29340 -9295 29385 -9175
rect 29505 -9295 29560 -9175
rect 29680 -9295 29705 -9175
rect 24175 -9340 29705 -9295
rect 24175 -9460 24200 -9340
rect 24320 -9460 24365 -9340
rect 24485 -9460 24530 -9340
rect 24650 -9460 24695 -9340
rect 24815 -9460 24870 -9340
rect 24990 -9460 25035 -9340
rect 25155 -9460 25200 -9340
rect 25320 -9460 25365 -9340
rect 25485 -9460 25540 -9340
rect 25660 -9460 25705 -9340
rect 25825 -9460 25870 -9340
rect 25990 -9460 26035 -9340
rect 26155 -9460 26210 -9340
rect 26330 -9460 26375 -9340
rect 26495 -9460 26540 -9340
rect 26660 -9460 26705 -9340
rect 26825 -9460 26880 -9340
rect 27000 -9460 27045 -9340
rect 27165 -9460 27210 -9340
rect 27330 -9460 27375 -9340
rect 27495 -9460 27550 -9340
rect 27670 -9460 27715 -9340
rect 27835 -9460 27880 -9340
rect 28000 -9460 28045 -9340
rect 28165 -9460 28220 -9340
rect 28340 -9460 28385 -9340
rect 28505 -9460 28550 -9340
rect 28670 -9460 28715 -9340
rect 28835 -9460 28890 -9340
rect 29010 -9460 29055 -9340
rect 29175 -9460 29220 -9340
rect 29340 -9460 29385 -9340
rect 29505 -9460 29560 -9340
rect 29680 -9460 29705 -9340
rect 24175 -9505 29705 -9460
rect 24175 -9625 24200 -9505
rect 24320 -9625 24365 -9505
rect 24485 -9625 24530 -9505
rect 24650 -9625 24695 -9505
rect 24815 -9625 24870 -9505
rect 24990 -9625 25035 -9505
rect 25155 -9625 25200 -9505
rect 25320 -9625 25365 -9505
rect 25485 -9625 25540 -9505
rect 25660 -9625 25705 -9505
rect 25825 -9625 25870 -9505
rect 25990 -9625 26035 -9505
rect 26155 -9625 26210 -9505
rect 26330 -9625 26375 -9505
rect 26495 -9625 26540 -9505
rect 26660 -9625 26705 -9505
rect 26825 -9625 26880 -9505
rect 27000 -9625 27045 -9505
rect 27165 -9625 27210 -9505
rect 27330 -9625 27375 -9505
rect 27495 -9625 27550 -9505
rect 27670 -9625 27715 -9505
rect 27835 -9625 27880 -9505
rect 28000 -9625 28045 -9505
rect 28165 -9625 28220 -9505
rect 28340 -9625 28385 -9505
rect 28505 -9625 28550 -9505
rect 28670 -9625 28715 -9505
rect 28835 -9625 28890 -9505
rect 29010 -9625 29055 -9505
rect 29175 -9625 29220 -9505
rect 29340 -9625 29385 -9505
rect 29505 -9625 29560 -9505
rect 29680 -9625 29705 -9505
rect 24175 -9670 29705 -9625
rect 24175 -9790 24200 -9670
rect 24320 -9790 24365 -9670
rect 24485 -9790 24530 -9670
rect 24650 -9790 24695 -9670
rect 24815 -9790 24870 -9670
rect 24990 -9790 25035 -9670
rect 25155 -9790 25200 -9670
rect 25320 -9790 25365 -9670
rect 25485 -9790 25540 -9670
rect 25660 -9790 25705 -9670
rect 25825 -9790 25870 -9670
rect 25990 -9790 26035 -9670
rect 26155 -9790 26210 -9670
rect 26330 -9790 26375 -9670
rect 26495 -9790 26540 -9670
rect 26660 -9790 26705 -9670
rect 26825 -9790 26880 -9670
rect 27000 -9790 27045 -9670
rect 27165 -9790 27210 -9670
rect 27330 -9790 27375 -9670
rect 27495 -9790 27550 -9670
rect 27670 -9790 27715 -9670
rect 27835 -9790 27880 -9670
rect 28000 -9790 28045 -9670
rect 28165 -9790 28220 -9670
rect 28340 -9790 28385 -9670
rect 28505 -9790 28550 -9670
rect 28670 -9790 28715 -9670
rect 28835 -9790 28890 -9670
rect 29010 -9790 29055 -9670
rect 29175 -9790 29220 -9670
rect 29340 -9790 29385 -9670
rect 29505 -9790 29560 -9670
rect 29680 -9790 29705 -9670
rect 24175 -9860 29705 -9790
rect 7105 -9880 29705 -9860
rect 7105 -10000 7170 -9880
rect 7290 -10000 7335 -9880
rect 7455 -10000 7500 -9880
rect 7620 -10000 7665 -9880
rect 7785 -10000 7830 -9880
rect 7950 -10000 7995 -9880
rect 8115 -10000 8160 -9880
rect 8280 -10000 8325 -9880
rect 8445 -10000 8490 -9880
rect 8610 -10000 8655 -9880
rect 8775 -10000 8820 -9880
rect 8940 -10000 8985 -9880
rect 9105 -10000 9150 -9880
rect 9270 -10000 9315 -9880
rect 9435 -10000 9480 -9880
rect 9600 -10000 9645 -9880
rect 9765 -10000 9810 -9880
rect 9930 -10000 9975 -9880
rect 10095 -10000 10140 -9880
rect 10260 -10000 10305 -9880
rect 10425 -10000 10470 -9880
rect 10590 -10000 10635 -9880
rect 10755 -10000 10800 -9880
rect 10920 -10000 10965 -9880
rect 11085 -10000 11130 -9880
rect 11250 -10000 11295 -9880
rect 11415 -10000 11460 -9880
rect 11580 -10000 11625 -9880
rect 11745 -10000 11790 -9880
rect 11910 -10000 11955 -9880
rect 12075 -10000 12120 -9880
rect 12240 -10000 12285 -9880
rect 12405 -10000 12450 -9880
rect 12570 -10000 12860 -9880
rect 12980 -10000 13025 -9880
rect 13145 -10000 13190 -9880
rect 13310 -10000 13355 -9880
rect 13475 -10000 13520 -9880
rect 13640 -10000 13685 -9880
rect 13805 -10000 13850 -9880
rect 13970 -10000 14015 -9880
rect 14135 -10000 14180 -9880
rect 14300 -10000 14345 -9880
rect 14465 -10000 14510 -9880
rect 14630 -10000 14675 -9880
rect 14795 -10000 14840 -9880
rect 14960 -10000 15005 -9880
rect 15125 -10000 15170 -9880
rect 15290 -10000 15335 -9880
rect 15455 -10000 15500 -9880
rect 15620 -10000 15665 -9880
rect 15785 -10000 15830 -9880
rect 15950 -10000 15995 -9880
rect 16115 -10000 16160 -9880
rect 16280 -10000 16325 -9880
rect 16445 -10000 16490 -9880
rect 16610 -10000 16655 -9880
rect 16775 -10000 16820 -9880
rect 16940 -10000 16985 -9880
rect 17105 -10000 17150 -9880
rect 17270 -10000 17315 -9880
rect 17435 -10000 17480 -9880
rect 17600 -10000 17645 -9880
rect 17765 -10000 17810 -9880
rect 17930 -10000 17975 -9880
rect 18095 -10000 18140 -9880
rect 18260 -10000 18550 -9880
rect 18670 -10000 18715 -9880
rect 18835 -10000 18880 -9880
rect 19000 -10000 19045 -9880
rect 19165 -10000 19210 -9880
rect 19330 -10000 19375 -9880
rect 19495 -10000 19540 -9880
rect 19660 -10000 19705 -9880
rect 19825 -10000 19870 -9880
rect 19990 -10000 20035 -9880
rect 20155 -10000 20200 -9880
rect 20320 -10000 20365 -9880
rect 20485 -10000 20530 -9880
rect 20650 -10000 20695 -9880
rect 20815 -10000 20860 -9880
rect 20980 -10000 21025 -9880
rect 21145 -10000 21190 -9880
rect 21310 -10000 21355 -9880
rect 21475 -10000 21520 -9880
rect 21640 -10000 21685 -9880
rect 21805 -10000 21850 -9880
rect 21970 -10000 22015 -9880
rect 22135 -10000 22180 -9880
rect 22300 -10000 22345 -9880
rect 22465 -10000 22510 -9880
rect 22630 -10000 22675 -9880
rect 22795 -10000 22840 -9880
rect 22960 -10000 23005 -9880
rect 23125 -10000 23170 -9880
rect 23290 -10000 23335 -9880
rect 23455 -10000 23500 -9880
rect 23620 -10000 23665 -9880
rect 23785 -10000 23830 -9880
rect 23950 -10000 24240 -9880
rect 24360 -10000 24405 -9880
rect 24525 -10000 24570 -9880
rect 24690 -10000 24735 -9880
rect 24855 -10000 24900 -9880
rect 25020 -10000 25065 -9880
rect 25185 -10000 25230 -9880
rect 25350 -10000 25395 -9880
rect 25515 -10000 25560 -9880
rect 25680 -10000 25725 -9880
rect 25845 -10000 25890 -9880
rect 26010 -10000 26055 -9880
rect 26175 -10000 26220 -9880
rect 26340 -10000 26385 -9880
rect 26505 -10000 26550 -9880
rect 26670 -10000 26715 -9880
rect 26835 -10000 26880 -9880
rect 27000 -10000 27045 -9880
rect 27165 -10000 27210 -9880
rect 27330 -10000 27375 -9880
rect 27495 -10000 27540 -9880
rect 27660 -10000 27705 -9880
rect 27825 -10000 27870 -9880
rect 27990 -10000 28035 -9880
rect 28155 -10000 28200 -9880
rect 28320 -10000 28365 -9880
rect 28485 -10000 28530 -9880
rect 28650 -10000 28695 -9880
rect 28815 -10000 28860 -9880
rect 28980 -10000 29025 -9880
rect 29145 -10000 29190 -9880
rect 29310 -10000 29355 -9880
rect 29475 -10000 29520 -9880
rect 29640 -10000 29705 -9880
rect 7105 -10020 29705 -10000
rect 7105 -10090 12635 -10020
rect 7105 -10210 7130 -10090
rect 7250 -10210 7305 -10090
rect 7425 -10210 7470 -10090
rect 7590 -10210 7635 -10090
rect 7755 -10210 7800 -10090
rect 7920 -10210 7975 -10090
rect 8095 -10210 8140 -10090
rect 8260 -10210 8305 -10090
rect 8425 -10210 8470 -10090
rect 8590 -10210 8645 -10090
rect 8765 -10210 8810 -10090
rect 8930 -10210 8975 -10090
rect 9095 -10210 9140 -10090
rect 9260 -10210 9315 -10090
rect 9435 -10210 9480 -10090
rect 9600 -10210 9645 -10090
rect 9765 -10210 9810 -10090
rect 9930 -10210 9985 -10090
rect 10105 -10210 10150 -10090
rect 10270 -10210 10315 -10090
rect 10435 -10210 10480 -10090
rect 10600 -10210 10655 -10090
rect 10775 -10210 10820 -10090
rect 10940 -10210 10985 -10090
rect 11105 -10210 11150 -10090
rect 11270 -10210 11325 -10090
rect 11445 -10210 11490 -10090
rect 11610 -10210 11655 -10090
rect 11775 -10210 11820 -10090
rect 11940 -10210 11995 -10090
rect 12115 -10210 12160 -10090
rect 12280 -10210 12325 -10090
rect 12445 -10210 12490 -10090
rect 12610 -10210 12635 -10090
rect 7105 -10255 12635 -10210
rect 7105 -10375 7130 -10255
rect 7250 -10375 7305 -10255
rect 7425 -10375 7470 -10255
rect 7590 -10375 7635 -10255
rect 7755 -10375 7800 -10255
rect 7920 -10375 7975 -10255
rect 8095 -10375 8140 -10255
rect 8260 -10375 8305 -10255
rect 8425 -10375 8470 -10255
rect 8590 -10375 8645 -10255
rect 8765 -10375 8810 -10255
rect 8930 -10375 8975 -10255
rect 9095 -10375 9140 -10255
rect 9260 -10375 9315 -10255
rect 9435 -10375 9480 -10255
rect 9600 -10375 9645 -10255
rect 9765 -10375 9810 -10255
rect 9930 -10375 9985 -10255
rect 10105 -10375 10150 -10255
rect 10270 -10375 10315 -10255
rect 10435 -10375 10480 -10255
rect 10600 -10375 10655 -10255
rect 10775 -10375 10820 -10255
rect 10940 -10375 10985 -10255
rect 11105 -10375 11150 -10255
rect 11270 -10375 11325 -10255
rect 11445 -10375 11490 -10255
rect 11610 -10375 11655 -10255
rect 11775 -10375 11820 -10255
rect 11940 -10375 11995 -10255
rect 12115 -10375 12160 -10255
rect 12280 -10375 12325 -10255
rect 12445 -10375 12490 -10255
rect 12610 -10375 12635 -10255
rect 7105 -10420 12635 -10375
rect 7105 -10540 7130 -10420
rect 7250 -10540 7305 -10420
rect 7425 -10540 7470 -10420
rect 7590 -10540 7635 -10420
rect 7755 -10540 7800 -10420
rect 7920 -10540 7975 -10420
rect 8095 -10540 8140 -10420
rect 8260 -10540 8305 -10420
rect 8425 -10540 8470 -10420
rect 8590 -10540 8645 -10420
rect 8765 -10540 8810 -10420
rect 8930 -10540 8975 -10420
rect 9095 -10540 9140 -10420
rect 9260 -10540 9315 -10420
rect 9435 -10540 9480 -10420
rect 9600 -10540 9645 -10420
rect 9765 -10540 9810 -10420
rect 9930 -10540 9985 -10420
rect 10105 -10540 10150 -10420
rect 10270 -10540 10315 -10420
rect 10435 -10540 10480 -10420
rect 10600 -10540 10655 -10420
rect 10775 -10540 10820 -10420
rect 10940 -10540 10985 -10420
rect 11105 -10540 11150 -10420
rect 11270 -10540 11325 -10420
rect 11445 -10540 11490 -10420
rect 11610 -10540 11655 -10420
rect 11775 -10540 11820 -10420
rect 11940 -10540 11995 -10420
rect 12115 -10540 12160 -10420
rect 12280 -10540 12325 -10420
rect 12445 -10540 12490 -10420
rect 12610 -10540 12635 -10420
rect 7105 -10585 12635 -10540
rect 7105 -10705 7130 -10585
rect 7250 -10705 7305 -10585
rect 7425 -10705 7470 -10585
rect 7590 -10705 7635 -10585
rect 7755 -10705 7800 -10585
rect 7920 -10705 7975 -10585
rect 8095 -10705 8140 -10585
rect 8260 -10705 8305 -10585
rect 8425 -10705 8470 -10585
rect 8590 -10705 8645 -10585
rect 8765 -10705 8810 -10585
rect 8930 -10705 8975 -10585
rect 9095 -10705 9140 -10585
rect 9260 -10705 9315 -10585
rect 9435 -10705 9480 -10585
rect 9600 -10705 9645 -10585
rect 9765 -10705 9810 -10585
rect 9930 -10705 9985 -10585
rect 10105 -10705 10150 -10585
rect 10270 -10705 10315 -10585
rect 10435 -10705 10480 -10585
rect 10600 -10705 10655 -10585
rect 10775 -10705 10820 -10585
rect 10940 -10705 10985 -10585
rect 11105 -10705 11150 -10585
rect 11270 -10705 11325 -10585
rect 11445 -10705 11490 -10585
rect 11610 -10705 11655 -10585
rect 11775 -10705 11820 -10585
rect 11940 -10705 11995 -10585
rect 12115 -10705 12160 -10585
rect 12280 -10705 12325 -10585
rect 12445 -10705 12490 -10585
rect 12610 -10705 12635 -10585
rect 7105 -10760 12635 -10705
rect 7105 -10880 7130 -10760
rect 7250 -10880 7305 -10760
rect 7425 -10880 7470 -10760
rect 7590 -10880 7635 -10760
rect 7755 -10880 7800 -10760
rect 7920 -10880 7975 -10760
rect 8095 -10880 8140 -10760
rect 8260 -10880 8305 -10760
rect 8425 -10880 8470 -10760
rect 8590 -10880 8645 -10760
rect 8765 -10880 8810 -10760
rect 8930 -10880 8975 -10760
rect 9095 -10880 9140 -10760
rect 9260 -10880 9315 -10760
rect 9435 -10880 9480 -10760
rect 9600 -10880 9645 -10760
rect 9765 -10880 9810 -10760
rect 9930 -10880 9985 -10760
rect 10105 -10880 10150 -10760
rect 10270 -10880 10315 -10760
rect 10435 -10880 10480 -10760
rect 10600 -10880 10655 -10760
rect 10775 -10880 10820 -10760
rect 10940 -10880 10985 -10760
rect 11105 -10880 11150 -10760
rect 11270 -10880 11325 -10760
rect 11445 -10880 11490 -10760
rect 11610 -10880 11655 -10760
rect 11775 -10880 11820 -10760
rect 11940 -10880 11995 -10760
rect 12115 -10880 12160 -10760
rect 12280 -10880 12325 -10760
rect 12445 -10880 12490 -10760
rect 12610 -10880 12635 -10760
rect 7105 -10925 12635 -10880
rect 7105 -11045 7130 -10925
rect 7250 -11045 7305 -10925
rect 7425 -11045 7470 -10925
rect 7590 -11045 7635 -10925
rect 7755 -11045 7800 -10925
rect 7920 -11045 7975 -10925
rect 8095 -11045 8140 -10925
rect 8260 -11045 8305 -10925
rect 8425 -11045 8470 -10925
rect 8590 -11045 8645 -10925
rect 8765 -11045 8810 -10925
rect 8930 -11045 8975 -10925
rect 9095 -11045 9140 -10925
rect 9260 -11045 9315 -10925
rect 9435 -11045 9480 -10925
rect 9600 -11045 9645 -10925
rect 9765 -11045 9810 -10925
rect 9930 -11045 9985 -10925
rect 10105 -11045 10150 -10925
rect 10270 -11045 10315 -10925
rect 10435 -11045 10480 -10925
rect 10600 -11045 10655 -10925
rect 10775 -11045 10820 -10925
rect 10940 -11045 10985 -10925
rect 11105 -11045 11150 -10925
rect 11270 -11045 11325 -10925
rect 11445 -11045 11490 -10925
rect 11610 -11045 11655 -10925
rect 11775 -11045 11820 -10925
rect 11940 -11045 11995 -10925
rect 12115 -11045 12160 -10925
rect 12280 -11045 12325 -10925
rect 12445 -11045 12490 -10925
rect 12610 -11045 12635 -10925
rect 7105 -11090 12635 -11045
rect 7105 -11210 7130 -11090
rect 7250 -11210 7305 -11090
rect 7425 -11210 7470 -11090
rect 7590 -11210 7635 -11090
rect 7755 -11210 7800 -11090
rect 7920 -11210 7975 -11090
rect 8095 -11210 8140 -11090
rect 8260 -11210 8305 -11090
rect 8425 -11210 8470 -11090
rect 8590 -11210 8645 -11090
rect 8765 -11210 8810 -11090
rect 8930 -11210 8975 -11090
rect 9095 -11210 9140 -11090
rect 9260 -11210 9315 -11090
rect 9435 -11210 9480 -11090
rect 9600 -11210 9645 -11090
rect 9765 -11210 9810 -11090
rect 9930 -11210 9985 -11090
rect 10105 -11210 10150 -11090
rect 10270 -11210 10315 -11090
rect 10435 -11210 10480 -11090
rect 10600 -11210 10655 -11090
rect 10775 -11210 10820 -11090
rect 10940 -11210 10985 -11090
rect 11105 -11210 11150 -11090
rect 11270 -11210 11325 -11090
rect 11445 -11210 11490 -11090
rect 11610 -11210 11655 -11090
rect 11775 -11210 11820 -11090
rect 11940 -11210 11995 -11090
rect 12115 -11210 12160 -11090
rect 12280 -11210 12325 -11090
rect 12445 -11210 12490 -11090
rect 12610 -11210 12635 -11090
rect 7105 -11255 12635 -11210
rect 7105 -11375 7130 -11255
rect 7250 -11375 7305 -11255
rect 7425 -11375 7470 -11255
rect 7590 -11375 7635 -11255
rect 7755 -11375 7800 -11255
rect 7920 -11375 7975 -11255
rect 8095 -11375 8140 -11255
rect 8260 -11375 8305 -11255
rect 8425 -11375 8470 -11255
rect 8590 -11375 8645 -11255
rect 8765 -11375 8810 -11255
rect 8930 -11375 8975 -11255
rect 9095 -11375 9140 -11255
rect 9260 -11375 9315 -11255
rect 9435 -11375 9480 -11255
rect 9600 -11375 9645 -11255
rect 9765 -11375 9810 -11255
rect 9930 -11375 9985 -11255
rect 10105 -11375 10150 -11255
rect 10270 -11375 10315 -11255
rect 10435 -11375 10480 -11255
rect 10600 -11375 10655 -11255
rect 10775 -11375 10820 -11255
rect 10940 -11375 10985 -11255
rect 11105 -11375 11150 -11255
rect 11270 -11375 11325 -11255
rect 11445 -11375 11490 -11255
rect 11610 -11375 11655 -11255
rect 11775 -11375 11820 -11255
rect 11940 -11375 11995 -11255
rect 12115 -11375 12160 -11255
rect 12280 -11375 12325 -11255
rect 12445 -11375 12490 -11255
rect 12610 -11375 12635 -11255
rect 7105 -11430 12635 -11375
rect 7105 -11550 7130 -11430
rect 7250 -11550 7305 -11430
rect 7425 -11550 7470 -11430
rect 7590 -11550 7635 -11430
rect 7755 -11550 7800 -11430
rect 7920 -11550 7975 -11430
rect 8095 -11550 8140 -11430
rect 8260 -11550 8305 -11430
rect 8425 -11550 8470 -11430
rect 8590 -11550 8645 -11430
rect 8765 -11550 8810 -11430
rect 8930 -11550 8975 -11430
rect 9095 -11550 9140 -11430
rect 9260 -11550 9315 -11430
rect 9435 -11550 9480 -11430
rect 9600 -11550 9645 -11430
rect 9765 -11550 9810 -11430
rect 9930 -11550 9985 -11430
rect 10105 -11550 10150 -11430
rect 10270 -11550 10315 -11430
rect 10435 -11550 10480 -11430
rect 10600 -11550 10655 -11430
rect 10775 -11550 10820 -11430
rect 10940 -11550 10985 -11430
rect 11105 -11550 11150 -11430
rect 11270 -11550 11325 -11430
rect 11445 -11550 11490 -11430
rect 11610 -11550 11655 -11430
rect 11775 -11550 11820 -11430
rect 11940 -11550 11995 -11430
rect 12115 -11550 12160 -11430
rect 12280 -11550 12325 -11430
rect 12445 -11550 12490 -11430
rect 12610 -11550 12635 -11430
rect 7105 -11595 12635 -11550
rect 7105 -11715 7130 -11595
rect 7250 -11715 7305 -11595
rect 7425 -11715 7470 -11595
rect 7590 -11715 7635 -11595
rect 7755 -11715 7800 -11595
rect 7920 -11715 7975 -11595
rect 8095 -11715 8140 -11595
rect 8260 -11715 8305 -11595
rect 8425 -11715 8470 -11595
rect 8590 -11715 8645 -11595
rect 8765 -11715 8810 -11595
rect 8930 -11715 8975 -11595
rect 9095 -11715 9140 -11595
rect 9260 -11715 9315 -11595
rect 9435 -11715 9480 -11595
rect 9600 -11715 9645 -11595
rect 9765 -11715 9810 -11595
rect 9930 -11715 9985 -11595
rect 10105 -11715 10150 -11595
rect 10270 -11715 10315 -11595
rect 10435 -11715 10480 -11595
rect 10600 -11715 10655 -11595
rect 10775 -11715 10820 -11595
rect 10940 -11715 10985 -11595
rect 11105 -11715 11150 -11595
rect 11270 -11715 11325 -11595
rect 11445 -11715 11490 -11595
rect 11610 -11715 11655 -11595
rect 11775 -11715 11820 -11595
rect 11940 -11715 11995 -11595
rect 12115 -11715 12160 -11595
rect 12280 -11715 12325 -11595
rect 12445 -11715 12490 -11595
rect 12610 -11715 12635 -11595
rect 7105 -11760 12635 -11715
rect 7105 -11880 7130 -11760
rect 7250 -11880 7305 -11760
rect 7425 -11880 7470 -11760
rect 7590 -11880 7635 -11760
rect 7755 -11880 7800 -11760
rect 7920 -11880 7975 -11760
rect 8095 -11880 8140 -11760
rect 8260 -11880 8305 -11760
rect 8425 -11880 8470 -11760
rect 8590 -11880 8645 -11760
rect 8765 -11880 8810 -11760
rect 8930 -11880 8975 -11760
rect 9095 -11880 9140 -11760
rect 9260 -11880 9315 -11760
rect 9435 -11880 9480 -11760
rect 9600 -11880 9645 -11760
rect 9765 -11880 9810 -11760
rect 9930 -11880 9985 -11760
rect 10105 -11880 10150 -11760
rect 10270 -11880 10315 -11760
rect 10435 -11880 10480 -11760
rect 10600 -11880 10655 -11760
rect 10775 -11880 10820 -11760
rect 10940 -11880 10985 -11760
rect 11105 -11880 11150 -11760
rect 11270 -11880 11325 -11760
rect 11445 -11880 11490 -11760
rect 11610 -11880 11655 -11760
rect 11775 -11880 11820 -11760
rect 11940 -11880 11995 -11760
rect 12115 -11880 12160 -11760
rect 12280 -11880 12325 -11760
rect 12445 -11880 12490 -11760
rect 12610 -11880 12635 -11760
rect 7105 -11925 12635 -11880
rect 7105 -12045 7130 -11925
rect 7250 -12045 7305 -11925
rect 7425 -12045 7470 -11925
rect 7590 -12045 7635 -11925
rect 7755 -12045 7800 -11925
rect 7920 -12045 7975 -11925
rect 8095 -12045 8140 -11925
rect 8260 -12045 8305 -11925
rect 8425 -12045 8470 -11925
rect 8590 -12045 8645 -11925
rect 8765 -12045 8810 -11925
rect 8930 -12045 8975 -11925
rect 9095 -12045 9140 -11925
rect 9260 -12045 9315 -11925
rect 9435 -12045 9480 -11925
rect 9600 -12045 9645 -11925
rect 9765 -12045 9810 -11925
rect 9930 -12045 9985 -11925
rect 10105 -12045 10150 -11925
rect 10270 -12045 10315 -11925
rect 10435 -12045 10480 -11925
rect 10600 -12045 10655 -11925
rect 10775 -12045 10820 -11925
rect 10940 -12045 10985 -11925
rect 11105 -12045 11150 -11925
rect 11270 -12045 11325 -11925
rect 11445 -12045 11490 -11925
rect 11610 -12045 11655 -11925
rect 11775 -12045 11820 -11925
rect 11940 -12045 11995 -11925
rect 12115 -12045 12160 -11925
rect 12280 -12045 12325 -11925
rect 12445 -12045 12490 -11925
rect 12610 -12045 12635 -11925
rect 7105 -12100 12635 -12045
rect 7105 -12220 7130 -12100
rect 7250 -12220 7305 -12100
rect 7425 -12220 7470 -12100
rect 7590 -12220 7635 -12100
rect 7755 -12220 7800 -12100
rect 7920 -12220 7975 -12100
rect 8095 -12220 8140 -12100
rect 8260 -12220 8305 -12100
rect 8425 -12220 8470 -12100
rect 8590 -12220 8645 -12100
rect 8765 -12220 8810 -12100
rect 8930 -12220 8975 -12100
rect 9095 -12220 9140 -12100
rect 9260 -12220 9315 -12100
rect 9435 -12220 9480 -12100
rect 9600 -12220 9645 -12100
rect 9765 -12220 9810 -12100
rect 9930 -12220 9985 -12100
rect 10105 -12220 10150 -12100
rect 10270 -12220 10315 -12100
rect 10435 -12220 10480 -12100
rect 10600 -12220 10655 -12100
rect 10775 -12220 10820 -12100
rect 10940 -12220 10985 -12100
rect 11105 -12220 11150 -12100
rect 11270 -12220 11325 -12100
rect 11445 -12220 11490 -12100
rect 11610 -12220 11655 -12100
rect 11775 -12220 11820 -12100
rect 11940 -12220 11995 -12100
rect 12115 -12220 12160 -12100
rect 12280 -12220 12325 -12100
rect 12445 -12220 12490 -12100
rect 12610 -12220 12635 -12100
rect 7105 -12265 12635 -12220
rect 7105 -12385 7130 -12265
rect 7250 -12385 7305 -12265
rect 7425 -12385 7470 -12265
rect 7590 -12385 7635 -12265
rect 7755 -12385 7800 -12265
rect 7920 -12385 7975 -12265
rect 8095 -12385 8140 -12265
rect 8260 -12385 8305 -12265
rect 8425 -12385 8470 -12265
rect 8590 -12385 8645 -12265
rect 8765 -12385 8810 -12265
rect 8930 -12385 8975 -12265
rect 9095 -12385 9140 -12265
rect 9260 -12385 9315 -12265
rect 9435 -12385 9480 -12265
rect 9600 -12385 9645 -12265
rect 9765 -12385 9810 -12265
rect 9930 -12385 9985 -12265
rect 10105 -12385 10150 -12265
rect 10270 -12385 10315 -12265
rect 10435 -12385 10480 -12265
rect 10600 -12385 10655 -12265
rect 10775 -12385 10820 -12265
rect 10940 -12385 10985 -12265
rect 11105 -12385 11150 -12265
rect 11270 -12385 11325 -12265
rect 11445 -12385 11490 -12265
rect 11610 -12385 11655 -12265
rect 11775 -12385 11820 -12265
rect 11940 -12385 11995 -12265
rect 12115 -12385 12160 -12265
rect 12280 -12385 12325 -12265
rect 12445 -12385 12490 -12265
rect 12610 -12385 12635 -12265
rect 7105 -12430 12635 -12385
rect 7105 -12550 7130 -12430
rect 7250 -12550 7305 -12430
rect 7425 -12550 7470 -12430
rect 7590 -12550 7635 -12430
rect 7755 -12550 7800 -12430
rect 7920 -12550 7975 -12430
rect 8095 -12550 8140 -12430
rect 8260 -12550 8305 -12430
rect 8425 -12550 8470 -12430
rect 8590 -12550 8645 -12430
rect 8765 -12550 8810 -12430
rect 8930 -12550 8975 -12430
rect 9095 -12550 9140 -12430
rect 9260 -12550 9315 -12430
rect 9435 -12550 9480 -12430
rect 9600 -12550 9645 -12430
rect 9765 -12550 9810 -12430
rect 9930 -12550 9985 -12430
rect 10105 -12550 10150 -12430
rect 10270 -12550 10315 -12430
rect 10435 -12550 10480 -12430
rect 10600 -12550 10655 -12430
rect 10775 -12550 10820 -12430
rect 10940 -12550 10985 -12430
rect 11105 -12550 11150 -12430
rect 11270 -12550 11325 -12430
rect 11445 -12550 11490 -12430
rect 11610 -12550 11655 -12430
rect 11775 -12550 11820 -12430
rect 11940 -12550 11995 -12430
rect 12115 -12550 12160 -12430
rect 12280 -12550 12325 -12430
rect 12445 -12550 12490 -12430
rect 12610 -12550 12635 -12430
rect 7105 -12595 12635 -12550
rect 7105 -12715 7130 -12595
rect 7250 -12715 7305 -12595
rect 7425 -12715 7470 -12595
rect 7590 -12715 7635 -12595
rect 7755 -12715 7800 -12595
rect 7920 -12715 7975 -12595
rect 8095 -12715 8140 -12595
rect 8260 -12715 8305 -12595
rect 8425 -12715 8470 -12595
rect 8590 -12715 8645 -12595
rect 8765 -12715 8810 -12595
rect 8930 -12715 8975 -12595
rect 9095 -12715 9140 -12595
rect 9260 -12715 9315 -12595
rect 9435 -12715 9480 -12595
rect 9600 -12715 9645 -12595
rect 9765 -12715 9810 -12595
rect 9930 -12715 9985 -12595
rect 10105 -12715 10150 -12595
rect 10270 -12715 10315 -12595
rect 10435 -12715 10480 -12595
rect 10600 -12715 10655 -12595
rect 10775 -12715 10820 -12595
rect 10940 -12715 10985 -12595
rect 11105 -12715 11150 -12595
rect 11270 -12715 11325 -12595
rect 11445 -12715 11490 -12595
rect 11610 -12715 11655 -12595
rect 11775 -12715 11820 -12595
rect 11940 -12715 11995 -12595
rect 12115 -12715 12160 -12595
rect 12280 -12715 12325 -12595
rect 12445 -12715 12490 -12595
rect 12610 -12715 12635 -12595
rect 7105 -12770 12635 -12715
rect 7105 -12890 7130 -12770
rect 7250 -12890 7305 -12770
rect 7425 -12890 7470 -12770
rect 7590 -12890 7635 -12770
rect 7755 -12890 7800 -12770
rect 7920 -12890 7975 -12770
rect 8095 -12890 8140 -12770
rect 8260 -12890 8305 -12770
rect 8425 -12890 8470 -12770
rect 8590 -12890 8645 -12770
rect 8765 -12890 8810 -12770
rect 8930 -12890 8975 -12770
rect 9095 -12890 9140 -12770
rect 9260 -12890 9315 -12770
rect 9435 -12890 9480 -12770
rect 9600 -12890 9645 -12770
rect 9765 -12890 9810 -12770
rect 9930 -12890 9985 -12770
rect 10105 -12890 10150 -12770
rect 10270 -12890 10315 -12770
rect 10435 -12890 10480 -12770
rect 10600 -12890 10655 -12770
rect 10775 -12890 10820 -12770
rect 10940 -12890 10985 -12770
rect 11105 -12890 11150 -12770
rect 11270 -12890 11325 -12770
rect 11445 -12890 11490 -12770
rect 11610 -12890 11655 -12770
rect 11775 -12890 11820 -12770
rect 11940 -12890 11995 -12770
rect 12115 -12890 12160 -12770
rect 12280 -12890 12325 -12770
rect 12445 -12890 12490 -12770
rect 12610 -12890 12635 -12770
rect 7105 -12935 12635 -12890
rect 7105 -13055 7130 -12935
rect 7250 -13055 7305 -12935
rect 7425 -13055 7470 -12935
rect 7590 -13055 7635 -12935
rect 7755 -13055 7800 -12935
rect 7920 -13055 7975 -12935
rect 8095 -13055 8140 -12935
rect 8260 -13055 8305 -12935
rect 8425 -13055 8470 -12935
rect 8590 -13055 8645 -12935
rect 8765 -13055 8810 -12935
rect 8930 -13055 8975 -12935
rect 9095 -13055 9140 -12935
rect 9260 -13055 9315 -12935
rect 9435 -13055 9480 -12935
rect 9600 -13055 9645 -12935
rect 9765 -13055 9810 -12935
rect 9930 -13055 9985 -12935
rect 10105 -13055 10150 -12935
rect 10270 -13055 10315 -12935
rect 10435 -13055 10480 -12935
rect 10600 -13055 10655 -12935
rect 10775 -13055 10820 -12935
rect 10940 -13055 10985 -12935
rect 11105 -13055 11150 -12935
rect 11270 -13055 11325 -12935
rect 11445 -13055 11490 -12935
rect 11610 -13055 11655 -12935
rect 11775 -13055 11820 -12935
rect 11940 -13055 11995 -12935
rect 12115 -13055 12160 -12935
rect 12280 -13055 12325 -12935
rect 12445 -13055 12490 -12935
rect 12610 -13055 12635 -12935
rect 7105 -13100 12635 -13055
rect 7105 -13220 7130 -13100
rect 7250 -13220 7305 -13100
rect 7425 -13220 7470 -13100
rect 7590 -13220 7635 -13100
rect 7755 -13220 7800 -13100
rect 7920 -13220 7975 -13100
rect 8095 -13220 8140 -13100
rect 8260 -13220 8305 -13100
rect 8425 -13220 8470 -13100
rect 8590 -13220 8645 -13100
rect 8765 -13220 8810 -13100
rect 8930 -13220 8975 -13100
rect 9095 -13220 9140 -13100
rect 9260 -13220 9315 -13100
rect 9435 -13220 9480 -13100
rect 9600 -13220 9645 -13100
rect 9765 -13220 9810 -13100
rect 9930 -13220 9985 -13100
rect 10105 -13220 10150 -13100
rect 10270 -13220 10315 -13100
rect 10435 -13220 10480 -13100
rect 10600 -13220 10655 -13100
rect 10775 -13220 10820 -13100
rect 10940 -13220 10985 -13100
rect 11105 -13220 11150 -13100
rect 11270 -13220 11325 -13100
rect 11445 -13220 11490 -13100
rect 11610 -13220 11655 -13100
rect 11775 -13220 11820 -13100
rect 11940 -13220 11995 -13100
rect 12115 -13220 12160 -13100
rect 12280 -13220 12325 -13100
rect 12445 -13220 12490 -13100
rect 12610 -13220 12635 -13100
rect 7105 -13265 12635 -13220
rect 7105 -13385 7130 -13265
rect 7250 -13385 7305 -13265
rect 7425 -13385 7470 -13265
rect 7590 -13385 7635 -13265
rect 7755 -13385 7800 -13265
rect 7920 -13385 7975 -13265
rect 8095 -13385 8140 -13265
rect 8260 -13385 8305 -13265
rect 8425 -13385 8470 -13265
rect 8590 -13385 8645 -13265
rect 8765 -13385 8810 -13265
rect 8930 -13385 8975 -13265
rect 9095 -13385 9140 -13265
rect 9260 -13385 9315 -13265
rect 9435 -13385 9480 -13265
rect 9600 -13385 9645 -13265
rect 9765 -13385 9810 -13265
rect 9930 -13385 9985 -13265
rect 10105 -13385 10150 -13265
rect 10270 -13385 10315 -13265
rect 10435 -13385 10480 -13265
rect 10600 -13385 10655 -13265
rect 10775 -13385 10820 -13265
rect 10940 -13385 10985 -13265
rect 11105 -13385 11150 -13265
rect 11270 -13385 11325 -13265
rect 11445 -13385 11490 -13265
rect 11610 -13385 11655 -13265
rect 11775 -13385 11820 -13265
rect 11940 -13385 11995 -13265
rect 12115 -13385 12160 -13265
rect 12280 -13385 12325 -13265
rect 12445 -13385 12490 -13265
rect 12610 -13385 12635 -13265
rect 7105 -13440 12635 -13385
rect 7105 -13560 7130 -13440
rect 7250 -13560 7305 -13440
rect 7425 -13560 7470 -13440
rect 7590 -13560 7635 -13440
rect 7755 -13560 7800 -13440
rect 7920 -13560 7975 -13440
rect 8095 -13560 8140 -13440
rect 8260 -13560 8305 -13440
rect 8425 -13560 8470 -13440
rect 8590 -13560 8645 -13440
rect 8765 -13560 8810 -13440
rect 8930 -13560 8975 -13440
rect 9095 -13560 9140 -13440
rect 9260 -13560 9315 -13440
rect 9435 -13560 9480 -13440
rect 9600 -13560 9645 -13440
rect 9765 -13560 9810 -13440
rect 9930 -13560 9985 -13440
rect 10105 -13560 10150 -13440
rect 10270 -13560 10315 -13440
rect 10435 -13560 10480 -13440
rect 10600 -13560 10655 -13440
rect 10775 -13560 10820 -13440
rect 10940 -13560 10985 -13440
rect 11105 -13560 11150 -13440
rect 11270 -13560 11325 -13440
rect 11445 -13560 11490 -13440
rect 11610 -13560 11655 -13440
rect 11775 -13560 11820 -13440
rect 11940 -13560 11995 -13440
rect 12115 -13560 12160 -13440
rect 12280 -13560 12325 -13440
rect 12445 -13560 12490 -13440
rect 12610 -13560 12635 -13440
rect 7105 -13605 12635 -13560
rect 7105 -13725 7130 -13605
rect 7250 -13725 7305 -13605
rect 7425 -13725 7470 -13605
rect 7590 -13725 7635 -13605
rect 7755 -13725 7800 -13605
rect 7920 -13725 7975 -13605
rect 8095 -13725 8140 -13605
rect 8260 -13725 8305 -13605
rect 8425 -13725 8470 -13605
rect 8590 -13725 8645 -13605
rect 8765 -13725 8810 -13605
rect 8930 -13725 8975 -13605
rect 9095 -13725 9140 -13605
rect 9260 -13725 9315 -13605
rect 9435 -13725 9480 -13605
rect 9600 -13725 9645 -13605
rect 9765 -13725 9810 -13605
rect 9930 -13725 9985 -13605
rect 10105 -13725 10150 -13605
rect 10270 -13725 10315 -13605
rect 10435 -13725 10480 -13605
rect 10600 -13725 10655 -13605
rect 10775 -13725 10820 -13605
rect 10940 -13725 10985 -13605
rect 11105 -13725 11150 -13605
rect 11270 -13725 11325 -13605
rect 11445 -13725 11490 -13605
rect 11610 -13725 11655 -13605
rect 11775 -13725 11820 -13605
rect 11940 -13725 11995 -13605
rect 12115 -13725 12160 -13605
rect 12280 -13725 12325 -13605
rect 12445 -13725 12490 -13605
rect 12610 -13725 12635 -13605
rect 7105 -13770 12635 -13725
rect 7105 -13890 7130 -13770
rect 7250 -13890 7305 -13770
rect 7425 -13890 7470 -13770
rect 7590 -13890 7635 -13770
rect 7755 -13890 7800 -13770
rect 7920 -13890 7975 -13770
rect 8095 -13890 8140 -13770
rect 8260 -13890 8305 -13770
rect 8425 -13890 8470 -13770
rect 8590 -13890 8645 -13770
rect 8765 -13890 8810 -13770
rect 8930 -13890 8975 -13770
rect 9095 -13890 9140 -13770
rect 9260 -13890 9315 -13770
rect 9435 -13890 9480 -13770
rect 9600 -13890 9645 -13770
rect 9765 -13890 9810 -13770
rect 9930 -13890 9985 -13770
rect 10105 -13890 10150 -13770
rect 10270 -13890 10315 -13770
rect 10435 -13890 10480 -13770
rect 10600 -13890 10655 -13770
rect 10775 -13890 10820 -13770
rect 10940 -13890 10985 -13770
rect 11105 -13890 11150 -13770
rect 11270 -13890 11325 -13770
rect 11445 -13890 11490 -13770
rect 11610 -13890 11655 -13770
rect 11775 -13890 11820 -13770
rect 11940 -13890 11995 -13770
rect 12115 -13890 12160 -13770
rect 12280 -13890 12325 -13770
rect 12445 -13890 12490 -13770
rect 12610 -13890 12635 -13770
rect 7105 -13935 12635 -13890
rect 7105 -14055 7130 -13935
rect 7250 -14055 7305 -13935
rect 7425 -14055 7470 -13935
rect 7590 -14055 7635 -13935
rect 7755 -14055 7800 -13935
rect 7920 -14055 7975 -13935
rect 8095 -14055 8140 -13935
rect 8260 -14055 8305 -13935
rect 8425 -14055 8470 -13935
rect 8590 -14055 8645 -13935
rect 8765 -14055 8810 -13935
rect 8930 -14055 8975 -13935
rect 9095 -14055 9140 -13935
rect 9260 -14055 9315 -13935
rect 9435 -14055 9480 -13935
rect 9600 -14055 9645 -13935
rect 9765 -14055 9810 -13935
rect 9930 -14055 9985 -13935
rect 10105 -14055 10150 -13935
rect 10270 -14055 10315 -13935
rect 10435 -14055 10480 -13935
rect 10600 -14055 10655 -13935
rect 10775 -14055 10820 -13935
rect 10940 -14055 10985 -13935
rect 11105 -14055 11150 -13935
rect 11270 -14055 11325 -13935
rect 11445 -14055 11490 -13935
rect 11610 -14055 11655 -13935
rect 11775 -14055 11820 -13935
rect 11940 -14055 11995 -13935
rect 12115 -14055 12160 -13935
rect 12280 -14055 12325 -13935
rect 12445 -14055 12490 -13935
rect 12610 -14055 12635 -13935
rect 7105 -14110 12635 -14055
rect 7105 -14230 7130 -14110
rect 7250 -14230 7305 -14110
rect 7425 -14230 7470 -14110
rect 7590 -14230 7635 -14110
rect 7755 -14230 7800 -14110
rect 7920 -14230 7975 -14110
rect 8095 -14230 8140 -14110
rect 8260 -14230 8305 -14110
rect 8425 -14230 8470 -14110
rect 8590 -14230 8645 -14110
rect 8765 -14230 8810 -14110
rect 8930 -14230 8975 -14110
rect 9095 -14230 9140 -14110
rect 9260 -14230 9315 -14110
rect 9435 -14230 9480 -14110
rect 9600 -14230 9645 -14110
rect 9765 -14230 9810 -14110
rect 9930 -14230 9985 -14110
rect 10105 -14230 10150 -14110
rect 10270 -14230 10315 -14110
rect 10435 -14230 10480 -14110
rect 10600 -14230 10655 -14110
rect 10775 -14230 10820 -14110
rect 10940 -14230 10985 -14110
rect 11105 -14230 11150 -14110
rect 11270 -14230 11325 -14110
rect 11445 -14230 11490 -14110
rect 11610 -14230 11655 -14110
rect 11775 -14230 11820 -14110
rect 11940 -14230 11995 -14110
rect 12115 -14230 12160 -14110
rect 12280 -14230 12325 -14110
rect 12445 -14230 12490 -14110
rect 12610 -14230 12635 -14110
rect 7105 -14275 12635 -14230
rect 7105 -14395 7130 -14275
rect 7250 -14395 7305 -14275
rect 7425 -14395 7470 -14275
rect 7590 -14395 7635 -14275
rect 7755 -14395 7800 -14275
rect 7920 -14395 7975 -14275
rect 8095 -14395 8140 -14275
rect 8260 -14395 8305 -14275
rect 8425 -14395 8470 -14275
rect 8590 -14395 8645 -14275
rect 8765 -14395 8810 -14275
rect 8930 -14395 8975 -14275
rect 9095 -14395 9140 -14275
rect 9260 -14395 9315 -14275
rect 9435 -14395 9480 -14275
rect 9600 -14395 9645 -14275
rect 9765 -14395 9810 -14275
rect 9930 -14395 9985 -14275
rect 10105 -14395 10150 -14275
rect 10270 -14395 10315 -14275
rect 10435 -14395 10480 -14275
rect 10600 -14395 10655 -14275
rect 10775 -14395 10820 -14275
rect 10940 -14395 10985 -14275
rect 11105 -14395 11150 -14275
rect 11270 -14395 11325 -14275
rect 11445 -14395 11490 -14275
rect 11610 -14395 11655 -14275
rect 11775 -14395 11820 -14275
rect 11940 -14395 11995 -14275
rect 12115 -14395 12160 -14275
rect 12280 -14395 12325 -14275
rect 12445 -14395 12490 -14275
rect 12610 -14395 12635 -14275
rect 7105 -14440 12635 -14395
rect 7105 -14560 7130 -14440
rect 7250 -14560 7305 -14440
rect 7425 -14560 7470 -14440
rect 7590 -14560 7635 -14440
rect 7755 -14560 7800 -14440
rect 7920 -14560 7975 -14440
rect 8095 -14560 8140 -14440
rect 8260 -14560 8305 -14440
rect 8425 -14560 8470 -14440
rect 8590 -14560 8645 -14440
rect 8765 -14560 8810 -14440
rect 8930 -14560 8975 -14440
rect 9095 -14560 9140 -14440
rect 9260 -14560 9315 -14440
rect 9435 -14560 9480 -14440
rect 9600 -14560 9645 -14440
rect 9765 -14560 9810 -14440
rect 9930 -14560 9985 -14440
rect 10105 -14560 10150 -14440
rect 10270 -14560 10315 -14440
rect 10435 -14560 10480 -14440
rect 10600 -14560 10655 -14440
rect 10775 -14560 10820 -14440
rect 10940 -14560 10985 -14440
rect 11105 -14560 11150 -14440
rect 11270 -14560 11325 -14440
rect 11445 -14560 11490 -14440
rect 11610 -14560 11655 -14440
rect 11775 -14560 11820 -14440
rect 11940 -14560 11995 -14440
rect 12115 -14560 12160 -14440
rect 12280 -14560 12325 -14440
rect 12445 -14560 12490 -14440
rect 12610 -14560 12635 -14440
rect 7105 -14605 12635 -14560
rect 7105 -14725 7130 -14605
rect 7250 -14725 7305 -14605
rect 7425 -14725 7470 -14605
rect 7590 -14725 7635 -14605
rect 7755 -14725 7800 -14605
rect 7920 -14725 7975 -14605
rect 8095 -14725 8140 -14605
rect 8260 -14725 8305 -14605
rect 8425 -14725 8470 -14605
rect 8590 -14725 8645 -14605
rect 8765 -14725 8810 -14605
rect 8930 -14725 8975 -14605
rect 9095 -14725 9140 -14605
rect 9260 -14725 9315 -14605
rect 9435 -14725 9480 -14605
rect 9600 -14725 9645 -14605
rect 9765 -14725 9810 -14605
rect 9930 -14725 9985 -14605
rect 10105 -14725 10150 -14605
rect 10270 -14725 10315 -14605
rect 10435 -14725 10480 -14605
rect 10600 -14725 10655 -14605
rect 10775 -14725 10820 -14605
rect 10940 -14725 10985 -14605
rect 11105 -14725 11150 -14605
rect 11270 -14725 11325 -14605
rect 11445 -14725 11490 -14605
rect 11610 -14725 11655 -14605
rect 11775 -14725 11820 -14605
rect 11940 -14725 11995 -14605
rect 12115 -14725 12160 -14605
rect 12280 -14725 12325 -14605
rect 12445 -14725 12490 -14605
rect 12610 -14725 12635 -14605
rect 7105 -14780 12635 -14725
rect 7105 -14900 7130 -14780
rect 7250 -14900 7305 -14780
rect 7425 -14900 7470 -14780
rect 7590 -14900 7635 -14780
rect 7755 -14900 7800 -14780
rect 7920 -14900 7975 -14780
rect 8095 -14900 8140 -14780
rect 8260 -14900 8305 -14780
rect 8425 -14900 8470 -14780
rect 8590 -14900 8645 -14780
rect 8765 -14900 8810 -14780
rect 8930 -14900 8975 -14780
rect 9095 -14900 9140 -14780
rect 9260 -14900 9315 -14780
rect 9435 -14900 9480 -14780
rect 9600 -14900 9645 -14780
rect 9765 -14900 9810 -14780
rect 9930 -14900 9985 -14780
rect 10105 -14900 10150 -14780
rect 10270 -14900 10315 -14780
rect 10435 -14900 10480 -14780
rect 10600 -14900 10655 -14780
rect 10775 -14900 10820 -14780
rect 10940 -14900 10985 -14780
rect 11105 -14900 11150 -14780
rect 11270 -14900 11325 -14780
rect 11445 -14900 11490 -14780
rect 11610 -14900 11655 -14780
rect 11775 -14900 11820 -14780
rect 11940 -14900 11995 -14780
rect 12115 -14900 12160 -14780
rect 12280 -14900 12325 -14780
rect 12445 -14900 12490 -14780
rect 12610 -14900 12635 -14780
rect 7105 -14945 12635 -14900
rect 7105 -15065 7130 -14945
rect 7250 -15065 7305 -14945
rect 7425 -15065 7470 -14945
rect 7590 -15065 7635 -14945
rect 7755 -15065 7800 -14945
rect 7920 -15065 7975 -14945
rect 8095 -15065 8140 -14945
rect 8260 -15065 8305 -14945
rect 8425 -15065 8470 -14945
rect 8590 -15065 8645 -14945
rect 8765 -15065 8810 -14945
rect 8930 -15065 8975 -14945
rect 9095 -15065 9140 -14945
rect 9260 -15065 9315 -14945
rect 9435 -15065 9480 -14945
rect 9600 -15065 9645 -14945
rect 9765 -15065 9810 -14945
rect 9930 -15065 9985 -14945
rect 10105 -15065 10150 -14945
rect 10270 -15065 10315 -14945
rect 10435 -15065 10480 -14945
rect 10600 -15065 10655 -14945
rect 10775 -15065 10820 -14945
rect 10940 -15065 10985 -14945
rect 11105 -15065 11150 -14945
rect 11270 -15065 11325 -14945
rect 11445 -15065 11490 -14945
rect 11610 -15065 11655 -14945
rect 11775 -15065 11820 -14945
rect 11940 -15065 11995 -14945
rect 12115 -15065 12160 -14945
rect 12280 -15065 12325 -14945
rect 12445 -15065 12490 -14945
rect 12610 -15065 12635 -14945
rect 7105 -15110 12635 -15065
rect 7105 -15230 7130 -15110
rect 7250 -15230 7305 -15110
rect 7425 -15230 7470 -15110
rect 7590 -15230 7635 -15110
rect 7755 -15230 7800 -15110
rect 7920 -15230 7975 -15110
rect 8095 -15230 8140 -15110
rect 8260 -15230 8305 -15110
rect 8425 -15230 8470 -15110
rect 8590 -15230 8645 -15110
rect 8765 -15230 8810 -15110
rect 8930 -15230 8975 -15110
rect 9095 -15230 9140 -15110
rect 9260 -15230 9315 -15110
rect 9435 -15230 9480 -15110
rect 9600 -15230 9645 -15110
rect 9765 -15230 9810 -15110
rect 9930 -15230 9985 -15110
rect 10105 -15230 10150 -15110
rect 10270 -15230 10315 -15110
rect 10435 -15230 10480 -15110
rect 10600 -15230 10655 -15110
rect 10775 -15230 10820 -15110
rect 10940 -15230 10985 -15110
rect 11105 -15230 11150 -15110
rect 11270 -15230 11325 -15110
rect 11445 -15230 11490 -15110
rect 11610 -15230 11655 -15110
rect 11775 -15230 11820 -15110
rect 11940 -15230 11995 -15110
rect 12115 -15230 12160 -15110
rect 12280 -15230 12325 -15110
rect 12445 -15230 12490 -15110
rect 12610 -15230 12635 -15110
rect 7105 -15275 12635 -15230
rect 7105 -15395 7130 -15275
rect 7250 -15395 7305 -15275
rect 7425 -15395 7470 -15275
rect 7590 -15395 7635 -15275
rect 7755 -15395 7800 -15275
rect 7920 -15395 7975 -15275
rect 8095 -15395 8140 -15275
rect 8260 -15395 8305 -15275
rect 8425 -15395 8470 -15275
rect 8590 -15395 8645 -15275
rect 8765 -15395 8810 -15275
rect 8930 -15395 8975 -15275
rect 9095 -15395 9140 -15275
rect 9260 -15395 9315 -15275
rect 9435 -15395 9480 -15275
rect 9600 -15395 9645 -15275
rect 9765 -15395 9810 -15275
rect 9930 -15395 9985 -15275
rect 10105 -15395 10150 -15275
rect 10270 -15395 10315 -15275
rect 10435 -15395 10480 -15275
rect 10600 -15395 10655 -15275
rect 10775 -15395 10820 -15275
rect 10940 -15395 10985 -15275
rect 11105 -15395 11150 -15275
rect 11270 -15395 11325 -15275
rect 11445 -15395 11490 -15275
rect 11610 -15395 11655 -15275
rect 11775 -15395 11820 -15275
rect 11940 -15395 11995 -15275
rect 12115 -15395 12160 -15275
rect 12280 -15395 12325 -15275
rect 12445 -15395 12490 -15275
rect 12610 -15395 12635 -15275
rect 7105 -15450 12635 -15395
rect 7105 -15570 7130 -15450
rect 7250 -15570 7305 -15450
rect 7425 -15570 7470 -15450
rect 7590 -15570 7635 -15450
rect 7755 -15570 7800 -15450
rect 7920 -15570 7975 -15450
rect 8095 -15570 8140 -15450
rect 8260 -15570 8305 -15450
rect 8425 -15570 8470 -15450
rect 8590 -15570 8645 -15450
rect 8765 -15570 8810 -15450
rect 8930 -15570 8975 -15450
rect 9095 -15570 9140 -15450
rect 9260 -15570 9315 -15450
rect 9435 -15570 9480 -15450
rect 9600 -15570 9645 -15450
rect 9765 -15570 9810 -15450
rect 9930 -15570 9985 -15450
rect 10105 -15570 10150 -15450
rect 10270 -15570 10315 -15450
rect 10435 -15570 10480 -15450
rect 10600 -15570 10655 -15450
rect 10775 -15570 10820 -15450
rect 10940 -15570 10985 -15450
rect 11105 -15570 11150 -15450
rect 11270 -15570 11325 -15450
rect 11445 -15570 11490 -15450
rect 11610 -15570 11655 -15450
rect 11775 -15570 11820 -15450
rect 11940 -15570 11995 -15450
rect 12115 -15570 12160 -15450
rect 12280 -15570 12325 -15450
rect 12445 -15570 12490 -15450
rect 12610 -15570 12635 -15450
rect 7105 -15595 12635 -15570
rect 12795 -10090 18325 -10020
rect 12795 -10210 12820 -10090
rect 12940 -10210 12995 -10090
rect 13115 -10210 13160 -10090
rect 13280 -10210 13325 -10090
rect 13445 -10210 13490 -10090
rect 13610 -10210 13665 -10090
rect 13785 -10210 13830 -10090
rect 13950 -10210 13995 -10090
rect 14115 -10210 14160 -10090
rect 14280 -10210 14335 -10090
rect 14455 -10210 14500 -10090
rect 14620 -10210 14665 -10090
rect 14785 -10210 14830 -10090
rect 14950 -10210 15005 -10090
rect 15125 -10210 15170 -10090
rect 15290 -10210 15335 -10090
rect 15455 -10210 15500 -10090
rect 15620 -10210 15675 -10090
rect 15795 -10210 15840 -10090
rect 15960 -10210 16005 -10090
rect 16125 -10210 16170 -10090
rect 16290 -10210 16345 -10090
rect 16465 -10210 16510 -10090
rect 16630 -10210 16675 -10090
rect 16795 -10210 16840 -10090
rect 16960 -10210 17015 -10090
rect 17135 -10210 17180 -10090
rect 17300 -10210 17345 -10090
rect 17465 -10210 17510 -10090
rect 17630 -10210 17685 -10090
rect 17805 -10210 17850 -10090
rect 17970 -10210 18015 -10090
rect 18135 -10210 18180 -10090
rect 18300 -10210 18325 -10090
rect 12795 -10255 18325 -10210
rect 12795 -10375 12820 -10255
rect 12940 -10375 12995 -10255
rect 13115 -10375 13160 -10255
rect 13280 -10375 13325 -10255
rect 13445 -10375 13490 -10255
rect 13610 -10375 13665 -10255
rect 13785 -10375 13830 -10255
rect 13950 -10375 13995 -10255
rect 14115 -10375 14160 -10255
rect 14280 -10375 14335 -10255
rect 14455 -10375 14500 -10255
rect 14620 -10375 14665 -10255
rect 14785 -10375 14830 -10255
rect 14950 -10375 15005 -10255
rect 15125 -10375 15170 -10255
rect 15290 -10375 15335 -10255
rect 15455 -10375 15500 -10255
rect 15620 -10375 15675 -10255
rect 15795 -10375 15840 -10255
rect 15960 -10375 16005 -10255
rect 16125 -10375 16170 -10255
rect 16290 -10375 16345 -10255
rect 16465 -10375 16510 -10255
rect 16630 -10375 16675 -10255
rect 16795 -10375 16840 -10255
rect 16960 -10375 17015 -10255
rect 17135 -10375 17180 -10255
rect 17300 -10375 17345 -10255
rect 17465 -10375 17510 -10255
rect 17630 -10375 17685 -10255
rect 17805 -10375 17850 -10255
rect 17970 -10375 18015 -10255
rect 18135 -10375 18180 -10255
rect 18300 -10375 18325 -10255
rect 12795 -10420 18325 -10375
rect 12795 -10540 12820 -10420
rect 12940 -10540 12995 -10420
rect 13115 -10540 13160 -10420
rect 13280 -10540 13325 -10420
rect 13445 -10540 13490 -10420
rect 13610 -10540 13665 -10420
rect 13785 -10540 13830 -10420
rect 13950 -10540 13995 -10420
rect 14115 -10540 14160 -10420
rect 14280 -10540 14335 -10420
rect 14455 -10540 14500 -10420
rect 14620 -10540 14665 -10420
rect 14785 -10540 14830 -10420
rect 14950 -10540 15005 -10420
rect 15125 -10540 15170 -10420
rect 15290 -10540 15335 -10420
rect 15455 -10540 15500 -10420
rect 15620 -10540 15675 -10420
rect 15795 -10540 15840 -10420
rect 15960 -10540 16005 -10420
rect 16125 -10540 16170 -10420
rect 16290 -10540 16345 -10420
rect 16465 -10540 16510 -10420
rect 16630 -10540 16675 -10420
rect 16795 -10540 16840 -10420
rect 16960 -10540 17015 -10420
rect 17135 -10540 17180 -10420
rect 17300 -10540 17345 -10420
rect 17465 -10540 17510 -10420
rect 17630 -10540 17685 -10420
rect 17805 -10540 17850 -10420
rect 17970 -10540 18015 -10420
rect 18135 -10540 18180 -10420
rect 18300 -10540 18325 -10420
rect 12795 -10585 18325 -10540
rect 12795 -10705 12820 -10585
rect 12940 -10705 12995 -10585
rect 13115 -10705 13160 -10585
rect 13280 -10705 13325 -10585
rect 13445 -10705 13490 -10585
rect 13610 -10705 13665 -10585
rect 13785 -10705 13830 -10585
rect 13950 -10705 13995 -10585
rect 14115 -10705 14160 -10585
rect 14280 -10705 14335 -10585
rect 14455 -10705 14500 -10585
rect 14620 -10705 14665 -10585
rect 14785 -10705 14830 -10585
rect 14950 -10705 15005 -10585
rect 15125 -10705 15170 -10585
rect 15290 -10705 15335 -10585
rect 15455 -10705 15500 -10585
rect 15620 -10705 15675 -10585
rect 15795 -10705 15840 -10585
rect 15960 -10705 16005 -10585
rect 16125 -10705 16170 -10585
rect 16290 -10705 16345 -10585
rect 16465 -10705 16510 -10585
rect 16630 -10705 16675 -10585
rect 16795 -10705 16840 -10585
rect 16960 -10705 17015 -10585
rect 17135 -10705 17180 -10585
rect 17300 -10705 17345 -10585
rect 17465 -10705 17510 -10585
rect 17630 -10705 17685 -10585
rect 17805 -10705 17850 -10585
rect 17970 -10705 18015 -10585
rect 18135 -10705 18180 -10585
rect 18300 -10705 18325 -10585
rect 12795 -10760 18325 -10705
rect 12795 -10880 12820 -10760
rect 12940 -10880 12995 -10760
rect 13115 -10880 13160 -10760
rect 13280 -10880 13325 -10760
rect 13445 -10880 13490 -10760
rect 13610 -10880 13665 -10760
rect 13785 -10880 13830 -10760
rect 13950 -10880 13995 -10760
rect 14115 -10880 14160 -10760
rect 14280 -10880 14335 -10760
rect 14455 -10880 14500 -10760
rect 14620 -10880 14665 -10760
rect 14785 -10880 14830 -10760
rect 14950 -10880 15005 -10760
rect 15125 -10880 15170 -10760
rect 15290 -10880 15335 -10760
rect 15455 -10880 15500 -10760
rect 15620 -10880 15675 -10760
rect 15795 -10880 15840 -10760
rect 15960 -10880 16005 -10760
rect 16125 -10880 16170 -10760
rect 16290 -10880 16345 -10760
rect 16465 -10880 16510 -10760
rect 16630 -10880 16675 -10760
rect 16795 -10880 16840 -10760
rect 16960 -10880 17015 -10760
rect 17135 -10880 17180 -10760
rect 17300 -10880 17345 -10760
rect 17465 -10880 17510 -10760
rect 17630 -10880 17685 -10760
rect 17805 -10880 17850 -10760
rect 17970 -10880 18015 -10760
rect 18135 -10880 18180 -10760
rect 18300 -10880 18325 -10760
rect 12795 -10925 18325 -10880
rect 12795 -11045 12820 -10925
rect 12940 -11045 12995 -10925
rect 13115 -11045 13160 -10925
rect 13280 -11045 13325 -10925
rect 13445 -11045 13490 -10925
rect 13610 -11045 13665 -10925
rect 13785 -11045 13830 -10925
rect 13950 -11045 13995 -10925
rect 14115 -11045 14160 -10925
rect 14280 -11045 14335 -10925
rect 14455 -11045 14500 -10925
rect 14620 -11045 14665 -10925
rect 14785 -11045 14830 -10925
rect 14950 -11045 15005 -10925
rect 15125 -11045 15170 -10925
rect 15290 -11045 15335 -10925
rect 15455 -11045 15500 -10925
rect 15620 -11045 15675 -10925
rect 15795 -11045 15840 -10925
rect 15960 -11045 16005 -10925
rect 16125 -11045 16170 -10925
rect 16290 -11045 16345 -10925
rect 16465 -11045 16510 -10925
rect 16630 -11045 16675 -10925
rect 16795 -11045 16840 -10925
rect 16960 -11045 17015 -10925
rect 17135 -11045 17180 -10925
rect 17300 -11045 17345 -10925
rect 17465 -11045 17510 -10925
rect 17630 -11045 17685 -10925
rect 17805 -11045 17850 -10925
rect 17970 -11045 18015 -10925
rect 18135 -11045 18180 -10925
rect 18300 -11045 18325 -10925
rect 12795 -11090 18325 -11045
rect 12795 -11210 12820 -11090
rect 12940 -11210 12995 -11090
rect 13115 -11210 13160 -11090
rect 13280 -11210 13325 -11090
rect 13445 -11210 13490 -11090
rect 13610 -11210 13665 -11090
rect 13785 -11210 13830 -11090
rect 13950 -11210 13995 -11090
rect 14115 -11210 14160 -11090
rect 14280 -11210 14335 -11090
rect 14455 -11210 14500 -11090
rect 14620 -11210 14665 -11090
rect 14785 -11210 14830 -11090
rect 14950 -11210 15005 -11090
rect 15125 -11210 15170 -11090
rect 15290 -11210 15335 -11090
rect 15455 -11210 15500 -11090
rect 15620 -11210 15675 -11090
rect 15795 -11210 15840 -11090
rect 15960 -11210 16005 -11090
rect 16125 -11210 16170 -11090
rect 16290 -11210 16345 -11090
rect 16465 -11210 16510 -11090
rect 16630 -11210 16675 -11090
rect 16795 -11210 16840 -11090
rect 16960 -11210 17015 -11090
rect 17135 -11210 17180 -11090
rect 17300 -11210 17345 -11090
rect 17465 -11210 17510 -11090
rect 17630 -11210 17685 -11090
rect 17805 -11210 17850 -11090
rect 17970 -11210 18015 -11090
rect 18135 -11210 18180 -11090
rect 18300 -11210 18325 -11090
rect 12795 -11255 18325 -11210
rect 12795 -11375 12820 -11255
rect 12940 -11375 12995 -11255
rect 13115 -11375 13160 -11255
rect 13280 -11375 13325 -11255
rect 13445 -11375 13490 -11255
rect 13610 -11375 13665 -11255
rect 13785 -11375 13830 -11255
rect 13950 -11375 13995 -11255
rect 14115 -11375 14160 -11255
rect 14280 -11375 14335 -11255
rect 14455 -11375 14500 -11255
rect 14620 -11375 14665 -11255
rect 14785 -11375 14830 -11255
rect 14950 -11375 15005 -11255
rect 15125 -11375 15170 -11255
rect 15290 -11375 15335 -11255
rect 15455 -11375 15500 -11255
rect 15620 -11375 15675 -11255
rect 15795 -11375 15840 -11255
rect 15960 -11375 16005 -11255
rect 16125 -11375 16170 -11255
rect 16290 -11375 16345 -11255
rect 16465 -11375 16510 -11255
rect 16630 -11375 16675 -11255
rect 16795 -11375 16840 -11255
rect 16960 -11375 17015 -11255
rect 17135 -11375 17180 -11255
rect 17300 -11375 17345 -11255
rect 17465 -11375 17510 -11255
rect 17630 -11375 17685 -11255
rect 17805 -11375 17850 -11255
rect 17970 -11375 18015 -11255
rect 18135 -11375 18180 -11255
rect 18300 -11375 18325 -11255
rect 12795 -11430 18325 -11375
rect 12795 -11550 12820 -11430
rect 12940 -11550 12995 -11430
rect 13115 -11550 13160 -11430
rect 13280 -11550 13325 -11430
rect 13445 -11550 13490 -11430
rect 13610 -11550 13665 -11430
rect 13785 -11550 13830 -11430
rect 13950 -11550 13995 -11430
rect 14115 -11550 14160 -11430
rect 14280 -11550 14335 -11430
rect 14455 -11550 14500 -11430
rect 14620 -11550 14665 -11430
rect 14785 -11550 14830 -11430
rect 14950 -11550 15005 -11430
rect 15125 -11550 15170 -11430
rect 15290 -11550 15335 -11430
rect 15455 -11550 15500 -11430
rect 15620 -11550 15675 -11430
rect 15795 -11550 15840 -11430
rect 15960 -11550 16005 -11430
rect 16125 -11550 16170 -11430
rect 16290 -11550 16345 -11430
rect 16465 -11550 16510 -11430
rect 16630 -11550 16675 -11430
rect 16795 -11550 16840 -11430
rect 16960 -11550 17015 -11430
rect 17135 -11550 17180 -11430
rect 17300 -11550 17345 -11430
rect 17465 -11550 17510 -11430
rect 17630 -11550 17685 -11430
rect 17805 -11550 17850 -11430
rect 17970 -11550 18015 -11430
rect 18135 -11550 18180 -11430
rect 18300 -11550 18325 -11430
rect 12795 -11595 18325 -11550
rect 12795 -11715 12820 -11595
rect 12940 -11715 12995 -11595
rect 13115 -11715 13160 -11595
rect 13280 -11715 13325 -11595
rect 13445 -11715 13490 -11595
rect 13610 -11715 13665 -11595
rect 13785 -11715 13830 -11595
rect 13950 -11715 13995 -11595
rect 14115 -11715 14160 -11595
rect 14280 -11715 14335 -11595
rect 14455 -11715 14500 -11595
rect 14620 -11715 14665 -11595
rect 14785 -11715 14830 -11595
rect 14950 -11715 15005 -11595
rect 15125 -11715 15170 -11595
rect 15290 -11715 15335 -11595
rect 15455 -11715 15500 -11595
rect 15620 -11715 15675 -11595
rect 15795 -11715 15840 -11595
rect 15960 -11715 16005 -11595
rect 16125 -11715 16170 -11595
rect 16290 -11715 16345 -11595
rect 16465 -11715 16510 -11595
rect 16630 -11715 16675 -11595
rect 16795 -11715 16840 -11595
rect 16960 -11715 17015 -11595
rect 17135 -11715 17180 -11595
rect 17300 -11715 17345 -11595
rect 17465 -11715 17510 -11595
rect 17630 -11715 17685 -11595
rect 17805 -11715 17850 -11595
rect 17970 -11715 18015 -11595
rect 18135 -11715 18180 -11595
rect 18300 -11715 18325 -11595
rect 12795 -11760 18325 -11715
rect 12795 -11880 12820 -11760
rect 12940 -11880 12995 -11760
rect 13115 -11880 13160 -11760
rect 13280 -11880 13325 -11760
rect 13445 -11880 13490 -11760
rect 13610 -11880 13665 -11760
rect 13785 -11880 13830 -11760
rect 13950 -11880 13995 -11760
rect 14115 -11880 14160 -11760
rect 14280 -11880 14335 -11760
rect 14455 -11880 14500 -11760
rect 14620 -11880 14665 -11760
rect 14785 -11880 14830 -11760
rect 14950 -11880 15005 -11760
rect 15125 -11880 15170 -11760
rect 15290 -11880 15335 -11760
rect 15455 -11880 15500 -11760
rect 15620 -11880 15675 -11760
rect 15795 -11880 15840 -11760
rect 15960 -11880 16005 -11760
rect 16125 -11880 16170 -11760
rect 16290 -11880 16345 -11760
rect 16465 -11880 16510 -11760
rect 16630 -11880 16675 -11760
rect 16795 -11880 16840 -11760
rect 16960 -11880 17015 -11760
rect 17135 -11880 17180 -11760
rect 17300 -11880 17345 -11760
rect 17465 -11880 17510 -11760
rect 17630 -11880 17685 -11760
rect 17805 -11880 17850 -11760
rect 17970 -11880 18015 -11760
rect 18135 -11880 18180 -11760
rect 18300 -11880 18325 -11760
rect 12795 -11925 18325 -11880
rect 12795 -12045 12820 -11925
rect 12940 -12045 12995 -11925
rect 13115 -12045 13160 -11925
rect 13280 -12045 13325 -11925
rect 13445 -12045 13490 -11925
rect 13610 -12045 13665 -11925
rect 13785 -12045 13830 -11925
rect 13950 -12045 13995 -11925
rect 14115 -12045 14160 -11925
rect 14280 -12045 14335 -11925
rect 14455 -12045 14500 -11925
rect 14620 -12045 14665 -11925
rect 14785 -12045 14830 -11925
rect 14950 -12045 15005 -11925
rect 15125 -12045 15170 -11925
rect 15290 -12045 15335 -11925
rect 15455 -12045 15500 -11925
rect 15620 -12045 15675 -11925
rect 15795 -12045 15840 -11925
rect 15960 -12045 16005 -11925
rect 16125 -12045 16170 -11925
rect 16290 -12045 16345 -11925
rect 16465 -12045 16510 -11925
rect 16630 -12045 16675 -11925
rect 16795 -12045 16840 -11925
rect 16960 -12045 17015 -11925
rect 17135 -12045 17180 -11925
rect 17300 -12045 17345 -11925
rect 17465 -12045 17510 -11925
rect 17630 -12045 17685 -11925
rect 17805 -12045 17850 -11925
rect 17970 -12045 18015 -11925
rect 18135 -12045 18180 -11925
rect 18300 -12045 18325 -11925
rect 12795 -12100 18325 -12045
rect 12795 -12220 12820 -12100
rect 12940 -12220 12995 -12100
rect 13115 -12220 13160 -12100
rect 13280 -12220 13325 -12100
rect 13445 -12220 13490 -12100
rect 13610 -12220 13665 -12100
rect 13785 -12220 13830 -12100
rect 13950 -12220 13995 -12100
rect 14115 -12220 14160 -12100
rect 14280 -12220 14335 -12100
rect 14455 -12220 14500 -12100
rect 14620 -12220 14665 -12100
rect 14785 -12220 14830 -12100
rect 14950 -12220 15005 -12100
rect 15125 -12220 15170 -12100
rect 15290 -12220 15335 -12100
rect 15455 -12220 15500 -12100
rect 15620 -12220 15675 -12100
rect 15795 -12220 15840 -12100
rect 15960 -12220 16005 -12100
rect 16125 -12220 16170 -12100
rect 16290 -12220 16345 -12100
rect 16465 -12220 16510 -12100
rect 16630 -12220 16675 -12100
rect 16795 -12220 16840 -12100
rect 16960 -12220 17015 -12100
rect 17135 -12220 17180 -12100
rect 17300 -12220 17345 -12100
rect 17465 -12220 17510 -12100
rect 17630 -12220 17685 -12100
rect 17805 -12220 17850 -12100
rect 17970 -12220 18015 -12100
rect 18135 -12220 18180 -12100
rect 18300 -12220 18325 -12100
rect 12795 -12265 18325 -12220
rect 12795 -12385 12820 -12265
rect 12940 -12385 12995 -12265
rect 13115 -12385 13160 -12265
rect 13280 -12385 13325 -12265
rect 13445 -12385 13490 -12265
rect 13610 -12385 13665 -12265
rect 13785 -12385 13830 -12265
rect 13950 -12385 13995 -12265
rect 14115 -12385 14160 -12265
rect 14280 -12385 14335 -12265
rect 14455 -12385 14500 -12265
rect 14620 -12385 14665 -12265
rect 14785 -12385 14830 -12265
rect 14950 -12385 15005 -12265
rect 15125 -12385 15170 -12265
rect 15290 -12385 15335 -12265
rect 15455 -12385 15500 -12265
rect 15620 -12385 15675 -12265
rect 15795 -12385 15840 -12265
rect 15960 -12385 16005 -12265
rect 16125 -12385 16170 -12265
rect 16290 -12385 16345 -12265
rect 16465 -12385 16510 -12265
rect 16630 -12385 16675 -12265
rect 16795 -12385 16840 -12265
rect 16960 -12385 17015 -12265
rect 17135 -12385 17180 -12265
rect 17300 -12385 17345 -12265
rect 17465 -12385 17510 -12265
rect 17630 -12385 17685 -12265
rect 17805 -12385 17850 -12265
rect 17970 -12385 18015 -12265
rect 18135 -12385 18180 -12265
rect 18300 -12385 18325 -12265
rect 12795 -12430 18325 -12385
rect 12795 -12550 12820 -12430
rect 12940 -12550 12995 -12430
rect 13115 -12550 13160 -12430
rect 13280 -12550 13325 -12430
rect 13445 -12550 13490 -12430
rect 13610 -12550 13665 -12430
rect 13785 -12550 13830 -12430
rect 13950 -12550 13995 -12430
rect 14115 -12550 14160 -12430
rect 14280 -12550 14335 -12430
rect 14455 -12550 14500 -12430
rect 14620 -12550 14665 -12430
rect 14785 -12550 14830 -12430
rect 14950 -12550 15005 -12430
rect 15125 -12550 15170 -12430
rect 15290 -12550 15335 -12430
rect 15455 -12550 15500 -12430
rect 15620 -12550 15675 -12430
rect 15795 -12550 15840 -12430
rect 15960 -12550 16005 -12430
rect 16125 -12550 16170 -12430
rect 16290 -12550 16345 -12430
rect 16465 -12550 16510 -12430
rect 16630 -12550 16675 -12430
rect 16795 -12550 16840 -12430
rect 16960 -12550 17015 -12430
rect 17135 -12550 17180 -12430
rect 17300 -12550 17345 -12430
rect 17465 -12550 17510 -12430
rect 17630 -12550 17685 -12430
rect 17805 -12550 17850 -12430
rect 17970 -12550 18015 -12430
rect 18135 -12550 18180 -12430
rect 18300 -12550 18325 -12430
rect 12795 -12595 18325 -12550
rect 12795 -12715 12820 -12595
rect 12940 -12715 12995 -12595
rect 13115 -12715 13160 -12595
rect 13280 -12715 13325 -12595
rect 13445 -12715 13490 -12595
rect 13610 -12715 13665 -12595
rect 13785 -12715 13830 -12595
rect 13950 -12715 13995 -12595
rect 14115 -12715 14160 -12595
rect 14280 -12715 14335 -12595
rect 14455 -12715 14500 -12595
rect 14620 -12715 14665 -12595
rect 14785 -12715 14830 -12595
rect 14950 -12715 15005 -12595
rect 15125 -12715 15170 -12595
rect 15290 -12715 15335 -12595
rect 15455 -12715 15500 -12595
rect 15620 -12715 15675 -12595
rect 15795 -12715 15840 -12595
rect 15960 -12715 16005 -12595
rect 16125 -12715 16170 -12595
rect 16290 -12715 16345 -12595
rect 16465 -12715 16510 -12595
rect 16630 -12715 16675 -12595
rect 16795 -12715 16840 -12595
rect 16960 -12715 17015 -12595
rect 17135 -12715 17180 -12595
rect 17300 -12715 17345 -12595
rect 17465 -12715 17510 -12595
rect 17630 -12715 17685 -12595
rect 17805 -12715 17850 -12595
rect 17970 -12715 18015 -12595
rect 18135 -12715 18180 -12595
rect 18300 -12715 18325 -12595
rect 12795 -12770 18325 -12715
rect 12795 -12890 12820 -12770
rect 12940 -12890 12995 -12770
rect 13115 -12890 13160 -12770
rect 13280 -12890 13325 -12770
rect 13445 -12890 13490 -12770
rect 13610 -12890 13665 -12770
rect 13785 -12890 13830 -12770
rect 13950 -12890 13995 -12770
rect 14115 -12890 14160 -12770
rect 14280 -12890 14335 -12770
rect 14455 -12890 14500 -12770
rect 14620 -12890 14665 -12770
rect 14785 -12890 14830 -12770
rect 14950 -12890 15005 -12770
rect 15125 -12890 15170 -12770
rect 15290 -12890 15335 -12770
rect 15455 -12890 15500 -12770
rect 15620 -12890 15675 -12770
rect 15795 -12890 15840 -12770
rect 15960 -12890 16005 -12770
rect 16125 -12890 16170 -12770
rect 16290 -12890 16345 -12770
rect 16465 -12890 16510 -12770
rect 16630 -12890 16675 -12770
rect 16795 -12890 16840 -12770
rect 16960 -12890 17015 -12770
rect 17135 -12890 17180 -12770
rect 17300 -12890 17345 -12770
rect 17465 -12890 17510 -12770
rect 17630 -12890 17685 -12770
rect 17805 -12890 17850 -12770
rect 17970 -12890 18015 -12770
rect 18135 -12890 18180 -12770
rect 18300 -12890 18325 -12770
rect 12795 -12935 18325 -12890
rect 12795 -13055 12820 -12935
rect 12940 -13055 12995 -12935
rect 13115 -13055 13160 -12935
rect 13280 -13055 13325 -12935
rect 13445 -13055 13490 -12935
rect 13610 -13055 13665 -12935
rect 13785 -13055 13830 -12935
rect 13950 -13055 13995 -12935
rect 14115 -13055 14160 -12935
rect 14280 -13055 14335 -12935
rect 14455 -13055 14500 -12935
rect 14620 -13055 14665 -12935
rect 14785 -13055 14830 -12935
rect 14950 -13055 15005 -12935
rect 15125 -13055 15170 -12935
rect 15290 -13055 15335 -12935
rect 15455 -13055 15500 -12935
rect 15620 -13055 15675 -12935
rect 15795 -13055 15840 -12935
rect 15960 -13055 16005 -12935
rect 16125 -13055 16170 -12935
rect 16290 -13055 16345 -12935
rect 16465 -13055 16510 -12935
rect 16630 -13055 16675 -12935
rect 16795 -13055 16840 -12935
rect 16960 -13055 17015 -12935
rect 17135 -13055 17180 -12935
rect 17300 -13055 17345 -12935
rect 17465 -13055 17510 -12935
rect 17630 -13055 17685 -12935
rect 17805 -13055 17850 -12935
rect 17970 -13055 18015 -12935
rect 18135 -13055 18180 -12935
rect 18300 -13055 18325 -12935
rect 12795 -13100 18325 -13055
rect 12795 -13220 12820 -13100
rect 12940 -13220 12995 -13100
rect 13115 -13220 13160 -13100
rect 13280 -13220 13325 -13100
rect 13445 -13220 13490 -13100
rect 13610 -13220 13665 -13100
rect 13785 -13220 13830 -13100
rect 13950 -13220 13995 -13100
rect 14115 -13220 14160 -13100
rect 14280 -13220 14335 -13100
rect 14455 -13220 14500 -13100
rect 14620 -13220 14665 -13100
rect 14785 -13220 14830 -13100
rect 14950 -13220 15005 -13100
rect 15125 -13220 15170 -13100
rect 15290 -13220 15335 -13100
rect 15455 -13220 15500 -13100
rect 15620 -13220 15675 -13100
rect 15795 -13220 15840 -13100
rect 15960 -13220 16005 -13100
rect 16125 -13220 16170 -13100
rect 16290 -13220 16345 -13100
rect 16465 -13220 16510 -13100
rect 16630 -13220 16675 -13100
rect 16795 -13220 16840 -13100
rect 16960 -13220 17015 -13100
rect 17135 -13220 17180 -13100
rect 17300 -13220 17345 -13100
rect 17465 -13220 17510 -13100
rect 17630 -13220 17685 -13100
rect 17805 -13220 17850 -13100
rect 17970 -13220 18015 -13100
rect 18135 -13220 18180 -13100
rect 18300 -13220 18325 -13100
rect 12795 -13265 18325 -13220
rect 12795 -13385 12820 -13265
rect 12940 -13385 12995 -13265
rect 13115 -13385 13160 -13265
rect 13280 -13385 13325 -13265
rect 13445 -13385 13490 -13265
rect 13610 -13385 13665 -13265
rect 13785 -13385 13830 -13265
rect 13950 -13385 13995 -13265
rect 14115 -13385 14160 -13265
rect 14280 -13385 14335 -13265
rect 14455 -13385 14500 -13265
rect 14620 -13385 14665 -13265
rect 14785 -13385 14830 -13265
rect 14950 -13385 15005 -13265
rect 15125 -13385 15170 -13265
rect 15290 -13385 15335 -13265
rect 15455 -13385 15500 -13265
rect 15620 -13385 15675 -13265
rect 15795 -13385 15840 -13265
rect 15960 -13385 16005 -13265
rect 16125 -13385 16170 -13265
rect 16290 -13385 16345 -13265
rect 16465 -13385 16510 -13265
rect 16630 -13385 16675 -13265
rect 16795 -13385 16840 -13265
rect 16960 -13385 17015 -13265
rect 17135 -13385 17180 -13265
rect 17300 -13385 17345 -13265
rect 17465 -13385 17510 -13265
rect 17630 -13385 17685 -13265
rect 17805 -13385 17850 -13265
rect 17970 -13385 18015 -13265
rect 18135 -13385 18180 -13265
rect 18300 -13385 18325 -13265
rect 12795 -13440 18325 -13385
rect 12795 -13560 12820 -13440
rect 12940 -13560 12995 -13440
rect 13115 -13560 13160 -13440
rect 13280 -13560 13325 -13440
rect 13445 -13560 13490 -13440
rect 13610 -13560 13665 -13440
rect 13785 -13560 13830 -13440
rect 13950 -13560 13995 -13440
rect 14115 -13560 14160 -13440
rect 14280 -13560 14335 -13440
rect 14455 -13560 14500 -13440
rect 14620 -13560 14665 -13440
rect 14785 -13560 14830 -13440
rect 14950 -13560 15005 -13440
rect 15125 -13560 15170 -13440
rect 15290 -13560 15335 -13440
rect 15455 -13560 15500 -13440
rect 15620 -13560 15675 -13440
rect 15795 -13560 15840 -13440
rect 15960 -13560 16005 -13440
rect 16125 -13560 16170 -13440
rect 16290 -13560 16345 -13440
rect 16465 -13560 16510 -13440
rect 16630 -13560 16675 -13440
rect 16795 -13560 16840 -13440
rect 16960 -13560 17015 -13440
rect 17135 -13560 17180 -13440
rect 17300 -13560 17345 -13440
rect 17465 -13560 17510 -13440
rect 17630 -13560 17685 -13440
rect 17805 -13560 17850 -13440
rect 17970 -13560 18015 -13440
rect 18135 -13560 18180 -13440
rect 18300 -13560 18325 -13440
rect 12795 -13605 18325 -13560
rect 12795 -13725 12820 -13605
rect 12940 -13725 12995 -13605
rect 13115 -13725 13160 -13605
rect 13280 -13725 13325 -13605
rect 13445 -13725 13490 -13605
rect 13610 -13725 13665 -13605
rect 13785 -13725 13830 -13605
rect 13950 -13725 13995 -13605
rect 14115 -13725 14160 -13605
rect 14280 -13725 14335 -13605
rect 14455 -13725 14500 -13605
rect 14620 -13725 14665 -13605
rect 14785 -13725 14830 -13605
rect 14950 -13725 15005 -13605
rect 15125 -13725 15170 -13605
rect 15290 -13725 15335 -13605
rect 15455 -13725 15500 -13605
rect 15620 -13725 15675 -13605
rect 15795 -13725 15840 -13605
rect 15960 -13725 16005 -13605
rect 16125 -13725 16170 -13605
rect 16290 -13725 16345 -13605
rect 16465 -13725 16510 -13605
rect 16630 -13725 16675 -13605
rect 16795 -13725 16840 -13605
rect 16960 -13725 17015 -13605
rect 17135 -13725 17180 -13605
rect 17300 -13725 17345 -13605
rect 17465 -13725 17510 -13605
rect 17630 -13725 17685 -13605
rect 17805 -13725 17850 -13605
rect 17970 -13725 18015 -13605
rect 18135 -13725 18180 -13605
rect 18300 -13725 18325 -13605
rect 12795 -13770 18325 -13725
rect 12795 -13890 12820 -13770
rect 12940 -13890 12995 -13770
rect 13115 -13890 13160 -13770
rect 13280 -13890 13325 -13770
rect 13445 -13890 13490 -13770
rect 13610 -13890 13665 -13770
rect 13785 -13890 13830 -13770
rect 13950 -13890 13995 -13770
rect 14115 -13890 14160 -13770
rect 14280 -13890 14335 -13770
rect 14455 -13890 14500 -13770
rect 14620 -13890 14665 -13770
rect 14785 -13890 14830 -13770
rect 14950 -13890 15005 -13770
rect 15125 -13890 15170 -13770
rect 15290 -13890 15335 -13770
rect 15455 -13890 15500 -13770
rect 15620 -13890 15675 -13770
rect 15795 -13890 15840 -13770
rect 15960 -13890 16005 -13770
rect 16125 -13890 16170 -13770
rect 16290 -13890 16345 -13770
rect 16465 -13890 16510 -13770
rect 16630 -13890 16675 -13770
rect 16795 -13890 16840 -13770
rect 16960 -13890 17015 -13770
rect 17135 -13890 17180 -13770
rect 17300 -13890 17345 -13770
rect 17465 -13890 17510 -13770
rect 17630 -13890 17685 -13770
rect 17805 -13890 17850 -13770
rect 17970 -13890 18015 -13770
rect 18135 -13890 18180 -13770
rect 18300 -13890 18325 -13770
rect 12795 -13935 18325 -13890
rect 12795 -14055 12820 -13935
rect 12940 -14055 12995 -13935
rect 13115 -14055 13160 -13935
rect 13280 -14055 13325 -13935
rect 13445 -14055 13490 -13935
rect 13610 -14055 13665 -13935
rect 13785 -14055 13830 -13935
rect 13950 -14055 13995 -13935
rect 14115 -14055 14160 -13935
rect 14280 -14055 14335 -13935
rect 14455 -14055 14500 -13935
rect 14620 -14055 14665 -13935
rect 14785 -14055 14830 -13935
rect 14950 -14055 15005 -13935
rect 15125 -14055 15170 -13935
rect 15290 -14055 15335 -13935
rect 15455 -14055 15500 -13935
rect 15620 -14055 15675 -13935
rect 15795 -14055 15840 -13935
rect 15960 -14055 16005 -13935
rect 16125 -14055 16170 -13935
rect 16290 -14055 16345 -13935
rect 16465 -14055 16510 -13935
rect 16630 -14055 16675 -13935
rect 16795 -14055 16840 -13935
rect 16960 -14055 17015 -13935
rect 17135 -14055 17180 -13935
rect 17300 -14055 17345 -13935
rect 17465 -14055 17510 -13935
rect 17630 -14055 17685 -13935
rect 17805 -14055 17850 -13935
rect 17970 -14055 18015 -13935
rect 18135 -14055 18180 -13935
rect 18300 -14055 18325 -13935
rect 12795 -14110 18325 -14055
rect 12795 -14230 12820 -14110
rect 12940 -14230 12995 -14110
rect 13115 -14230 13160 -14110
rect 13280 -14230 13325 -14110
rect 13445 -14230 13490 -14110
rect 13610 -14230 13665 -14110
rect 13785 -14230 13830 -14110
rect 13950 -14230 13995 -14110
rect 14115 -14230 14160 -14110
rect 14280 -14230 14335 -14110
rect 14455 -14230 14500 -14110
rect 14620 -14230 14665 -14110
rect 14785 -14230 14830 -14110
rect 14950 -14230 15005 -14110
rect 15125 -14230 15170 -14110
rect 15290 -14230 15335 -14110
rect 15455 -14230 15500 -14110
rect 15620 -14230 15675 -14110
rect 15795 -14230 15840 -14110
rect 15960 -14230 16005 -14110
rect 16125 -14230 16170 -14110
rect 16290 -14230 16345 -14110
rect 16465 -14230 16510 -14110
rect 16630 -14230 16675 -14110
rect 16795 -14230 16840 -14110
rect 16960 -14230 17015 -14110
rect 17135 -14230 17180 -14110
rect 17300 -14230 17345 -14110
rect 17465 -14230 17510 -14110
rect 17630 -14230 17685 -14110
rect 17805 -14230 17850 -14110
rect 17970 -14230 18015 -14110
rect 18135 -14230 18180 -14110
rect 18300 -14230 18325 -14110
rect 12795 -14275 18325 -14230
rect 12795 -14395 12820 -14275
rect 12940 -14395 12995 -14275
rect 13115 -14395 13160 -14275
rect 13280 -14395 13325 -14275
rect 13445 -14395 13490 -14275
rect 13610 -14395 13665 -14275
rect 13785 -14395 13830 -14275
rect 13950 -14395 13995 -14275
rect 14115 -14395 14160 -14275
rect 14280 -14395 14335 -14275
rect 14455 -14395 14500 -14275
rect 14620 -14395 14665 -14275
rect 14785 -14395 14830 -14275
rect 14950 -14395 15005 -14275
rect 15125 -14395 15170 -14275
rect 15290 -14395 15335 -14275
rect 15455 -14395 15500 -14275
rect 15620 -14395 15675 -14275
rect 15795 -14395 15840 -14275
rect 15960 -14395 16005 -14275
rect 16125 -14395 16170 -14275
rect 16290 -14395 16345 -14275
rect 16465 -14395 16510 -14275
rect 16630 -14395 16675 -14275
rect 16795 -14395 16840 -14275
rect 16960 -14395 17015 -14275
rect 17135 -14395 17180 -14275
rect 17300 -14395 17345 -14275
rect 17465 -14395 17510 -14275
rect 17630 -14395 17685 -14275
rect 17805 -14395 17850 -14275
rect 17970 -14395 18015 -14275
rect 18135 -14395 18180 -14275
rect 18300 -14395 18325 -14275
rect 12795 -14440 18325 -14395
rect 12795 -14560 12820 -14440
rect 12940 -14560 12995 -14440
rect 13115 -14560 13160 -14440
rect 13280 -14560 13325 -14440
rect 13445 -14560 13490 -14440
rect 13610 -14560 13665 -14440
rect 13785 -14560 13830 -14440
rect 13950 -14560 13995 -14440
rect 14115 -14560 14160 -14440
rect 14280 -14560 14335 -14440
rect 14455 -14560 14500 -14440
rect 14620 -14560 14665 -14440
rect 14785 -14560 14830 -14440
rect 14950 -14560 15005 -14440
rect 15125 -14560 15170 -14440
rect 15290 -14560 15335 -14440
rect 15455 -14560 15500 -14440
rect 15620 -14560 15675 -14440
rect 15795 -14560 15840 -14440
rect 15960 -14560 16005 -14440
rect 16125 -14560 16170 -14440
rect 16290 -14560 16345 -14440
rect 16465 -14560 16510 -14440
rect 16630 -14560 16675 -14440
rect 16795 -14560 16840 -14440
rect 16960 -14560 17015 -14440
rect 17135 -14560 17180 -14440
rect 17300 -14560 17345 -14440
rect 17465 -14560 17510 -14440
rect 17630 -14560 17685 -14440
rect 17805 -14560 17850 -14440
rect 17970 -14560 18015 -14440
rect 18135 -14560 18180 -14440
rect 18300 -14560 18325 -14440
rect 12795 -14605 18325 -14560
rect 12795 -14725 12820 -14605
rect 12940 -14725 12995 -14605
rect 13115 -14725 13160 -14605
rect 13280 -14725 13325 -14605
rect 13445 -14725 13490 -14605
rect 13610 -14725 13665 -14605
rect 13785 -14725 13830 -14605
rect 13950 -14725 13995 -14605
rect 14115 -14725 14160 -14605
rect 14280 -14725 14335 -14605
rect 14455 -14725 14500 -14605
rect 14620 -14725 14665 -14605
rect 14785 -14725 14830 -14605
rect 14950 -14725 15005 -14605
rect 15125 -14725 15170 -14605
rect 15290 -14725 15335 -14605
rect 15455 -14725 15500 -14605
rect 15620 -14725 15675 -14605
rect 15795 -14725 15840 -14605
rect 15960 -14725 16005 -14605
rect 16125 -14725 16170 -14605
rect 16290 -14725 16345 -14605
rect 16465 -14725 16510 -14605
rect 16630 -14725 16675 -14605
rect 16795 -14725 16840 -14605
rect 16960 -14725 17015 -14605
rect 17135 -14725 17180 -14605
rect 17300 -14725 17345 -14605
rect 17465 -14725 17510 -14605
rect 17630 -14725 17685 -14605
rect 17805 -14725 17850 -14605
rect 17970 -14725 18015 -14605
rect 18135 -14725 18180 -14605
rect 18300 -14725 18325 -14605
rect 12795 -14780 18325 -14725
rect 12795 -14900 12820 -14780
rect 12940 -14900 12995 -14780
rect 13115 -14900 13160 -14780
rect 13280 -14900 13325 -14780
rect 13445 -14900 13490 -14780
rect 13610 -14900 13665 -14780
rect 13785 -14900 13830 -14780
rect 13950 -14900 13995 -14780
rect 14115 -14900 14160 -14780
rect 14280 -14900 14335 -14780
rect 14455 -14900 14500 -14780
rect 14620 -14900 14665 -14780
rect 14785 -14900 14830 -14780
rect 14950 -14900 15005 -14780
rect 15125 -14900 15170 -14780
rect 15290 -14900 15335 -14780
rect 15455 -14900 15500 -14780
rect 15620 -14900 15675 -14780
rect 15795 -14900 15840 -14780
rect 15960 -14900 16005 -14780
rect 16125 -14900 16170 -14780
rect 16290 -14900 16345 -14780
rect 16465 -14900 16510 -14780
rect 16630 -14900 16675 -14780
rect 16795 -14900 16840 -14780
rect 16960 -14900 17015 -14780
rect 17135 -14900 17180 -14780
rect 17300 -14900 17345 -14780
rect 17465 -14900 17510 -14780
rect 17630 -14900 17685 -14780
rect 17805 -14900 17850 -14780
rect 17970 -14900 18015 -14780
rect 18135 -14900 18180 -14780
rect 18300 -14900 18325 -14780
rect 12795 -14945 18325 -14900
rect 12795 -15065 12820 -14945
rect 12940 -15065 12995 -14945
rect 13115 -15065 13160 -14945
rect 13280 -15065 13325 -14945
rect 13445 -15065 13490 -14945
rect 13610 -15065 13665 -14945
rect 13785 -15065 13830 -14945
rect 13950 -15065 13995 -14945
rect 14115 -15065 14160 -14945
rect 14280 -15065 14335 -14945
rect 14455 -15065 14500 -14945
rect 14620 -15065 14665 -14945
rect 14785 -15065 14830 -14945
rect 14950 -15065 15005 -14945
rect 15125 -15065 15170 -14945
rect 15290 -15065 15335 -14945
rect 15455 -15065 15500 -14945
rect 15620 -15065 15675 -14945
rect 15795 -15065 15840 -14945
rect 15960 -15065 16005 -14945
rect 16125 -15065 16170 -14945
rect 16290 -15065 16345 -14945
rect 16465 -15065 16510 -14945
rect 16630 -15065 16675 -14945
rect 16795 -15065 16840 -14945
rect 16960 -15065 17015 -14945
rect 17135 -15065 17180 -14945
rect 17300 -15065 17345 -14945
rect 17465 -15065 17510 -14945
rect 17630 -15065 17685 -14945
rect 17805 -15065 17850 -14945
rect 17970 -15065 18015 -14945
rect 18135 -15065 18180 -14945
rect 18300 -15065 18325 -14945
rect 12795 -15110 18325 -15065
rect 12795 -15230 12820 -15110
rect 12940 -15230 12995 -15110
rect 13115 -15230 13160 -15110
rect 13280 -15230 13325 -15110
rect 13445 -15230 13490 -15110
rect 13610 -15230 13665 -15110
rect 13785 -15230 13830 -15110
rect 13950 -15230 13995 -15110
rect 14115 -15230 14160 -15110
rect 14280 -15230 14335 -15110
rect 14455 -15230 14500 -15110
rect 14620 -15230 14665 -15110
rect 14785 -15230 14830 -15110
rect 14950 -15230 15005 -15110
rect 15125 -15230 15170 -15110
rect 15290 -15230 15335 -15110
rect 15455 -15230 15500 -15110
rect 15620 -15230 15675 -15110
rect 15795 -15230 15840 -15110
rect 15960 -15230 16005 -15110
rect 16125 -15230 16170 -15110
rect 16290 -15230 16345 -15110
rect 16465 -15230 16510 -15110
rect 16630 -15230 16675 -15110
rect 16795 -15230 16840 -15110
rect 16960 -15230 17015 -15110
rect 17135 -15230 17180 -15110
rect 17300 -15230 17345 -15110
rect 17465 -15230 17510 -15110
rect 17630 -15230 17685 -15110
rect 17805 -15230 17850 -15110
rect 17970 -15230 18015 -15110
rect 18135 -15230 18180 -15110
rect 18300 -15230 18325 -15110
rect 12795 -15275 18325 -15230
rect 12795 -15395 12820 -15275
rect 12940 -15395 12995 -15275
rect 13115 -15395 13160 -15275
rect 13280 -15395 13325 -15275
rect 13445 -15395 13490 -15275
rect 13610 -15395 13665 -15275
rect 13785 -15395 13830 -15275
rect 13950 -15395 13995 -15275
rect 14115 -15395 14160 -15275
rect 14280 -15395 14335 -15275
rect 14455 -15395 14500 -15275
rect 14620 -15395 14665 -15275
rect 14785 -15395 14830 -15275
rect 14950 -15395 15005 -15275
rect 15125 -15395 15170 -15275
rect 15290 -15395 15335 -15275
rect 15455 -15395 15500 -15275
rect 15620 -15395 15675 -15275
rect 15795 -15395 15840 -15275
rect 15960 -15395 16005 -15275
rect 16125 -15395 16170 -15275
rect 16290 -15395 16345 -15275
rect 16465 -15395 16510 -15275
rect 16630 -15395 16675 -15275
rect 16795 -15395 16840 -15275
rect 16960 -15395 17015 -15275
rect 17135 -15395 17180 -15275
rect 17300 -15395 17345 -15275
rect 17465 -15395 17510 -15275
rect 17630 -15395 17685 -15275
rect 17805 -15395 17850 -15275
rect 17970 -15395 18015 -15275
rect 18135 -15395 18180 -15275
rect 18300 -15395 18325 -15275
rect 12795 -15450 18325 -15395
rect 12795 -15570 12820 -15450
rect 12940 -15570 12995 -15450
rect 13115 -15570 13160 -15450
rect 13280 -15570 13325 -15450
rect 13445 -15570 13490 -15450
rect 13610 -15570 13665 -15450
rect 13785 -15570 13830 -15450
rect 13950 -15570 13995 -15450
rect 14115 -15570 14160 -15450
rect 14280 -15570 14335 -15450
rect 14455 -15570 14500 -15450
rect 14620 -15570 14665 -15450
rect 14785 -15570 14830 -15450
rect 14950 -15570 15005 -15450
rect 15125 -15570 15170 -15450
rect 15290 -15570 15335 -15450
rect 15455 -15570 15500 -15450
rect 15620 -15570 15675 -15450
rect 15795 -15570 15840 -15450
rect 15960 -15570 16005 -15450
rect 16125 -15570 16170 -15450
rect 16290 -15570 16345 -15450
rect 16465 -15570 16510 -15450
rect 16630 -15570 16675 -15450
rect 16795 -15570 16840 -15450
rect 16960 -15570 17015 -15450
rect 17135 -15570 17180 -15450
rect 17300 -15570 17345 -15450
rect 17465 -15570 17510 -15450
rect 17630 -15570 17685 -15450
rect 17805 -15570 17850 -15450
rect 17970 -15570 18015 -15450
rect 18135 -15570 18180 -15450
rect 18300 -15570 18325 -15450
rect 12795 -15595 18325 -15570
rect 18485 -10090 24015 -10020
rect 18485 -10210 18510 -10090
rect 18630 -10210 18685 -10090
rect 18805 -10210 18850 -10090
rect 18970 -10210 19015 -10090
rect 19135 -10210 19180 -10090
rect 19300 -10210 19355 -10090
rect 19475 -10210 19520 -10090
rect 19640 -10210 19685 -10090
rect 19805 -10210 19850 -10090
rect 19970 -10210 20025 -10090
rect 20145 -10210 20190 -10090
rect 20310 -10210 20355 -10090
rect 20475 -10210 20520 -10090
rect 20640 -10210 20695 -10090
rect 20815 -10210 20860 -10090
rect 20980 -10210 21025 -10090
rect 21145 -10210 21190 -10090
rect 21310 -10210 21365 -10090
rect 21485 -10210 21530 -10090
rect 21650 -10210 21695 -10090
rect 21815 -10210 21860 -10090
rect 21980 -10210 22035 -10090
rect 22155 -10210 22200 -10090
rect 22320 -10210 22365 -10090
rect 22485 -10210 22530 -10090
rect 22650 -10210 22705 -10090
rect 22825 -10210 22870 -10090
rect 22990 -10210 23035 -10090
rect 23155 -10210 23200 -10090
rect 23320 -10210 23375 -10090
rect 23495 -10210 23540 -10090
rect 23660 -10210 23705 -10090
rect 23825 -10210 23870 -10090
rect 23990 -10210 24015 -10090
rect 18485 -10255 24015 -10210
rect 18485 -10375 18510 -10255
rect 18630 -10375 18685 -10255
rect 18805 -10375 18850 -10255
rect 18970 -10375 19015 -10255
rect 19135 -10375 19180 -10255
rect 19300 -10375 19355 -10255
rect 19475 -10375 19520 -10255
rect 19640 -10375 19685 -10255
rect 19805 -10375 19850 -10255
rect 19970 -10375 20025 -10255
rect 20145 -10375 20190 -10255
rect 20310 -10375 20355 -10255
rect 20475 -10375 20520 -10255
rect 20640 -10375 20695 -10255
rect 20815 -10375 20860 -10255
rect 20980 -10375 21025 -10255
rect 21145 -10375 21190 -10255
rect 21310 -10375 21365 -10255
rect 21485 -10375 21530 -10255
rect 21650 -10375 21695 -10255
rect 21815 -10375 21860 -10255
rect 21980 -10375 22035 -10255
rect 22155 -10375 22200 -10255
rect 22320 -10375 22365 -10255
rect 22485 -10375 22530 -10255
rect 22650 -10375 22705 -10255
rect 22825 -10375 22870 -10255
rect 22990 -10375 23035 -10255
rect 23155 -10375 23200 -10255
rect 23320 -10375 23375 -10255
rect 23495 -10375 23540 -10255
rect 23660 -10375 23705 -10255
rect 23825 -10375 23870 -10255
rect 23990 -10375 24015 -10255
rect 18485 -10420 24015 -10375
rect 18485 -10540 18510 -10420
rect 18630 -10540 18685 -10420
rect 18805 -10540 18850 -10420
rect 18970 -10540 19015 -10420
rect 19135 -10540 19180 -10420
rect 19300 -10540 19355 -10420
rect 19475 -10540 19520 -10420
rect 19640 -10540 19685 -10420
rect 19805 -10540 19850 -10420
rect 19970 -10540 20025 -10420
rect 20145 -10540 20190 -10420
rect 20310 -10540 20355 -10420
rect 20475 -10540 20520 -10420
rect 20640 -10540 20695 -10420
rect 20815 -10540 20860 -10420
rect 20980 -10540 21025 -10420
rect 21145 -10540 21190 -10420
rect 21310 -10540 21365 -10420
rect 21485 -10540 21530 -10420
rect 21650 -10540 21695 -10420
rect 21815 -10540 21860 -10420
rect 21980 -10540 22035 -10420
rect 22155 -10540 22200 -10420
rect 22320 -10540 22365 -10420
rect 22485 -10540 22530 -10420
rect 22650 -10540 22705 -10420
rect 22825 -10540 22870 -10420
rect 22990 -10540 23035 -10420
rect 23155 -10540 23200 -10420
rect 23320 -10540 23375 -10420
rect 23495 -10540 23540 -10420
rect 23660 -10540 23705 -10420
rect 23825 -10540 23870 -10420
rect 23990 -10540 24015 -10420
rect 18485 -10585 24015 -10540
rect 18485 -10705 18510 -10585
rect 18630 -10705 18685 -10585
rect 18805 -10705 18850 -10585
rect 18970 -10705 19015 -10585
rect 19135 -10705 19180 -10585
rect 19300 -10705 19355 -10585
rect 19475 -10705 19520 -10585
rect 19640 -10705 19685 -10585
rect 19805 -10705 19850 -10585
rect 19970 -10705 20025 -10585
rect 20145 -10705 20190 -10585
rect 20310 -10705 20355 -10585
rect 20475 -10705 20520 -10585
rect 20640 -10705 20695 -10585
rect 20815 -10705 20860 -10585
rect 20980 -10705 21025 -10585
rect 21145 -10705 21190 -10585
rect 21310 -10705 21365 -10585
rect 21485 -10705 21530 -10585
rect 21650 -10705 21695 -10585
rect 21815 -10705 21860 -10585
rect 21980 -10705 22035 -10585
rect 22155 -10705 22200 -10585
rect 22320 -10705 22365 -10585
rect 22485 -10705 22530 -10585
rect 22650 -10705 22705 -10585
rect 22825 -10705 22870 -10585
rect 22990 -10705 23035 -10585
rect 23155 -10705 23200 -10585
rect 23320 -10705 23375 -10585
rect 23495 -10705 23540 -10585
rect 23660 -10705 23705 -10585
rect 23825 -10705 23870 -10585
rect 23990 -10705 24015 -10585
rect 18485 -10760 24015 -10705
rect 18485 -10880 18510 -10760
rect 18630 -10880 18685 -10760
rect 18805 -10880 18850 -10760
rect 18970 -10880 19015 -10760
rect 19135 -10880 19180 -10760
rect 19300 -10880 19355 -10760
rect 19475 -10880 19520 -10760
rect 19640 -10880 19685 -10760
rect 19805 -10880 19850 -10760
rect 19970 -10880 20025 -10760
rect 20145 -10880 20190 -10760
rect 20310 -10880 20355 -10760
rect 20475 -10880 20520 -10760
rect 20640 -10880 20695 -10760
rect 20815 -10880 20860 -10760
rect 20980 -10880 21025 -10760
rect 21145 -10880 21190 -10760
rect 21310 -10880 21365 -10760
rect 21485 -10880 21530 -10760
rect 21650 -10880 21695 -10760
rect 21815 -10880 21860 -10760
rect 21980 -10880 22035 -10760
rect 22155 -10880 22200 -10760
rect 22320 -10880 22365 -10760
rect 22485 -10880 22530 -10760
rect 22650 -10880 22705 -10760
rect 22825 -10880 22870 -10760
rect 22990 -10880 23035 -10760
rect 23155 -10880 23200 -10760
rect 23320 -10880 23375 -10760
rect 23495 -10880 23540 -10760
rect 23660 -10880 23705 -10760
rect 23825 -10880 23870 -10760
rect 23990 -10880 24015 -10760
rect 18485 -10925 24015 -10880
rect 18485 -11045 18510 -10925
rect 18630 -11045 18685 -10925
rect 18805 -11045 18850 -10925
rect 18970 -11045 19015 -10925
rect 19135 -11045 19180 -10925
rect 19300 -11045 19355 -10925
rect 19475 -11045 19520 -10925
rect 19640 -11045 19685 -10925
rect 19805 -11045 19850 -10925
rect 19970 -11045 20025 -10925
rect 20145 -11045 20190 -10925
rect 20310 -11045 20355 -10925
rect 20475 -11045 20520 -10925
rect 20640 -11045 20695 -10925
rect 20815 -11045 20860 -10925
rect 20980 -11045 21025 -10925
rect 21145 -11045 21190 -10925
rect 21310 -11045 21365 -10925
rect 21485 -11045 21530 -10925
rect 21650 -11045 21695 -10925
rect 21815 -11045 21860 -10925
rect 21980 -11045 22035 -10925
rect 22155 -11045 22200 -10925
rect 22320 -11045 22365 -10925
rect 22485 -11045 22530 -10925
rect 22650 -11045 22705 -10925
rect 22825 -11045 22870 -10925
rect 22990 -11045 23035 -10925
rect 23155 -11045 23200 -10925
rect 23320 -11045 23375 -10925
rect 23495 -11045 23540 -10925
rect 23660 -11045 23705 -10925
rect 23825 -11045 23870 -10925
rect 23990 -11045 24015 -10925
rect 18485 -11090 24015 -11045
rect 18485 -11210 18510 -11090
rect 18630 -11210 18685 -11090
rect 18805 -11210 18850 -11090
rect 18970 -11210 19015 -11090
rect 19135 -11210 19180 -11090
rect 19300 -11210 19355 -11090
rect 19475 -11210 19520 -11090
rect 19640 -11210 19685 -11090
rect 19805 -11210 19850 -11090
rect 19970 -11210 20025 -11090
rect 20145 -11210 20190 -11090
rect 20310 -11210 20355 -11090
rect 20475 -11210 20520 -11090
rect 20640 -11210 20695 -11090
rect 20815 -11210 20860 -11090
rect 20980 -11210 21025 -11090
rect 21145 -11210 21190 -11090
rect 21310 -11210 21365 -11090
rect 21485 -11210 21530 -11090
rect 21650 -11210 21695 -11090
rect 21815 -11210 21860 -11090
rect 21980 -11210 22035 -11090
rect 22155 -11210 22200 -11090
rect 22320 -11210 22365 -11090
rect 22485 -11210 22530 -11090
rect 22650 -11210 22705 -11090
rect 22825 -11210 22870 -11090
rect 22990 -11210 23035 -11090
rect 23155 -11210 23200 -11090
rect 23320 -11210 23375 -11090
rect 23495 -11210 23540 -11090
rect 23660 -11210 23705 -11090
rect 23825 -11210 23870 -11090
rect 23990 -11210 24015 -11090
rect 18485 -11255 24015 -11210
rect 18485 -11375 18510 -11255
rect 18630 -11375 18685 -11255
rect 18805 -11375 18850 -11255
rect 18970 -11375 19015 -11255
rect 19135 -11375 19180 -11255
rect 19300 -11375 19355 -11255
rect 19475 -11375 19520 -11255
rect 19640 -11375 19685 -11255
rect 19805 -11375 19850 -11255
rect 19970 -11375 20025 -11255
rect 20145 -11375 20190 -11255
rect 20310 -11375 20355 -11255
rect 20475 -11375 20520 -11255
rect 20640 -11375 20695 -11255
rect 20815 -11375 20860 -11255
rect 20980 -11375 21025 -11255
rect 21145 -11375 21190 -11255
rect 21310 -11375 21365 -11255
rect 21485 -11375 21530 -11255
rect 21650 -11375 21695 -11255
rect 21815 -11375 21860 -11255
rect 21980 -11375 22035 -11255
rect 22155 -11375 22200 -11255
rect 22320 -11375 22365 -11255
rect 22485 -11375 22530 -11255
rect 22650 -11375 22705 -11255
rect 22825 -11375 22870 -11255
rect 22990 -11375 23035 -11255
rect 23155 -11375 23200 -11255
rect 23320 -11375 23375 -11255
rect 23495 -11375 23540 -11255
rect 23660 -11375 23705 -11255
rect 23825 -11375 23870 -11255
rect 23990 -11375 24015 -11255
rect 18485 -11430 24015 -11375
rect 18485 -11550 18510 -11430
rect 18630 -11550 18685 -11430
rect 18805 -11550 18850 -11430
rect 18970 -11550 19015 -11430
rect 19135 -11550 19180 -11430
rect 19300 -11550 19355 -11430
rect 19475 -11550 19520 -11430
rect 19640 -11550 19685 -11430
rect 19805 -11550 19850 -11430
rect 19970 -11550 20025 -11430
rect 20145 -11550 20190 -11430
rect 20310 -11550 20355 -11430
rect 20475 -11550 20520 -11430
rect 20640 -11550 20695 -11430
rect 20815 -11550 20860 -11430
rect 20980 -11550 21025 -11430
rect 21145 -11550 21190 -11430
rect 21310 -11550 21365 -11430
rect 21485 -11550 21530 -11430
rect 21650 -11550 21695 -11430
rect 21815 -11550 21860 -11430
rect 21980 -11550 22035 -11430
rect 22155 -11550 22200 -11430
rect 22320 -11550 22365 -11430
rect 22485 -11550 22530 -11430
rect 22650 -11550 22705 -11430
rect 22825 -11550 22870 -11430
rect 22990 -11550 23035 -11430
rect 23155 -11550 23200 -11430
rect 23320 -11550 23375 -11430
rect 23495 -11550 23540 -11430
rect 23660 -11550 23705 -11430
rect 23825 -11550 23870 -11430
rect 23990 -11550 24015 -11430
rect 18485 -11595 24015 -11550
rect 18485 -11715 18510 -11595
rect 18630 -11715 18685 -11595
rect 18805 -11715 18850 -11595
rect 18970 -11715 19015 -11595
rect 19135 -11715 19180 -11595
rect 19300 -11715 19355 -11595
rect 19475 -11715 19520 -11595
rect 19640 -11715 19685 -11595
rect 19805 -11715 19850 -11595
rect 19970 -11715 20025 -11595
rect 20145 -11715 20190 -11595
rect 20310 -11715 20355 -11595
rect 20475 -11715 20520 -11595
rect 20640 -11715 20695 -11595
rect 20815 -11715 20860 -11595
rect 20980 -11715 21025 -11595
rect 21145 -11715 21190 -11595
rect 21310 -11715 21365 -11595
rect 21485 -11715 21530 -11595
rect 21650 -11715 21695 -11595
rect 21815 -11715 21860 -11595
rect 21980 -11715 22035 -11595
rect 22155 -11715 22200 -11595
rect 22320 -11715 22365 -11595
rect 22485 -11715 22530 -11595
rect 22650 -11715 22705 -11595
rect 22825 -11715 22870 -11595
rect 22990 -11715 23035 -11595
rect 23155 -11715 23200 -11595
rect 23320 -11715 23375 -11595
rect 23495 -11715 23540 -11595
rect 23660 -11715 23705 -11595
rect 23825 -11715 23870 -11595
rect 23990 -11715 24015 -11595
rect 18485 -11760 24015 -11715
rect 18485 -11880 18510 -11760
rect 18630 -11880 18685 -11760
rect 18805 -11880 18850 -11760
rect 18970 -11880 19015 -11760
rect 19135 -11880 19180 -11760
rect 19300 -11880 19355 -11760
rect 19475 -11880 19520 -11760
rect 19640 -11880 19685 -11760
rect 19805 -11880 19850 -11760
rect 19970 -11880 20025 -11760
rect 20145 -11880 20190 -11760
rect 20310 -11880 20355 -11760
rect 20475 -11880 20520 -11760
rect 20640 -11880 20695 -11760
rect 20815 -11880 20860 -11760
rect 20980 -11880 21025 -11760
rect 21145 -11880 21190 -11760
rect 21310 -11880 21365 -11760
rect 21485 -11880 21530 -11760
rect 21650 -11880 21695 -11760
rect 21815 -11880 21860 -11760
rect 21980 -11880 22035 -11760
rect 22155 -11880 22200 -11760
rect 22320 -11880 22365 -11760
rect 22485 -11880 22530 -11760
rect 22650 -11880 22705 -11760
rect 22825 -11880 22870 -11760
rect 22990 -11880 23035 -11760
rect 23155 -11880 23200 -11760
rect 23320 -11880 23375 -11760
rect 23495 -11880 23540 -11760
rect 23660 -11880 23705 -11760
rect 23825 -11880 23870 -11760
rect 23990 -11880 24015 -11760
rect 18485 -11925 24015 -11880
rect 18485 -12045 18510 -11925
rect 18630 -12045 18685 -11925
rect 18805 -12045 18850 -11925
rect 18970 -12045 19015 -11925
rect 19135 -12045 19180 -11925
rect 19300 -12045 19355 -11925
rect 19475 -12045 19520 -11925
rect 19640 -12045 19685 -11925
rect 19805 -12045 19850 -11925
rect 19970 -12045 20025 -11925
rect 20145 -12045 20190 -11925
rect 20310 -12045 20355 -11925
rect 20475 -12045 20520 -11925
rect 20640 -12045 20695 -11925
rect 20815 -12045 20860 -11925
rect 20980 -12045 21025 -11925
rect 21145 -12045 21190 -11925
rect 21310 -12045 21365 -11925
rect 21485 -12045 21530 -11925
rect 21650 -12045 21695 -11925
rect 21815 -12045 21860 -11925
rect 21980 -12045 22035 -11925
rect 22155 -12045 22200 -11925
rect 22320 -12045 22365 -11925
rect 22485 -12045 22530 -11925
rect 22650 -12045 22705 -11925
rect 22825 -12045 22870 -11925
rect 22990 -12045 23035 -11925
rect 23155 -12045 23200 -11925
rect 23320 -12045 23375 -11925
rect 23495 -12045 23540 -11925
rect 23660 -12045 23705 -11925
rect 23825 -12045 23870 -11925
rect 23990 -12045 24015 -11925
rect 18485 -12100 24015 -12045
rect 18485 -12220 18510 -12100
rect 18630 -12220 18685 -12100
rect 18805 -12220 18850 -12100
rect 18970 -12220 19015 -12100
rect 19135 -12220 19180 -12100
rect 19300 -12220 19355 -12100
rect 19475 -12220 19520 -12100
rect 19640 -12220 19685 -12100
rect 19805 -12220 19850 -12100
rect 19970 -12220 20025 -12100
rect 20145 -12220 20190 -12100
rect 20310 -12220 20355 -12100
rect 20475 -12220 20520 -12100
rect 20640 -12220 20695 -12100
rect 20815 -12220 20860 -12100
rect 20980 -12220 21025 -12100
rect 21145 -12220 21190 -12100
rect 21310 -12220 21365 -12100
rect 21485 -12220 21530 -12100
rect 21650 -12220 21695 -12100
rect 21815 -12220 21860 -12100
rect 21980 -12220 22035 -12100
rect 22155 -12220 22200 -12100
rect 22320 -12220 22365 -12100
rect 22485 -12220 22530 -12100
rect 22650 -12220 22705 -12100
rect 22825 -12220 22870 -12100
rect 22990 -12220 23035 -12100
rect 23155 -12220 23200 -12100
rect 23320 -12220 23375 -12100
rect 23495 -12220 23540 -12100
rect 23660 -12220 23705 -12100
rect 23825 -12220 23870 -12100
rect 23990 -12220 24015 -12100
rect 18485 -12265 24015 -12220
rect 18485 -12385 18510 -12265
rect 18630 -12385 18685 -12265
rect 18805 -12385 18850 -12265
rect 18970 -12385 19015 -12265
rect 19135 -12385 19180 -12265
rect 19300 -12385 19355 -12265
rect 19475 -12385 19520 -12265
rect 19640 -12385 19685 -12265
rect 19805 -12385 19850 -12265
rect 19970 -12385 20025 -12265
rect 20145 -12385 20190 -12265
rect 20310 -12385 20355 -12265
rect 20475 -12385 20520 -12265
rect 20640 -12385 20695 -12265
rect 20815 -12385 20860 -12265
rect 20980 -12385 21025 -12265
rect 21145 -12385 21190 -12265
rect 21310 -12385 21365 -12265
rect 21485 -12385 21530 -12265
rect 21650 -12385 21695 -12265
rect 21815 -12385 21860 -12265
rect 21980 -12385 22035 -12265
rect 22155 -12385 22200 -12265
rect 22320 -12385 22365 -12265
rect 22485 -12385 22530 -12265
rect 22650 -12385 22705 -12265
rect 22825 -12385 22870 -12265
rect 22990 -12385 23035 -12265
rect 23155 -12385 23200 -12265
rect 23320 -12385 23375 -12265
rect 23495 -12385 23540 -12265
rect 23660 -12385 23705 -12265
rect 23825 -12385 23870 -12265
rect 23990 -12385 24015 -12265
rect 18485 -12430 24015 -12385
rect 18485 -12550 18510 -12430
rect 18630 -12550 18685 -12430
rect 18805 -12550 18850 -12430
rect 18970 -12550 19015 -12430
rect 19135 -12550 19180 -12430
rect 19300 -12550 19355 -12430
rect 19475 -12550 19520 -12430
rect 19640 -12550 19685 -12430
rect 19805 -12550 19850 -12430
rect 19970 -12550 20025 -12430
rect 20145 -12550 20190 -12430
rect 20310 -12550 20355 -12430
rect 20475 -12550 20520 -12430
rect 20640 -12550 20695 -12430
rect 20815 -12550 20860 -12430
rect 20980 -12550 21025 -12430
rect 21145 -12550 21190 -12430
rect 21310 -12550 21365 -12430
rect 21485 -12550 21530 -12430
rect 21650 -12550 21695 -12430
rect 21815 -12550 21860 -12430
rect 21980 -12550 22035 -12430
rect 22155 -12550 22200 -12430
rect 22320 -12550 22365 -12430
rect 22485 -12550 22530 -12430
rect 22650 -12550 22705 -12430
rect 22825 -12550 22870 -12430
rect 22990 -12550 23035 -12430
rect 23155 -12550 23200 -12430
rect 23320 -12550 23375 -12430
rect 23495 -12550 23540 -12430
rect 23660 -12550 23705 -12430
rect 23825 -12550 23870 -12430
rect 23990 -12550 24015 -12430
rect 18485 -12595 24015 -12550
rect 18485 -12715 18510 -12595
rect 18630 -12715 18685 -12595
rect 18805 -12715 18850 -12595
rect 18970 -12715 19015 -12595
rect 19135 -12715 19180 -12595
rect 19300 -12715 19355 -12595
rect 19475 -12715 19520 -12595
rect 19640 -12715 19685 -12595
rect 19805 -12715 19850 -12595
rect 19970 -12715 20025 -12595
rect 20145 -12715 20190 -12595
rect 20310 -12715 20355 -12595
rect 20475 -12715 20520 -12595
rect 20640 -12715 20695 -12595
rect 20815 -12715 20860 -12595
rect 20980 -12715 21025 -12595
rect 21145 -12715 21190 -12595
rect 21310 -12715 21365 -12595
rect 21485 -12715 21530 -12595
rect 21650 -12715 21695 -12595
rect 21815 -12715 21860 -12595
rect 21980 -12715 22035 -12595
rect 22155 -12715 22200 -12595
rect 22320 -12715 22365 -12595
rect 22485 -12715 22530 -12595
rect 22650 -12715 22705 -12595
rect 22825 -12715 22870 -12595
rect 22990 -12715 23035 -12595
rect 23155 -12715 23200 -12595
rect 23320 -12715 23375 -12595
rect 23495 -12715 23540 -12595
rect 23660 -12715 23705 -12595
rect 23825 -12715 23870 -12595
rect 23990 -12715 24015 -12595
rect 18485 -12770 24015 -12715
rect 18485 -12890 18510 -12770
rect 18630 -12890 18685 -12770
rect 18805 -12890 18850 -12770
rect 18970 -12890 19015 -12770
rect 19135 -12890 19180 -12770
rect 19300 -12890 19355 -12770
rect 19475 -12890 19520 -12770
rect 19640 -12890 19685 -12770
rect 19805 -12890 19850 -12770
rect 19970 -12890 20025 -12770
rect 20145 -12890 20190 -12770
rect 20310 -12890 20355 -12770
rect 20475 -12890 20520 -12770
rect 20640 -12890 20695 -12770
rect 20815 -12890 20860 -12770
rect 20980 -12890 21025 -12770
rect 21145 -12890 21190 -12770
rect 21310 -12890 21365 -12770
rect 21485 -12890 21530 -12770
rect 21650 -12890 21695 -12770
rect 21815 -12890 21860 -12770
rect 21980 -12890 22035 -12770
rect 22155 -12890 22200 -12770
rect 22320 -12890 22365 -12770
rect 22485 -12890 22530 -12770
rect 22650 -12890 22705 -12770
rect 22825 -12890 22870 -12770
rect 22990 -12890 23035 -12770
rect 23155 -12890 23200 -12770
rect 23320 -12890 23375 -12770
rect 23495 -12890 23540 -12770
rect 23660 -12890 23705 -12770
rect 23825 -12890 23870 -12770
rect 23990 -12890 24015 -12770
rect 18485 -12935 24015 -12890
rect 18485 -13055 18510 -12935
rect 18630 -13055 18685 -12935
rect 18805 -13055 18850 -12935
rect 18970 -13055 19015 -12935
rect 19135 -13055 19180 -12935
rect 19300 -13055 19355 -12935
rect 19475 -13055 19520 -12935
rect 19640 -13055 19685 -12935
rect 19805 -13055 19850 -12935
rect 19970 -13055 20025 -12935
rect 20145 -13055 20190 -12935
rect 20310 -13055 20355 -12935
rect 20475 -13055 20520 -12935
rect 20640 -13055 20695 -12935
rect 20815 -13055 20860 -12935
rect 20980 -13055 21025 -12935
rect 21145 -13055 21190 -12935
rect 21310 -13055 21365 -12935
rect 21485 -13055 21530 -12935
rect 21650 -13055 21695 -12935
rect 21815 -13055 21860 -12935
rect 21980 -13055 22035 -12935
rect 22155 -13055 22200 -12935
rect 22320 -13055 22365 -12935
rect 22485 -13055 22530 -12935
rect 22650 -13055 22705 -12935
rect 22825 -13055 22870 -12935
rect 22990 -13055 23035 -12935
rect 23155 -13055 23200 -12935
rect 23320 -13055 23375 -12935
rect 23495 -13055 23540 -12935
rect 23660 -13055 23705 -12935
rect 23825 -13055 23870 -12935
rect 23990 -13055 24015 -12935
rect 18485 -13100 24015 -13055
rect 18485 -13220 18510 -13100
rect 18630 -13220 18685 -13100
rect 18805 -13220 18850 -13100
rect 18970 -13220 19015 -13100
rect 19135 -13220 19180 -13100
rect 19300 -13220 19355 -13100
rect 19475 -13220 19520 -13100
rect 19640 -13220 19685 -13100
rect 19805 -13220 19850 -13100
rect 19970 -13220 20025 -13100
rect 20145 -13220 20190 -13100
rect 20310 -13220 20355 -13100
rect 20475 -13220 20520 -13100
rect 20640 -13220 20695 -13100
rect 20815 -13220 20860 -13100
rect 20980 -13220 21025 -13100
rect 21145 -13220 21190 -13100
rect 21310 -13220 21365 -13100
rect 21485 -13220 21530 -13100
rect 21650 -13220 21695 -13100
rect 21815 -13220 21860 -13100
rect 21980 -13220 22035 -13100
rect 22155 -13220 22200 -13100
rect 22320 -13220 22365 -13100
rect 22485 -13220 22530 -13100
rect 22650 -13220 22705 -13100
rect 22825 -13220 22870 -13100
rect 22990 -13220 23035 -13100
rect 23155 -13220 23200 -13100
rect 23320 -13220 23375 -13100
rect 23495 -13220 23540 -13100
rect 23660 -13220 23705 -13100
rect 23825 -13220 23870 -13100
rect 23990 -13220 24015 -13100
rect 18485 -13265 24015 -13220
rect 18485 -13385 18510 -13265
rect 18630 -13385 18685 -13265
rect 18805 -13385 18850 -13265
rect 18970 -13385 19015 -13265
rect 19135 -13385 19180 -13265
rect 19300 -13385 19355 -13265
rect 19475 -13385 19520 -13265
rect 19640 -13385 19685 -13265
rect 19805 -13385 19850 -13265
rect 19970 -13385 20025 -13265
rect 20145 -13385 20190 -13265
rect 20310 -13385 20355 -13265
rect 20475 -13385 20520 -13265
rect 20640 -13385 20695 -13265
rect 20815 -13385 20860 -13265
rect 20980 -13385 21025 -13265
rect 21145 -13385 21190 -13265
rect 21310 -13385 21365 -13265
rect 21485 -13385 21530 -13265
rect 21650 -13385 21695 -13265
rect 21815 -13385 21860 -13265
rect 21980 -13385 22035 -13265
rect 22155 -13385 22200 -13265
rect 22320 -13385 22365 -13265
rect 22485 -13385 22530 -13265
rect 22650 -13385 22705 -13265
rect 22825 -13385 22870 -13265
rect 22990 -13385 23035 -13265
rect 23155 -13385 23200 -13265
rect 23320 -13385 23375 -13265
rect 23495 -13385 23540 -13265
rect 23660 -13385 23705 -13265
rect 23825 -13385 23870 -13265
rect 23990 -13385 24015 -13265
rect 18485 -13440 24015 -13385
rect 18485 -13560 18510 -13440
rect 18630 -13560 18685 -13440
rect 18805 -13560 18850 -13440
rect 18970 -13560 19015 -13440
rect 19135 -13560 19180 -13440
rect 19300 -13560 19355 -13440
rect 19475 -13560 19520 -13440
rect 19640 -13560 19685 -13440
rect 19805 -13560 19850 -13440
rect 19970 -13560 20025 -13440
rect 20145 -13560 20190 -13440
rect 20310 -13560 20355 -13440
rect 20475 -13560 20520 -13440
rect 20640 -13560 20695 -13440
rect 20815 -13560 20860 -13440
rect 20980 -13560 21025 -13440
rect 21145 -13560 21190 -13440
rect 21310 -13560 21365 -13440
rect 21485 -13560 21530 -13440
rect 21650 -13560 21695 -13440
rect 21815 -13560 21860 -13440
rect 21980 -13560 22035 -13440
rect 22155 -13560 22200 -13440
rect 22320 -13560 22365 -13440
rect 22485 -13560 22530 -13440
rect 22650 -13560 22705 -13440
rect 22825 -13560 22870 -13440
rect 22990 -13560 23035 -13440
rect 23155 -13560 23200 -13440
rect 23320 -13560 23375 -13440
rect 23495 -13560 23540 -13440
rect 23660 -13560 23705 -13440
rect 23825 -13560 23870 -13440
rect 23990 -13560 24015 -13440
rect 18485 -13605 24015 -13560
rect 18485 -13725 18510 -13605
rect 18630 -13725 18685 -13605
rect 18805 -13725 18850 -13605
rect 18970 -13725 19015 -13605
rect 19135 -13725 19180 -13605
rect 19300 -13725 19355 -13605
rect 19475 -13725 19520 -13605
rect 19640 -13725 19685 -13605
rect 19805 -13725 19850 -13605
rect 19970 -13725 20025 -13605
rect 20145 -13725 20190 -13605
rect 20310 -13725 20355 -13605
rect 20475 -13725 20520 -13605
rect 20640 -13725 20695 -13605
rect 20815 -13725 20860 -13605
rect 20980 -13725 21025 -13605
rect 21145 -13725 21190 -13605
rect 21310 -13725 21365 -13605
rect 21485 -13725 21530 -13605
rect 21650 -13725 21695 -13605
rect 21815 -13725 21860 -13605
rect 21980 -13725 22035 -13605
rect 22155 -13725 22200 -13605
rect 22320 -13725 22365 -13605
rect 22485 -13725 22530 -13605
rect 22650 -13725 22705 -13605
rect 22825 -13725 22870 -13605
rect 22990 -13725 23035 -13605
rect 23155 -13725 23200 -13605
rect 23320 -13725 23375 -13605
rect 23495 -13725 23540 -13605
rect 23660 -13725 23705 -13605
rect 23825 -13725 23870 -13605
rect 23990 -13725 24015 -13605
rect 18485 -13770 24015 -13725
rect 18485 -13890 18510 -13770
rect 18630 -13890 18685 -13770
rect 18805 -13890 18850 -13770
rect 18970 -13890 19015 -13770
rect 19135 -13890 19180 -13770
rect 19300 -13890 19355 -13770
rect 19475 -13890 19520 -13770
rect 19640 -13890 19685 -13770
rect 19805 -13890 19850 -13770
rect 19970 -13890 20025 -13770
rect 20145 -13890 20190 -13770
rect 20310 -13890 20355 -13770
rect 20475 -13890 20520 -13770
rect 20640 -13890 20695 -13770
rect 20815 -13890 20860 -13770
rect 20980 -13890 21025 -13770
rect 21145 -13890 21190 -13770
rect 21310 -13890 21365 -13770
rect 21485 -13890 21530 -13770
rect 21650 -13890 21695 -13770
rect 21815 -13890 21860 -13770
rect 21980 -13890 22035 -13770
rect 22155 -13890 22200 -13770
rect 22320 -13890 22365 -13770
rect 22485 -13890 22530 -13770
rect 22650 -13890 22705 -13770
rect 22825 -13890 22870 -13770
rect 22990 -13890 23035 -13770
rect 23155 -13890 23200 -13770
rect 23320 -13890 23375 -13770
rect 23495 -13890 23540 -13770
rect 23660 -13890 23705 -13770
rect 23825 -13890 23870 -13770
rect 23990 -13890 24015 -13770
rect 18485 -13935 24015 -13890
rect 18485 -14055 18510 -13935
rect 18630 -14055 18685 -13935
rect 18805 -14055 18850 -13935
rect 18970 -14055 19015 -13935
rect 19135 -14055 19180 -13935
rect 19300 -14055 19355 -13935
rect 19475 -14055 19520 -13935
rect 19640 -14055 19685 -13935
rect 19805 -14055 19850 -13935
rect 19970 -14055 20025 -13935
rect 20145 -14055 20190 -13935
rect 20310 -14055 20355 -13935
rect 20475 -14055 20520 -13935
rect 20640 -14055 20695 -13935
rect 20815 -14055 20860 -13935
rect 20980 -14055 21025 -13935
rect 21145 -14055 21190 -13935
rect 21310 -14055 21365 -13935
rect 21485 -14055 21530 -13935
rect 21650 -14055 21695 -13935
rect 21815 -14055 21860 -13935
rect 21980 -14055 22035 -13935
rect 22155 -14055 22200 -13935
rect 22320 -14055 22365 -13935
rect 22485 -14055 22530 -13935
rect 22650 -14055 22705 -13935
rect 22825 -14055 22870 -13935
rect 22990 -14055 23035 -13935
rect 23155 -14055 23200 -13935
rect 23320 -14055 23375 -13935
rect 23495 -14055 23540 -13935
rect 23660 -14055 23705 -13935
rect 23825 -14055 23870 -13935
rect 23990 -14055 24015 -13935
rect 18485 -14110 24015 -14055
rect 18485 -14230 18510 -14110
rect 18630 -14230 18685 -14110
rect 18805 -14230 18850 -14110
rect 18970 -14230 19015 -14110
rect 19135 -14230 19180 -14110
rect 19300 -14230 19355 -14110
rect 19475 -14230 19520 -14110
rect 19640 -14230 19685 -14110
rect 19805 -14230 19850 -14110
rect 19970 -14230 20025 -14110
rect 20145 -14230 20190 -14110
rect 20310 -14230 20355 -14110
rect 20475 -14230 20520 -14110
rect 20640 -14230 20695 -14110
rect 20815 -14230 20860 -14110
rect 20980 -14230 21025 -14110
rect 21145 -14230 21190 -14110
rect 21310 -14230 21365 -14110
rect 21485 -14230 21530 -14110
rect 21650 -14230 21695 -14110
rect 21815 -14230 21860 -14110
rect 21980 -14230 22035 -14110
rect 22155 -14230 22200 -14110
rect 22320 -14230 22365 -14110
rect 22485 -14230 22530 -14110
rect 22650 -14230 22705 -14110
rect 22825 -14230 22870 -14110
rect 22990 -14230 23035 -14110
rect 23155 -14230 23200 -14110
rect 23320 -14230 23375 -14110
rect 23495 -14230 23540 -14110
rect 23660 -14230 23705 -14110
rect 23825 -14230 23870 -14110
rect 23990 -14230 24015 -14110
rect 18485 -14275 24015 -14230
rect 18485 -14395 18510 -14275
rect 18630 -14395 18685 -14275
rect 18805 -14395 18850 -14275
rect 18970 -14395 19015 -14275
rect 19135 -14395 19180 -14275
rect 19300 -14395 19355 -14275
rect 19475 -14395 19520 -14275
rect 19640 -14395 19685 -14275
rect 19805 -14395 19850 -14275
rect 19970 -14395 20025 -14275
rect 20145 -14395 20190 -14275
rect 20310 -14395 20355 -14275
rect 20475 -14395 20520 -14275
rect 20640 -14395 20695 -14275
rect 20815 -14395 20860 -14275
rect 20980 -14395 21025 -14275
rect 21145 -14395 21190 -14275
rect 21310 -14395 21365 -14275
rect 21485 -14395 21530 -14275
rect 21650 -14395 21695 -14275
rect 21815 -14395 21860 -14275
rect 21980 -14395 22035 -14275
rect 22155 -14395 22200 -14275
rect 22320 -14395 22365 -14275
rect 22485 -14395 22530 -14275
rect 22650 -14395 22705 -14275
rect 22825 -14395 22870 -14275
rect 22990 -14395 23035 -14275
rect 23155 -14395 23200 -14275
rect 23320 -14395 23375 -14275
rect 23495 -14395 23540 -14275
rect 23660 -14395 23705 -14275
rect 23825 -14395 23870 -14275
rect 23990 -14395 24015 -14275
rect 18485 -14440 24015 -14395
rect 18485 -14560 18510 -14440
rect 18630 -14560 18685 -14440
rect 18805 -14560 18850 -14440
rect 18970 -14560 19015 -14440
rect 19135 -14560 19180 -14440
rect 19300 -14560 19355 -14440
rect 19475 -14560 19520 -14440
rect 19640 -14560 19685 -14440
rect 19805 -14560 19850 -14440
rect 19970 -14560 20025 -14440
rect 20145 -14560 20190 -14440
rect 20310 -14560 20355 -14440
rect 20475 -14560 20520 -14440
rect 20640 -14560 20695 -14440
rect 20815 -14560 20860 -14440
rect 20980 -14560 21025 -14440
rect 21145 -14560 21190 -14440
rect 21310 -14560 21365 -14440
rect 21485 -14560 21530 -14440
rect 21650 -14560 21695 -14440
rect 21815 -14560 21860 -14440
rect 21980 -14560 22035 -14440
rect 22155 -14560 22200 -14440
rect 22320 -14560 22365 -14440
rect 22485 -14560 22530 -14440
rect 22650 -14560 22705 -14440
rect 22825 -14560 22870 -14440
rect 22990 -14560 23035 -14440
rect 23155 -14560 23200 -14440
rect 23320 -14560 23375 -14440
rect 23495 -14560 23540 -14440
rect 23660 -14560 23705 -14440
rect 23825 -14560 23870 -14440
rect 23990 -14560 24015 -14440
rect 18485 -14605 24015 -14560
rect 18485 -14725 18510 -14605
rect 18630 -14725 18685 -14605
rect 18805 -14725 18850 -14605
rect 18970 -14725 19015 -14605
rect 19135 -14725 19180 -14605
rect 19300 -14725 19355 -14605
rect 19475 -14725 19520 -14605
rect 19640 -14725 19685 -14605
rect 19805 -14725 19850 -14605
rect 19970 -14725 20025 -14605
rect 20145 -14725 20190 -14605
rect 20310 -14725 20355 -14605
rect 20475 -14725 20520 -14605
rect 20640 -14725 20695 -14605
rect 20815 -14725 20860 -14605
rect 20980 -14725 21025 -14605
rect 21145 -14725 21190 -14605
rect 21310 -14725 21365 -14605
rect 21485 -14725 21530 -14605
rect 21650 -14725 21695 -14605
rect 21815 -14725 21860 -14605
rect 21980 -14725 22035 -14605
rect 22155 -14725 22200 -14605
rect 22320 -14725 22365 -14605
rect 22485 -14725 22530 -14605
rect 22650 -14725 22705 -14605
rect 22825 -14725 22870 -14605
rect 22990 -14725 23035 -14605
rect 23155 -14725 23200 -14605
rect 23320 -14725 23375 -14605
rect 23495 -14725 23540 -14605
rect 23660 -14725 23705 -14605
rect 23825 -14725 23870 -14605
rect 23990 -14725 24015 -14605
rect 18485 -14780 24015 -14725
rect 18485 -14900 18510 -14780
rect 18630 -14900 18685 -14780
rect 18805 -14900 18850 -14780
rect 18970 -14900 19015 -14780
rect 19135 -14900 19180 -14780
rect 19300 -14900 19355 -14780
rect 19475 -14900 19520 -14780
rect 19640 -14900 19685 -14780
rect 19805 -14900 19850 -14780
rect 19970 -14900 20025 -14780
rect 20145 -14900 20190 -14780
rect 20310 -14900 20355 -14780
rect 20475 -14900 20520 -14780
rect 20640 -14900 20695 -14780
rect 20815 -14900 20860 -14780
rect 20980 -14900 21025 -14780
rect 21145 -14900 21190 -14780
rect 21310 -14900 21365 -14780
rect 21485 -14900 21530 -14780
rect 21650 -14900 21695 -14780
rect 21815 -14900 21860 -14780
rect 21980 -14900 22035 -14780
rect 22155 -14900 22200 -14780
rect 22320 -14900 22365 -14780
rect 22485 -14900 22530 -14780
rect 22650 -14900 22705 -14780
rect 22825 -14900 22870 -14780
rect 22990 -14900 23035 -14780
rect 23155 -14900 23200 -14780
rect 23320 -14900 23375 -14780
rect 23495 -14900 23540 -14780
rect 23660 -14900 23705 -14780
rect 23825 -14900 23870 -14780
rect 23990 -14900 24015 -14780
rect 18485 -14945 24015 -14900
rect 18485 -15065 18510 -14945
rect 18630 -15065 18685 -14945
rect 18805 -15065 18850 -14945
rect 18970 -15065 19015 -14945
rect 19135 -15065 19180 -14945
rect 19300 -15065 19355 -14945
rect 19475 -15065 19520 -14945
rect 19640 -15065 19685 -14945
rect 19805 -15065 19850 -14945
rect 19970 -15065 20025 -14945
rect 20145 -15065 20190 -14945
rect 20310 -15065 20355 -14945
rect 20475 -15065 20520 -14945
rect 20640 -15065 20695 -14945
rect 20815 -15065 20860 -14945
rect 20980 -15065 21025 -14945
rect 21145 -15065 21190 -14945
rect 21310 -15065 21365 -14945
rect 21485 -15065 21530 -14945
rect 21650 -15065 21695 -14945
rect 21815 -15065 21860 -14945
rect 21980 -15065 22035 -14945
rect 22155 -15065 22200 -14945
rect 22320 -15065 22365 -14945
rect 22485 -15065 22530 -14945
rect 22650 -15065 22705 -14945
rect 22825 -15065 22870 -14945
rect 22990 -15065 23035 -14945
rect 23155 -15065 23200 -14945
rect 23320 -15065 23375 -14945
rect 23495 -15065 23540 -14945
rect 23660 -15065 23705 -14945
rect 23825 -15065 23870 -14945
rect 23990 -15065 24015 -14945
rect 18485 -15110 24015 -15065
rect 18485 -15230 18510 -15110
rect 18630 -15230 18685 -15110
rect 18805 -15230 18850 -15110
rect 18970 -15230 19015 -15110
rect 19135 -15230 19180 -15110
rect 19300 -15230 19355 -15110
rect 19475 -15230 19520 -15110
rect 19640 -15230 19685 -15110
rect 19805 -15230 19850 -15110
rect 19970 -15230 20025 -15110
rect 20145 -15230 20190 -15110
rect 20310 -15230 20355 -15110
rect 20475 -15230 20520 -15110
rect 20640 -15230 20695 -15110
rect 20815 -15230 20860 -15110
rect 20980 -15230 21025 -15110
rect 21145 -15230 21190 -15110
rect 21310 -15230 21365 -15110
rect 21485 -15230 21530 -15110
rect 21650 -15230 21695 -15110
rect 21815 -15230 21860 -15110
rect 21980 -15230 22035 -15110
rect 22155 -15230 22200 -15110
rect 22320 -15230 22365 -15110
rect 22485 -15230 22530 -15110
rect 22650 -15230 22705 -15110
rect 22825 -15230 22870 -15110
rect 22990 -15230 23035 -15110
rect 23155 -15230 23200 -15110
rect 23320 -15230 23375 -15110
rect 23495 -15230 23540 -15110
rect 23660 -15230 23705 -15110
rect 23825 -15230 23870 -15110
rect 23990 -15230 24015 -15110
rect 18485 -15275 24015 -15230
rect 18485 -15395 18510 -15275
rect 18630 -15395 18685 -15275
rect 18805 -15395 18850 -15275
rect 18970 -15395 19015 -15275
rect 19135 -15395 19180 -15275
rect 19300 -15395 19355 -15275
rect 19475 -15395 19520 -15275
rect 19640 -15395 19685 -15275
rect 19805 -15395 19850 -15275
rect 19970 -15395 20025 -15275
rect 20145 -15395 20190 -15275
rect 20310 -15395 20355 -15275
rect 20475 -15395 20520 -15275
rect 20640 -15395 20695 -15275
rect 20815 -15395 20860 -15275
rect 20980 -15395 21025 -15275
rect 21145 -15395 21190 -15275
rect 21310 -15395 21365 -15275
rect 21485 -15395 21530 -15275
rect 21650 -15395 21695 -15275
rect 21815 -15395 21860 -15275
rect 21980 -15395 22035 -15275
rect 22155 -15395 22200 -15275
rect 22320 -15395 22365 -15275
rect 22485 -15395 22530 -15275
rect 22650 -15395 22705 -15275
rect 22825 -15395 22870 -15275
rect 22990 -15395 23035 -15275
rect 23155 -15395 23200 -15275
rect 23320 -15395 23375 -15275
rect 23495 -15395 23540 -15275
rect 23660 -15395 23705 -15275
rect 23825 -15395 23870 -15275
rect 23990 -15395 24015 -15275
rect 18485 -15450 24015 -15395
rect 18485 -15570 18510 -15450
rect 18630 -15570 18685 -15450
rect 18805 -15570 18850 -15450
rect 18970 -15570 19015 -15450
rect 19135 -15570 19180 -15450
rect 19300 -15570 19355 -15450
rect 19475 -15570 19520 -15450
rect 19640 -15570 19685 -15450
rect 19805 -15570 19850 -15450
rect 19970 -15570 20025 -15450
rect 20145 -15570 20190 -15450
rect 20310 -15570 20355 -15450
rect 20475 -15570 20520 -15450
rect 20640 -15570 20695 -15450
rect 20815 -15570 20860 -15450
rect 20980 -15570 21025 -15450
rect 21145 -15570 21190 -15450
rect 21310 -15570 21365 -15450
rect 21485 -15570 21530 -15450
rect 21650 -15570 21695 -15450
rect 21815 -15570 21860 -15450
rect 21980 -15570 22035 -15450
rect 22155 -15570 22200 -15450
rect 22320 -15570 22365 -15450
rect 22485 -15570 22530 -15450
rect 22650 -15570 22705 -15450
rect 22825 -15570 22870 -15450
rect 22990 -15570 23035 -15450
rect 23155 -15570 23200 -15450
rect 23320 -15570 23375 -15450
rect 23495 -15570 23540 -15450
rect 23660 -15570 23705 -15450
rect 23825 -15570 23870 -15450
rect 23990 -15570 24015 -15450
rect 18485 -15595 24015 -15570
rect 24175 -10090 29705 -10020
rect 24175 -10210 24200 -10090
rect 24320 -10210 24375 -10090
rect 24495 -10210 24540 -10090
rect 24660 -10210 24705 -10090
rect 24825 -10210 24870 -10090
rect 24990 -10210 25045 -10090
rect 25165 -10210 25210 -10090
rect 25330 -10210 25375 -10090
rect 25495 -10210 25540 -10090
rect 25660 -10210 25715 -10090
rect 25835 -10210 25880 -10090
rect 26000 -10210 26045 -10090
rect 26165 -10210 26210 -10090
rect 26330 -10210 26385 -10090
rect 26505 -10210 26550 -10090
rect 26670 -10210 26715 -10090
rect 26835 -10210 26880 -10090
rect 27000 -10210 27055 -10090
rect 27175 -10210 27220 -10090
rect 27340 -10210 27385 -10090
rect 27505 -10210 27550 -10090
rect 27670 -10210 27725 -10090
rect 27845 -10210 27890 -10090
rect 28010 -10210 28055 -10090
rect 28175 -10210 28220 -10090
rect 28340 -10210 28395 -10090
rect 28515 -10210 28560 -10090
rect 28680 -10210 28725 -10090
rect 28845 -10210 28890 -10090
rect 29010 -10210 29065 -10090
rect 29185 -10210 29230 -10090
rect 29350 -10210 29395 -10090
rect 29515 -10210 29560 -10090
rect 29680 -10210 29705 -10090
rect 24175 -10255 29705 -10210
rect 24175 -10375 24200 -10255
rect 24320 -10375 24375 -10255
rect 24495 -10375 24540 -10255
rect 24660 -10375 24705 -10255
rect 24825 -10375 24870 -10255
rect 24990 -10375 25045 -10255
rect 25165 -10375 25210 -10255
rect 25330 -10375 25375 -10255
rect 25495 -10375 25540 -10255
rect 25660 -10375 25715 -10255
rect 25835 -10375 25880 -10255
rect 26000 -10375 26045 -10255
rect 26165 -10375 26210 -10255
rect 26330 -10375 26385 -10255
rect 26505 -10375 26550 -10255
rect 26670 -10375 26715 -10255
rect 26835 -10375 26880 -10255
rect 27000 -10375 27055 -10255
rect 27175 -10375 27220 -10255
rect 27340 -10375 27385 -10255
rect 27505 -10375 27550 -10255
rect 27670 -10375 27725 -10255
rect 27845 -10375 27890 -10255
rect 28010 -10375 28055 -10255
rect 28175 -10375 28220 -10255
rect 28340 -10375 28395 -10255
rect 28515 -10375 28560 -10255
rect 28680 -10375 28725 -10255
rect 28845 -10375 28890 -10255
rect 29010 -10375 29065 -10255
rect 29185 -10375 29230 -10255
rect 29350 -10375 29395 -10255
rect 29515 -10375 29560 -10255
rect 29680 -10375 29705 -10255
rect 24175 -10420 29705 -10375
rect 24175 -10540 24200 -10420
rect 24320 -10540 24375 -10420
rect 24495 -10540 24540 -10420
rect 24660 -10540 24705 -10420
rect 24825 -10540 24870 -10420
rect 24990 -10540 25045 -10420
rect 25165 -10540 25210 -10420
rect 25330 -10540 25375 -10420
rect 25495 -10540 25540 -10420
rect 25660 -10540 25715 -10420
rect 25835 -10540 25880 -10420
rect 26000 -10540 26045 -10420
rect 26165 -10540 26210 -10420
rect 26330 -10540 26385 -10420
rect 26505 -10540 26550 -10420
rect 26670 -10540 26715 -10420
rect 26835 -10540 26880 -10420
rect 27000 -10540 27055 -10420
rect 27175 -10540 27220 -10420
rect 27340 -10540 27385 -10420
rect 27505 -10540 27550 -10420
rect 27670 -10540 27725 -10420
rect 27845 -10540 27890 -10420
rect 28010 -10540 28055 -10420
rect 28175 -10540 28220 -10420
rect 28340 -10540 28395 -10420
rect 28515 -10540 28560 -10420
rect 28680 -10540 28725 -10420
rect 28845 -10540 28890 -10420
rect 29010 -10540 29065 -10420
rect 29185 -10540 29230 -10420
rect 29350 -10540 29395 -10420
rect 29515 -10540 29560 -10420
rect 29680 -10540 29705 -10420
rect 24175 -10585 29705 -10540
rect 24175 -10705 24200 -10585
rect 24320 -10705 24375 -10585
rect 24495 -10705 24540 -10585
rect 24660 -10705 24705 -10585
rect 24825 -10705 24870 -10585
rect 24990 -10705 25045 -10585
rect 25165 -10705 25210 -10585
rect 25330 -10705 25375 -10585
rect 25495 -10705 25540 -10585
rect 25660 -10705 25715 -10585
rect 25835 -10705 25880 -10585
rect 26000 -10705 26045 -10585
rect 26165 -10705 26210 -10585
rect 26330 -10705 26385 -10585
rect 26505 -10705 26550 -10585
rect 26670 -10705 26715 -10585
rect 26835 -10705 26880 -10585
rect 27000 -10705 27055 -10585
rect 27175 -10705 27220 -10585
rect 27340 -10705 27385 -10585
rect 27505 -10705 27550 -10585
rect 27670 -10705 27725 -10585
rect 27845 -10705 27890 -10585
rect 28010 -10705 28055 -10585
rect 28175 -10705 28220 -10585
rect 28340 -10705 28395 -10585
rect 28515 -10705 28560 -10585
rect 28680 -10705 28725 -10585
rect 28845 -10705 28890 -10585
rect 29010 -10705 29065 -10585
rect 29185 -10705 29230 -10585
rect 29350 -10705 29395 -10585
rect 29515 -10705 29560 -10585
rect 29680 -10705 29705 -10585
rect 24175 -10760 29705 -10705
rect 24175 -10880 24200 -10760
rect 24320 -10880 24375 -10760
rect 24495 -10880 24540 -10760
rect 24660 -10880 24705 -10760
rect 24825 -10880 24870 -10760
rect 24990 -10880 25045 -10760
rect 25165 -10880 25210 -10760
rect 25330 -10880 25375 -10760
rect 25495 -10880 25540 -10760
rect 25660 -10880 25715 -10760
rect 25835 -10880 25880 -10760
rect 26000 -10880 26045 -10760
rect 26165 -10880 26210 -10760
rect 26330 -10880 26385 -10760
rect 26505 -10880 26550 -10760
rect 26670 -10880 26715 -10760
rect 26835 -10880 26880 -10760
rect 27000 -10880 27055 -10760
rect 27175 -10880 27220 -10760
rect 27340 -10880 27385 -10760
rect 27505 -10880 27550 -10760
rect 27670 -10880 27725 -10760
rect 27845 -10880 27890 -10760
rect 28010 -10880 28055 -10760
rect 28175 -10880 28220 -10760
rect 28340 -10880 28395 -10760
rect 28515 -10880 28560 -10760
rect 28680 -10880 28725 -10760
rect 28845 -10880 28890 -10760
rect 29010 -10880 29065 -10760
rect 29185 -10880 29230 -10760
rect 29350 -10880 29395 -10760
rect 29515 -10880 29560 -10760
rect 29680 -10880 29705 -10760
rect 24175 -10925 29705 -10880
rect 24175 -11045 24200 -10925
rect 24320 -11045 24375 -10925
rect 24495 -11045 24540 -10925
rect 24660 -11045 24705 -10925
rect 24825 -11045 24870 -10925
rect 24990 -11045 25045 -10925
rect 25165 -11045 25210 -10925
rect 25330 -11045 25375 -10925
rect 25495 -11045 25540 -10925
rect 25660 -11045 25715 -10925
rect 25835 -11045 25880 -10925
rect 26000 -11045 26045 -10925
rect 26165 -11045 26210 -10925
rect 26330 -11045 26385 -10925
rect 26505 -11045 26550 -10925
rect 26670 -11045 26715 -10925
rect 26835 -11045 26880 -10925
rect 27000 -11045 27055 -10925
rect 27175 -11045 27220 -10925
rect 27340 -11045 27385 -10925
rect 27505 -11045 27550 -10925
rect 27670 -11045 27725 -10925
rect 27845 -11045 27890 -10925
rect 28010 -11045 28055 -10925
rect 28175 -11045 28220 -10925
rect 28340 -11045 28395 -10925
rect 28515 -11045 28560 -10925
rect 28680 -11045 28725 -10925
rect 28845 -11045 28890 -10925
rect 29010 -11045 29065 -10925
rect 29185 -11045 29230 -10925
rect 29350 -11045 29395 -10925
rect 29515 -11045 29560 -10925
rect 29680 -11045 29705 -10925
rect 24175 -11090 29705 -11045
rect 24175 -11210 24200 -11090
rect 24320 -11210 24375 -11090
rect 24495 -11210 24540 -11090
rect 24660 -11210 24705 -11090
rect 24825 -11210 24870 -11090
rect 24990 -11210 25045 -11090
rect 25165 -11210 25210 -11090
rect 25330 -11210 25375 -11090
rect 25495 -11210 25540 -11090
rect 25660 -11210 25715 -11090
rect 25835 -11210 25880 -11090
rect 26000 -11210 26045 -11090
rect 26165 -11210 26210 -11090
rect 26330 -11210 26385 -11090
rect 26505 -11210 26550 -11090
rect 26670 -11210 26715 -11090
rect 26835 -11210 26880 -11090
rect 27000 -11210 27055 -11090
rect 27175 -11210 27220 -11090
rect 27340 -11210 27385 -11090
rect 27505 -11210 27550 -11090
rect 27670 -11210 27725 -11090
rect 27845 -11210 27890 -11090
rect 28010 -11210 28055 -11090
rect 28175 -11210 28220 -11090
rect 28340 -11210 28395 -11090
rect 28515 -11210 28560 -11090
rect 28680 -11210 28725 -11090
rect 28845 -11210 28890 -11090
rect 29010 -11210 29065 -11090
rect 29185 -11210 29230 -11090
rect 29350 -11210 29395 -11090
rect 29515 -11210 29560 -11090
rect 29680 -11210 29705 -11090
rect 24175 -11255 29705 -11210
rect 24175 -11375 24200 -11255
rect 24320 -11375 24375 -11255
rect 24495 -11375 24540 -11255
rect 24660 -11375 24705 -11255
rect 24825 -11375 24870 -11255
rect 24990 -11375 25045 -11255
rect 25165 -11375 25210 -11255
rect 25330 -11375 25375 -11255
rect 25495 -11375 25540 -11255
rect 25660 -11375 25715 -11255
rect 25835 -11375 25880 -11255
rect 26000 -11375 26045 -11255
rect 26165 -11375 26210 -11255
rect 26330 -11375 26385 -11255
rect 26505 -11375 26550 -11255
rect 26670 -11375 26715 -11255
rect 26835 -11375 26880 -11255
rect 27000 -11375 27055 -11255
rect 27175 -11375 27220 -11255
rect 27340 -11375 27385 -11255
rect 27505 -11375 27550 -11255
rect 27670 -11375 27725 -11255
rect 27845 -11375 27890 -11255
rect 28010 -11375 28055 -11255
rect 28175 -11375 28220 -11255
rect 28340 -11375 28395 -11255
rect 28515 -11375 28560 -11255
rect 28680 -11375 28725 -11255
rect 28845 -11375 28890 -11255
rect 29010 -11375 29065 -11255
rect 29185 -11375 29230 -11255
rect 29350 -11375 29395 -11255
rect 29515 -11375 29560 -11255
rect 29680 -11375 29705 -11255
rect 24175 -11430 29705 -11375
rect 24175 -11550 24200 -11430
rect 24320 -11550 24375 -11430
rect 24495 -11550 24540 -11430
rect 24660 -11550 24705 -11430
rect 24825 -11550 24870 -11430
rect 24990 -11550 25045 -11430
rect 25165 -11550 25210 -11430
rect 25330 -11550 25375 -11430
rect 25495 -11550 25540 -11430
rect 25660 -11550 25715 -11430
rect 25835 -11550 25880 -11430
rect 26000 -11550 26045 -11430
rect 26165 -11550 26210 -11430
rect 26330 -11550 26385 -11430
rect 26505 -11550 26550 -11430
rect 26670 -11550 26715 -11430
rect 26835 -11550 26880 -11430
rect 27000 -11550 27055 -11430
rect 27175 -11550 27220 -11430
rect 27340 -11550 27385 -11430
rect 27505 -11550 27550 -11430
rect 27670 -11550 27725 -11430
rect 27845 -11550 27890 -11430
rect 28010 -11550 28055 -11430
rect 28175 -11550 28220 -11430
rect 28340 -11550 28395 -11430
rect 28515 -11550 28560 -11430
rect 28680 -11550 28725 -11430
rect 28845 -11550 28890 -11430
rect 29010 -11550 29065 -11430
rect 29185 -11550 29230 -11430
rect 29350 -11550 29395 -11430
rect 29515 -11550 29560 -11430
rect 29680 -11550 29705 -11430
rect 24175 -11595 29705 -11550
rect 24175 -11715 24200 -11595
rect 24320 -11715 24375 -11595
rect 24495 -11715 24540 -11595
rect 24660 -11715 24705 -11595
rect 24825 -11715 24870 -11595
rect 24990 -11715 25045 -11595
rect 25165 -11715 25210 -11595
rect 25330 -11715 25375 -11595
rect 25495 -11715 25540 -11595
rect 25660 -11715 25715 -11595
rect 25835 -11715 25880 -11595
rect 26000 -11715 26045 -11595
rect 26165 -11715 26210 -11595
rect 26330 -11715 26385 -11595
rect 26505 -11715 26550 -11595
rect 26670 -11715 26715 -11595
rect 26835 -11715 26880 -11595
rect 27000 -11715 27055 -11595
rect 27175 -11715 27220 -11595
rect 27340 -11715 27385 -11595
rect 27505 -11715 27550 -11595
rect 27670 -11715 27725 -11595
rect 27845 -11715 27890 -11595
rect 28010 -11715 28055 -11595
rect 28175 -11715 28220 -11595
rect 28340 -11715 28395 -11595
rect 28515 -11715 28560 -11595
rect 28680 -11715 28725 -11595
rect 28845 -11715 28890 -11595
rect 29010 -11715 29065 -11595
rect 29185 -11715 29230 -11595
rect 29350 -11715 29395 -11595
rect 29515 -11715 29560 -11595
rect 29680 -11715 29705 -11595
rect 24175 -11760 29705 -11715
rect 24175 -11880 24200 -11760
rect 24320 -11880 24375 -11760
rect 24495 -11880 24540 -11760
rect 24660 -11880 24705 -11760
rect 24825 -11880 24870 -11760
rect 24990 -11880 25045 -11760
rect 25165 -11880 25210 -11760
rect 25330 -11880 25375 -11760
rect 25495 -11880 25540 -11760
rect 25660 -11880 25715 -11760
rect 25835 -11880 25880 -11760
rect 26000 -11880 26045 -11760
rect 26165 -11880 26210 -11760
rect 26330 -11880 26385 -11760
rect 26505 -11880 26550 -11760
rect 26670 -11880 26715 -11760
rect 26835 -11880 26880 -11760
rect 27000 -11880 27055 -11760
rect 27175 -11880 27220 -11760
rect 27340 -11880 27385 -11760
rect 27505 -11880 27550 -11760
rect 27670 -11880 27725 -11760
rect 27845 -11880 27890 -11760
rect 28010 -11880 28055 -11760
rect 28175 -11880 28220 -11760
rect 28340 -11880 28395 -11760
rect 28515 -11880 28560 -11760
rect 28680 -11880 28725 -11760
rect 28845 -11880 28890 -11760
rect 29010 -11880 29065 -11760
rect 29185 -11880 29230 -11760
rect 29350 -11880 29395 -11760
rect 29515 -11880 29560 -11760
rect 29680 -11880 29705 -11760
rect 24175 -11925 29705 -11880
rect 24175 -12045 24200 -11925
rect 24320 -12045 24375 -11925
rect 24495 -12045 24540 -11925
rect 24660 -12045 24705 -11925
rect 24825 -12045 24870 -11925
rect 24990 -12045 25045 -11925
rect 25165 -12045 25210 -11925
rect 25330 -12045 25375 -11925
rect 25495 -12045 25540 -11925
rect 25660 -12045 25715 -11925
rect 25835 -12045 25880 -11925
rect 26000 -12045 26045 -11925
rect 26165 -12045 26210 -11925
rect 26330 -12045 26385 -11925
rect 26505 -12045 26550 -11925
rect 26670 -12045 26715 -11925
rect 26835 -12045 26880 -11925
rect 27000 -12045 27055 -11925
rect 27175 -12045 27220 -11925
rect 27340 -12045 27385 -11925
rect 27505 -12045 27550 -11925
rect 27670 -12045 27725 -11925
rect 27845 -12045 27890 -11925
rect 28010 -12045 28055 -11925
rect 28175 -12045 28220 -11925
rect 28340 -12045 28395 -11925
rect 28515 -12045 28560 -11925
rect 28680 -12045 28725 -11925
rect 28845 -12045 28890 -11925
rect 29010 -12045 29065 -11925
rect 29185 -12045 29230 -11925
rect 29350 -12045 29395 -11925
rect 29515 -12045 29560 -11925
rect 29680 -12045 29705 -11925
rect 24175 -12100 29705 -12045
rect 24175 -12220 24200 -12100
rect 24320 -12220 24375 -12100
rect 24495 -12220 24540 -12100
rect 24660 -12220 24705 -12100
rect 24825 -12220 24870 -12100
rect 24990 -12220 25045 -12100
rect 25165 -12220 25210 -12100
rect 25330 -12220 25375 -12100
rect 25495 -12220 25540 -12100
rect 25660 -12220 25715 -12100
rect 25835 -12220 25880 -12100
rect 26000 -12220 26045 -12100
rect 26165 -12220 26210 -12100
rect 26330 -12220 26385 -12100
rect 26505 -12220 26550 -12100
rect 26670 -12220 26715 -12100
rect 26835 -12220 26880 -12100
rect 27000 -12220 27055 -12100
rect 27175 -12220 27220 -12100
rect 27340 -12220 27385 -12100
rect 27505 -12220 27550 -12100
rect 27670 -12220 27725 -12100
rect 27845 -12220 27890 -12100
rect 28010 -12220 28055 -12100
rect 28175 -12220 28220 -12100
rect 28340 -12220 28395 -12100
rect 28515 -12220 28560 -12100
rect 28680 -12220 28725 -12100
rect 28845 -12220 28890 -12100
rect 29010 -12220 29065 -12100
rect 29185 -12220 29230 -12100
rect 29350 -12220 29395 -12100
rect 29515 -12220 29560 -12100
rect 29680 -12220 29705 -12100
rect 24175 -12265 29705 -12220
rect 24175 -12385 24200 -12265
rect 24320 -12385 24375 -12265
rect 24495 -12385 24540 -12265
rect 24660 -12385 24705 -12265
rect 24825 -12385 24870 -12265
rect 24990 -12385 25045 -12265
rect 25165 -12385 25210 -12265
rect 25330 -12385 25375 -12265
rect 25495 -12385 25540 -12265
rect 25660 -12385 25715 -12265
rect 25835 -12385 25880 -12265
rect 26000 -12385 26045 -12265
rect 26165 -12385 26210 -12265
rect 26330 -12385 26385 -12265
rect 26505 -12385 26550 -12265
rect 26670 -12385 26715 -12265
rect 26835 -12385 26880 -12265
rect 27000 -12385 27055 -12265
rect 27175 -12385 27220 -12265
rect 27340 -12385 27385 -12265
rect 27505 -12385 27550 -12265
rect 27670 -12385 27725 -12265
rect 27845 -12385 27890 -12265
rect 28010 -12385 28055 -12265
rect 28175 -12385 28220 -12265
rect 28340 -12385 28395 -12265
rect 28515 -12385 28560 -12265
rect 28680 -12385 28725 -12265
rect 28845 -12385 28890 -12265
rect 29010 -12385 29065 -12265
rect 29185 -12385 29230 -12265
rect 29350 -12385 29395 -12265
rect 29515 -12385 29560 -12265
rect 29680 -12385 29705 -12265
rect 24175 -12430 29705 -12385
rect 24175 -12550 24200 -12430
rect 24320 -12550 24375 -12430
rect 24495 -12550 24540 -12430
rect 24660 -12550 24705 -12430
rect 24825 -12550 24870 -12430
rect 24990 -12550 25045 -12430
rect 25165 -12550 25210 -12430
rect 25330 -12550 25375 -12430
rect 25495 -12550 25540 -12430
rect 25660 -12550 25715 -12430
rect 25835 -12550 25880 -12430
rect 26000 -12550 26045 -12430
rect 26165 -12550 26210 -12430
rect 26330 -12550 26385 -12430
rect 26505 -12550 26550 -12430
rect 26670 -12550 26715 -12430
rect 26835 -12550 26880 -12430
rect 27000 -12550 27055 -12430
rect 27175 -12550 27220 -12430
rect 27340 -12550 27385 -12430
rect 27505 -12550 27550 -12430
rect 27670 -12550 27725 -12430
rect 27845 -12550 27890 -12430
rect 28010 -12550 28055 -12430
rect 28175 -12550 28220 -12430
rect 28340 -12550 28395 -12430
rect 28515 -12550 28560 -12430
rect 28680 -12550 28725 -12430
rect 28845 -12550 28890 -12430
rect 29010 -12550 29065 -12430
rect 29185 -12550 29230 -12430
rect 29350 -12550 29395 -12430
rect 29515 -12550 29560 -12430
rect 29680 -12550 29705 -12430
rect 24175 -12595 29705 -12550
rect 24175 -12715 24200 -12595
rect 24320 -12715 24375 -12595
rect 24495 -12715 24540 -12595
rect 24660 -12715 24705 -12595
rect 24825 -12715 24870 -12595
rect 24990 -12715 25045 -12595
rect 25165 -12715 25210 -12595
rect 25330 -12715 25375 -12595
rect 25495 -12715 25540 -12595
rect 25660 -12715 25715 -12595
rect 25835 -12715 25880 -12595
rect 26000 -12715 26045 -12595
rect 26165 -12715 26210 -12595
rect 26330 -12715 26385 -12595
rect 26505 -12715 26550 -12595
rect 26670 -12715 26715 -12595
rect 26835 -12715 26880 -12595
rect 27000 -12715 27055 -12595
rect 27175 -12715 27220 -12595
rect 27340 -12715 27385 -12595
rect 27505 -12715 27550 -12595
rect 27670 -12715 27725 -12595
rect 27845 -12715 27890 -12595
rect 28010 -12715 28055 -12595
rect 28175 -12715 28220 -12595
rect 28340 -12715 28395 -12595
rect 28515 -12715 28560 -12595
rect 28680 -12715 28725 -12595
rect 28845 -12715 28890 -12595
rect 29010 -12715 29065 -12595
rect 29185 -12715 29230 -12595
rect 29350 -12715 29395 -12595
rect 29515 -12715 29560 -12595
rect 29680 -12715 29705 -12595
rect 24175 -12770 29705 -12715
rect 24175 -12890 24200 -12770
rect 24320 -12890 24375 -12770
rect 24495 -12890 24540 -12770
rect 24660 -12890 24705 -12770
rect 24825 -12890 24870 -12770
rect 24990 -12890 25045 -12770
rect 25165 -12890 25210 -12770
rect 25330 -12890 25375 -12770
rect 25495 -12890 25540 -12770
rect 25660 -12890 25715 -12770
rect 25835 -12890 25880 -12770
rect 26000 -12890 26045 -12770
rect 26165 -12890 26210 -12770
rect 26330 -12890 26385 -12770
rect 26505 -12890 26550 -12770
rect 26670 -12890 26715 -12770
rect 26835 -12890 26880 -12770
rect 27000 -12890 27055 -12770
rect 27175 -12890 27220 -12770
rect 27340 -12890 27385 -12770
rect 27505 -12890 27550 -12770
rect 27670 -12890 27725 -12770
rect 27845 -12890 27890 -12770
rect 28010 -12890 28055 -12770
rect 28175 -12890 28220 -12770
rect 28340 -12890 28395 -12770
rect 28515 -12890 28560 -12770
rect 28680 -12890 28725 -12770
rect 28845 -12890 28890 -12770
rect 29010 -12890 29065 -12770
rect 29185 -12890 29230 -12770
rect 29350 -12890 29395 -12770
rect 29515 -12890 29560 -12770
rect 29680 -12890 29705 -12770
rect 24175 -12935 29705 -12890
rect 24175 -13055 24200 -12935
rect 24320 -13055 24375 -12935
rect 24495 -13055 24540 -12935
rect 24660 -13055 24705 -12935
rect 24825 -13055 24870 -12935
rect 24990 -13055 25045 -12935
rect 25165 -13055 25210 -12935
rect 25330 -13055 25375 -12935
rect 25495 -13055 25540 -12935
rect 25660 -13055 25715 -12935
rect 25835 -13055 25880 -12935
rect 26000 -13055 26045 -12935
rect 26165 -13055 26210 -12935
rect 26330 -13055 26385 -12935
rect 26505 -13055 26550 -12935
rect 26670 -13055 26715 -12935
rect 26835 -13055 26880 -12935
rect 27000 -13055 27055 -12935
rect 27175 -13055 27220 -12935
rect 27340 -13055 27385 -12935
rect 27505 -13055 27550 -12935
rect 27670 -13055 27725 -12935
rect 27845 -13055 27890 -12935
rect 28010 -13055 28055 -12935
rect 28175 -13055 28220 -12935
rect 28340 -13055 28395 -12935
rect 28515 -13055 28560 -12935
rect 28680 -13055 28725 -12935
rect 28845 -13055 28890 -12935
rect 29010 -13055 29065 -12935
rect 29185 -13055 29230 -12935
rect 29350 -13055 29395 -12935
rect 29515 -13055 29560 -12935
rect 29680 -13055 29705 -12935
rect 24175 -13100 29705 -13055
rect 24175 -13220 24200 -13100
rect 24320 -13220 24375 -13100
rect 24495 -13220 24540 -13100
rect 24660 -13220 24705 -13100
rect 24825 -13220 24870 -13100
rect 24990 -13220 25045 -13100
rect 25165 -13220 25210 -13100
rect 25330 -13220 25375 -13100
rect 25495 -13220 25540 -13100
rect 25660 -13220 25715 -13100
rect 25835 -13220 25880 -13100
rect 26000 -13220 26045 -13100
rect 26165 -13220 26210 -13100
rect 26330 -13220 26385 -13100
rect 26505 -13220 26550 -13100
rect 26670 -13220 26715 -13100
rect 26835 -13220 26880 -13100
rect 27000 -13220 27055 -13100
rect 27175 -13220 27220 -13100
rect 27340 -13220 27385 -13100
rect 27505 -13220 27550 -13100
rect 27670 -13220 27725 -13100
rect 27845 -13220 27890 -13100
rect 28010 -13220 28055 -13100
rect 28175 -13220 28220 -13100
rect 28340 -13220 28395 -13100
rect 28515 -13220 28560 -13100
rect 28680 -13220 28725 -13100
rect 28845 -13220 28890 -13100
rect 29010 -13220 29065 -13100
rect 29185 -13220 29230 -13100
rect 29350 -13220 29395 -13100
rect 29515 -13220 29560 -13100
rect 29680 -13220 29705 -13100
rect 24175 -13265 29705 -13220
rect 24175 -13385 24200 -13265
rect 24320 -13385 24375 -13265
rect 24495 -13385 24540 -13265
rect 24660 -13385 24705 -13265
rect 24825 -13385 24870 -13265
rect 24990 -13385 25045 -13265
rect 25165 -13385 25210 -13265
rect 25330 -13385 25375 -13265
rect 25495 -13385 25540 -13265
rect 25660 -13385 25715 -13265
rect 25835 -13385 25880 -13265
rect 26000 -13385 26045 -13265
rect 26165 -13385 26210 -13265
rect 26330 -13385 26385 -13265
rect 26505 -13385 26550 -13265
rect 26670 -13385 26715 -13265
rect 26835 -13385 26880 -13265
rect 27000 -13385 27055 -13265
rect 27175 -13385 27220 -13265
rect 27340 -13385 27385 -13265
rect 27505 -13385 27550 -13265
rect 27670 -13385 27725 -13265
rect 27845 -13385 27890 -13265
rect 28010 -13385 28055 -13265
rect 28175 -13385 28220 -13265
rect 28340 -13385 28395 -13265
rect 28515 -13385 28560 -13265
rect 28680 -13385 28725 -13265
rect 28845 -13385 28890 -13265
rect 29010 -13385 29065 -13265
rect 29185 -13385 29230 -13265
rect 29350 -13385 29395 -13265
rect 29515 -13385 29560 -13265
rect 29680 -13385 29705 -13265
rect 24175 -13440 29705 -13385
rect 24175 -13560 24200 -13440
rect 24320 -13560 24375 -13440
rect 24495 -13560 24540 -13440
rect 24660 -13560 24705 -13440
rect 24825 -13560 24870 -13440
rect 24990 -13560 25045 -13440
rect 25165 -13560 25210 -13440
rect 25330 -13560 25375 -13440
rect 25495 -13560 25540 -13440
rect 25660 -13560 25715 -13440
rect 25835 -13560 25880 -13440
rect 26000 -13560 26045 -13440
rect 26165 -13560 26210 -13440
rect 26330 -13560 26385 -13440
rect 26505 -13560 26550 -13440
rect 26670 -13560 26715 -13440
rect 26835 -13560 26880 -13440
rect 27000 -13560 27055 -13440
rect 27175 -13560 27220 -13440
rect 27340 -13560 27385 -13440
rect 27505 -13560 27550 -13440
rect 27670 -13560 27725 -13440
rect 27845 -13560 27890 -13440
rect 28010 -13560 28055 -13440
rect 28175 -13560 28220 -13440
rect 28340 -13560 28395 -13440
rect 28515 -13560 28560 -13440
rect 28680 -13560 28725 -13440
rect 28845 -13560 28890 -13440
rect 29010 -13560 29065 -13440
rect 29185 -13560 29230 -13440
rect 29350 -13560 29395 -13440
rect 29515 -13560 29560 -13440
rect 29680 -13560 29705 -13440
rect 24175 -13605 29705 -13560
rect 24175 -13725 24200 -13605
rect 24320 -13725 24375 -13605
rect 24495 -13725 24540 -13605
rect 24660 -13725 24705 -13605
rect 24825 -13725 24870 -13605
rect 24990 -13725 25045 -13605
rect 25165 -13725 25210 -13605
rect 25330 -13725 25375 -13605
rect 25495 -13725 25540 -13605
rect 25660 -13725 25715 -13605
rect 25835 -13725 25880 -13605
rect 26000 -13725 26045 -13605
rect 26165 -13725 26210 -13605
rect 26330 -13725 26385 -13605
rect 26505 -13725 26550 -13605
rect 26670 -13725 26715 -13605
rect 26835 -13725 26880 -13605
rect 27000 -13725 27055 -13605
rect 27175 -13725 27220 -13605
rect 27340 -13725 27385 -13605
rect 27505 -13725 27550 -13605
rect 27670 -13725 27725 -13605
rect 27845 -13725 27890 -13605
rect 28010 -13725 28055 -13605
rect 28175 -13725 28220 -13605
rect 28340 -13725 28395 -13605
rect 28515 -13725 28560 -13605
rect 28680 -13725 28725 -13605
rect 28845 -13725 28890 -13605
rect 29010 -13725 29065 -13605
rect 29185 -13725 29230 -13605
rect 29350 -13725 29395 -13605
rect 29515 -13725 29560 -13605
rect 29680 -13725 29705 -13605
rect 24175 -13770 29705 -13725
rect 24175 -13890 24200 -13770
rect 24320 -13890 24375 -13770
rect 24495 -13890 24540 -13770
rect 24660 -13890 24705 -13770
rect 24825 -13890 24870 -13770
rect 24990 -13890 25045 -13770
rect 25165 -13890 25210 -13770
rect 25330 -13890 25375 -13770
rect 25495 -13890 25540 -13770
rect 25660 -13890 25715 -13770
rect 25835 -13890 25880 -13770
rect 26000 -13890 26045 -13770
rect 26165 -13890 26210 -13770
rect 26330 -13890 26385 -13770
rect 26505 -13890 26550 -13770
rect 26670 -13890 26715 -13770
rect 26835 -13890 26880 -13770
rect 27000 -13890 27055 -13770
rect 27175 -13890 27220 -13770
rect 27340 -13890 27385 -13770
rect 27505 -13890 27550 -13770
rect 27670 -13890 27725 -13770
rect 27845 -13890 27890 -13770
rect 28010 -13890 28055 -13770
rect 28175 -13890 28220 -13770
rect 28340 -13890 28395 -13770
rect 28515 -13890 28560 -13770
rect 28680 -13890 28725 -13770
rect 28845 -13890 28890 -13770
rect 29010 -13890 29065 -13770
rect 29185 -13890 29230 -13770
rect 29350 -13890 29395 -13770
rect 29515 -13890 29560 -13770
rect 29680 -13890 29705 -13770
rect 24175 -13935 29705 -13890
rect 24175 -14055 24200 -13935
rect 24320 -14055 24375 -13935
rect 24495 -14055 24540 -13935
rect 24660 -14055 24705 -13935
rect 24825 -14055 24870 -13935
rect 24990 -14055 25045 -13935
rect 25165 -14055 25210 -13935
rect 25330 -14055 25375 -13935
rect 25495 -14055 25540 -13935
rect 25660 -14055 25715 -13935
rect 25835 -14055 25880 -13935
rect 26000 -14055 26045 -13935
rect 26165 -14055 26210 -13935
rect 26330 -14055 26385 -13935
rect 26505 -14055 26550 -13935
rect 26670 -14055 26715 -13935
rect 26835 -14055 26880 -13935
rect 27000 -14055 27055 -13935
rect 27175 -14055 27220 -13935
rect 27340 -14055 27385 -13935
rect 27505 -14055 27550 -13935
rect 27670 -14055 27725 -13935
rect 27845 -14055 27890 -13935
rect 28010 -14055 28055 -13935
rect 28175 -14055 28220 -13935
rect 28340 -14055 28395 -13935
rect 28515 -14055 28560 -13935
rect 28680 -14055 28725 -13935
rect 28845 -14055 28890 -13935
rect 29010 -14055 29065 -13935
rect 29185 -14055 29230 -13935
rect 29350 -14055 29395 -13935
rect 29515 -14055 29560 -13935
rect 29680 -14055 29705 -13935
rect 24175 -14110 29705 -14055
rect 24175 -14230 24200 -14110
rect 24320 -14230 24375 -14110
rect 24495 -14230 24540 -14110
rect 24660 -14230 24705 -14110
rect 24825 -14230 24870 -14110
rect 24990 -14230 25045 -14110
rect 25165 -14230 25210 -14110
rect 25330 -14230 25375 -14110
rect 25495 -14230 25540 -14110
rect 25660 -14230 25715 -14110
rect 25835 -14230 25880 -14110
rect 26000 -14230 26045 -14110
rect 26165 -14230 26210 -14110
rect 26330 -14230 26385 -14110
rect 26505 -14230 26550 -14110
rect 26670 -14230 26715 -14110
rect 26835 -14230 26880 -14110
rect 27000 -14230 27055 -14110
rect 27175 -14230 27220 -14110
rect 27340 -14230 27385 -14110
rect 27505 -14230 27550 -14110
rect 27670 -14230 27725 -14110
rect 27845 -14230 27890 -14110
rect 28010 -14230 28055 -14110
rect 28175 -14230 28220 -14110
rect 28340 -14230 28395 -14110
rect 28515 -14230 28560 -14110
rect 28680 -14230 28725 -14110
rect 28845 -14230 28890 -14110
rect 29010 -14230 29065 -14110
rect 29185 -14230 29230 -14110
rect 29350 -14230 29395 -14110
rect 29515 -14230 29560 -14110
rect 29680 -14230 29705 -14110
rect 24175 -14275 29705 -14230
rect 24175 -14395 24200 -14275
rect 24320 -14395 24375 -14275
rect 24495 -14395 24540 -14275
rect 24660 -14395 24705 -14275
rect 24825 -14395 24870 -14275
rect 24990 -14395 25045 -14275
rect 25165 -14395 25210 -14275
rect 25330 -14395 25375 -14275
rect 25495 -14395 25540 -14275
rect 25660 -14395 25715 -14275
rect 25835 -14395 25880 -14275
rect 26000 -14395 26045 -14275
rect 26165 -14395 26210 -14275
rect 26330 -14395 26385 -14275
rect 26505 -14395 26550 -14275
rect 26670 -14395 26715 -14275
rect 26835 -14395 26880 -14275
rect 27000 -14395 27055 -14275
rect 27175 -14395 27220 -14275
rect 27340 -14395 27385 -14275
rect 27505 -14395 27550 -14275
rect 27670 -14395 27725 -14275
rect 27845 -14395 27890 -14275
rect 28010 -14395 28055 -14275
rect 28175 -14395 28220 -14275
rect 28340 -14395 28395 -14275
rect 28515 -14395 28560 -14275
rect 28680 -14395 28725 -14275
rect 28845 -14395 28890 -14275
rect 29010 -14395 29065 -14275
rect 29185 -14395 29230 -14275
rect 29350 -14395 29395 -14275
rect 29515 -14395 29560 -14275
rect 29680 -14395 29705 -14275
rect 24175 -14440 29705 -14395
rect 24175 -14560 24200 -14440
rect 24320 -14560 24375 -14440
rect 24495 -14560 24540 -14440
rect 24660 -14560 24705 -14440
rect 24825 -14560 24870 -14440
rect 24990 -14560 25045 -14440
rect 25165 -14560 25210 -14440
rect 25330 -14560 25375 -14440
rect 25495 -14560 25540 -14440
rect 25660 -14560 25715 -14440
rect 25835 -14560 25880 -14440
rect 26000 -14560 26045 -14440
rect 26165 -14560 26210 -14440
rect 26330 -14560 26385 -14440
rect 26505 -14560 26550 -14440
rect 26670 -14560 26715 -14440
rect 26835 -14560 26880 -14440
rect 27000 -14560 27055 -14440
rect 27175 -14560 27220 -14440
rect 27340 -14560 27385 -14440
rect 27505 -14560 27550 -14440
rect 27670 -14560 27725 -14440
rect 27845 -14560 27890 -14440
rect 28010 -14560 28055 -14440
rect 28175 -14560 28220 -14440
rect 28340 -14560 28395 -14440
rect 28515 -14560 28560 -14440
rect 28680 -14560 28725 -14440
rect 28845 -14560 28890 -14440
rect 29010 -14560 29065 -14440
rect 29185 -14560 29230 -14440
rect 29350 -14560 29395 -14440
rect 29515 -14560 29560 -14440
rect 29680 -14560 29705 -14440
rect 24175 -14605 29705 -14560
rect 24175 -14725 24200 -14605
rect 24320 -14725 24375 -14605
rect 24495 -14725 24540 -14605
rect 24660 -14725 24705 -14605
rect 24825 -14725 24870 -14605
rect 24990 -14725 25045 -14605
rect 25165 -14725 25210 -14605
rect 25330 -14725 25375 -14605
rect 25495 -14725 25540 -14605
rect 25660 -14725 25715 -14605
rect 25835 -14725 25880 -14605
rect 26000 -14725 26045 -14605
rect 26165 -14725 26210 -14605
rect 26330 -14725 26385 -14605
rect 26505 -14725 26550 -14605
rect 26670 -14725 26715 -14605
rect 26835 -14725 26880 -14605
rect 27000 -14725 27055 -14605
rect 27175 -14725 27220 -14605
rect 27340 -14725 27385 -14605
rect 27505 -14725 27550 -14605
rect 27670 -14725 27725 -14605
rect 27845 -14725 27890 -14605
rect 28010 -14725 28055 -14605
rect 28175 -14725 28220 -14605
rect 28340 -14725 28395 -14605
rect 28515 -14725 28560 -14605
rect 28680 -14725 28725 -14605
rect 28845 -14725 28890 -14605
rect 29010 -14725 29065 -14605
rect 29185 -14725 29230 -14605
rect 29350 -14725 29395 -14605
rect 29515 -14725 29560 -14605
rect 29680 -14725 29705 -14605
rect 24175 -14780 29705 -14725
rect 24175 -14900 24200 -14780
rect 24320 -14900 24375 -14780
rect 24495 -14900 24540 -14780
rect 24660 -14900 24705 -14780
rect 24825 -14900 24870 -14780
rect 24990 -14900 25045 -14780
rect 25165 -14900 25210 -14780
rect 25330 -14900 25375 -14780
rect 25495 -14900 25540 -14780
rect 25660 -14900 25715 -14780
rect 25835 -14900 25880 -14780
rect 26000 -14900 26045 -14780
rect 26165 -14900 26210 -14780
rect 26330 -14900 26385 -14780
rect 26505 -14900 26550 -14780
rect 26670 -14900 26715 -14780
rect 26835 -14900 26880 -14780
rect 27000 -14900 27055 -14780
rect 27175 -14900 27220 -14780
rect 27340 -14900 27385 -14780
rect 27505 -14900 27550 -14780
rect 27670 -14900 27725 -14780
rect 27845 -14900 27890 -14780
rect 28010 -14900 28055 -14780
rect 28175 -14900 28220 -14780
rect 28340 -14900 28395 -14780
rect 28515 -14900 28560 -14780
rect 28680 -14900 28725 -14780
rect 28845 -14900 28890 -14780
rect 29010 -14900 29065 -14780
rect 29185 -14900 29230 -14780
rect 29350 -14900 29395 -14780
rect 29515 -14900 29560 -14780
rect 29680 -14900 29705 -14780
rect 24175 -14945 29705 -14900
rect 24175 -15065 24200 -14945
rect 24320 -15065 24375 -14945
rect 24495 -15065 24540 -14945
rect 24660 -15065 24705 -14945
rect 24825 -15065 24870 -14945
rect 24990 -15065 25045 -14945
rect 25165 -15065 25210 -14945
rect 25330 -15065 25375 -14945
rect 25495 -15065 25540 -14945
rect 25660 -15065 25715 -14945
rect 25835 -15065 25880 -14945
rect 26000 -15065 26045 -14945
rect 26165 -15065 26210 -14945
rect 26330 -15065 26385 -14945
rect 26505 -15065 26550 -14945
rect 26670 -15065 26715 -14945
rect 26835 -15065 26880 -14945
rect 27000 -15065 27055 -14945
rect 27175 -15065 27220 -14945
rect 27340 -15065 27385 -14945
rect 27505 -15065 27550 -14945
rect 27670 -15065 27725 -14945
rect 27845 -15065 27890 -14945
rect 28010 -15065 28055 -14945
rect 28175 -15065 28220 -14945
rect 28340 -15065 28395 -14945
rect 28515 -15065 28560 -14945
rect 28680 -15065 28725 -14945
rect 28845 -15065 28890 -14945
rect 29010 -15065 29065 -14945
rect 29185 -15065 29230 -14945
rect 29350 -15065 29395 -14945
rect 29515 -15065 29560 -14945
rect 29680 -15065 29705 -14945
rect 24175 -15110 29705 -15065
rect 24175 -15230 24200 -15110
rect 24320 -15230 24375 -15110
rect 24495 -15230 24540 -15110
rect 24660 -15230 24705 -15110
rect 24825 -15230 24870 -15110
rect 24990 -15230 25045 -15110
rect 25165 -15230 25210 -15110
rect 25330 -15230 25375 -15110
rect 25495 -15230 25540 -15110
rect 25660 -15230 25715 -15110
rect 25835 -15230 25880 -15110
rect 26000 -15230 26045 -15110
rect 26165 -15230 26210 -15110
rect 26330 -15230 26385 -15110
rect 26505 -15230 26550 -15110
rect 26670 -15230 26715 -15110
rect 26835 -15230 26880 -15110
rect 27000 -15230 27055 -15110
rect 27175 -15230 27220 -15110
rect 27340 -15230 27385 -15110
rect 27505 -15230 27550 -15110
rect 27670 -15230 27725 -15110
rect 27845 -15230 27890 -15110
rect 28010 -15230 28055 -15110
rect 28175 -15230 28220 -15110
rect 28340 -15230 28395 -15110
rect 28515 -15230 28560 -15110
rect 28680 -15230 28725 -15110
rect 28845 -15230 28890 -15110
rect 29010 -15230 29065 -15110
rect 29185 -15230 29230 -15110
rect 29350 -15230 29395 -15110
rect 29515 -15230 29560 -15110
rect 29680 -15230 29705 -15110
rect 24175 -15275 29705 -15230
rect 24175 -15395 24200 -15275
rect 24320 -15395 24375 -15275
rect 24495 -15395 24540 -15275
rect 24660 -15395 24705 -15275
rect 24825 -15395 24870 -15275
rect 24990 -15395 25045 -15275
rect 25165 -15395 25210 -15275
rect 25330 -15395 25375 -15275
rect 25495 -15395 25540 -15275
rect 25660 -15395 25715 -15275
rect 25835 -15395 25880 -15275
rect 26000 -15395 26045 -15275
rect 26165 -15395 26210 -15275
rect 26330 -15395 26385 -15275
rect 26505 -15395 26550 -15275
rect 26670 -15395 26715 -15275
rect 26835 -15395 26880 -15275
rect 27000 -15395 27055 -15275
rect 27175 -15395 27220 -15275
rect 27340 -15395 27385 -15275
rect 27505 -15395 27550 -15275
rect 27670 -15395 27725 -15275
rect 27845 -15395 27890 -15275
rect 28010 -15395 28055 -15275
rect 28175 -15395 28220 -15275
rect 28340 -15395 28395 -15275
rect 28515 -15395 28560 -15275
rect 28680 -15395 28725 -15275
rect 28845 -15395 28890 -15275
rect 29010 -15395 29065 -15275
rect 29185 -15395 29230 -15275
rect 29350 -15395 29395 -15275
rect 29515 -15395 29560 -15275
rect 29680 -15395 29705 -15275
rect 24175 -15450 29705 -15395
rect 24175 -15570 24200 -15450
rect 24320 -15570 24375 -15450
rect 24495 -15570 24540 -15450
rect 24660 -15570 24705 -15450
rect 24825 -15570 24870 -15450
rect 24990 -15570 25045 -15450
rect 25165 -15570 25210 -15450
rect 25330 -15570 25375 -15450
rect 25495 -15570 25540 -15450
rect 25660 -15570 25715 -15450
rect 25835 -15570 25880 -15450
rect 26000 -15570 26045 -15450
rect 26165 -15570 26210 -15450
rect 26330 -15570 26385 -15450
rect 26505 -15570 26550 -15450
rect 26670 -15570 26715 -15450
rect 26835 -15570 26880 -15450
rect 27000 -15570 27055 -15450
rect 27175 -15570 27220 -15450
rect 27340 -15570 27385 -15450
rect 27505 -15570 27550 -15450
rect 27670 -15570 27725 -15450
rect 27845 -15570 27890 -15450
rect 28010 -15570 28055 -15450
rect 28175 -15570 28220 -15450
rect 28340 -15570 28395 -15450
rect 28515 -15570 28560 -15450
rect 28680 -15570 28725 -15450
rect 28845 -15570 28890 -15450
rect 29010 -15570 29065 -15450
rect 29185 -15570 29230 -15450
rect 29350 -15570 29395 -15450
rect 29515 -15570 29560 -15450
rect 29680 -15570 29705 -15450
rect 24175 -15595 29705 -15570
<< end >>
