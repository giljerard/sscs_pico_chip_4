.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31]
+ wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23]
+ wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7]
+ wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31]
+ wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23]
+ wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7]
+ wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24]
+ wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8]
+ wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107]
+ la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100]
+ la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79]
+ la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72]
+ la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58]
+ la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51]
+ la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37]
+ la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16]
+ la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9]
+ la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123]
+ la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111]
+ la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98]
+ la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63]
+ la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35]
+ la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17] io_in[16] io_in[15]
+ io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4]
+ io_in[3] io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14]
+ io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6]
+ io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5]
+ io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22]
+ io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12]
+ io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] gpio_noesd[17]
+ gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10]
+ gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1]
+ io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127]
+ la_oenb[126] la_oenb[125] la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119]
+ la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94]
+ la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85]
+ la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68] la_oenb[67]
+ la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58]
+ la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49]
+ la_oenb[48] la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31]
+ la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22]
+ la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0]
*.iopin vdda1
*.iopin vdda2
*.iopin vssa1
*.iopin vssa2
*.iopin vccd1
*.iopin vccd2
*.iopin vssd1
*.iopin vssd2
*.ipin wb_clk_i
*.ipin wb_rst_i
*.ipin wbs_stb_i
*.ipin wbs_cyc_i
*.ipin wbs_we_i
*.ipin wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
*.ipin
*+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
*.ipin
*+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0]
*.opin wbs_ack_o
*.opin
*+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
*.ipin
*+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
*.opin
*+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
*.ipin
*+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
*.ipin
*+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0]
*.ipin user_clock2
*.opin
*+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
*.opin
*+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
*.iopin
*+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
*.iopin
*+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
*.iopin
*+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0]
*.iopin io_clamp_high[2],io_clamp_high[1],io_clamp_high[0]
*.iopin io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
*.opin user_irq[2],user_irq[1],user_irq[0]
*.ipin
*+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
x1 io_analog[6] io_analog[5] io_analog[2] io_analog[4] io_analog[1] io_analog[0] io_analog[3]
+ io_analog[9] io_analog[10] io_analog[8] io_analog[7] top
x2 io_analog[9] io_analog[10] big_cap
.ends

* expanding   symbol:  sscs_pico_chip_4/xschem/top.sym # of pins=11
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/top.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/top.sch
.subckt top  Iin_p Iin_n Vb1_ Vb2 Vb3_ Vb4_ Vb5 VDD GND Vout_n Vout_p
*.iopin VDD
*.iopin GND
*.opin Vout_n
*.ipin Iin_n
*.ipin Iin_p
*.ipin Vb1_
*.opin Vout_p
*.ipin Vb2
*.ipin Vb3_
*.ipin Vb4_
*.ipin Vb5
XR6 Vinn pre_Vout_p GND sky130_fd_pr__res_xhigh_po W=1.41 L=53 mult=1 m=1
XR1 pre_Vout_n Vinp GND sky130_fd_pr__res_xhigh_po W=1.41 L=53 mult=1 m=1
XR3 Vcm2 pre_Vout_p GND sky130_fd_pr__res_xhigh_po W=1.41 L=35 mult=1 m=1
XR5 pre_Vout_n Vcm2 GND sky130_fd_pr__res_xhigh_po W=1.41 L=35 mult=1 m=1
XR4 Vop net1 GND sky130_fd_pr__res_xhigh_po W=1.41 L=1.41 mult=1 m=1
XR10 Von net2 GND sky130_fd_pr__res_xhigh_po W=1.41 L=1.41 mult=1 m=1
XR17 Vcm1 Von GND sky130_fd_pr__res_xhigh_po W=1.41 L=35 mult=1 m=1
XR18 Vop Vcm1 GND sky130_fd_pr__res_xhigh_po W=1.41 L=35 mult=1 m=1
x1 Vinn Vinp Vb2 Vb1 Vcmfb1 VDD GND Vop Von core
x2 Vop Von Vb2 Vb1 Vcmfb2 VDD GND pre_Vout_n pre_Vout_p core
X1 VDD GND pre_Vout_n pre_Vout_p Vout_n Vout_p Vb4 sf
x3 Vcm1 Vb5 Vb3 VDD GND Vcmfb1 cmfb
x4 Vcm2 Vb5 Vb3 VDD GND Vcmfb2 cmfb
x5 Vb1 Vb1_ GND mirror_1
x6 Vb3 Vb3_ GND mirror_3
x7 Vb4 Vb4_ GND mirror_4
XC3 net1 pre_Vout_n sky130_fd_pr__cap_mim_m3_1 W=7.75 L=7.75 MF=1 m=1
XC4 pre_Vout_n net1 sky130_fd_pr__cap_mim_m3_2 W=7.75 L=7.75 MF=1 m=1
XC1 net2 pre_Vout_p sky130_fd_pr__cap_mim_m3_1 W=7.75 L=7.75 MF=1 m=1
XC2 pre_Vout_p net2 sky130_fd_pr__cap_mim_m3_2 W=7.75 L=7.75 MF=1 m=1
XC5 Vinn Iin_n sky130_fd_pr__cap_mim_m3_1 W=61.2 L=61.2 MF=1 m=1
XC6 Iin_n Vinn sky130_fd_pr__cap_mim_m3_2 W=61.2 L=61.2 MF=1 m=1
XC7 Vinp Iin_p sky130_fd_pr__cap_mim_m3_1 W=61.2 L=61.2 MF=1 m=1
XC8 Iin_p Vinp sky130_fd_pr__cap_mim_m3_2 W=61.2 L=61.2 MF=1 m=1
XC9 Vcmfb1 GND sky130_fd_pr__cap_mim_m3_1 W=33.5 L=33.5 MF=1 m=1
XC10 GND Vcmfb1 sky130_fd_pr__cap_mim_m3_2 W=33.5 L=33.5 MF=1 m=1
XC11 Vcmfb2 GND sky130_fd_pr__cap_mim_m3_1 W=33.5 L=33.5 MF=1 m=1
XC12 GND Vcmfb2 sky130_fd_pr__cap_mim_m3_2 W=33.5 L=33.5 MF=1 m=1
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/big_cap.sym # of pins=2
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/big_cap.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/big_cap.sch
.subckt big_cap  VDD GND
*.iopin VDD
*.iopin GND
XC5 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC6 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC1 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC2 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC3 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC4 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC7 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC8 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC9 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC10 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC11 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC12 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC13 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC14 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC15 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC16 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC17 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC18 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC19 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC20 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC21 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC22 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC23 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC24 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC25 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC26 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC27 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC28 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC29 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC30 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
XC31 VDD GND sky130_fd_pr__cap_mim_m3_1 W=55 L=55 MF=1 m=1
XC32 GND VDD sky130_fd_pr__cap_mim_m3_2 W=55 L=55 MF=1 m=1
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/core.sym # of pins=9
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/core.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/core.sch
.subckt core  Vin_n Vin_p Vb2 Vb1 Vcmfb VDD GND Vout_p Vout_n
*.ipin Vb2
*.ipin Vcmfb
*.iopin VDD
*.iopin GND
*.opin Vout_p
*.ipin Vin_p
*.ipin Vin_n
*.opin Vout_n
*.ipin Vb1
XM1 net1 Vb1 GND GND sky130_fd_pr__nfet_01v8 L=.5 W=710 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x1 Vin_p Vb2 Vcmfb VDD GND Vout_n net1 core_half
x2 Vin_n Vb2 Vcmfb VDD GND Vout_p net1 core_half
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/sf.sym # of pins=7
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/sf.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/sf.sch
.subckt sf  VDD GND Vin_p Vin_n Vout_p Vout_n Vb4
*.ipin Vin_n
*.iopin VDD
*.iopin GND
*.ipin Vin_p
*.opin Vout_n
*.opin Vout_p
*.iopin Vb4
X1 VDD Vb4 Vout_p Vin_p GND sf_half
X2 VDD Vb4 Vout_n Vin_n GND sf_half
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/cmfb.sym # of pins=6
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/cmfb.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/cmfb.sch
.subckt cmfb  Vcm Vref Vb3 VDD GND Vcmfb
*.iopin VDD
*.iopin GND
*.opin Vcmfb
*.ipin Vref
*.iopin Vb3
*.ipin Vcm
x1 Vref net2 VDD GND Vb3 net3 Vcmfb cmfb_half
x2 Vcm net1 VDD GND Vb3 net3 net3 cmfb_half
XR20 net2 net1 GND sky130_fd_pr__res_xhigh_po W=1.41 L=1.41 mult=1 m=1
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/mirror_1.sym # of pins=3
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/mirror_1.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/mirror_1.sch
.subckt mirror_1  Vb1 Vb1_ GND
*.iopin GND
*.iopin Vb1_
*.opin Vb1
XM27 Vb1_ Vb1_ GND GND sky130_fd_pr__nfet_01v8 L=.5 W=3.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC1 Vb1 GND sky130_fd_pr__cap_mim_m3_1 W=15.8 L=15.8 MF=1 m=1
XC2 GND Vb1 sky130_fd_pr__cap_mim_m3_2 W=15.8 L=15.8 MF=1 m=1
XR11 V10 Vb1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR1 Vb1_ V1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR2 V10 V9 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR3 V2 V1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR4 V8 V9 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR5 V2 V3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR6 V8 V7 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR7 V4 V3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR8 V6 V7 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR9 V4 V5 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR10 V6 V5 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XM1 GND GND Vb1_ GND sky130_fd_pr__nfet_01v8 L=.5 W=3.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 GND GND GND GND sky130_fd_pr__nfet_01v8 L=.5 W=3.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/mirror_3.sym # of pins=3
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/mirror_3.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/mirror_3.sch
.subckt mirror_3  Vb3 Vb3_ GND
*.iopin GND
*.iopin Vb3_
*.opin Vb3
XM27 Vb3_ Vb3_ GND GND sky130_fd_pr__nfet_01v8 L=.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XR11 V10 Vb3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XC1 Vb3 GND sky130_fd_pr__cap_mim_m3_1 W=15.8 L=15.8 MF=1 m=1
XC2 GND Vb3 sky130_fd_pr__cap_mim_m3_2 W=15.8 L=15.8 MF=1 m=1
XR1 Vb3_ V1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR2 V10 V9 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR3 V2 V1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR4 V8 V9 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR5 V2 V3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR6 V8 V7 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR7 V4 V3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR8 V6 V7 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR9 V4 V5 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR10 V6 V5 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XM1 GND GND GND GND sky130_fd_pr__nfet_01v8 L=.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 GND GND GND GND sky130_fd_pr__nfet_01v8 L=.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/mirror_4.sym # of pins=3
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/mirror_4.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/mirror_4.sch
.subckt mirror_4  Vb4 Vb4_ GND
*.iopin GND
*.iopin Vb4_
*.opin Vb4
XM27 Vb4_ Vb4_ GND GND sky130_fd_pr__nfet_01v8 L=.45 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC1 Vb4 GND sky130_fd_pr__cap_mim_m3_1 W=15.8 L=15.8 MF=1 m=1
XC2 GND Vb4 sky130_fd_pr__cap_mim_m3_2 W=15.8 L=15.8 MF=1 m=1
XR11 V10 Vb4 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR1 Vb4_ V1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR2 V10 V9 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR3 V2 V1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR4 V8 V9 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR5 V2 V3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR6 V8 V7 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR7 V4 V3 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR8 V6 V7 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR9 V4 V5 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XR10 V6 V5 GND sky130_fd_pr__res_xhigh_po W=0.35 L=16 mult=1 m=1
XM1 GND GND Vb4_ GND sky130_fd_pr__nfet_01v8 L=.45 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 GND GND GND GND sky130_fd_pr__nfet_01v8 L=.45 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/core_half.sym # of pins=7
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/core_half.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/core_half.sch
.subckt core_half  Vin Vb2 Vcmfb VDD GND Vout s
*.ipin Vb2
*.ipin Vcmfb
*.iopin VDD
*.iopin GND
*.opin Vout
*.iopin s
*.ipin Vin
XM3 Vout Vin s GND sky130_fd_pr__nfet_01v8 L=0.15 W=150 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 Vout Vcmfb VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=112 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM25 Vout Vb2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=448 nf=15 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/sf_half.sym # of pins=5
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/sf_half.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/sf_half.sch
.subckt sf_half  VDD g_d Vout g_u GND
*.iopin VDD
*.iopin g_u
*.iopin GND
*.iopin Vout
*.iopin g_d
XM17 VDD g_u Vout GND sky130_fd_pr__nfet_01v8_lvt L=0.32 W=650 nf=26 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM19 Vout g_d GND GND sky130_fd_pr__nfet_01v8 L=.45 W=650 nf=26 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sscs_pico_chip_4/xschem/cmfb_half.sym # of pins=7
* sym_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/cmfb_half.sym
* sch_path: /home/jared/Documents/GS_Design/sscs_pico_chip_4/xschem/cmfb_half.sch
.subckt cmfb_half  Vin res VDD GND Vb3 diode Vout
*.iopin VDD
*.iopin GND
*.opin Vout
*.ipin Vin
*.iopin diode
*.iopin Vb3
*.iopin res
XM11 Vout Vin res GND sky130_fd_pr__nfet_01v8 L=0.20 W=150 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM14 Vout diode VDD VDD sky130_fd_pr__pfet_01v8 L=0.2 W=42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 res Vb3 GND GND sky130_fd_pr__nfet_01v8 L=.5 W=65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
