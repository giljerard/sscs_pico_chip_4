magic
tech sky130A
timestamp 1636159292
<< nwell >>
rect -3670 -55 -660 1470
<< nmos >>
rect -3485 -200 -985 -185
rect -3485 -265 -985 -250
rect -3485 -330 -985 -315
rect -3485 -395 -985 -380
rect -3485 -460 -985 -445
rect -3485 -525 -985 -510
<< pmos >>
rect -3485 1342 -685 1360
rect -3485 1274 -685 1292
rect -3485 1206 -685 1224
rect -3485 1138 -685 1156
rect -3485 1070 -685 1088
rect -3485 1002 -685 1020
rect -3485 934 -685 952
rect -3485 866 -685 884
rect -3485 798 -685 816
rect -3485 730 -685 748
rect -3485 662 -685 680
rect -3485 594 -685 612
rect -3485 526 -685 544
rect -3485 458 -685 476
rect -3485 390 -685 408
rect -3485 322 -685 340
rect -3485 254 -685 272
rect -3485 186 -685 204
rect -3485 118 -685 136
rect -3485 50 -685 68
<< ndiff >>
rect -3485 -150 -985 -140
rect -3485 -170 -3470 -150
rect -3450 -170 -3430 -150
rect -3410 -170 -3390 -150
rect -3370 -170 -3350 -150
rect -3330 -170 -3310 -150
rect -3290 -170 -3270 -150
rect -3250 -170 -3230 -150
rect -3210 -170 -3190 -150
rect -3170 -170 -3150 -150
rect -3130 -170 -3110 -150
rect -3090 -170 -3070 -150
rect -3050 -170 -3030 -150
rect -3010 -170 -2990 -150
rect -2970 -170 -2950 -150
rect -2930 -170 -2910 -150
rect -2890 -170 -2870 -150
rect -2850 -170 -2830 -150
rect -2810 -170 -2790 -150
rect -2770 -170 -2750 -150
rect -2730 -170 -2710 -150
rect -2690 -170 -2670 -150
rect -2650 -170 -2630 -150
rect -2610 -170 -2590 -150
rect -2570 -170 -2550 -150
rect -2530 -170 -2510 -150
rect -2490 -170 -2470 -150
rect -2450 -170 -2430 -150
rect -2410 -170 -2390 -150
rect -2370 -170 -2350 -150
rect -2330 -170 -2310 -150
rect -2290 -170 -2270 -150
rect -2250 -170 -2230 -150
rect -2210 -170 -2190 -150
rect -2170 -170 -2150 -150
rect -2130 -170 -2110 -150
rect -2090 -170 -2070 -150
rect -2050 -170 -2030 -150
rect -2010 -170 -1990 -150
rect -1970 -170 -1950 -150
rect -1930 -170 -1910 -150
rect -1890 -170 -1870 -150
rect -1850 -170 -1830 -150
rect -1810 -170 -1790 -150
rect -1770 -170 -1750 -150
rect -1730 -170 -1710 -150
rect -1690 -170 -1670 -150
rect -1650 -170 -1630 -150
rect -1610 -170 -1590 -150
rect -1570 -170 -1550 -150
rect -1530 -170 -1510 -150
rect -1490 -170 -1470 -150
rect -1450 -170 -1430 -150
rect -1410 -170 -1390 -150
rect -1370 -170 -1350 -150
rect -1330 -170 -1310 -150
rect -1290 -170 -1270 -150
rect -1250 -170 -1230 -150
rect -1210 -170 -1190 -150
rect -1170 -170 -1150 -150
rect -1130 -170 -1110 -150
rect -1090 -170 -1070 -150
rect -1050 -170 -1030 -150
rect -1005 -170 -985 -150
rect -3485 -185 -985 -170
rect -3485 -215 -985 -200
rect -3485 -235 -3470 -215
rect -3450 -235 -3430 -215
rect -3410 -235 -3390 -215
rect -3370 -235 -3350 -215
rect -3330 -235 -3310 -215
rect -3290 -235 -3270 -215
rect -3250 -235 -3230 -215
rect -3210 -235 -3190 -215
rect -3170 -235 -3150 -215
rect -3130 -235 -3110 -215
rect -3090 -235 -3070 -215
rect -3050 -235 -3030 -215
rect -3010 -235 -2990 -215
rect -2970 -235 -2950 -215
rect -2930 -235 -2910 -215
rect -2890 -235 -2870 -215
rect -2850 -235 -2830 -215
rect -2810 -235 -2790 -215
rect -2770 -235 -2750 -215
rect -2730 -235 -2710 -215
rect -2690 -235 -2670 -215
rect -2650 -235 -2630 -215
rect -2610 -235 -2590 -215
rect -2570 -235 -2550 -215
rect -2530 -235 -2510 -215
rect -2490 -235 -2470 -215
rect -2450 -235 -2430 -215
rect -2410 -235 -2390 -215
rect -2370 -235 -2350 -215
rect -2330 -235 -2310 -215
rect -2290 -235 -2270 -215
rect -2250 -235 -2230 -215
rect -2210 -235 -2190 -215
rect -2170 -235 -2150 -215
rect -2130 -235 -2110 -215
rect -2090 -235 -2070 -215
rect -2050 -235 -2030 -215
rect -2010 -235 -1990 -215
rect -1970 -235 -1950 -215
rect -1930 -235 -1910 -215
rect -1890 -235 -1870 -215
rect -1850 -235 -1830 -215
rect -1810 -235 -1790 -215
rect -1770 -235 -1750 -215
rect -1730 -235 -1710 -215
rect -1690 -235 -1670 -215
rect -1650 -235 -1630 -215
rect -1610 -235 -1590 -215
rect -1570 -235 -1550 -215
rect -1530 -235 -1510 -215
rect -1490 -235 -1470 -215
rect -1450 -235 -1430 -215
rect -1410 -235 -1390 -215
rect -1370 -235 -1350 -215
rect -1330 -235 -1310 -215
rect -1290 -235 -1270 -215
rect -1250 -235 -1230 -215
rect -1210 -235 -1190 -215
rect -1170 -235 -1150 -215
rect -1130 -235 -1110 -215
rect -1090 -235 -1070 -215
rect -1050 -235 -1030 -215
rect -1005 -235 -985 -215
rect -3485 -250 -985 -235
rect -3485 -280 -985 -265
rect -3485 -300 -3470 -280
rect -3450 -300 -3430 -280
rect -3410 -300 -3390 -280
rect -3370 -300 -3350 -280
rect -3330 -300 -3310 -280
rect -3290 -300 -3270 -280
rect -3250 -300 -3230 -280
rect -3210 -300 -3190 -280
rect -3170 -300 -3150 -280
rect -3130 -300 -3110 -280
rect -3090 -300 -3070 -280
rect -3050 -300 -3030 -280
rect -3010 -300 -2990 -280
rect -2970 -300 -2950 -280
rect -2930 -300 -2910 -280
rect -2890 -300 -2870 -280
rect -2850 -300 -2830 -280
rect -2810 -300 -2790 -280
rect -2770 -300 -2750 -280
rect -2730 -300 -2710 -280
rect -2690 -300 -2670 -280
rect -2650 -300 -2630 -280
rect -2610 -300 -2590 -280
rect -2570 -300 -2550 -280
rect -2530 -300 -2510 -280
rect -2490 -300 -2470 -280
rect -2450 -300 -2430 -280
rect -2410 -300 -2390 -280
rect -2370 -300 -2350 -280
rect -2330 -300 -2310 -280
rect -2290 -300 -2270 -280
rect -2250 -300 -2230 -280
rect -2210 -300 -2190 -280
rect -2170 -300 -2150 -280
rect -2130 -300 -2110 -280
rect -2090 -300 -2070 -280
rect -2050 -300 -2030 -280
rect -2010 -300 -1990 -280
rect -1970 -300 -1950 -280
rect -1930 -300 -1910 -280
rect -1890 -300 -1870 -280
rect -1850 -300 -1830 -280
rect -1810 -300 -1790 -280
rect -1770 -300 -1750 -280
rect -1730 -300 -1710 -280
rect -1690 -300 -1670 -280
rect -1650 -300 -1630 -280
rect -1610 -300 -1590 -280
rect -1570 -300 -1550 -280
rect -1530 -300 -1510 -280
rect -1490 -300 -1470 -280
rect -1450 -300 -1430 -280
rect -1410 -300 -1390 -280
rect -1370 -300 -1350 -280
rect -1330 -300 -1310 -280
rect -1290 -300 -1270 -280
rect -1250 -300 -1230 -280
rect -1210 -300 -1190 -280
rect -1170 -300 -1150 -280
rect -1130 -300 -1110 -280
rect -1090 -300 -1070 -280
rect -1050 -300 -1030 -280
rect -1005 -300 -985 -280
rect -3485 -315 -985 -300
rect -3485 -345 -985 -330
rect -3485 -365 -3470 -345
rect -3450 -365 -3430 -345
rect -3410 -365 -3390 -345
rect -3370 -365 -3350 -345
rect -3330 -365 -3310 -345
rect -3290 -365 -3270 -345
rect -3250 -365 -3230 -345
rect -3210 -365 -3190 -345
rect -3170 -365 -3150 -345
rect -3130 -365 -3110 -345
rect -3090 -365 -3070 -345
rect -3050 -365 -3030 -345
rect -3010 -365 -2990 -345
rect -2970 -365 -2950 -345
rect -2930 -365 -2910 -345
rect -2890 -365 -2870 -345
rect -2850 -365 -2830 -345
rect -2810 -365 -2790 -345
rect -2770 -365 -2750 -345
rect -2730 -365 -2710 -345
rect -2690 -365 -2670 -345
rect -2650 -365 -2630 -345
rect -2610 -365 -2590 -345
rect -2570 -365 -2550 -345
rect -2530 -365 -2510 -345
rect -2490 -365 -2470 -345
rect -2450 -365 -2430 -345
rect -2410 -365 -2390 -345
rect -2370 -365 -2350 -345
rect -2330 -365 -2310 -345
rect -2290 -365 -2270 -345
rect -2250 -365 -2230 -345
rect -2210 -365 -2190 -345
rect -2170 -365 -2150 -345
rect -2130 -365 -2110 -345
rect -2090 -365 -2070 -345
rect -2050 -365 -2030 -345
rect -2010 -365 -1990 -345
rect -1970 -365 -1950 -345
rect -1930 -365 -1910 -345
rect -1890 -365 -1870 -345
rect -1850 -365 -1830 -345
rect -1810 -365 -1790 -345
rect -1770 -365 -1750 -345
rect -1730 -365 -1710 -345
rect -1690 -365 -1670 -345
rect -1650 -365 -1630 -345
rect -1610 -365 -1590 -345
rect -1570 -365 -1550 -345
rect -1530 -365 -1510 -345
rect -1490 -365 -1470 -345
rect -1450 -365 -1430 -345
rect -1410 -365 -1390 -345
rect -1370 -365 -1350 -345
rect -1330 -365 -1310 -345
rect -1290 -365 -1270 -345
rect -1250 -365 -1230 -345
rect -1210 -365 -1190 -345
rect -1170 -365 -1150 -345
rect -1130 -365 -1110 -345
rect -1090 -365 -1070 -345
rect -1050 -365 -1030 -345
rect -1005 -365 -985 -345
rect -3485 -380 -985 -365
rect -3485 -410 -985 -395
rect -3485 -430 -3470 -410
rect -3450 -430 -3430 -410
rect -3410 -430 -3390 -410
rect -3370 -430 -3350 -410
rect -3330 -430 -3310 -410
rect -3290 -430 -3270 -410
rect -3250 -430 -3230 -410
rect -3210 -430 -3190 -410
rect -3170 -430 -3150 -410
rect -3130 -430 -3110 -410
rect -3090 -430 -3070 -410
rect -3050 -430 -3030 -410
rect -3010 -430 -2990 -410
rect -2970 -430 -2950 -410
rect -2930 -430 -2910 -410
rect -2890 -430 -2870 -410
rect -2850 -430 -2830 -410
rect -2810 -430 -2790 -410
rect -2770 -430 -2750 -410
rect -2730 -430 -2710 -410
rect -2690 -430 -2670 -410
rect -2650 -430 -2630 -410
rect -2610 -430 -2590 -410
rect -2570 -430 -2550 -410
rect -2530 -430 -2510 -410
rect -2490 -430 -2470 -410
rect -2450 -430 -2430 -410
rect -2410 -430 -2390 -410
rect -2370 -430 -2350 -410
rect -2330 -430 -2310 -410
rect -2290 -430 -2270 -410
rect -2250 -430 -2230 -410
rect -2210 -430 -2190 -410
rect -2170 -430 -2150 -410
rect -2130 -430 -2110 -410
rect -2090 -430 -2070 -410
rect -2050 -430 -2030 -410
rect -2010 -430 -1990 -410
rect -1970 -430 -1950 -410
rect -1930 -430 -1910 -410
rect -1890 -430 -1870 -410
rect -1850 -430 -1830 -410
rect -1810 -430 -1790 -410
rect -1770 -430 -1750 -410
rect -1730 -430 -1710 -410
rect -1690 -430 -1670 -410
rect -1650 -430 -1630 -410
rect -1610 -430 -1590 -410
rect -1570 -430 -1550 -410
rect -1530 -430 -1510 -410
rect -1490 -430 -1470 -410
rect -1450 -430 -1430 -410
rect -1410 -430 -1390 -410
rect -1370 -430 -1350 -410
rect -1330 -430 -1310 -410
rect -1290 -430 -1270 -410
rect -1250 -430 -1230 -410
rect -1210 -430 -1190 -410
rect -1170 -430 -1150 -410
rect -1130 -430 -1110 -410
rect -1090 -430 -1070 -410
rect -1050 -430 -1030 -410
rect -1005 -430 -985 -410
rect -3485 -445 -985 -430
rect -3485 -475 -985 -460
rect -3485 -495 -3470 -475
rect -3450 -495 -3430 -475
rect -3410 -495 -3390 -475
rect -3370 -495 -3350 -475
rect -3330 -495 -3310 -475
rect -3290 -495 -3270 -475
rect -3250 -495 -3230 -475
rect -3210 -495 -3190 -475
rect -3170 -495 -3150 -475
rect -3130 -495 -3110 -475
rect -3090 -495 -3070 -475
rect -3050 -495 -3030 -475
rect -3010 -495 -2990 -475
rect -2970 -495 -2950 -475
rect -2930 -495 -2910 -475
rect -2890 -495 -2870 -475
rect -2850 -495 -2830 -475
rect -2810 -495 -2790 -475
rect -2770 -495 -2750 -475
rect -2730 -495 -2710 -475
rect -2690 -495 -2670 -475
rect -2650 -495 -2630 -475
rect -2610 -495 -2590 -475
rect -2570 -495 -2550 -475
rect -2530 -495 -2510 -475
rect -2490 -495 -2470 -475
rect -2450 -495 -2430 -475
rect -2410 -495 -2390 -475
rect -2370 -495 -2350 -475
rect -2330 -495 -2310 -475
rect -2290 -495 -2270 -475
rect -2250 -495 -2230 -475
rect -2210 -495 -2190 -475
rect -2170 -495 -2150 -475
rect -2130 -495 -2110 -475
rect -2090 -495 -2070 -475
rect -2050 -495 -2030 -475
rect -2010 -495 -1990 -475
rect -1970 -495 -1950 -475
rect -1930 -495 -1910 -475
rect -1890 -495 -1870 -475
rect -1850 -495 -1830 -475
rect -1810 -495 -1790 -475
rect -1770 -495 -1750 -475
rect -1730 -495 -1710 -475
rect -1690 -495 -1670 -475
rect -1650 -495 -1630 -475
rect -1610 -495 -1590 -475
rect -1570 -495 -1550 -475
rect -1530 -495 -1510 -475
rect -1490 -495 -1470 -475
rect -1450 -495 -1430 -475
rect -1410 -495 -1390 -475
rect -1370 -495 -1350 -475
rect -1330 -495 -1310 -475
rect -1290 -495 -1270 -475
rect -1250 -495 -1230 -475
rect -1210 -495 -1190 -475
rect -1170 -495 -1150 -475
rect -1130 -495 -1110 -475
rect -1090 -495 -1070 -475
rect -1050 -495 -1030 -475
rect -1005 -495 -985 -475
rect -3485 -510 -985 -495
rect -3485 -540 -985 -525
rect -3485 -560 -3470 -540
rect -3450 -560 -3430 -540
rect -3410 -560 -3390 -540
rect -3370 -560 -3350 -540
rect -3330 -560 -3310 -540
rect -3290 -560 -3270 -540
rect -3250 -560 -3230 -540
rect -3210 -560 -3190 -540
rect -3170 -560 -3150 -540
rect -3130 -560 -3110 -540
rect -3090 -560 -3070 -540
rect -3050 -560 -3030 -540
rect -3010 -560 -2990 -540
rect -2970 -560 -2950 -540
rect -2930 -560 -2910 -540
rect -2890 -560 -2870 -540
rect -2850 -560 -2830 -540
rect -2810 -560 -2790 -540
rect -2770 -560 -2750 -540
rect -2730 -560 -2710 -540
rect -2690 -560 -2670 -540
rect -2650 -560 -2630 -540
rect -2610 -560 -2590 -540
rect -2570 -560 -2550 -540
rect -2530 -560 -2510 -540
rect -2490 -560 -2470 -540
rect -2450 -560 -2430 -540
rect -2410 -560 -2390 -540
rect -2370 -560 -2350 -540
rect -2330 -560 -2310 -540
rect -2290 -560 -2270 -540
rect -2250 -560 -2230 -540
rect -2210 -560 -2190 -540
rect -2170 -560 -2150 -540
rect -2130 -560 -2110 -540
rect -2090 -560 -2070 -540
rect -2050 -560 -2030 -540
rect -2010 -560 -1990 -540
rect -1970 -560 -1950 -540
rect -1930 -560 -1910 -540
rect -1890 -560 -1870 -540
rect -1850 -560 -1830 -540
rect -1810 -560 -1790 -540
rect -1770 -560 -1750 -540
rect -1730 -560 -1710 -540
rect -1690 -560 -1670 -540
rect -1650 -560 -1630 -540
rect -1610 -560 -1590 -540
rect -1570 -560 -1550 -540
rect -1530 -560 -1510 -540
rect -1490 -560 -1470 -540
rect -1450 -560 -1430 -540
rect -1410 -560 -1390 -540
rect -1370 -560 -1350 -540
rect -1330 -560 -1310 -540
rect -1290 -560 -1270 -540
rect -1250 -560 -1230 -540
rect -1210 -560 -1190 -540
rect -1170 -560 -1150 -540
rect -1130 -560 -1110 -540
rect -1090 -560 -1070 -540
rect -1050 -560 -1030 -540
rect -1005 -560 -985 -540
rect -3485 -570 -985 -560
<< pdiff >>
rect -3485 1395 -685 1405
rect -3485 1375 -3470 1395
rect -3450 1375 -3430 1395
rect -3410 1375 -3390 1395
rect -3370 1375 -3350 1395
rect -3330 1375 -3310 1395
rect -3290 1375 -3270 1395
rect -3250 1375 -3230 1395
rect -3210 1375 -3190 1395
rect -3170 1375 -3150 1395
rect -3130 1375 -3110 1395
rect -3090 1375 -3070 1395
rect -3050 1375 -3030 1395
rect -3010 1375 -2990 1395
rect -2970 1375 -2950 1395
rect -2930 1375 -2910 1395
rect -2890 1375 -2870 1395
rect -2850 1375 -2830 1395
rect -2810 1375 -2790 1395
rect -2770 1375 -2750 1395
rect -2730 1375 -2710 1395
rect -2690 1375 -2670 1395
rect -2650 1375 -2630 1395
rect -2610 1375 -2590 1395
rect -2570 1375 -2550 1395
rect -2530 1375 -2510 1395
rect -2490 1375 -2470 1395
rect -2450 1375 -2430 1395
rect -2410 1375 -2390 1395
rect -2370 1375 -2350 1395
rect -2330 1375 -2310 1395
rect -2290 1375 -2270 1395
rect -2250 1375 -2230 1395
rect -2210 1375 -2190 1395
rect -2170 1375 -2150 1395
rect -2130 1375 -2110 1395
rect -2090 1375 -2070 1395
rect -2050 1375 -2030 1395
rect -2010 1375 -1990 1395
rect -1970 1375 -1950 1395
rect -1930 1375 -1910 1395
rect -1890 1375 -1870 1395
rect -1850 1375 -1830 1395
rect -1810 1375 -1790 1395
rect -1770 1375 -1750 1395
rect -1730 1375 -1710 1395
rect -1690 1375 -1670 1395
rect -1650 1375 -1630 1395
rect -1610 1375 -1590 1395
rect -1570 1375 -1550 1395
rect -1530 1375 -1510 1395
rect -1490 1375 -1470 1395
rect -1450 1375 -1430 1395
rect -1410 1375 -1390 1395
rect -1370 1375 -1350 1395
rect -1330 1375 -1310 1395
rect -1290 1375 -1270 1395
rect -1250 1375 -1230 1395
rect -1210 1375 -1190 1395
rect -1170 1375 -1150 1395
rect -1130 1375 -1110 1395
rect -1090 1375 -1070 1395
rect -1050 1375 -1030 1395
rect -1010 1375 -990 1395
rect -970 1375 -950 1395
rect -930 1375 -910 1395
rect -890 1375 -870 1395
rect -850 1375 -830 1395
rect -810 1375 -790 1395
rect -770 1375 -740 1395
rect -710 1375 -685 1395
rect -3485 1360 -685 1375
rect -3485 1327 -685 1342
rect -3485 1307 -3470 1327
rect -3450 1307 -3430 1327
rect -3410 1307 -3390 1327
rect -3370 1307 -3350 1327
rect -3330 1307 -3310 1327
rect -3290 1307 -3270 1327
rect -3250 1307 -3230 1327
rect -3210 1307 -3190 1327
rect -3170 1307 -3150 1327
rect -3130 1307 -3110 1327
rect -3090 1307 -3070 1327
rect -3050 1307 -3030 1327
rect -3010 1307 -2990 1327
rect -2970 1307 -2950 1327
rect -2930 1307 -2910 1327
rect -2890 1307 -2870 1327
rect -2850 1307 -2830 1327
rect -2810 1307 -2790 1327
rect -2770 1307 -2750 1327
rect -2730 1307 -2710 1327
rect -2690 1307 -2670 1327
rect -2650 1307 -2630 1327
rect -2610 1307 -2590 1327
rect -2570 1307 -2550 1327
rect -2530 1307 -2510 1327
rect -2490 1307 -2470 1327
rect -2450 1307 -2430 1327
rect -2410 1307 -2390 1327
rect -2370 1307 -2350 1327
rect -2330 1307 -2310 1327
rect -2290 1307 -2270 1327
rect -2250 1307 -2230 1327
rect -2210 1307 -2190 1327
rect -2170 1307 -2150 1327
rect -2130 1307 -2110 1327
rect -2090 1307 -2070 1327
rect -2050 1307 -2030 1327
rect -2010 1307 -1990 1327
rect -1970 1307 -1950 1327
rect -1930 1307 -1910 1327
rect -1890 1307 -1870 1327
rect -1850 1307 -1830 1327
rect -1810 1307 -1790 1327
rect -1770 1307 -1750 1327
rect -1730 1307 -1710 1327
rect -1690 1307 -1670 1327
rect -1650 1307 -1630 1327
rect -1610 1307 -1590 1327
rect -1570 1307 -1550 1327
rect -1530 1307 -1510 1327
rect -1490 1307 -1470 1327
rect -1450 1307 -1430 1327
rect -1410 1307 -1390 1327
rect -1370 1307 -1350 1327
rect -1330 1307 -1310 1327
rect -1290 1307 -1270 1327
rect -1250 1307 -1230 1327
rect -1210 1307 -1190 1327
rect -1170 1307 -1150 1327
rect -1130 1307 -1110 1327
rect -1090 1307 -1070 1327
rect -1050 1307 -1030 1327
rect -1010 1307 -990 1327
rect -970 1307 -950 1327
rect -930 1307 -910 1327
rect -890 1307 -870 1327
rect -850 1307 -830 1327
rect -810 1307 -790 1327
rect -770 1307 -740 1327
rect -710 1307 -685 1327
rect -3485 1292 -685 1307
rect -3485 1259 -685 1274
rect -3485 1239 -3470 1259
rect -3450 1239 -3430 1259
rect -3410 1239 -3390 1259
rect -3370 1239 -3350 1259
rect -3330 1239 -3310 1259
rect -3290 1239 -3270 1259
rect -3250 1239 -3230 1259
rect -3210 1239 -3190 1259
rect -3170 1239 -3150 1259
rect -3130 1239 -3110 1259
rect -3090 1239 -3070 1259
rect -3050 1239 -3030 1259
rect -3010 1239 -2990 1259
rect -2970 1239 -2950 1259
rect -2930 1239 -2910 1259
rect -2890 1239 -2870 1259
rect -2850 1239 -2830 1259
rect -2810 1239 -2790 1259
rect -2770 1239 -2750 1259
rect -2730 1239 -2710 1259
rect -2690 1239 -2670 1259
rect -2650 1239 -2630 1259
rect -2610 1239 -2590 1259
rect -2570 1239 -2550 1259
rect -2530 1239 -2510 1259
rect -2490 1239 -2470 1259
rect -2450 1239 -2430 1259
rect -2410 1239 -2390 1259
rect -2370 1239 -2350 1259
rect -2330 1239 -2310 1259
rect -2290 1239 -2270 1259
rect -2250 1239 -2230 1259
rect -2210 1239 -2190 1259
rect -2170 1239 -2150 1259
rect -2130 1239 -2110 1259
rect -2090 1239 -2070 1259
rect -2050 1239 -2030 1259
rect -2010 1239 -1990 1259
rect -1970 1239 -1950 1259
rect -1930 1239 -1910 1259
rect -1890 1239 -1870 1259
rect -1850 1239 -1830 1259
rect -1810 1239 -1790 1259
rect -1770 1239 -1750 1259
rect -1730 1239 -1710 1259
rect -1690 1239 -1670 1259
rect -1650 1239 -1630 1259
rect -1610 1239 -1590 1259
rect -1570 1239 -1550 1259
rect -1530 1239 -1510 1259
rect -1490 1239 -1470 1259
rect -1450 1239 -1430 1259
rect -1410 1239 -1390 1259
rect -1370 1239 -1350 1259
rect -1330 1239 -1310 1259
rect -1290 1239 -1270 1259
rect -1250 1239 -1230 1259
rect -1210 1239 -1190 1259
rect -1170 1239 -1150 1259
rect -1130 1239 -1110 1259
rect -1090 1239 -1070 1259
rect -1050 1239 -1030 1259
rect -1010 1239 -990 1259
rect -970 1239 -950 1259
rect -930 1239 -910 1259
rect -890 1239 -870 1259
rect -850 1239 -830 1259
rect -810 1239 -790 1259
rect -770 1239 -740 1259
rect -710 1239 -685 1259
rect -3485 1224 -685 1239
rect -3485 1191 -685 1206
rect -3485 1171 -3470 1191
rect -3450 1171 -3430 1191
rect -3410 1171 -3390 1191
rect -3370 1171 -3350 1191
rect -3330 1171 -3310 1191
rect -3290 1171 -3270 1191
rect -3250 1171 -3230 1191
rect -3210 1171 -3190 1191
rect -3170 1171 -3150 1191
rect -3130 1171 -3110 1191
rect -3090 1171 -3070 1191
rect -3050 1171 -3030 1191
rect -3010 1171 -2990 1191
rect -2970 1171 -2950 1191
rect -2930 1171 -2910 1191
rect -2890 1171 -2870 1191
rect -2850 1171 -2830 1191
rect -2810 1171 -2790 1191
rect -2770 1171 -2750 1191
rect -2730 1171 -2710 1191
rect -2690 1171 -2670 1191
rect -2650 1171 -2630 1191
rect -2610 1171 -2590 1191
rect -2570 1171 -2550 1191
rect -2530 1171 -2510 1191
rect -2490 1171 -2470 1191
rect -2450 1171 -2430 1191
rect -2410 1171 -2390 1191
rect -2370 1171 -2350 1191
rect -2330 1171 -2310 1191
rect -2290 1171 -2270 1191
rect -2250 1171 -2230 1191
rect -2210 1171 -2190 1191
rect -2170 1171 -2150 1191
rect -2130 1171 -2110 1191
rect -2090 1171 -2070 1191
rect -2050 1171 -2030 1191
rect -2010 1171 -1990 1191
rect -1970 1171 -1950 1191
rect -1930 1171 -1910 1191
rect -1890 1171 -1870 1191
rect -1850 1171 -1830 1191
rect -1810 1171 -1790 1191
rect -1770 1171 -1750 1191
rect -1730 1171 -1710 1191
rect -1690 1171 -1670 1191
rect -1650 1171 -1630 1191
rect -1610 1171 -1590 1191
rect -1570 1171 -1550 1191
rect -1530 1171 -1510 1191
rect -1490 1171 -1470 1191
rect -1450 1171 -1430 1191
rect -1410 1171 -1390 1191
rect -1370 1171 -1350 1191
rect -1330 1171 -1310 1191
rect -1290 1171 -1270 1191
rect -1250 1171 -1230 1191
rect -1210 1171 -1190 1191
rect -1170 1171 -1150 1191
rect -1130 1171 -1110 1191
rect -1090 1171 -1070 1191
rect -1050 1171 -1030 1191
rect -1010 1171 -990 1191
rect -970 1171 -950 1191
rect -930 1171 -910 1191
rect -890 1171 -870 1191
rect -850 1171 -830 1191
rect -810 1171 -790 1191
rect -770 1171 -740 1191
rect -710 1171 -685 1191
rect -3485 1156 -685 1171
rect -3485 1123 -685 1138
rect -3485 1103 -3470 1123
rect -3450 1103 -3430 1123
rect -3410 1103 -3390 1123
rect -3370 1103 -3350 1123
rect -3330 1103 -3310 1123
rect -3290 1103 -3270 1123
rect -3250 1103 -3230 1123
rect -3210 1103 -3190 1123
rect -3170 1103 -3150 1123
rect -3130 1103 -3110 1123
rect -3090 1103 -3070 1123
rect -3050 1103 -3030 1123
rect -3010 1103 -2990 1123
rect -2970 1103 -2950 1123
rect -2930 1103 -2910 1123
rect -2890 1103 -2870 1123
rect -2850 1103 -2830 1123
rect -2810 1103 -2790 1123
rect -2770 1103 -2750 1123
rect -2730 1103 -2710 1123
rect -2690 1103 -2670 1123
rect -2650 1103 -2630 1123
rect -2610 1103 -2590 1123
rect -2570 1103 -2550 1123
rect -2530 1103 -2510 1123
rect -2490 1103 -2470 1123
rect -2450 1103 -2430 1123
rect -2410 1103 -2390 1123
rect -2370 1103 -2350 1123
rect -2330 1103 -2310 1123
rect -2290 1103 -2270 1123
rect -2250 1103 -2230 1123
rect -2210 1103 -2190 1123
rect -2170 1103 -2150 1123
rect -2130 1103 -2110 1123
rect -2090 1103 -2070 1123
rect -2050 1103 -2030 1123
rect -2010 1103 -1990 1123
rect -1970 1103 -1950 1123
rect -1930 1103 -1910 1123
rect -1890 1103 -1870 1123
rect -1850 1103 -1830 1123
rect -1810 1103 -1790 1123
rect -1770 1103 -1750 1123
rect -1730 1103 -1710 1123
rect -1690 1103 -1670 1123
rect -1650 1103 -1630 1123
rect -1610 1103 -1590 1123
rect -1570 1103 -1550 1123
rect -1530 1103 -1510 1123
rect -1490 1103 -1470 1123
rect -1450 1103 -1430 1123
rect -1410 1103 -1390 1123
rect -1370 1103 -1350 1123
rect -1330 1103 -1310 1123
rect -1290 1103 -1270 1123
rect -1250 1103 -1230 1123
rect -1210 1103 -1190 1123
rect -1170 1103 -1150 1123
rect -1130 1103 -1110 1123
rect -1090 1103 -1070 1123
rect -1050 1103 -1030 1123
rect -1010 1103 -990 1123
rect -970 1103 -950 1123
rect -930 1103 -910 1123
rect -890 1103 -870 1123
rect -850 1103 -830 1123
rect -810 1103 -790 1123
rect -770 1103 -740 1123
rect -710 1103 -685 1123
rect -3485 1088 -685 1103
rect -3485 1055 -685 1070
rect -3485 1035 -3470 1055
rect -3450 1035 -3430 1055
rect -3410 1035 -3390 1055
rect -3370 1035 -3350 1055
rect -3330 1035 -3310 1055
rect -3290 1035 -3270 1055
rect -3250 1035 -3230 1055
rect -3210 1035 -3190 1055
rect -3170 1035 -3150 1055
rect -3130 1035 -3110 1055
rect -3090 1035 -3070 1055
rect -3050 1035 -3030 1055
rect -3010 1035 -2990 1055
rect -2970 1035 -2950 1055
rect -2930 1035 -2910 1055
rect -2890 1035 -2870 1055
rect -2850 1035 -2830 1055
rect -2810 1035 -2790 1055
rect -2770 1035 -2750 1055
rect -2730 1035 -2710 1055
rect -2690 1035 -2670 1055
rect -2650 1035 -2630 1055
rect -2610 1035 -2590 1055
rect -2570 1035 -2550 1055
rect -2530 1035 -2510 1055
rect -2490 1035 -2470 1055
rect -2450 1035 -2430 1055
rect -2410 1035 -2390 1055
rect -2370 1035 -2350 1055
rect -2330 1035 -2310 1055
rect -2290 1035 -2270 1055
rect -2250 1035 -2230 1055
rect -2210 1035 -2190 1055
rect -2170 1035 -2150 1055
rect -2130 1035 -2110 1055
rect -2090 1035 -2070 1055
rect -2050 1035 -2030 1055
rect -2010 1035 -1990 1055
rect -1970 1035 -1950 1055
rect -1930 1035 -1910 1055
rect -1890 1035 -1870 1055
rect -1850 1035 -1830 1055
rect -1810 1035 -1790 1055
rect -1770 1035 -1750 1055
rect -1730 1035 -1710 1055
rect -1690 1035 -1670 1055
rect -1650 1035 -1630 1055
rect -1610 1035 -1590 1055
rect -1570 1035 -1550 1055
rect -1530 1035 -1510 1055
rect -1490 1035 -1470 1055
rect -1450 1035 -1430 1055
rect -1410 1035 -1390 1055
rect -1370 1035 -1350 1055
rect -1330 1035 -1310 1055
rect -1290 1035 -1270 1055
rect -1250 1035 -1230 1055
rect -1210 1035 -1190 1055
rect -1170 1035 -1150 1055
rect -1130 1035 -1110 1055
rect -1090 1035 -1070 1055
rect -1050 1035 -1030 1055
rect -1010 1035 -990 1055
rect -970 1035 -950 1055
rect -930 1035 -910 1055
rect -890 1035 -870 1055
rect -850 1035 -830 1055
rect -810 1035 -790 1055
rect -770 1035 -740 1055
rect -710 1035 -685 1055
rect -3485 1020 -685 1035
rect -3485 987 -685 1002
rect -3485 967 -3470 987
rect -3450 967 -3430 987
rect -3410 967 -3390 987
rect -3370 967 -3350 987
rect -3330 967 -3310 987
rect -3290 967 -3270 987
rect -3250 967 -3230 987
rect -3210 967 -3190 987
rect -3170 967 -3150 987
rect -3130 967 -3110 987
rect -3090 967 -3070 987
rect -3050 967 -3030 987
rect -3010 967 -2990 987
rect -2970 967 -2950 987
rect -2930 967 -2910 987
rect -2890 967 -2870 987
rect -2850 967 -2830 987
rect -2810 967 -2790 987
rect -2770 967 -2750 987
rect -2730 967 -2710 987
rect -2690 967 -2670 987
rect -2650 967 -2630 987
rect -2610 967 -2590 987
rect -2570 967 -2550 987
rect -2530 967 -2510 987
rect -2490 967 -2470 987
rect -2450 967 -2430 987
rect -2410 967 -2390 987
rect -2370 967 -2350 987
rect -2330 967 -2310 987
rect -2290 967 -2270 987
rect -2250 967 -2230 987
rect -2210 967 -2190 987
rect -2170 967 -2150 987
rect -2130 967 -2110 987
rect -2090 967 -2070 987
rect -2050 967 -2030 987
rect -2010 967 -1990 987
rect -1970 967 -1950 987
rect -1930 967 -1910 987
rect -1890 967 -1870 987
rect -1850 967 -1830 987
rect -1810 967 -1790 987
rect -1770 967 -1750 987
rect -1730 967 -1710 987
rect -1690 967 -1670 987
rect -1650 967 -1630 987
rect -1610 967 -1590 987
rect -1570 967 -1550 987
rect -1530 967 -1510 987
rect -1490 967 -1470 987
rect -1450 967 -1430 987
rect -1410 967 -1390 987
rect -1370 967 -1350 987
rect -1330 967 -1310 987
rect -1290 967 -1270 987
rect -1250 967 -1230 987
rect -1210 967 -1190 987
rect -1170 967 -1150 987
rect -1130 967 -1110 987
rect -1090 967 -1070 987
rect -1050 967 -1030 987
rect -1010 967 -990 987
rect -970 967 -950 987
rect -930 967 -910 987
rect -890 967 -870 987
rect -850 967 -830 987
rect -810 967 -790 987
rect -770 967 -740 987
rect -710 967 -685 987
rect -3485 952 -685 967
rect -3485 919 -685 934
rect -3485 899 -3470 919
rect -3450 899 -3430 919
rect -3410 899 -3390 919
rect -3370 899 -3350 919
rect -3330 899 -3310 919
rect -3290 899 -3270 919
rect -3250 899 -3230 919
rect -3210 899 -3190 919
rect -3170 899 -3150 919
rect -3130 899 -3110 919
rect -3090 899 -3070 919
rect -3050 899 -3030 919
rect -3010 899 -2990 919
rect -2970 899 -2950 919
rect -2930 899 -2910 919
rect -2890 899 -2870 919
rect -2850 899 -2830 919
rect -2810 899 -2790 919
rect -2770 899 -2750 919
rect -2730 899 -2710 919
rect -2690 899 -2670 919
rect -2650 899 -2630 919
rect -2610 899 -2590 919
rect -2570 899 -2550 919
rect -2530 899 -2510 919
rect -2490 899 -2470 919
rect -2450 899 -2430 919
rect -2410 899 -2390 919
rect -2370 899 -2350 919
rect -2330 899 -2310 919
rect -2290 899 -2270 919
rect -2250 899 -2230 919
rect -2210 899 -2190 919
rect -2170 899 -2150 919
rect -2130 899 -2110 919
rect -2090 899 -2070 919
rect -2050 899 -2030 919
rect -2010 899 -1990 919
rect -1970 899 -1950 919
rect -1930 899 -1910 919
rect -1890 899 -1870 919
rect -1850 899 -1830 919
rect -1810 899 -1790 919
rect -1770 899 -1750 919
rect -1730 899 -1710 919
rect -1690 899 -1670 919
rect -1650 899 -1630 919
rect -1610 899 -1590 919
rect -1570 899 -1550 919
rect -1530 899 -1510 919
rect -1490 899 -1470 919
rect -1450 899 -1430 919
rect -1410 899 -1390 919
rect -1370 899 -1350 919
rect -1330 899 -1310 919
rect -1290 899 -1270 919
rect -1250 899 -1230 919
rect -1210 899 -1190 919
rect -1170 899 -1150 919
rect -1130 899 -1110 919
rect -1090 899 -1070 919
rect -1050 899 -1030 919
rect -1010 899 -990 919
rect -970 899 -950 919
rect -930 899 -910 919
rect -890 899 -870 919
rect -850 899 -830 919
rect -810 899 -790 919
rect -770 899 -740 919
rect -710 899 -685 919
rect -3485 884 -685 899
rect -3485 851 -685 866
rect -3485 831 -3470 851
rect -3450 831 -3430 851
rect -3410 831 -3390 851
rect -3370 831 -3350 851
rect -3330 831 -3310 851
rect -3290 831 -3270 851
rect -3250 831 -3230 851
rect -3210 831 -3190 851
rect -3170 831 -3150 851
rect -3130 831 -3110 851
rect -3090 831 -3070 851
rect -3050 831 -3030 851
rect -3010 831 -2990 851
rect -2970 831 -2950 851
rect -2930 831 -2910 851
rect -2890 831 -2870 851
rect -2850 831 -2830 851
rect -2810 831 -2790 851
rect -2770 831 -2750 851
rect -2730 831 -2710 851
rect -2690 831 -2670 851
rect -2650 831 -2630 851
rect -2610 831 -2590 851
rect -2570 831 -2550 851
rect -2530 831 -2510 851
rect -2490 831 -2470 851
rect -2450 831 -2430 851
rect -2410 831 -2390 851
rect -2370 831 -2350 851
rect -2330 831 -2310 851
rect -2290 831 -2270 851
rect -2250 831 -2230 851
rect -2210 831 -2190 851
rect -2170 831 -2150 851
rect -2130 831 -2110 851
rect -2090 831 -2070 851
rect -2050 831 -2030 851
rect -2010 831 -1990 851
rect -1970 831 -1950 851
rect -1930 831 -1910 851
rect -1890 831 -1870 851
rect -1850 831 -1830 851
rect -1810 831 -1790 851
rect -1770 831 -1750 851
rect -1730 831 -1710 851
rect -1690 831 -1670 851
rect -1650 831 -1630 851
rect -1610 831 -1590 851
rect -1570 831 -1550 851
rect -1530 831 -1510 851
rect -1490 831 -1470 851
rect -1450 831 -1430 851
rect -1410 831 -1390 851
rect -1370 831 -1350 851
rect -1330 831 -1310 851
rect -1290 831 -1270 851
rect -1250 831 -1230 851
rect -1210 831 -1190 851
rect -1170 831 -1150 851
rect -1130 831 -1110 851
rect -1090 831 -1070 851
rect -1050 831 -1030 851
rect -1010 831 -990 851
rect -970 831 -950 851
rect -930 831 -910 851
rect -890 831 -870 851
rect -850 831 -830 851
rect -810 831 -790 851
rect -770 831 -740 851
rect -710 831 -685 851
rect -3485 816 -685 831
rect -3485 783 -685 798
rect -3485 763 -3470 783
rect -3450 763 -3430 783
rect -3410 763 -3390 783
rect -3370 763 -3350 783
rect -3330 763 -3310 783
rect -3290 763 -3270 783
rect -3250 763 -3230 783
rect -3210 763 -3190 783
rect -3170 763 -3150 783
rect -3130 763 -3110 783
rect -3090 763 -3070 783
rect -3050 763 -3030 783
rect -3010 763 -2990 783
rect -2970 763 -2950 783
rect -2930 763 -2910 783
rect -2890 763 -2870 783
rect -2850 763 -2830 783
rect -2810 763 -2790 783
rect -2770 763 -2750 783
rect -2730 763 -2710 783
rect -2690 763 -2670 783
rect -2650 763 -2630 783
rect -2610 763 -2590 783
rect -2570 763 -2550 783
rect -2530 763 -2510 783
rect -2490 763 -2470 783
rect -2450 763 -2430 783
rect -2410 763 -2390 783
rect -2370 763 -2350 783
rect -2330 763 -2310 783
rect -2290 763 -2270 783
rect -2250 763 -2230 783
rect -2210 763 -2190 783
rect -2170 763 -2150 783
rect -2130 763 -2110 783
rect -2090 763 -2070 783
rect -2050 763 -2030 783
rect -2010 763 -1990 783
rect -1970 763 -1950 783
rect -1930 763 -1910 783
rect -1890 763 -1870 783
rect -1850 763 -1830 783
rect -1810 763 -1790 783
rect -1770 763 -1750 783
rect -1730 763 -1710 783
rect -1690 763 -1670 783
rect -1650 763 -1630 783
rect -1610 763 -1590 783
rect -1570 763 -1550 783
rect -1530 763 -1510 783
rect -1490 763 -1470 783
rect -1450 763 -1430 783
rect -1410 763 -1390 783
rect -1370 763 -1350 783
rect -1330 763 -1310 783
rect -1290 763 -1270 783
rect -1250 763 -1230 783
rect -1210 763 -1190 783
rect -1170 763 -1150 783
rect -1130 763 -1110 783
rect -1090 763 -1070 783
rect -1050 763 -1030 783
rect -1010 763 -990 783
rect -970 763 -950 783
rect -930 763 -910 783
rect -890 763 -870 783
rect -850 763 -830 783
rect -810 763 -790 783
rect -770 763 -740 783
rect -710 763 -685 783
rect -3485 748 -685 763
rect -3485 715 -685 730
rect -3485 695 -3470 715
rect -3450 695 -3430 715
rect -3410 695 -3390 715
rect -3370 695 -3350 715
rect -3330 695 -3310 715
rect -3290 695 -3270 715
rect -3250 695 -3230 715
rect -3210 695 -3190 715
rect -3170 695 -3150 715
rect -3130 695 -3110 715
rect -3090 695 -3070 715
rect -3050 695 -3030 715
rect -3010 695 -2990 715
rect -2970 695 -2950 715
rect -2930 695 -2910 715
rect -2890 695 -2870 715
rect -2850 695 -2830 715
rect -2810 695 -2790 715
rect -2770 695 -2750 715
rect -2730 695 -2710 715
rect -2690 695 -2670 715
rect -2650 695 -2630 715
rect -2610 695 -2590 715
rect -2570 695 -2550 715
rect -2530 695 -2510 715
rect -2490 695 -2470 715
rect -2450 695 -2430 715
rect -2410 695 -2390 715
rect -2370 695 -2350 715
rect -2330 695 -2310 715
rect -2290 695 -2270 715
rect -2250 695 -2230 715
rect -2210 695 -2190 715
rect -2170 695 -2150 715
rect -2130 695 -2110 715
rect -2090 695 -2070 715
rect -2050 695 -2030 715
rect -2010 695 -1990 715
rect -1970 695 -1950 715
rect -1930 695 -1910 715
rect -1890 695 -1870 715
rect -1850 695 -1830 715
rect -1810 695 -1790 715
rect -1770 695 -1750 715
rect -1730 695 -1710 715
rect -1690 695 -1670 715
rect -1650 695 -1630 715
rect -1610 695 -1590 715
rect -1570 695 -1550 715
rect -1530 695 -1510 715
rect -1490 695 -1470 715
rect -1450 695 -1430 715
rect -1410 695 -1390 715
rect -1370 695 -1350 715
rect -1330 695 -1310 715
rect -1290 695 -1270 715
rect -1250 695 -1230 715
rect -1210 695 -1190 715
rect -1170 695 -1150 715
rect -1130 695 -1110 715
rect -1090 695 -1070 715
rect -1050 695 -1030 715
rect -1010 695 -990 715
rect -970 695 -950 715
rect -930 695 -910 715
rect -890 695 -870 715
rect -850 695 -830 715
rect -810 695 -790 715
rect -770 695 -740 715
rect -710 695 -685 715
rect -3485 680 -685 695
rect -3485 647 -685 662
rect -3485 627 -3470 647
rect -3450 627 -3430 647
rect -3410 627 -3390 647
rect -3370 627 -3350 647
rect -3330 627 -3310 647
rect -3290 627 -3270 647
rect -3250 627 -3230 647
rect -3210 627 -3190 647
rect -3170 627 -3150 647
rect -3130 627 -3110 647
rect -3090 627 -3070 647
rect -3050 627 -3030 647
rect -3010 627 -2990 647
rect -2970 627 -2950 647
rect -2930 627 -2910 647
rect -2890 627 -2870 647
rect -2850 627 -2830 647
rect -2810 627 -2790 647
rect -2770 627 -2750 647
rect -2730 627 -2710 647
rect -2690 627 -2670 647
rect -2650 627 -2630 647
rect -2610 627 -2590 647
rect -2570 627 -2550 647
rect -2530 627 -2510 647
rect -2490 627 -2470 647
rect -2450 627 -2430 647
rect -2410 627 -2390 647
rect -2370 627 -2350 647
rect -2330 627 -2310 647
rect -2290 627 -2270 647
rect -2250 627 -2230 647
rect -2210 627 -2190 647
rect -2170 627 -2150 647
rect -2130 627 -2110 647
rect -2090 627 -2070 647
rect -2050 627 -2030 647
rect -2010 627 -1990 647
rect -1970 627 -1950 647
rect -1930 627 -1910 647
rect -1890 627 -1870 647
rect -1850 627 -1830 647
rect -1810 627 -1790 647
rect -1770 627 -1750 647
rect -1730 627 -1710 647
rect -1690 627 -1670 647
rect -1650 627 -1630 647
rect -1610 627 -1590 647
rect -1570 627 -1550 647
rect -1530 627 -1510 647
rect -1490 627 -1470 647
rect -1450 627 -1430 647
rect -1410 627 -1390 647
rect -1370 627 -1350 647
rect -1330 627 -1310 647
rect -1290 627 -1270 647
rect -1250 627 -1230 647
rect -1210 627 -1190 647
rect -1170 627 -1150 647
rect -1130 627 -1110 647
rect -1090 627 -1070 647
rect -1050 627 -1030 647
rect -1010 627 -990 647
rect -970 627 -950 647
rect -930 627 -910 647
rect -890 627 -870 647
rect -850 627 -830 647
rect -810 627 -790 647
rect -770 627 -740 647
rect -710 627 -685 647
rect -3485 612 -685 627
rect -3485 579 -685 594
rect -3485 559 -3470 579
rect -3450 559 -3430 579
rect -3410 559 -3390 579
rect -3370 559 -3350 579
rect -3330 559 -3310 579
rect -3290 559 -3270 579
rect -3250 559 -3230 579
rect -3210 559 -3190 579
rect -3170 559 -3150 579
rect -3130 559 -3110 579
rect -3090 559 -3070 579
rect -3050 559 -3030 579
rect -3010 559 -2990 579
rect -2970 559 -2950 579
rect -2930 559 -2910 579
rect -2890 559 -2870 579
rect -2850 559 -2830 579
rect -2810 559 -2790 579
rect -2770 559 -2750 579
rect -2730 559 -2710 579
rect -2690 559 -2670 579
rect -2650 559 -2630 579
rect -2610 559 -2590 579
rect -2570 559 -2550 579
rect -2530 559 -2510 579
rect -2490 559 -2470 579
rect -2450 559 -2430 579
rect -2410 559 -2390 579
rect -2370 559 -2350 579
rect -2330 559 -2310 579
rect -2290 559 -2270 579
rect -2250 559 -2230 579
rect -2210 559 -2190 579
rect -2170 559 -2150 579
rect -2130 559 -2110 579
rect -2090 559 -2070 579
rect -2050 559 -2030 579
rect -2010 559 -1990 579
rect -1970 559 -1950 579
rect -1930 559 -1910 579
rect -1890 559 -1870 579
rect -1850 559 -1830 579
rect -1810 559 -1790 579
rect -1770 559 -1750 579
rect -1730 559 -1710 579
rect -1690 559 -1670 579
rect -1650 559 -1630 579
rect -1610 559 -1590 579
rect -1570 559 -1550 579
rect -1530 559 -1510 579
rect -1490 559 -1470 579
rect -1450 559 -1430 579
rect -1410 559 -1390 579
rect -1370 559 -1350 579
rect -1330 559 -1310 579
rect -1290 559 -1270 579
rect -1250 559 -1230 579
rect -1210 559 -1190 579
rect -1170 559 -1150 579
rect -1130 559 -1110 579
rect -1090 559 -1070 579
rect -1050 559 -1030 579
rect -1010 559 -990 579
rect -970 559 -950 579
rect -930 559 -910 579
rect -890 559 -870 579
rect -850 559 -830 579
rect -810 559 -790 579
rect -770 559 -740 579
rect -710 559 -685 579
rect -3485 544 -685 559
rect -3485 511 -685 526
rect -3485 491 -3470 511
rect -3450 491 -3430 511
rect -3410 491 -3390 511
rect -3370 491 -3350 511
rect -3330 491 -3310 511
rect -3290 491 -3270 511
rect -3250 491 -3230 511
rect -3210 491 -3190 511
rect -3170 491 -3150 511
rect -3130 491 -3110 511
rect -3090 491 -3070 511
rect -3050 491 -3030 511
rect -3010 491 -2990 511
rect -2970 491 -2950 511
rect -2930 491 -2910 511
rect -2890 491 -2870 511
rect -2850 491 -2830 511
rect -2810 491 -2790 511
rect -2770 491 -2750 511
rect -2730 491 -2710 511
rect -2690 491 -2670 511
rect -2650 491 -2630 511
rect -2610 491 -2590 511
rect -2570 491 -2550 511
rect -2530 491 -2510 511
rect -2490 491 -2470 511
rect -2450 491 -2430 511
rect -2410 491 -2390 511
rect -2370 491 -2350 511
rect -2330 491 -2310 511
rect -2290 491 -2270 511
rect -2250 491 -2230 511
rect -2210 491 -2190 511
rect -2170 491 -2150 511
rect -2130 491 -2110 511
rect -2090 491 -2070 511
rect -2050 491 -2030 511
rect -2010 491 -1990 511
rect -1970 491 -1950 511
rect -1930 491 -1910 511
rect -1890 491 -1870 511
rect -1850 491 -1830 511
rect -1810 491 -1790 511
rect -1770 491 -1750 511
rect -1730 491 -1710 511
rect -1690 491 -1670 511
rect -1650 491 -1630 511
rect -1610 491 -1590 511
rect -1570 491 -1550 511
rect -1530 491 -1510 511
rect -1490 491 -1470 511
rect -1450 491 -1430 511
rect -1410 491 -1390 511
rect -1370 491 -1350 511
rect -1330 491 -1310 511
rect -1290 491 -1270 511
rect -1250 491 -1230 511
rect -1210 491 -1190 511
rect -1170 491 -1150 511
rect -1130 491 -1110 511
rect -1090 491 -1070 511
rect -1050 491 -1030 511
rect -1010 491 -990 511
rect -970 491 -950 511
rect -930 491 -910 511
rect -890 491 -870 511
rect -850 491 -830 511
rect -810 491 -790 511
rect -770 491 -740 511
rect -710 491 -685 511
rect -3485 476 -685 491
rect -3485 443 -685 458
rect -3485 423 -3470 443
rect -3450 423 -3430 443
rect -3410 423 -3390 443
rect -3370 423 -3350 443
rect -3330 423 -3310 443
rect -3290 423 -3270 443
rect -3250 423 -3230 443
rect -3210 423 -3190 443
rect -3170 423 -3150 443
rect -3130 423 -3110 443
rect -3090 423 -3070 443
rect -3050 423 -3030 443
rect -3010 423 -2990 443
rect -2970 423 -2950 443
rect -2930 423 -2910 443
rect -2890 423 -2870 443
rect -2850 423 -2830 443
rect -2810 423 -2790 443
rect -2770 423 -2750 443
rect -2730 423 -2710 443
rect -2690 423 -2670 443
rect -2650 423 -2630 443
rect -2610 423 -2590 443
rect -2570 423 -2550 443
rect -2530 423 -2510 443
rect -2490 423 -2470 443
rect -2450 423 -2430 443
rect -2410 423 -2390 443
rect -2370 423 -2350 443
rect -2330 423 -2310 443
rect -2290 423 -2270 443
rect -2250 423 -2230 443
rect -2210 423 -2190 443
rect -2170 423 -2150 443
rect -2130 423 -2110 443
rect -2090 423 -2070 443
rect -2050 423 -2030 443
rect -2010 423 -1990 443
rect -1970 423 -1950 443
rect -1930 423 -1910 443
rect -1890 423 -1870 443
rect -1850 423 -1830 443
rect -1810 423 -1790 443
rect -1770 423 -1750 443
rect -1730 423 -1710 443
rect -1690 423 -1670 443
rect -1650 423 -1630 443
rect -1610 423 -1590 443
rect -1570 423 -1550 443
rect -1530 423 -1510 443
rect -1490 423 -1470 443
rect -1450 423 -1430 443
rect -1410 423 -1390 443
rect -1370 423 -1350 443
rect -1330 423 -1310 443
rect -1290 423 -1270 443
rect -1250 423 -1230 443
rect -1210 423 -1190 443
rect -1170 423 -1150 443
rect -1130 423 -1110 443
rect -1090 423 -1070 443
rect -1050 423 -1030 443
rect -1010 423 -990 443
rect -970 423 -950 443
rect -930 423 -910 443
rect -890 423 -870 443
rect -850 423 -830 443
rect -810 423 -790 443
rect -770 423 -740 443
rect -710 423 -685 443
rect -3485 408 -685 423
rect -3485 375 -685 390
rect -3485 355 -3470 375
rect -3450 355 -3430 375
rect -3410 355 -3390 375
rect -3370 355 -3350 375
rect -3330 355 -3310 375
rect -3290 355 -3270 375
rect -3250 355 -3230 375
rect -3210 355 -3190 375
rect -3170 355 -3150 375
rect -3130 355 -3110 375
rect -3090 355 -3070 375
rect -3050 355 -3030 375
rect -3010 355 -2990 375
rect -2970 355 -2950 375
rect -2930 355 -2910 375
rect -2890 355 -2870 375
rect -2850 355 -2830 375
rect -2810 355 -2790 375
rect -2770 355 -2750 375
rect -2730 355 -2710 375
rect -2690 355 -2670 375
rect -2650 355 -2630 375
rect -2610 355 -2590 375
rect -2570 355 -2550 375
rect -2530 355 -2510 375
rect -2490 355 -2470 375
rect -2450 355 -2430 375
rect -2410 355 -2390 375
rect -2370 355 -2350 375
rect -2330 355 -2310 375
rect -2290 355 -2270 375
rect -2250 355 -2230 375
rect -2210 355 -2190 375
rect -2170 355 -2150 375
rect -2130 355 -2110 375
rect -2090 355 -2070 375
rect -2050 355 -2030 375
rect -2010 355 -1990 375
rect -1970 355 -1950 375
rect -1930 355 -1910 375
rect -1890 355 -1870 375
rect -1850 355 -1830 375
rect -1810 355 -1790 375
rect -1770 355 -1750 375
rect -1730 355 -1710 375
rect -1690 355 -1670 375
rect -1650 355 -1630 375
rect -1610 355 -1590 375
rect -1570 355 -1550 375
rect -1530 355 -1510 375
rect -1490 355 -1470 375
rect -1450 355 -1430 375
rect -1410 355 -1390 375
rect -1370 355 -1350 375
rect -1330 355 -1310 375
rect -1290 355 -1270 375
rect -1250 355 -1230 375
rect -1210 355 -1190 375
rect -1170 355 -1150 375
rect -1130 355 -1110 375
rect -1090 355 -1070 375
rect -1050 355 -1030 375
rect -1010 355 -990 375
rect -970 355 -950 375
rect -930 355 -910 375
rect -890 355 -870 375
rect -850 355 -830 375
rect -810 355 -790 375
rect -770 355 -740 375
rect -710 355 -685 375
rect -3485 340 -685 355
rect -3485 307 -685 322
rect -3485 287 -3470 307
rect -3450 287 -3430 307
rect -3410 287 -3390 307
rect -3370 287 -3350 307
rect -3330 287 -3310 307
rect -3290 287 -3270 307
rect -3250 287 -3230 307
rect -3210 287 -3190 307
rect -3170 287 -3150 307
rect -3130 287 -3110 307
rect -3090 287 -3070 307
rect -3050 287 -3030 307
rect -3010 287 -2990 307
rect -2970 287 -2950 307
rect -2930 287 -2910 307
rect -2890 287 -2870 307
rect -2850 287 -2830 307
rect -2810 287 -2790 307
rect -2770 287 -2750 307
rect -2730 287 -2710 307
rect -2690 287 -2670 307
rect -2650 287 -2630 307
rect -2610 287 -2590 307
rect -2570 287 -2550 307
rect -2530 287 -2510 307
rect -2490 287 -2470 307
rect -2450 287 -2430 307
rect -2410 287 -2390 307
rect -2370 287 -2350 307
rect -2330 287 -2310 307
rect -2290 287 -2270 307
rect -2250 287 -2230 307
rect -2210 287 -2190 307
rect -2170 287 -2150 307
rect -2130 287 -2110 307
rect -2090 287 -2070 307
rect -2050 287 -2030 307
rect -2010 287 -1990 307
rect -1970 287 -1950 307
rect -1930 287 -1910 307
rect -1890 287 -1870 307
rect -1850 287 -1830 307
rect -1810 287 -1790 307
rect -1770 287 -1750 307
rect -1730 287 -1710 307
rect -1690 287 -1670 307
rect -1650 287 -1630 307
rect -1610 287 -1590 307
rect -1570 287 -1550 307
rect -1530 287 -1510 307
rect -1490 287 -1470 307
rect -1450 287 -1430 307
rect -1410 287 -1390 307
rect -1370 287 -1350 307
rect -1330 287 -1310 307
rect -1290 287 -1270 307
rect -1250 287 -1230 307
rect -1210 287 -1190 307
rect -1170 287 -1150 307
rect -1130 287 -1110 307
rect -1090 287 -1070 307
rect -1050 287 -1030 307
rect -1010 287 -990 307
rect -970 287 -950 307
rect -930 287 -910 307
rect -890 287 -870 307
rect -850 287 -830 307
rect -810 287 -790 307
rect -770 287 -740 307
rect -710 287 -685 307
rect -3485 272 -685 287
rect -3485 239 -685 254
rect -3485 219 -3470 239
rect -3450 219 -3430 239
rect -3410 219 -3390 239
rect -3370 219 -3350 239
rect -3330 219 -3310 239
rect -3290 219 -3270 239
rect -3250 219 -3230 239
rect -3210 219 -3190 239
rect -3170 219 -3150 239
rect -3130 219 -3110 239
rect -3090 219 -3070 239
rect -3050 219 -3030 239
rect -3010 219 -2990 239
rect -2970 219 -2950 239
rect -2930 219 -2910 239
rect -2890 219 -2870 239
rect -2850 219 -2830 239
rect -2810 219 -2790 239
rect -2770 219 -2750 239
rect -2730 219 -2710 239
rect -2690 219 -2670 239
rect -2650 219 -2630 239
rect -2610 219 -2590 239
rect -2570 219 -2550 239
rect -2530 219 -2510 239
rect -2490 219 -2470 239
rect -2450 219 -2430 239
rect -2410 219 -2390 239
rect -2370 219 -2350 239
rect -2330 219 -2310 239
rect -2290 219 -2270 239
rect -2250 219 -2230 239
rect -2210 219 -2190 239
rect -2170 219 -2150 239
rect -2130 219 -2110 239
rect -2090 219 -2070 239
rect -2050 219 -2030 239
rect -2010 219 -1990 239
rect -1970 219 -1950 239
rect -1930 219 -1910 239
rect -1890 219 -1870 239
rect -1850 219 -1830 239
rect -1810 219 -1790 239
rect -1770 219 -1750 239
rect -1730 219 -1710 239
rect -1690 219 -1670 239
rect -1650 219 -1630 239
rect -1610 219 -1590 239
rect -1570 219 -1550 239
rect -1530 219 -1510 239
rect -1490 219 -1470 239
rect -1450 219 -1430 239
rect -1410 219 -1390 239
rect -1370 219 -1350 239
rect -1330 219 -1310 239
rect -1290 219 -1270 239
rect -1250 219 -1230 239
rect -1210 219 -1190 239
rect -1170 219 -1150 239
rect -1130 219 -1110 239
rect -1090 219 -1070 239
rect -1050 219 -1030 239
rect -1010 219 -990 239
rect -970 219 -950 239
rect -930 219 -910 239
rect -890 219 -870 239
rect -850 219 -830 239
rect -810 219 -790 239
rect -770 219 -740 239
rect -710 219 -685 239
rect -3485 204 -685 219
rect -3485 171 -685 186
rect -3485 151 -3470 171
rect -3450 151 -3430 171
rect -3410 151 -3390 171
rect -3370 151 -3350 171
rect -3330 151 -3310 171
rect -3290 151 -3270 171
rect -3250 151 -3230 171
rect -3210 151 -3190 171
rect -3170 151 -3150 171
rect -3130 151 -3110 171
rect -3090 151 -3070 171
rect -3050 151 -3030 171
rect -3010 151 -2990 171
rect -2970 151 -2950 171
rect -2930 151 -2910 171
rect -2890 151 -2870 171
rect -2850 151 -2830 171
rect -2810 151 -2790 171
rect -2770 151 -2750 171
rect -2730 151 -2710 171
rect -2690 151 -2670 171
rect -2650 151 -2630 171
rect -2610 151 -2590 171
rect -2570 151 -2550 171
rect -2530 151 -2510 171
rect -2490 151 -2470 171
rect -2450 151 -2430 171
rect -2410 151 -2390 171
rect -2370 151 -2350 171
rect -2330 151 -2310 171
rect -2290 151 -2270 171
rect -2250 151 -2230 171
rect -2210 151 -2190 171
rect -2170 151 -2150 171
rect -2130 151 -2110 171
rect -2090 151 -2070 171
rect -2050 151 -2030 171
rect -2010 151 -1990 171
rect -1970 151 -1950 171
rect -1930 151 -1910 171
rect -1890 151 -1870 171
rect -1850 151 -1830 171
rect -1810 151 -1790 171
rect -1770 151 -1750 171
rect -1730 151 -1710 171
rect -1690 151 -1670 171
rect -1650 151 -1630 171
rect -1610 151 -1590 171
rect -1570 151 -1550 171
rect -1530 151 -1510 171
rect -1490 151 -1470 171
rect -1450 151 -1430 171
rect -1410 151 -1390 171
rect -1370 151 -1350 171
rect -1330 151 -1310 171
rect -1290 151 -1270 171
rect -1250 151 -1230 171
rect -1210 151 -1190 171
rect -1170 151 -1150 171
rect -1130 151 -1110 171
rect -1090 151 -1070 171
rect -1050 151 -1030 171
rect -1010 151 -990 171
rect -970 151 -950 171
rect -930 151 -910 171
rect -890 151 -870 171
rect -850 151 -830 171
rect -810 151 -790 171
rect -770 151 -740 171
rect -710 151 -685 171
rect -3485 136 -685 151
rect -3485 103 -685 118
rect -3485 83 -3470 103
rect -3450 83 -3430 103
rect -3410 83 -3390 103
rect -3370 83 -3350 103
rect -3330 83 -3310 103
rect -3290 83 -3270 103
rect -3250 83 -3230 103
rect -3210 83 -3190 103
rect -3170 83 -3150 103
rect -3130 83 -3110 103
rect -3090 83 -3070 103
rect -3050 83 -3030 103
rect -3010 83 -2990 103
rect -2970 83 -2950 103
rect -2930 83 -2910 103
rect -2890 83 -2870 103
rect -2850 83 -2830 103
rect -2810 83 -2790 103
rect -2770 83 -2750 103
rect -2730 83 -2710 103
rect -2690 83 -2670 103
rect -2650 83 -2630 103
rect -2610 83 -2590 103
rect -2570 83 -2550 103
rect -2530 83 -2510 103
rect -2490 83 -2470 103
rect -2450 83 -2430 103
rect -2410 83 -2390 103
rect -2370 83 -2350 103
rect -2330 83 -2310 103
rect -2290 83 -2270 103
rect -2250 83 -2230 103
rect -2210 83 -2190 103
rect -2170 83 -2150 103
rect -2130 83 -2110 103
rect -2090 83 -2070 103
rect -2050 83 -2030 103
rect -2010 83 -1990 103
rect -1970 83 -1950 103
rect -1930 83 -1910 103
rect -1890 83 -1870 103
rect -1850 83 -1830 103
rect -1810 83 -1790 103
rect -1770 83 -1750 103
rect -1730 83 -1710 103
rect -1690 83 -1670 103
rect -1650 83 -1630 103
rect -1610 83 -1590 103
rect -1570 83 -1550 103
rect -1530 83 -1510 103
rect -1490 83 -1470 103
rect -1450 83 -1430 103
rect -1410 83 -1390 103
rect -1370 83 -1350 103
rect -1330 83 -1310 103
rect -1290 83 -1270 103
rect -1250 83 -1230 103
rect -1210 83 -1190 103
rect -1170 83 -1150 103
rect -1130 83 -1110 103
rect -1090 83 -1070 103
rect -1050 83 -1030 103
rect -1010 83 -990 103
rect -970 83 -950 103
rect -930 83 -910 103
rect -890 83 -870 103
rect -850 83 -830 103
rect -810 83 -790 103
rect -770 83 -740 103
rect -710 83 -685 103
rect -3485 68 -685 83
rect -3485 35 -685 50
rect -3485 15 -3470 35
rect -3450 15 -3430 35
rect -3410 15 -3390 35
rect -3370 15 -3350 35
rect -3330 15 -3310 35
rect -3290 15 -3270 35
rect -3250 15 -3230 35
rect -3210 15 -3190 35
rect -3170 15 -3150 35
rect -3130 15 -3110 35
rect -3090 15 -3070 35
rect -3050 15 -3030 35
rect -3010 15 -2990 35
rect -2970 15 -2950 35
rect -2930 15 -2910 35
rect -2890 15 -2870 35
rect -2850 15 -2830 35
rect -2810 15 -2790 35
rect -2770 15 -2750 35
rect -2730 15 -2710 35
rect -2690 15 -2670 35
rect -2650 15 -2630 35
rect -2610 15 -2590 35
rect -2570 15 -2550 35
rect -2530 15 -2510 35
rect -2490 15 -2470 35
rect -2450 15 -2430 35
rect -2410 15 -2390 35
rect -2370 15 -2350 35
rect -2330 15 -2310 35
rect -2290 15 -2270 35
rect -2250 15 -2230 35
rect -2210 15 -2190 35
rect -2170 15 -2150 35
rect -2130 15 -2110 35
rect -2090 15 -2070 35
rect -2050 15 -2030 35
rect -2010 15 -1990 35
rect -1970 15 -1950 35
rect -1930 15 -1910 35
rect -1890 15 -1870 35
rect -1850 15 -1830 35
rect -1810 15 -1790 35
rect -1770 15 -1750 35
rect -1730 15 -1710 35
rect -1690 15 -1670 35
rect -1650 15 -1630 35
rect -1610 15 -1590 35
rect -1570 15 -1550 35
rect -1530 15 -1510 35
rect -1490 15 -1470 35
rect -1450 15 -1430 35
rect -1410 15 -1390 35
rect -1370 15 -1350 35
rect -1330 15 -1310 35
rect -1290 15 -1270 35
rect -1250 15 -1230 35
rect -1210 15 -1190 35
rect -1170 15 -1150 35
rect -1130 15 -1110 35
rect -1090 15 -1070 35
rect -1050 15 -1030 35
rect -1010 15 -990 35
rect -970 15 -950 35
rect -930 15 -910 35
rect -890 15 -870 35
rect -850 15 -830 35
rect -810 15 -790 35
rect -770 15 -740 35
rect -710 15 -685 35
rect -3485 5 -685 15
<< ndiffc >>
rect -3470 -170 -3450 -150
rect -3430 -170 -3410 -150
rect -3390 -170 -3370 -150
rect -3350 -170 -3330 -150
rect -3310 -170 -3290 -150
rect -3270 -170 -3250 -150
rect -3230 -170 -3210 -150
rect -3190 -170 -3170 -150
rect -3150 -170 -3130 -150
rect -3110 -170 -3090 -150
rect -3070 -170 -3050 -150
rect -3030 -170 -3010 -150
rect -2990 -170 -2970 -150
rect -2950 -170 -2930 -150
rect -2910 -170 -2890 -150
rect -2870 -170 -2850 -150
rect -2830 -170 -2810 -150
rect -2790 -170 -2770 -150
rect -2750 -170 -2730 -150
rect -2710 -170 -2690 -150
rect -2670 -170 -2650 -150
rect -2630 -170 -2610 -150
rect -2590 -170 -2570 -150
rect -2550 -170 -2530 -150
rect -2510 -170 -2490 -150
rect -2470 -170 -2450 -150
rect -2430 -170 -2410 -150
rect -2390 -170 -2370 -150
rect -2350 -170 -2330 -150
rect -2310 -170 -2290 -150
rect -2270 -170 -2250 -150
rect -2230 -170 -2210 -150
rect -2190 -170 -2170 -150
rect -2150 -170 -2130 -150
rect -2110 -170 -2090 -150
rect -2070 -170 -2050 -150
rect -2030 -170 -2010 -150
rect -1990 -170 -1970 -150
rect -1950 -170 -1930 -150
rect -1910 -170 -1890 -150
rect -1870 -170 -1850 -150
rect -1830 -170 -1810 -150
rect -1790 -170 -1770 -150
rect -1750 -170 -1730 -150
rect -1710 -170 -1690 -150
rect -1670 -170 -1650 -150
rect -1630 -170 -1610 -150
rect -1590 -170 -1570 -150
rect -1550 -170 -1530 -150
rect -1510 -170 -1490 -150
rect -1470 -170 -1450 -150
rect -1430 -170 -1410 -150
rect -1390 -170 -1370 -150
rect -1350 -170 -1330 -150
rect -1310 -170 -1290 -150
rect -1270 -170 -1250 -150
rect -1230 -170 -1210 -150
rect -1190 -170 -1170 -150
rect -1150 -170 -1130 -150
rect -1110 -170 -1090 -150
rect -1070 -170 -1050 -150
rect -1030 -170 -1005 -150
rect -3470 -235 -3450 -215
rect -3430 -235 -3410 -215
rect -3390 -235 -3370 -215
rect -3350 -235 -3330 -215
rect -3310 -235 -3290 -215
rect -3270 -235 -3250 -215
rect -3230 -235 -3210 -215
rect -3190 -235 -3170 -215
rect -3150 -235 -3130 -215
rect -3110 -235 -3090 -215
rect -3070 -235 -3050 -215
rect -3030 -235 -3010 -215
rect -2990 -235 -2970 -215
rect -2950 -235 -2930 -215
rect -2910 -235 -2890 -215
rect -2870 -235 -2850 -215
rect -2830 -235 -2810 -215
rect -2790 -235 -2770 -215
rect -2750 -235 -2730 -215
rect -2710 -235 -2690 -215
rect -2670 -235 -2650 -215
rect -2630 -235 -2610 -215
rect -2590 -235 -2570 -215
rect -2550 -235 -2530 -215
rect -2510 -235 -2490 -215
rect -2470 -235 -2450 -215
rect -2430 -235 -2410 -215
rect -2390 -235 -2370 -215
rect -2350 -235 -2330 -215
rect -2310 -235 -2290 -215
rect -2270 -235 -2250 -215
rect -2230 -235 -2210 -215
rect -2190 -235 -2170 -215
rect -2150 -235 -2130 -215
rect -2110 -235 -2090 -215
rect -2070 -235 -2050 -215
rect -2030 -235 -2010 -215
rect -1990 -235 -1970 -215
rect -1950 -235 -1930 -215
rect -1910 -235 -1890 -215
rect -1870 -235 -1850 -215
rect -1830 -235 -1810 -215
rect -1790 -235 -1770 -215
rect -1750 -235 -1730 -215
rect -1710 -235 -1690 -215
rect -1670 -235 -1650 -215
rect -1630 -235 -1610 -215
rect -1590 -235 -1570 -215
rect -1550 -235 -1530 -215
rect -1510 -235 -1490 -215
rect -1470 -235 -1450 -215
rect -1430 -235 -1410 -215
rect -1390 -235 -1370 -215
rect -1350 -235 -1330 -215
rect -1310 -235 -1290 -215
rect -1270 -235 -1250 -215
rect -1230 -235 -1210 -215
rect -1190 -235 -1170 -215
rect -1150 -235 -1130 -215
rect -1110 -235 -1090 -215
rect -1070 -235 -1050 -215
rect -1030 -235 -1005 -215
rect -3470 -300 -3450 -280
rect -3430 -300 -3410 -280
rect -3390 -300 -3370 -280
rect -3350 -300 -3330 -280
rect -3310 -300 -3290 -280
rect -3270 -300 -3250 -280
rect -3230 -300 -3210 -280
rect -3190 -300 -3170 -280
rect -3150 -300 -3130 -280
rect -3110 -300 -3090 -280
rect -3070 -300 -3050 -280
rect -3030 -300 -3010 -280
rect -2990 -300 -2970 -280
rect -2950 -300 -2930 -280
rect -2910 -300 -2890 -280
rect -2870 -300 -2850 -280
rect -2830 -300 -2810 -280
rect -2790 -300 -2770 -280
rect -2750 -300 -2730 -280
rect -2710 -300 -2690 -280
rect -2670 -300 -2650 -280
rect -2630 -300 -2610 -280
rect -2590 -300 -2570 -280
rect -2550 -300 -2530 -280
rect -2510 -300 -2490 -280
rect -2470 -300 -2450 -280
rect -2430 -300 -2410 -280
rect -2390 -300 -2370 -280
rect -2350 -300 -2330 -280
rect -2310 -300 -2290 -280
rect -2270 -300 -2250 -280
rect -2230 -300 -2210 -280
rect -2190 -300 -2170 -280
rect -2150 -300 -2130 -280
rect -2110 -300 -2090 -280
rect -2070 -300 -2050 -280
rect -2030 -300 -2010 -280
rect -1990 -300 -1970 -280
rect -1950 -300 -1930 -280
rect -1910 -300 -1890 -280
rect -1870 -300 -1850 -280
rect -1830 -300 -1810 -280
rect -1790 -300 -1770 -280
rect -1750 -300 -1730 -280
rect -1710 -300 -1690 -280
rect -1670 -300 -1650 -280
rect -1630 -300 -1610 -280
rect -1590 -300 -1570 -280
rect -1550 -300 -1530 -280
rect -1510 -300 -1490 -280
rect -1470 -300 -1450 -280
rect -1430 -300 -1410 -280
rect -1390 -300 -1370 -280
rect -1350 -300 -1330 -280
rect -1310 -300 -1290 -280
rect -1270 -300 -1250 -280
rect -1230 -300 -1210 -280
rect -1190 -300 -1170 -280
rect -1150 -300 -1130 -280
rect -1110 -300 -1090 -280
rect -1070 -300 -1050 -280
rect -1030 -300 -1005 -280
rect -3470 -365 -3450 -345
rect -3430 -365 -3410 -345
rect -3390 -365 -3370 -345
rect -3350 -365 -3330 -345
rect -3310 -365 -3290 -345
rect -3270 -365 -3250 -345
rect -3230 -365 -3210 -345
rect -3190 -365 -3170 -345
rect -3150 -365 -3130 -345
rect -3110 -365 -3090 -345
rect -3070 -365 -3050 -345
rect -3030 -365 -3010 -345
rect -2990 -365 -2970 -345
rect -2950 -365 -2930 -345
rect -2910 -365 -2890 -345
rect -2870 -365 -2850 -345
rect -2830 -365 -2810 -345
rect -2790 -365 -2770 -345
rect -2750 -365 -2730 -345
rect -2710 -365 -2690 -345
rect -2670 -365 -2650 -345
rect -2630 -365 -2610 -345
rect -2590 -365 -2570 -345
rect -2550 -365 -2530 -345
rect -2510 -365 -2490 -345
rect -2470 -365 -2450 -345
rect -2430 -365 -2410 -345
rect -2390 -365 -2370 -345
rect -2350 -365 -2330 -345
rect -2310 -365 -2290 -345
rect -2270 -365 -2250 -345
rect -2230 -365 -2210 -345
rect -2190 -365 -2170 -345
rect -2150 -365 -2130 -345
rect -2110 -365 -2090 -345
rect -2070 -365 -2050 -345
rect -2030 -365 -2010 -345
rect -1990 -365 -1970 -345
rect -1950 -365 -1930 -345
rect -1910 -365 -1890 -345
rect -1870 -365 -1850 -345
rect -1830 -365 -1810 -345
rect -1790 -365 -1770 -345
rect -1750 -365 -1730 -345
rect -1710 -365 -1690 -345
rect -1670 -365 -1650 -345
rect -1630 -365 -1610 -345
rect -1590 -365 -1570 -345
rect -1550 -365 -1530 -345
rect -1510 -365 -1490 -345
rect -1470 -365 -1450 -345
rect -1430 -365 -1410 -345
rect -1390 -365 -1370 -345
rect -1350 -365 -1330 -345
rect -1310 -365 -1290 -345
rect -1270 -365 -1250 -345
rect -1230 -365 -1210 -345
rect -1190 -365 -1170 -345
rect -1150 -365 -1130 -345
rect -1110 -365 -1090 -345
rect -1070 -365 -1050 -345
rect -1030 -365 -1005 -345
rect -3470 -430 -3450 -410
rect -3430 -430 -3410 -410
rect -3390 -430 -3370 -410
rect -3350 -430 -3330 -410
rect -3310 -430 -3290 -410
rect -3270 -430 -3250 -410
rect -3230 -430 -3210 -410
rect -3190 -430 -3170 -410
rect -3150 -430 -3130 -410
rect -3110 -430 -3090 -410
rect -3070 -430 -3050 -410
rect -3030 -430 -3010 -410
rect -2990 -430 -2970 -410
rect -2950 -430 -2930 -410
rect -2910 -430 -2890 -410
rect -2870 -430 -2850 -410
rect -2830 -430 -2810 -410
rect -2790 -430 -2770 -410
rect -2750 -430 -2730 -410
rect -2710 -430 -2690 -410
rect -2670 -430 -2650 -410
rect -2630 -430 -2610 -410
rect -2590 -430 -2570 -410
rect -2550 -430 -2530 -410
rect -2510 -430 -2490 -410
rect -2470 -430 -2450 -410
rect -2430 -430 -2410 -410
rect -2390 -430 -2370 -410
rect -2350 -430 -2330 -410
rect -2310 -430 -2290 -410
rect -2270 -430 -2250 -410
rect -2230 -430 -2210 -410
rect -2190 -430 -2170 -410
rect -2150 -430 -2130 -410
rect -2110 -430 -2090 -410
rect -2070 -430 -2050 -410
rect -2030 -430 -2010 -410
rect -1990 -430 -1970 -410
rect -1950 -430 -1930 -410
rect -1910 -430 -1890 -410
rect -1870 -430 -1850 -410
rect -1830 -430 -1810 -410
rect -1790 -430 -1770 -410
rect -1750 -430 -1730 -410
rect -1710 -430 -1690 -410
rect -1670 -430 -1650 -410
rect -1630 -430 -1610 -410
rect -1590 -430 -1570 -410
rect -1550 -430 -1530 -410
rect -1510 -430 -1490 -410
rect -1470 -430 -1450 -410
rect -1430 -430 -1410 -410
rect -1390 -430 -1370 -410
rect -1350 -430 -1330 -410
rect -1310 -430 -1290 -410
rect -1270 -430 -1250 -410
rect -1230 -430 -1210 -410
rect -1190 -430 -1170 -410
rect -1150 -430 -1130 -410
rect -1110 -430 -1090 -410
rect -1070 -430 -1050 -410
rect -1030 -430 -1005 -410
rect -3470 -495 -3450 -475
rect -3430 -495 -3410 -475
rect -3390 -495 -3370 -475
rect -3350 -495 -3330 -475
rect -3310 -495 -3290 -475
rect -3270 -495 -3250 -475
rect -3230 -495 -3210 -475
rect -3190 -495 -3170 -475
rect -3150 -495 -3130 -475
rect -3110 -495 -3090 -475
rect -3070 -495 -3050 -475
rect -3030 -495 -3010 -475
rect -2990 -495 -2970 -475
rect -2950 -495 -2930 -475
rect -2910 -495 -2890 -475
rect -2870 -495 -2850 -475
rect -2830 -495 -2810 -475
rect -2790 -495 -2770 -475
rect -2750 -495 -2730 -475
rect -2710 -495 -2690 -475
rect -2670 -495 -2650 -475
rect -2630 -495 -2610 -475
rect -2590 -495 -2570 -475
rect -2550 -495 -2530 -475
rect -2510 -495 -2490 -475
rect -2470 -495 -2450 -475
rect -2430 -495 -2410 -475
rect -2390 -495 -2370 -475
rect -2350 -495 -2330 -475
rect -2310 -495 -2290 -475
rect -2270 -495 -2250 -475
rect -2230 -495 -2210 -475
rect -2190 -495 -2170 -475
rect -2150 -495 -2130 -475
rect -2110 -495 -2090 -475
rect -2070 -495 -2050 -475
rect -2030 -495 -2010 -475
rect -1990 -495 -1970 -475
rect -1950 -495 -1930 -475
rect -1910 -495 -1890 -475
rect -1870 -495 -1850 -475
rect -1830 -495 -1810 -475
rect -1790 -495 -1770 -475
rect -1750 -495 -1730 -475
rect -1710 -495 -1690 -475
rect -1670 -495 -1650 -475
rect -1630 -495 -1610 -475
rect -1590 -495 -1570 -475
rect -1550 -495 -1530 -475
rect -1510 -495 -1490 -475
rect -1470 -495 -1450 -475
rect -1430 -495 -1410 -475
rect -1390 -495 -1370 -475
rect -1350 -495 -1330 -475
rect -1310 -495 -1290 -475
rect -1270 -495 -1250 -475
rect -1230 -495 -1210 -475
rect -1190 -495 -1170 -475
rect -1150 -495 -1130 -475
rect -1110 -495 -1090 -475
rect -1070 -495 -1050 -475
rect -1030 -495 -1005 -475
rect -3470 -560 -3450 -540
rect -3430 -560 -3410 -540
rect -3390 -560 -3370 -540
rect -3350 -560 -3330 -540
rect -3310 -560 -3290 -540
rect -3270 -560 -3250 -540
rect -3230 -560 -3210 -540
rect -3190 -560 -3170 -540
rect -3150 -560 -3130 -540
rect -3110 -560 -3090 -540
rect -3070 -560 -3050 -540
rect -3030 -560 -3010 -540
rect -2990 -560 -2970 -540
rect -2950 -560 -2930 -540
rect -2910 -560 -2890 -540
rect -2870 -560 -2850 -540
rect -2830 -560 -2810 -540
rect -2790 -560 -2770 -540
rect -2750 -560 -2730 -540
rect -2710 -560 -2690 -540
rect -2670 -560 -2650 -540
rect -2630 -560 -2610 -540
rect -2590 -560 -2570 -540
rect -2550 -560 -2530 -540
rect -2510 -560 -2490 -540
rect -2470 -560 -2450 -540
rect -2430 -560 -2410 -540
rect -2390 -560 -2370 -540
rect -2350 -560 -2330 -540
rect -2310 -560 -2290 -540
rect -2270 -560 -2250 -540
rect -2230 -560 -2210 -540
rect -2190 -560 -2170 -540
rect -2150 -560 -2130 -540
rect -2110 -560 -2090 -540
rect -2070 -560 -2050 -540
rect -2030 -560 -2010 -540
rect -1990 -560 -1970 -540
rect -1950 -560 -1930 -540
rect -1910 -560 -1890 -540
rect -1870 -560 -1850 -540
rect -1830 -560 -1810 -540
rect -1790 -560 -1770 -540
rect -1750 -560 -1730 -540
rect -1710 -560 -1690 -540
rect -1670 -560 -1650 -540
rect -1630 -560 -1610 -540
rect -1590 -560 -1570 -540
rect -1550 -560 -1530 -540
rect -1510 -560 -1490 -540
rect -1470 -560 -1450 -540
rect -1430 -560 -1410 -540
rect -1390 -560 -1370 -540
rect -1350 -560 -1330 -540
rect -1310 -560 -1290 -540
rect -1270 -560 -1250 -540
rect -1230 -560 -1210 -540
rect -1190 -560 -1170 -540
rect -1150 -560 -1130 -540
rect -1110 -560 -1090 -540
rect -1070 -560 -1050 -540
rect -1030 -560 -1005 -540
<< pdiffc >>
rect -3470 1375 -3450 1395
rect -3430 1375 -3410 1395
rect -3390 1375 -3370 1395
rect -3350 1375 -3330 1395
rect -3310 1375 -3290 1395
rect -3270 1375 -3250 1395
rect -3230 1375 -3210 1395
rect -3190 1375 -3170 1395
rect -3150 1375 -3130 1395
rect -3110 1375 -3090 1395
rect -3070 1375 -3050 1395
rect -3030 1375 -3010 1395
rect -2990 1375 -2970 1395
rect -2950 1375 -2930 1395
rect -2910 1375 -2890 1395
rect -2870 1375 -2850 1395
rect -2830 1375 -2810 1395
rect -2790 1375 -2770 1395
rect -2750 1375 -2730 1395
rect -2710 1375 -2690 1395
rect -2670 1375 -2650 1395
rect -2630 1375 -2610 1395
rect -2590 1375 -2570 1395
rect -2550 1375 -2530 1395
rect -2510 1375 -2490 1395
rect -2470 1375 -2450 1395
rect -2430 1375 -2410 1395
rect -2390 1375 -2370 1395
rect -2350 1375 -2330 1395
rect -2310 1375 -2290 1395
rect -2270 1375 -2250 1395
rect -2230 1375 -2210 1395
rect -2190 1375 -2170 1395
rect -2150 1375 -2130 1395
rect -2110 1375 -2090 1395
rect -2070 1375 -2050 1395
rect -2030 1375 -2010 1395
rect -1990 1375 -1970 1395
rect -1950 1375 -1930 1395
rect -1910 1375 -1890 1395
rect -1870 1375 -1850 1395
rect -1830 1375 -1810 1395
rect -1790 1375 -1770 1395
rect -1750 1375 -1730 1395
rect -1710 1375 -1690 1395
rect -1670 1375 -1650 1395
rect -1630 1375 -1610 1395
rect -1590 1375 -1570 1395
rect -1550 1375 -1530 1395
rect -1510 1375 -1490 1395
rect -1470 1375 -1450 1395
rect -1430 1375 -1410 1395
rect -1390 1375 -1370 1395
rect -1350 1375 -1330 1395
rect -1310 1375 -1290 1395
rect -1270 1375 -1250 1395
rect -1230 1375 -1210 1395
rect -1190 1375 -1170 1395
rect -1150 1375 -1130 1395
rect -1110 1375 -1090 1395
rect -1070 1375 -1050 1395
rect -1030 1375 -1010 1395
rect -990 1375 -970 1395
rect -950 1375 -930 1395
rect -910 1375 -890 1395
rect -870 1375 -850 1395
rect -830 1375 -810 1395
rect -790 1375 -770 1395
rect -740 1375 -710 1395
rect -3470 1307 -3450 1327
rect -3430 1307 -3410 1327
rect -3390 1307 -3370 1327
rect -3350 1307 -3330 1327
rect -3310 1307 -3290 1327
rect -3270 1307 -3250 1327
rect -3230 1307 -3210 1327
rect -3190 1307 -3170 1327
rect -3150 1307 -3130 1327
rect -3110 1307 -3090 1327
rect -3070 1307 -3050 1327
rect -3030 1307 -3010 1327
rect -2990 1307 -2970 1327
rect -2950 1307 -2930 1327
rect -2910 1307 -2890 1327
rect -2870 1307 -2850 1327
rect -2830 1307 -2810 1327
rect -2790 1307 -2770 1327
rect -2750 1307 -2730 1327
rect -2710 1307 -2690 1327
rect -2670 1307 -2650 1327
rect -2630 1307 -2610 1327
rect -2590 1307 -2570 1327
rect -2550 1307 -2530 1327
rect -2510 1307 -2490 1327
rect -2470 1307 -2450 1327
rect -2430 1307 -2410 1327
rect -2390 1307 -2370 1327
rect -2350 1307 -2330 1327
rect -2310 1307 -2290 1327
rect -2270 1307 -2250 1327
rect -2230 1307 -2210 1327
rect -2190 1307 -2170 1327
rect -2150 1307 -2130 1327
rect -2110 1307 -2090 1327
rect -2070 1307 -2050 1327
rect -2030 1307 -2010 1327
rect -1990 1307 -1970 1327
rect -1950 1307 -1930 1327
rect -1910 1307 -1890 1327
rect -1870 1307 -1850 1327
rect -1830 1307 -1810 1327
rect -1790 1307 -1770 1327
rect -1750 1307 -1730 1327
rect -1710 1307 -1690 1327
rect -1670 1307 -1650 1327
rect -1630 1307 -1610 1327
rect -1590 1307 -1570 1327
rect -1550 1307 -1530 1327
rect -1510 1307 -1490 1327
rect -1470 1307 -1450 1327
rect -1430 1307 -1410 1327
rect -1390 1307 -1370 1327
rect -1350 1307 -1330 1327
rect -1310 1307 -1290 1327
rect -1270 1307 -1250 1327
rect -1230 1307 -1210 1327
rect -1190 1307 -1170 1327
rect -1150 1307 -1130 1327
rect -1110 1307 -1090 1327
rect -1070 1307 -1050 1327
rect -1030 1307 -1010 1327
rect -990 1307 -970 1327
rect -950 1307 -930 1327
rect -910 1307 -890 1327
rect -870 1307 -850 1327
rect -830 1307 -810 1327
rect -790 1307 -770 1327
rect -740 1307 -710 1327
rect -3470 1239 -3450 1259
rect -3430 1239 -3410 1259
rect -3390 1239 -3370 1259
rect -3350 1239 -3330 1259
rect -3310 1239 -3290 1259
rect -3270 1239 -3250 1259
rect -3230 1239 -3210 1259
rect -3190 1239 -3170 1259
rect -3150 1239 -3130 1259
rect -3110 1239 -3090 1259
rect -3070 1239 -3050 1259
rect -3030 1239 -3010 1259
rect -2990 1239 -2970 1259
rect -2950 1239 -2930 1259
rect -2910 1239 -2890 1259
rect -2870 1239 -2850 1259
rect -2830 1239 -2810 1259
rect -2790 1239 -2770 1259
rect -2750 1239 -2730 1259
rect -2710 1239 -2690 1259
rect -2670 1239 -2650 1259
rect -2630 1239 -2610 1259
rect -2590 1239 -2570 1259
rect -2550 1239 -2530 1259
rect -2510 1239 -2490 1259
rect -2470 1239 -2450 1259
rect -2430 1239 -2410 1259
rect -2390 1239 -2370 1259
rect -2350 1239 -2330 1259
rect -2310 1239 -2290 1259
rect -2270 1239 -2250 1259
rect -2230 1239 -2210 1259
rect -2190 1239 -2170 1259
rect -2150 1239 -2130 1259
rect -2110 1239 -2090 1259
rect -2070 1239 -2050 1259
rect -2030 1239 -2010 1259
rect -1990 1239 -1970 1259
rect -1950 1239 -1930 1259
rect -1910 1239 -1890 1259
rect -1870 1239 -1850 1259
rect -1830 1239 -1810 1259
rect -1790 1239 -1770 1259
rect -1750 1239 -1730 1259
rect -1710 1239 -1690 1259
rect -1670 1239 -1650 1259
rect -1630 1239 -1610 1259
rect -1590 1239 -1570 1259
rect -1550 1239 -1530 1259
rect -1510 1239 -1490 1259
rect -1470 1239 -1450 1259
rect -1430 1239 -1410 1259
rect -1390 1239 -1370 1259
rect -1350 1239 -1330 1259
rect -1310 1239 -1290 1259
rect -1270 1239 -1250 1259
rect -1230 1239 -1210 1259
rect -1190 1239 -1170 1259
rect -1150 1239 -1130 1259
rect -1110 1239 -1090 1259
rect -1070 1239 -1050 1259
rect -1030 1239 -1010 1259
rect -990 1239 -970 1259
rect -950 1239 -930 1259
rect -910 1239 -890 1259
rect -870 1239 -850 1259
rect -830 1239 -810 1259
rect -790 1239 -770 1259
rect -740 1239 -710 1259
rect -3470 1171 -3450 1191
rect -3430 1171 -3410 1191
rect -3390 1171 -3370 1191
rect -3350 1171 -3330 1191
rect -3310 1171 -3290 1191
rect -3270 1171 -3250 1191
rect -3230 1171 -3210 1191
rect -3190 1171 -3170 1191
rect -3150 1171 -3130 1191
rect -3110 1171 -3090 1191
rect -3070 1171 -3050 1191
rect -3030 1171 -3010 1191
rect -2990 1171 -2970 1191
rect -2950 1171 -2930 1191
rect -2910 1171 -2890 1191
rect -2870 1171 -2850 1191
rect -2830 1171 -2810 1191
rect -2790 1171 -2770 1191
rect -2750 1171 -2730 1191
rect -2710 1171 -2690 1191
rect -2670 1171 -2650 1191
rect -2630 1171 -2610 1191
rect -2590 1171 -2570 1191
rect -2550 1171 -2530 1191
rect -2510 1171 -2490 1191
rect -2470 1171 -2450 1191
rect -2430 1171 -2410 1191
rect -2390 1171 -2370 1191
rect -2350 1171 -2330 1191
rect -2310 1171 -2290 1191
rect -2270 1171 -2250 1191
rect -2230 1171 -2210 1191
rect -2190 1171 -2170 1191
rect -2150 1171 -2130 1191
rect -2110 1171 -2090 1191
rect -2070 1171 -2050 1191
rect -2030 1171 -2010 1191
rect -1990 1171 -1970 1191
rect -1950 1171 -1930 1191
rect -1910 1171 -1890 1191
rect -1870 1171 -1850 1191
rect -1830 1171 -1810 1191
rect -1790 1171 -1770 1191
rect -1750 1171 -1730 1191
rect -1710 1171 -1690 1191
rect -1670 1171 -1650 1191
rect -1630 1171 -1610 1191
rect -1590 1171 -1570 1191
rect -1550 1171 -1530 1191
rect -1510 1171 -1490 1191
rect -1470 1171 -1450 1191
rect -1430 1171 -1410 1191
rect -1390 1171 -1370 1191
rect -1350 1171 -1330 1191
rect -1310 1171 -1290 1191
rect -1270 1171 -1250 1191
rect -1230 1171 -1210 1191
rect -1190 1171 -1170 1191
rect -1150 1171 -1130 1191
rect -1110 1171 -1090 1191
rect -1070 1171 -1050 1191
rect -1030 1171 -1010 1191
rect -990 1171 -970 1191
rect -950 1171 -930 1191
rect -910 1171 -890 1191
rect -870 1171 -850 1191
rect -830 1171 -810 1191
rect -790 1171 -770 1191
rect -740 1171 -710 1191
rect -3470 1103 -3450 1123
rect -3430 1103 -3410 1123
rect -3390 1103 -3370 1123
rect -3350 1103 -3330 1123
rect -3310 1103 -3290 1123
rect -3270 1103 -3250 1123
rect -3230 1103 -3210 1123
rect -3190 1103 -3170 1123
rect -3150 1103 -3130 1123
rect -3110 1103 -3090 1123
rect -3070 1103 -3050 1123
rect -3030 1103 -3010 1123
rect -2990 1103 -2970 1123
rect -2950 1103 -2930 1123
rect -2910 1103 -2890 1123
rect -2870 1103 -2850 1123
rect -2830 1103 -2810 1123
rect -2790 1103 -2770 1123
rect -2750 1103 -2730 1123
rect -2710 1103 -2690 1123
rect -2670 1103 -2650 1123
rect -2630 1103 -2610 1123
rect -2590 1103 -2570 1123
rect -2550 1103 -2530 1123
rect -2510 1103 -2490 1123
rect -2470 1103 -2450 1123
rect -2430 1103 -2410 1123
rect -2390 1103 -2370 1123
rect -2350 1103 -2330 1123
rect -2310 1103 -2290 1123
rect -2270 1103 -2250 1123
rect -2230 1103 -2210 1123
rect -2190 1103 -2170 1123
rect -2150 1103 -2130 1123
rect -2110 1103 -2090 1123
rect -2070 1103 -2050 1123
rect -2030 1103 -2010 1123
rect -1990 1103 -1970 1123
rect -1950 1103 -1930 1123
rect -1910 1103 -1890 1123
rect -1870 1103 -1850 1123
rect -1830 1103 -1810 1123
rect -1790 1103 -1770 1123
rect -1750 1103 -1730 1123
rect -1710 1103 -1690 1123
rect -1670 1103 -1650 1123
rect -1630 1103 -1610 1123
rect -1590 1103 -1570 1123
rect -1550 1103 -1530 1123
rect -1510 1103 -1490 1123
rect -1470 1103 -1450 1123
rect -1430 1103 -1410 1123
rect -1390 1103 -1370 1123
rect -1350 1103 -1330 1123
rect -1310 1103 -1290 1123
rect -1270 1103 -1250 1123
rect -1230 1103 -1210 1123
rect -1190 1103 -1170 1123
rect -1150 1103 -1130 1123
rect -1110 1103 -1090 1123
rect -1070 1103 -1050 1123
rect -1030 1103 -1010 1123
rect -990 1103 -970 1123
rect -950 1103 -930 1123
rect -910 1103 -890 1123
rect -870 1103 -850 1123
rect -830 1103 -810 1123
rect -790 1103 -770 1123
rect -740 1103 -710 1123
rect -3470 1035 -3450 1055
rect -3430 1035 -3410 1055
rect -3390 1035 -3370 1055
rect -3350 1035 -3330 1055
rect -3310 1035 -3290 1055
rect -3270 1035 -3250 1055
rect -3230 1035 -3210 1055
rect -3190 1035 -3170 1055
rect -3150 1035 -3130 1055
rect -3110 1035 -3090 1055
rect -3070 1035 -3050 1055
rect -3030 1035 -3010 1055
rect -2990 1035 -2970 1055
rect -2950 1035 -2930 1055
rect -2910 1035 -2890 1055
rect -2870 1035 -2850 1055
rect -2830 1035 -2810 1055
rect -2790 1035 -2770 1055
rect -2750 1035 -2730 1055
rect -2710 1035 -2690 1055
rect -2670 1035 -2650 1055
rect -2630 1035 -2610 1055
rect -2590 1035 -2570 1055
rect -2550 1035 -2530 1055
rect -2510 1035 -2490 1055
rect -2470 1035 -2450 1055
rect -2430 1035 -2410 1055
rect -2390 1035 -2370 1055
rect -2350 1035 -2330 1055
rect -2310 1035 -2290 1055
rect -2270 1035 -2250 1055
rect -2230 1035 -2210 1055
rect -2190 1035 -2170 1055
rect -2150 1035 -2130 1055
rect -2110 1035 -2090 1055
rect -2070 1035 -2050 1055
rect -2030 1035 -2010 1055
rect -1990 1035 -1970 1055
rect -1950 1035 -1930 1055
rect -1910 1035 -1890 1055
rect -1870 1035 -1850 1055
rect -1830 1035 -1810 1055
rect -1790 1035 -1770 1055
rect -1750 1035 -1730 1055
rect -1710 1035 -1690 1055
rect -1670 1035 -1650 1055
rect -1630 1035 -1610 1055
rect -1590 1035 -1570 1055
rect -1550 1035 -1530 1055
rect -1510 1035 -1490 1055
rect -1470 1035 -1450 1055
rect -1430 1035 -1410 1055
rect -1390 1035 -1370 1055
rect -1350 1035 -1330 1055
rect -1310 1035 -1290 1055
rect -1270 1035 -1250 1055
rect -1230 1035 -1210 1055
rect -1190 1035 -1170 1055
rect -1150 1035 -1130 1055
rect -1110 1035 -1090 1055
rect -1070 1035 -1050 1055
rect -1030 1035 -1010 1055
rect -990 1035 -970 1055
rect -950 1035 -930 1055
rect -910 1035 -890 1055
rect -870 1035 -850 1055
rect -830 1035 -810 1055
rect -790 1035 -770 1055
rect -740 1035 -710 1055
rect -3470 967 -3450 987
rect -3430 967 -3410 987
rect -3390 967 -3370 987
rect -3350 967 -3330 987
rect -3310 967 -3290 987
rect -3270 967 -3250 987
rect -3230 967 -3210 987
rect -3190 967 -3170 987
rect -3150 967 -3130 987
rect -3110 967 -3090 987
rect -3070 967 -3050 987
rect -3030 967 -3010 987
rect -2990 967 -2970 987
rect -2950 967 -2930 987
rect -2910 967 -2890 987
rect -2870 967 -2850 987
rect -2830 967 -2810 987
rect -2790 967 -2770 987
rect -2750 967 -2730 987
rect -2710 967 -2690 987
rect -2670 967 -2650 987
rect -2630 967 -2610 987
rect -2590 967 -2570 987
rect -2550 967 -2530 987
rect -2510 967 -2490 987
rect -2470 967 -2450 987
rect -2430 967 -2410 987
rect -2390 967 -2370 987
rect -2350 967 -2330 987
rect -2310 967 -2290 987
rect -2270 967 -2250 987
rect -2230 967 -2210 987
rect -2190 967 -2170 987
rect -2150 967 -2130 987
rect -2110 967 -2090 987
rect -2070 967 -2050 987
rect -2030 967 -2010 987
rect -1990 967 -1970 987
rect -1950 967 -1930 987
rect -1910 967 -1890 987
rect -1870 967 -1850 987
rect -1830 967 -1810 987
rect -1790 967 -1770 987
rect -1750 967 -1730 987
rect -1710 967 -1690 987
rect -1670 967 -1650 987
rect -1630 967 -1610 987
rect -1590 967 -1570 987
rect -1550 967 -1530 987
rect -1510 967 -1490 987
rect -1470 967 -1450 987
rect -1430 967 -1410 987
rect -1390 967 -1370 987
rect -1350 967 -1330 987
rect -1310 967 -1290 987
rect -1270 967 -1250 987
rect -1230 967 -1210 987
rect -1190 967 -1170 987
rect -1150 967 -1130 987
rect -1110 967 -1090 987
rect -1070 967 -1050 987
rect -1030 967 -1010 987
rect -990 967 -970 987
rect -950 967 -930 987
rect -910 967 -890 987
rect -870 967 -850 987
rect -830 967 -810 987
rect -790 967 -770 987
rect -740 967 -710 987
rect -3470 899 -3450 919
rect -3430 899 -3410 919
rect -3390 899 -3370 919
rect -3350 899 -3330 919
rect -3310 899 -3290 919
rect -3270 899 -3250 919
rect -3230 899 -3210 919
rect -3190 899 -3170 919
rect -3150 899 -3130 919
rect -3110 899 -3090 919
rect -3070 899 -3050 919
rect -3030 899 -3010 919
rect -2990 899 -2970 919
rect -2950 899 -2930 919
rect -2910 899 -2890 919
rect -2870 899 -2850 919
rect -2830 899 -2810 919
rect -2790 899 -2770 919
rect -2750 899 -2730 919
rect -2710 899 -2690 919
rect -2670 899 -2650 919
rect -2630 899 -2610 919
rect -2590 899 -2570 919
rect -2550 899 -2530 919
rect -2510 899 -2490 919
rect -2470 899 -2450 919
rect -2430 899 -2410 919
rect -2390 899 -2370 919
rect -2350 899 -2330 919
rect -2310 899 -2290 919
rect -2270 899 -2250 919
rect -2230 899 -2210 919
rect -2190 899 -2170 919
rect -2150 899 -2130 919
rect -2110 899 -2090 919
rect -2070 899 -2050 919
rect -2030 899 -2010 919
rect -1990 899 -1970 919
rect -1950 899 -1930 919
rect -1910 899 -1890 919
rect -1870 899 -1850 919
rect -1830 899 -1810 919
rect -1790 899 -1770 919
rect -1750 899 -1730 919
rect -1710 899 -1690 919
rect -1670 899 -1650 919
rect -1630 899 -1610 919
rect -1590 899 -1570 919
rect -1550 899 -1530 919
rect -1510 899 -1490 919
rect -1470 899 -1450 919
rect -1430 899 -1410 919
rect -1390 899 -1370 919
rect -1350 899 -1330 919
rect -1310 899 -1290 919
rect -1270 899 -1250 919
rect -1230 899 -1210 919
rect -1190 899 -1170 919
rect -1150 899 -1130 919
rect -1110 899 -1090 919
rect -1070 899 -1050 919
rect -1030 899 -1010 919
rect -990 899 -970 919
rect -950 899 -930 919
rect -910 899 -890 919
rect -870 899 -850 919
rect -830 899 -810 919
rect -790 899 -770 919
rect -740 899 -710 919
rect -3470 831 -3450 851
rect -3430 831 -3410 851
rect -3390 831 -3370 851
rect -3350 831 -3330 851
rect -3310 831 -3290 851
rect -3270 831 -3250 851
rect -3230 831 -3210 851
rect -3190 831 -3170 851
rect -3150 831 -3130 851
rect -3110 831 -3090 851
rect -3070 831 -3050 851
rect -3030 831 -3010 851
rect -2990 831 -2970 851
rect -2950 831 -2930 851
rect -2910 831 -2890 851
rect -2870 831 -2850 851
rect -2830 831 -2810 851
rect -2790 831 -2770 851
rect -2750 831 -2730 851
rect -2710 831 -2690 851
rect -2670 831 -2650 851
rect -2630 831 -2610 851
rect -2590 831 -2570 851
rect -2550 831 -2530 851
rect -2510 831 -2490 851
rect -2470 831 -2450 851
rect -2430 831 -2410 851
rect -2390 831 -2370 851
rect -2350 831 -2330 851
rect -2310 831 -2290 851
rect -2270 831 -2250 851
rect -2230 831 -2210 851
rect -2190 831 -2170 851
rect -2150 831 -2130 851
rect -2110 831 -2090 851
rect -2070 831 -2050 851
rect -2030 831 -2010 851
rect -1990 831 -1970 851
rect -1950 831 -1930 851
rect -1910 831 -1890 851
rect -1870 831 -1850 851
rect -1830 831 -1810 851
rect -1790 831 -1770 851
rect -1750 831 -1730 851
rect -1710 831 -1690 851
rect -1670 831 -1650 851
rect -1630 831 -1610 851
rect -1590 831 -1570 851
rect -1550 831 -1530 851
rect -1510 831 -1490 851
rect -1470 831 -1450 851
rect -1430 831 -1410 851
rect -1390 831 -1370 851
rect -1350 831 -1330 851
rect -1310 831 -1290 851
rect -1270 831 -1250 851
rect -1230 831 -1210 851
rect -1190 831 -1170 851
rect -1150 831 -1130 851
rect -1110 831 -1090 851
rect -1070 831 -1050 851
rect -1030 831 -1010 851
rect -990 831 -970 851
rect -950 831 -930 851
rect -910 831 -890 851
rect -870 831 -850 851
rect -830 831 -810 851
rect -790 831 -770 851
rect -740 831 -710 851
rect -3470 763 -3450 783
rect -3430 763 -3410 783
rect -3390 763 -3370 783
rect -3350 763 -3330 783
rect -3310 763 -3290 783
rect -3270 763 -3250 783
rect -3230 763 -3210 783
rect -3190 763 -3170 783
rect -3150 763 -3130 783
rect -3110 763 -3090 783
rect -3070 763 -3050 783
rect -3030 763 -3010 783
rect -2990 763 -2970 783
rect -2950 763 -2930 783
rect -2910 763 -2890 783
rect -2870 763 -2850 783
rect -2830 763 -2810 783
rect -2790 763 -2770 783
rect -2750 763 -2730 783
rect -2710 763 -2690 783
rect -2670 763 -2650 783
rect -2630 763 -2610 783
rect -2590 763 -2570 783
rect -2550 763 -2530 783
rect -2510 763 -2490 783
rect -2470 763 -2450 783
rect -2430 763 -2410 783
rect -2390 763 -2370 783
rect -2350 763 -2330 783
rect -2310 763 -2290 783
rect -2270 763 -2250 783
rect -2230 763 -2210 783
rect -2190 763 -2170 783
rect -2150 763 -2130 783
rect -2110 763 -2090 783
rect -2070 763 -2050 783
rect -2030 763 -2010 783
rect -1990 763 -1970 783
rect -1950 763 -1930 783
rect -1910 763 -1890 783
rect -1870 763 -1850 783
rect -1830 763 -1810 783
rect -1790 763 -1770 783
rect -1750 763 -1730 783
rect -1710 763 -1690 783
rect -1670 763 -1650 783
rect -1630 763 -1610 783
rect -1590 763 -1570 783
rect -1550 763 -1530 783
rect -1510 763 -1490 783
rect -1470 763 -1450 783
rect -1430 763 -1410 783
rect -1390 763 -1370 783
rect -1350 763 -1330 783
rect -1310 763 -1290 783
rect -1270 763 -1250 783
rect -1230 763 -1210 783
rect -1190 763 -1170 783
rect -1150 763 -1130 783
rect -1110 763 -1090 783
rect -1070 763 -1050 783
rect -1030 763 -1010 783
rect -990 763 -970 783
rect -950 763 -930 783
rect -910 763 -890 783
rect -870 763 -850 783
rect -830 763 -810 783
rect -790 763 -770 783
rect -740 763 -710 783
rect -3470 695 -3450 715
rect -3430 695 -3410 715
rect -3390 695 -3370 715
rect -3350 695 -3330 715
rect -3310 695 -3290 715
rect -3270 695 -3250 715
rect -3230 695 -3210 715
rect -3190 695 -3170 715
rect -3150 695 -3130 715
rect -3110 695 -3090 715
rect -3070 695 -3050 715
rect -3030 695 -3010 715
rect -2990 695 -2970 715
rect -2950 695 -2930 715
rect -2910 695 -2890 715
rect -2870 695 -2850 715
rect -2830 695 -2810 715
rect -2790 695 -2770 715
rect -2750 695 -2730 715
rect -2710 695 -2690 715
rect -2670 695 -2650 715
rect -2630 695 -2610 715
rect -2590 695 -2570 715
rect -2550 695 -2530 715
rect -2510 695 -2490 715
rect -2470 695 -2450 715
rect -2430 695 -2410 715
rect -2390 695 -2370 715
rect -2350 695 -2330 715
rect -2310 695 -2290 715
rect -2270 695 -2250 715
rect -2230 695 -2210 715
rect -2190 695 -2170 715
rect -2150 695 -2130 715
rect -2110 695 -2090 715
rect -2070 695 -2050 715
rect -2030 695 -2010 715
rect -1990 695 -1970 715
rect -1950 695 -1930 715
rect -1910 695 -1890 715
rect -1870 695 -1850 715
rect -1830 695 -1810 715
rect -1790 695 -1770 715
rect -1750 695 -1730 715
rect -1710 695 -1690 715
rect -1670 695 -1650 715
rect -1630 695 -1610 715
rect -1590 695 -1570 715
rect -1550 695 -1530 715
rect -1510 695 -1490 715
rect -1470 695 -1450 715
rect -1430 695 -1410 715
rect -1390 695 -1370 715
rect -1350 695 -1330 715
rect -1310 695 -1290 715
rect -1270 695 -1250 715
rect -1230 695 -1210 715
rect -1190 695 -1170 715
rect -1150 695 -1130 715
rect -1110 695 -1090 715
rect -1070 695 -1050 715
rect -1030 695 -1010 715
rect -990 695 -970 715
rect -950 695 -930 715
rect -910 695 -890 715
rect -870 695 -850 715
rect -830 695 -810 715
rect -790 695 -770 715
rect -740 695 -710 715
rect -3470 627 -3450 647
rect -3430 627 -3410 647
rect -3390 627 -3370 647
rect -3350 627 -3330 647
rect -3310 627 -3290 647
rect -3270 627 -3250 647
rect -3230 627 -3210 647
rect -3190 627 -3170 647
rect -3150 627 -3130 647
rect -3110 627 -3090 647
rect -3070 627 -3050 647
rect -3030 627 -3010 647
rect -2990 627 -2970 647
rect -2950 627 -2930 647
rect -2910 627 -2890 647
rect -2870 627 -2850 647
rect -2830 627 -2810 647
rect -2790 627 -2770 647
rect -2750 627 -2730 647
rect -2710 627 -2690 647
rect -2670 627 -2650 647
rect -2630 627 -2610 647
rect -2590 627 -2570 647
rect -2550 627 -2530 647
rect -2510 627 -2490 647
rect -2470 627 -2450 647
rect -2430 627 -2410 647
rect -2390 627 -2370 647
rect -2350 627 -2330 647
rect -2310 627 -2290 647
rect -2270 627 -2250 647
rect -2230 627 -2210 647
rect -2190 627 -2170 647
rect -2150 627 -2130 647
rect -2110 627 -2090 647
rect -2070 627 -2050 647
rect -2030 627 -2010 647
rect -1990 627 -1970 647
rect -1950 627 -1930 647
rect -1910 627 -1890 647
rect -1870 627 -1850 647
rect -1830 627 -1810 647
rect -1790 627 -1770 647
rect -1750 627 -1730 647
rect -1710 627 -1690 647
rect -1670 627 -1650 647
rect -1630 627 -1610 647
rect -1590 627 -1570 647
rect -1550 627 -1530 647
rect -1510 627 -1490 647
rect -1470 627 -1450 647
rect -1430 627 -1410 647
rect -1390 627 -1370 647
rect -1350 627 -1330 647
rect -1310 627 -1290 647
rect -1270 627 -1250 647
rect -1230 627 -1210 647
rect -1190 627 -1170 647
rect -1150 627 -1130 647
rect -1110 627 -1090 647
rect -1070 627 -1050 647
rect -1030 627 -1010 647
rect -990 627 -970 647
rect -950 627 -930 647
rect -910 627 -890 647
rect -870 627 -850 647
rect -830 627 -810 647
rect -790 627 -770 647
rect -740 627 -710 647
rect -3470 559 -3450 579
rect -3430 559 -3410 579
rect -3390 559 -3370 579
rect -3350 559 -3330 579
rect -3310 559 -3290 579
rect -3270 559 -3250 579
rect -3230 559 -3210 579
rect -3190 559 -3170 579
rect -3150 559 -3130 579
rect -3110 559 -3090 579
rect -3070 559 -3050 579
rect -3030 559 -3010 579
rect -2990 559 -2970 579
rect -2950 559 -2930 579
rect -2910 559 -2890 579
rect -2870 559 -2850 579
rect -2830 559 -2810 579
rect -2790 559 -2770 579
rect -2750 559 -2730 579
rect -2710 559 -2690 579
rect -2670 559 -2650 579
rect -2630 559 -2610 579
rect -2590 559 -2570 579
rect -2550 559 -2530 579
rect -2510 559 -2490 579
rect -2470 559 -2450 579
rect -2430 559 -2410 579
rect -2390 559 -2370 579
rect -2350 559 -2330 579
rect -2310 559 -2290 579
rect -2270 559 -2250 579
rect -2230 559 -2210 579
rect -2190 559 -2170 579
rect -2150 559 -2130 579
rect -2110 559 -2090 579
rect -2070 559 -2050 579
rect -2030 559 -2010 579
rect -1990 559 -1970 579
rect -1950 559 -1930 579
rect -1910 559 -1890 579
rect -1870 559 -1850 579
rect -1830 559 -1810 579
rect -1790 559 -1770 579
rect -1750 559 -1730 579
rect -1710 559 -1690 579
rect -1670 559 -1650 579
rect -1630 559 -1610 579
rect -1590 559 -1570 579
rect -1550 559 -1530 579
rect -1510 559 -1490 579
rect -1470 559 -1450 579
rect -1430 559 -1410 579
rect -1390 559 -1370 579
rect -1350 559 -1330 579
rect -1310 559 -1290 579
rect -1270 559 -1250 579
rect -1230 559 -1210 579
rect -1190 559 -1170 579
rect -1150 559 -1130 579
rect -1110 559 -1090 579
rect -1070 559 -1050 579
rect -1030 559 -1010 579
rect -990 559 -970 579
rect -950 559 -930 579
rect -910 559 -890 579
rect -870 559 -850 579
rect -830 559 -810 579
rect -790 559 -770 579
rect -740 559 -710 579
rect -3470 491 -3450 511
rect -3430 491 -3410 511
rect -3390 491 -3370 511
rect -3350 491 -3330 511
rect -3310 491 -3290 511
rect -3270 491 -3250 511
rect -3230 491 -3210 511
rect -3190 491 -3170 511
rect -3150 491 -3130 511
rect -3110 491 -3090 511
rect -3070 491 -3050 511
rect -3030 491 -3010 511
rect -2990 491 -2970 511
rect -2950 491 -2930 511
rect -2910 491 -2890 511
rect -2870 491 -2850 511
rect -2830 491 -2810 511
rect -2790 491 -2770 511
rect -2750 491 -2730 511
rect -2710 491 -2690 511
rect -2670 491 -2650 511
rect -2630 491 -2610 511
rect -2590 491 -2570 511
rect -2550 491 -2530 511
rect -2510 491 -2490 511
rect -2470 491 -2450 511
rect -2430 491 -2410 511
rect -2390 491 -2370 511
rect -2350 491 -2330 511
rect -2310 491 -2290 511
rect -2270 491 -2250 511
rect -2230 491 -2210 511
rect -2190 491 -2170 511
rect -2150 491 -2130 511
rect -2110 491 -2090 511
rect -2070 491 -2050 511
rect -2030 491 -2010 511
rect -1990 491 -1970 511
rect -1950 491 -1930 511
rect -1910 491 -1890 511
rect -1870 491 -1850 511
rect -1830 491 -1810 511
rect -1790 491 -1770 511
rect -1750 491 -1730 511
rect -1710 491 -1690 511
rect -1670 491 -1650 511
rect -1630 491 -1610 511
rect -1590 491 -1570 511
rect -1550 491 -1530 511
rect -1510 491 -1490 511
rect -1470 491 -1450 511
rect -1430 491 -1410 511
rect -1390 491 -1370 511
rect -1350 491 -1330 511
rect -1310 491 -1290 511
rect -1270 491 -1250 511
rect -1230 491 -1210 511
rect -1190 491 -1170 511
rect -1150 491 -1130 511
rect -1110 491 -1090 511
rect -1070 491 -1050 511
rect -1030 491 -1010 511
rect -990 491 -970 511
rect -950 491 -930 511
rect -910 491 -890 511
rect -870 491 -850 511
rect -830 491 -810 511
rect -790 491 -770 511
rect -740 491 -710 511
rect -3470 423 -3450 443
rect -3430 423 -3410 443
rect -3390 423 -3370 443
rect -3350 423 -3330 443
rect -3310 423 -3290 443
rect -3270 423 -3250 443
rect -3230 423 -3210 443
rect -3190 423 -3170 443
rect -3150 423 -3130 443
rect -3110 423 -3090 443
rect -3070 423 -3050 443
rect -3030 423 -3010 443
rect -2990 423 -2970 443
rect -2950 423 -2930 443
rect -2910 423 -2890 443
rect -2870 423 -2850 443
rect -2830 423 -2810 443
rect -2790 423 -2770 443
rect -2750 423 -2730 443
rect -2710 423 -2690 443
rect -2670 423 -2650 443
rect -2630 423 -2610 443
rect -2590 423 -2570 443
rect -2550 423 -2530 443
rect -2510 423 -2490 443
rect -2470 423 -2450 443
rect -2430 423 -2410 443
rect -2390 423 -2370 443
rect -2350 423 -2330 443
rect -2310 423 -2290 443
rect -2270 423 -2250 443
rect -2230 423 -2210 443
rect -2190 423 -2170 443
rect -2150 423 -2130 443
rect -2110 423 -2090 443
rect -2070 423 -2050 443
rect -2030 423 -2010 443
rect -1990 423 -1970 443
rect -1950 423 -1930 443
rect -1910 423 -1890 443
rect -1870 423 -1850 443
rect -1830 423 -1810 443
rect -1790 423 -1770 443
rect -1750 423 -1730 443
rect -1710 423 -1690 443
rect -1670 423 -1650 443
rect -1630 423 -1610 443
rect -1590 423 -1570 443
rect -1550 423 -1530 443
rect -1510 423 -1490 443
rect -1470 423 -1450 443
rect -1430 423 -1410 443
rect -1390 423 -1370 443
rect -1350 423 -1330 443
rect -1310 423 -1290 443
rect -1270 423 -1250 443
rect -1230 423 -1210 443
rect -1190 423 -1170 443
rect -1150 423 -1130 443
rect -1110 423 -1090 443
rect -1070 423 -1050 443
rect -1030 423 -1010 443
rect -990 423 -970 443
rect -950 423 -930 443
rect -910 423 -890 443
rect -870 423 -850 443
rect -830 423 -810 443
rect -790 423 -770 443
rect -740 423 -710 443
rect -3470 355 -3450 375
rect -3430 355 -3410 375
rect -3390 355 -3370 375
rect -3350 355 -3330 375
rect -3310 355 -3290 375
rect -3270 355 -3250 375
rect -3230 355 -3210 375
rect -3190 355 -3170 375
rect -3150 355 -3130 375
rect -3110 355 -3090 375
rect -3070 355 -3050 375
rect -3030 355 -3010 375
rect -2990 355 -2970 375
rect -2950 355 -2930 375
rect -2910 355 -2890 375
rect -2870 355 -2850 375
rect -2830 355 -2810 375
rect -2790 355 -2770 375
rect -2750 355 -2730 375
rect -2710 355 -2690 375
rect -2670 355 -2650 375
rect -2630 355 -2610 375
rect -2590 355 -2570 375
rect -2550 355 -2530 375
rect -2510 355 -2490 375
rect -2470 355 -2450 375
rect -2430 355 -2410 375
rect -2390 355 -2370 375
rect -2350 355 -2330 375
rect -2310 355 -2290 375
rect -2270 355 -2250 375
rect -2230 355 -2210 375
rect -2190 355 -2170 375
rect -2150 355 -2130 375
rect -2110 355 -2090 375
rect -2070 355 -2050 375
rect -2030 355 -2010 375
rect -1990 355 -1970 375
rect -1950 355 -1930 375
rect -1910 355 -1890 375
rect -1870 355 -1850 375
rect -1830 355 -1810 375
rect -1790 355 -1770 375
rect -1750 355 -1730 375
rect -1710 355 -1690 375
rect -1670 355 -1650 375
rect -1630 355 -1610 375
rect -1590 355 -1570 375
rect -1550 355 -1530 375
rect -1510 355 -1490 375
rect -1470 355 -1450 375
rect -1430 355 -1410 375
rect -1390 355 -1370 375
rect -1350 355 -1330 375
rect -1310 355 -1290 375
rect -1270 355 -1250 375
rect -1230 355 -1210 375
rect -1190 355 -1170 375
rect -1150 355 -1130 375
rect -1110 355 -1090 375
rect -1070 355 -1050 375
rect -1030 355 -1010 375
rect -990 355 -970 375
rect -950 355 -930 375
rect -910 355 -890 375
rect -870 355 -850 375
rect -830 355 -810 375
rect -790 355 -770 375
rect -740 355 -710 375
rect -3470 287 -3450 307
rect -3430 287 -3410 307
rect -3390 287 -3370 307
rect -3350 287 -3330 307
rect -3310 287 -3290 307
rect -3270 287 -3250 307
rect -3230 287 -3210 307
rect -3190 287 -3170 307
rect -3150 287 -3130 307
rect -3110 287 -3090 307
rect -3070 287 -3050 307
rect -3030 287 -3010 307
rect -2990 287 -2970 307
rect -2950 287 -2930 307
rect -2910 287 -2890 307
rect -2870 287 -2850 307
rect -2830 287 -2810 307
rect -2790 287 -2770 307
rect -2750 287 -2730 307
rect -2710 287 -2690 307
rect -2670 287 -2650 307
rect -2630 287 -2610 307
rect -2590 287 -2570 307
rect -2550 287 -2530 307
rect -2510 287 -2490 307
rect -2470 287 -2450 307
rect -2430 287 -2410 307
rect -2390 287 -2370 307
rect -2350 287 -2330 307
rect -2310 287 -2290 307
rect -2270 287 -2250 307
rect -2230 287 -2210 307
rect -2190 287 -2170 307
rect -2150 287 -2130 307
rect -2110 287 -2090 307
rect -2070 287 -2050 307
rect -2030 287 -2010 307
rect -1990 287 -1970 307
rect -1950 287 -1930 307
rect -1910 287 -1890 307
rect -1870 287 -1850 307
rect -1830 287 -1810 307
rect -1790 287 -1770 307
rect -1750 287 -1730 307
rect -1710 287 -1690 307
rect -1670 287 -1650 307
rect -1630 287 -1610 307
rect -1590 287 -1570 307
rect -1550 287 -1530 307
rect -1510 287 -1490 307
rect -1470 287 -1450 307
rect -1430 287 -1410 307
rect -1390 287 -1370 307
rect -1350 287 -1330 307
rect -1310 287 -1290 307
rect -1270 287 -1250 307
rect -1230 287 -1210 307
rect -1190 287 -1170 307
rect -1150 287 -1130 307
rect -1110 287 -1090 307
rect -1070 287 -1050 307
rect -1030 287 -1010 307
rect -990 287 -970 307
rect -950 287 -930 307
rect -910 287 -890 307
rect -870 287 -850 307
rect -830 287 -810 307
rect -790 287 -770 307
rect -740 287 -710 307
rect -3470 219 -3450 239
rect -3430 219 -3410 239
rect -3390 219 -3370 239
rect -3350 219 -3330 239
rect -3310 219 -3290 239
rect -3270 219 -3250 239
rect -3230 219 -3210 239
rect -3190 219 -3170 239
rect -3150 219 -3130 239
rect -3110 219 -3090 239
rect -3070 219 -3050 239
rect -3030 219 -3010 239
rect -2990 219 -2970 239
rect -2950 219 -2930 239
rect -2910 219 -2890 239
rect -2870 219 -2850 239
rect -2830 219 -2810 239
rect -2790 219 -2770 239
rect -2750 219 -2730 239
rect -2710 219 -2690 239
rect -2670 219 -2650 239
rect -2630 219 -2610 239
rect -2590 219 -2570 239
rect -2550 219 -2530 239
rect -2510 219 -2490 239
rect -2470 219 -2450 239
rect -2430 219 -2410 239
rect -2390 219 -2370 239
rect -2350 219 -2330 239
rect -2310 219 -2290 239
rect -2270 219 -2250 239
rect -2230 219 -2210 239
rect -2190 219 -2170 239
rect -2150 219 -2130 239
rect -2110 219 -2090 239
rect -2070 219 -2050 239
rect -2030 219 -2010 239
rect -1990 219 -1970 239
rect -1950 219 -1930 239
rect -1910 219 -1890 239
rect -1870 219 -1850 239
rect -1830 219 -1810 239
rect -1790 219 -1770 239
rect -1750 219 -1730 239
rect -1710 219 -1690 239
rect -1670 219 -1650 239
rect -1630 219 -1610 239
rect -1590 219 -1570 239
rect -1550 219 -1530 239
rect -1510 219 -1490 239
rect -1470 219 -1450 239
rect -1430 219 -1410 239
rect -1390 219 -1370 239
rect -1350 219 -1330 239
rect -1310 219 -1290 239
rect -1270 219 -1250 239
rect -1230 219 -1210 239
rect -1190 219 -1170 239
rect -1150 219 -1130 239
rect -1110 219 -1090 239
rect -1070 219 -1050 239
rect -1030 219 -1010 239
rect -990 219 -970 239
rect -950 219 -930 239
rect -910 219 -890 239
rect -870 219 -850 239
rect -830 219 -810 239
rect -790 219 -770 239
rect -740 219 -710 239
rect -3470 151 -3450 171
rect -3430 151 -3410 171
rect -3390 151 -3370 171
rect -3350 151 -3330 171
rect -3310 151 -3290 171
rect -3270 151 -3250 171
rect -3230 151 -3210 171
rect -3190 151 -3170 171
rect -3150 151 -3130 171
rect -3110 151 -3090 171
rect -3070 151 -3050 171
rect -3030 151 -3010 171
rect -2990 151 -2970 171
rect -2950 151 -2930 171
rect -2910 151 -2890 171
rect -2870 151 -2850 171
rect -2830 151 -2810 171
rect -2790 151 -2770 171
rect -2750 151 -2730 171
rect -2710 151 -2690 171
rect -2670 151 -2650 171
rect -2630 151 -2610 171
rect -2590 151 -2570 171
rect -2550 151 -2530 171
rect -2510 151 -2490 171
rect -2470 151 -2450 171
rect -2430 151 -2410 171
rect -2390 151 -2370 171
rect -2350 151 -2330 171
rect -2310 151 -2290 171
rect -2270 151 -2250 171
rect -2230 151 -2210 171
rect -2190 151 -2170 171
rect -2150 151 -2130 171
rect -2110 151 -2090 171
rect -2070 151 -2050 171
rect -2030 151 -2010 171
rect -1990 151 -1970 171
rect -1950 151 -1930 171
rect -1910 151 -1890 171
rect -1870 151 -1850 171
rect -1830 151 -1810 171
rect -1790 151 -1770 171
rect -1750 151 -1730 171
rect -1710 151 -1690 171
rect -1670 151 -1650 171
rect -1630 151 -1610 171
rect -1590 151 -1570 171
rect -1550 151 -1530 171
rect -1510 151 -1490 171
rect -1470 151 -1450 171
rect -1430 151 -1410 171
rect -1390 151 -1370 171
rect -1350 151 -1330 171
rect -1310 151 -1290 171
rect -1270 151 -1250 171
rect -1230 151 -1210 171
rect -1190 151 -1170 171
rect -1150 151 -1130 171
rect -1110 151 -1090 171
rect -1070 151 -1050 171
rect -1030 151 -1010 171
rect -990 151 -970 171
rect -950 151 -930 171
rect -910 151 -890 171
rect -870 151 -850 171
rect -830 151 -810 171
rect -790 151 -770 171
rect -740 151 -710 171
rect -3470 83 -3450 103
rect -3430 83 -3410 103
rect -3390 83 -3370 103
rect -3350 83 -3330 103
rect -3310 83 -3290 103
rect -3270 83 -3250 103
rect -3230 83 -3210 103
rect -3190 83 -3170 103
rect -3150 83 -3130 103
rect -3110 83 -3090 103
rect -3070 83 -3050 103
rect -3030 83 -3010 103
rect -2990 83 -2970 103
rect -2950 83 -2930 103
rect -2910 83 -2890 103
rect -2870 83 -2850 103
rect -2830 83 -2810 103
rect -2790 83 -2770 103
rect -2750 83 -2730 103
rect -2710 83 -2690 103
rect -2670 83 -2650 103
rect -2630 83 -2610 103
rect -2590 83 -2570 103
rect -2550 83 -2530 103
rect -2510 83 -2490 103
rect -2470 83 -2450 103
rect -2430 83 -2410 103
rect -2390 83 -2370 103
rect -2350 83 -2330 103
rect -2310 83 -2290 103
rect -2270 83 -2250 103
rect -2230 83 -2210 103
rect -2190 83 -2170 103
rect -2150 83 -2130 103
rect -2110 83 -2090 103
rect -2070 83 -2050 103
rect -2030 83 -2010 103
rect -1990 83 -1970 103
rect -1950 83 -1930 103
rect -1910 83 -1890 103
rect -1870 83 -1850 103
rect -1830 83 -1810 103
rect -1790 83 -1770 103
rect -1750 83 -1730 103
rect -1710 83 -1690 103
rect -1670 83 -1650 103
rect -1630 83 -1610 103
rect -1590 83 -1570 103
rect -1550 83 -1530 103
rect -1510 83 -1490 103
rect -1470 83 -1450 103
rect -1430 83 -1410 103
rect -1390 83 -1370 103
rect -1350 83 -1330 103
rect -1310 83 -1290 103
rect -1270 83 -1250 103
rect -1230 83 -1210 103
rect -1190 83 -1170 103
rect -1150 83 -1130 103
rect -1110 83 -1090 103
rect -1070 83 -1050 103
rect -1030 83 -1010 103
rect -990 83 -970 103
rect -950 83 -930 103
rect -910 83 -890 103
rect -870 83 -850 103
rect -830 83 -810 103
rect -790 83 -770 103
rect -740 83 -710 103
rect -3470 15 -3450 35
rect -3430 15 -3410 35
rect -3390 15 -3370 35
rect -3350 15 -3330 35
rect -3310 15 -3290 35
rect -3270 15 -3250 35
rect -3230 15 -3210 35
rect -3190 15 -3170 35
rect -3150 15 -3130 35
rect -3110 15 -3090 35
rect -3070 15 -3050 35
rect -3030 15 -3010 35
rect -2990 15 -2970 35
rect -2950 15 -2930 35
rect -2910 15 -2890 35
rect -2870 15 -2850 35
rect -2830 15 -2810 35
rect -2790 15 -2770 35
rect -2750 15 -2730 35
rect -2710 15 -2690 35
rect -2670 15 -2650 35
rect -2630 15 -2610 35
rect -2590 15 -2570 35
rect -2550 15 -2530 35
rect -2510 15 -2490 35
rect -2470 15 -2450 35
rect -2430 15 -2410 35
rect -2390 15 -2370 35
rect -2350 15 -2330 35
rect -2310 15 -2290 35
rect -2270 15 -2250 35
rect -2230 15 -2210 35
rect -2190 15 -2170 35
rect -2150 15 -2130 35
rect -2110 15 -2090 35
rect -2070 15 -2050 35
rect -2030 15 -2010 35
rect -1990 15 -1970 35
rect -1950 15 -1930 35
rect -1910 15 -1890 35
rect -1870 15 -1850 35
rect -1830 15 -1810 35
rect -1790 15 -1770 35
rect -1750 15 -1730 35
rect -1710 15 -1690 35
rect -1670 15 -1650 35
rect -1630 15 -1610 35
rect -1590 15 -1570 35
rect -1550 15 -1530 35
rect -1510 15 -1490 35
rect -1470 15 -1450 35
rect -1430 15 -1410 35
rect -1390 15 -1370 35
rect -1350 15 -1330 35
rect -1310 15 -1290 35
rect -1270 15 -1250 35
rect -1230 15 -1210 35
rect -1190 15 -1170 35
rect -1150 15 -1130 35
rect -1110 15 -1090 35
rect -1070 15 -1050 35
rect -1030 15 -1010 35
rect -990 15 -970 35
rect -950 15 -930 35
rect -910 15 -890 35
rect -870 15 -850 35
rect -830 15 -810 35
rect -790 15 -770 35
rect -740 15 -710 35
<< psubdiff >>
rect -3485 -80 -985 -70
rect -3485 -100 -3470 -80
rect -3450 -100 -3430 -80
rect -3410 -100 -3390 -80
rect -3370 -100 -3350 -80
rect -3330 -100 -3310 -80
rect -3290 -100 -3270 -80
rect -3250 -100 -3230 -80
rect -3210 -100 -3190 -80
rect -3170 -100 -3150 -80
rect -3130 -100 -3110 -80
rect -3090 -100 -3070 -80
rect -3050 -100 -3030 -80
rect -3010 -100 -2990 -80
rect -2970 -100 -2950 -80
rect -2930 -100 -2910 -80
rect -2890 -100 -2870 -80
rect -2850 -100 -2830 -80
rect -2810 -100 -2790 -80
rect -2770 -100 -2750 -80
rect -2730 -100 -2710 -80
rect -2690 -100 -2670 -80
rect -2650 -100 -2630 -80
rect -2610 -100 -2590 -80
rect -2570 -100 -2550 -80
rect -2530 -100 -2510 -80
rect -2490 -100 -2470 -80
rect -2450 -100 -2430 -80
rect -2410 -100 -2390 -80
rect -2370 -100 -2350 -80
rect -2330 -100 -2310 -80
rect -2290 -100 -2270 -80
rect -2250 -100 -2230 -80
rect -2210 -100 -2190 -80
rect -2170 -100 -2150 -80
rect -2130 -100 -2110 -80
rect -2090 -100 -2070 -80
rect -2050 -100 -2030 -80
rect -2010 -100 -1990 -80
rect -1970 -100 -1950 -80
rect -1930 -100 -1910 -80
rect -1890 -100 -1870 -80
rect -1850 -100 -1830 -80
rect -1810 -100 -1790 -80
rect -1770 -100 -1750 -80
rect -1730 -100 -1710 -80
rect -1690 -100 -1670 -80
rect -1650 -100 -1630 -80
rect -1610 -100 -1590 -80
rect -1570 -100 -1550 -80
rect -1530 -100 -1510 -80
rect -1490 -100 -1470 -80
rect -1450 -100 -1430 -80
rect -1410 -100 -1390 -80
rect -1370 -100 -1350 -80
rect -1330 -100 -1310 -80
rect -1290 -100 -1270 -80
rect -1250 -100 -1230 -80
rect -1210 -100 -1190 -80
rect -1170 -100 -1150 -80
rect -1130 -100 -1110 -80
rect -1090 -100 -1070 -80
rect -1050 -100 -1030 -80
rect -1005 -100 -985 -80
rect -3485 -110 -985 -100
rect -3485 -610 -985 -600
rect -3485 -630 -3470 -610
rect -3450 -630 -3430 -610
rect -3410 -630 -3390 -610
rect -3370 -630 -3350 -610
rect -3330 -630 -3310 -610
rect -3290 -630 -3270 -610
rect -3250 -630 -3230 -610
rect -3210 -630 -3190 -610
rect -3170 -630 -3150 -610
rect -3130 -630 -3110 -610
rect -3090 -630 -3070 -610
rect -3050 -630 -3030 -610
rect -3010 -630 -2990 -610
rect -2970 -630 -2950 -610
rect -2930 -630 -2910 -610
rect -2890 -630 -2870 -610
rect -2850 -630 -2830 -610
rect -2810 -630 -2790 -610
rect -2770 -630 -2750 -610
rect -2730 -630 -2710 -610
rect -2690 -630 -2670 -610
rect -2650 -630 -2630 -610
rect -2610 -630 -2590 -610
rect -2570 -630 -2550 -610
rect -2530 -630 -2510 -610
rect -2490 -630 -2470 -610
rect -2450 -630 -2430 -610
rect -2410 -630 -2390 -610
rect -2370 -630 -2350 -610
rect -2330 -630 -2310 -610
rect -2290 -630 -2270 -610
rect -2250 -630 -2230 -610
rect -2210 -630 -2190 -610
rect -2170 -630 -2150 -610
rect -2130 -630 -2110 -610
rect -2090 -630 -2070 -610
rect -2050 -630 -2030 -610
rect -2010 -630 -1990 -610
rect -1970 -630 -1950 -610
rect -1930 -630 -1910 -610
rect -1890 -630 -1870 -610
rect -1850 -630 -1830 -610
rect -1810 -630 -1790 -610
rect -1770 -630 -1750 -610
rect -1730 -630 -1710 -610
rect -1690 -630 -1670 -610
rect -1650 -630 -1630 -610
rect -1610 -630 -1590 -610
rect -1570 -630 -1550 -610
rect -1530 -630 -1510 -610
rect -1490 -630 -1470 -610
rect -1450 -630 -1430 -610
rect -1410 -630 -1390 -610
rect -1370 -630 -1350 -610
rect -1330 -630 -1310 -610
rect -1290 -630 -1270 -610
rect -1250 -630 -1230 -610
rect -1210 -630 -1190 -610
rect -1170 -630 -1150 -610
rect -1130 -630 -1110 -610
rect -1090 -630 -1070 -610
rect -1050 -630 -1030 -610
rect -1005 -630 -985 -610
rect -3485 -640 -985 -630
<< nsubdiff >>
rect -3485 1435 -685 1445
rect -3485 1415 -3470 1435
rect -3450 1415 -3430 1435
rect -3410 1415 -3390 1435
rect -3370 1415 -3350 1435
rect -3330 1415 -3310 1435
rect -3290 1415 -3270 1435
rect -3250 1415 -3230 1435
rect -3210 1415 -3190 1435
rect -3170 1415 -3150 1435
rect -3130 1415 -3110 1435
rect -3090 1415 -3070 1435
rect -3050 1415 -3030 1435
rect -3010 1415 -2990 1435
rect -2970 1415 -2950 1435
rect -2930 1415 -2910 1435
rect -2890 1415 -2870 1435
rect -2850 1415 -2830 1435
rect -2810 1415 -2790 1435
rect -2770 1415 -2750 1435
rect -2730 1415 -2710 1435
rect -2690 1415 -2670 1435
rect -2650 1415 -2630 1435
rect -2610 1415 -2590 1435
rect -2570 1415 -2550 1435
rect -2530 1415 -2510 1435
rect -2490 1415 -2470 1435
rect -2450 1415 -2430 1435
rect -2410 1415 -2390 1435
rect -2370 1415 -2350 1435
rect -2330 1415 -2310 1435
rect -2290 1415 -2270 1435
rect -2250 1415 -2230 1435
rect -2210 1415 -2190 1435
rect -2170 1415 -2150 1435
rect -2130 1415 -2110 1435
rect -2090 1415 -2070 1435
rect -2050 1415 -2030 1435
rect -2010 1415 -1990 1435
rect -1970 1415 -1950 1435
rect -1930 1415 -1910 1435
rect -1890 1415 -1870 1435
rect -1850 1415 -1830 1435
rect -1810 1415 -1790 1435
rect -1770 1415 -1750 1435
rect -1730 1415 -1710 1435
rect -1690 1415 -1670 1435
rect -1650 1415 -1630 1435
rect -1610 1415 -1590 1435
rect -1570 1415 -1550 1435
rect -1530 1415 -1510 1435
rect -1490 1415 -1470 1435
rect -1450 1415 -1430 1435
rect -1410 1415 -1390 1435
rect -1370 1415 -1350 1435
rect -1330 1415 -1310 1435
rect -1290 1415 -1270 1435
rect -1250 1415 -1230 1435
rect -1210 1415 -1190 1435
rect -1170 1415 -1150 1435
rect -1130 1415 -1110 1435
rect -1090 1415 -1070 1435
rect -1050 1415 -1030 1435
rect -1010 1415 -990 1435
rect -970 1415 -950 1435
rect -930 1415 -910 1435
rect -890 1415 -870 1435
rect -850 1415 -830 1435
rect -810 1415 -790 1435
rect -770 1415 -740 1435
rect -710 1415 -685 1435
rect -3485 1405 -685 1415
rect -3485 -5 -685 5
rect -3485 -25 -3470 -5
rect -3450 -25 -3430 -5
rect -3410 -25 -3390 -5
rect -3370 -25 -3350 -5
rect -3330 -25 -3310 -5
rect -3290 -25 -3270 -5
rect -3250 -25 -3230 -5
rect -3210 -25 -3190 -5
rect -3170 -25 -3150 -5
rect -3130 -25 -3110 -5
rect -3090 -25 -3070 -5
rect -3050 -25 -3030 -5
rect -3010 -25 -2990 -5
rect -2970 -25 -2950 -5
rect -2930 -25 -2910 -5
rect -2890 -25 -2870 -5
rect -2850 -25 -2830 -5
rect -2810 -25 -2790 -5
rect -2770 -25 -2750 -5
rect -2730 -25 -2710 -5
rect -2690 -25 -2670 -5
rect -2650 -25 -2630 -5
rect -2610 -25 -2590 -5
rect -2570 -25 -2550 -5
rect -2530 -25 -2510 -5
rect -2490 -25 -2470 -5
rect -2450 -25 -2430 -5
rect -2410 -25 -2390 -5
rect -2370 -25 -2350 -5
rect -2330 -25 -2310 -5
rect -2290 -25 -2270 -5
rect -2250 -25 -2230 -5
rect -2210 -25 -2190 -5
rect -2170 -25 -2150 -5
rect -2130 -25 -2110 -5
rect -2090 -25 -2070 -5
rect -2050 -25 -2030 -5
rect -2010 -25 -1990 -5
rect -1970 -25 -1950 -5
rect -1930 -25 -1910 -5
rect -1890 -25 -1870 -5
rect -1850 -25 -1830 -5
rect -1810 -25 -1790 -5
rect -1770 -25 -1750 -5
rect -1730 -25 -1710 -5
rect -1690 -25 -1670 -5
rect -1650 -25 -1630 -5
rect -1610 -25 -1590 -5
rect -1570 -25 -1550 -5
rect -1530 -25 -1510 -5
rect -1490 -25 -1470 -5
rect -1450 -25 -1430 -5
rect -1410 -25 -1390 -5
rect -1370 -25 -1350 -5
rect -1330 -25 -1310 -5
rect -1290 -25 -1270 -5
rect -1250 -25 -1230 -5
rect -1210 -25 -1190 -5
rect -1170 -25 -1150 -5
rect -1130 -25 -1110 -5
rect -1090 -25 -1070 -5
rect -1050 -25 -1030 -5
rect -1010 -25 -990 -5
rect -970 -25 -950 -5
rect -930 -25 -910 -5
rect -890 -25 -870 -5
rect -850 -25 -830 -5
rect -810 -25 -790 -5
rect -770 -25 -740 -5
rect -710 -25 -685 -5
rect -3485 -35 -685 -25
<< psubdiffcont >>
rect -3470 -100 -3450 -80
rect -3430 -100 -3410 -80
rect -3390 -100 -3370 -80
rect -3350 -100 -3330 -80
rect -3310 -100 -3290 -80
rect -3270 -100 -3250 -80
rect -3230 -100 -3210 -80
rect -3190 -100 -3170 -80
rect -3150 -100 -3130 -80
rect -3110 -100 -3090 -80
rect -3070 -100 -3050 -80
rect -3030 -100 -3010 -80
rect -2990 -100 -2970 -80
rect -2950 -100 -2930 -80
rect -2910 -100 -2890 -80
rect -2870 -100 -2850 -80
rect -2830 -100 -2810 -80
rect -2790 -100 -2770 -80
rect -2750 -100 -2730 -80
rect -2710 -100 -2690 -80
rect -2670 -100 -2650 -80
rect -2630 -100 -2610 -80
rect -2590 -100 -2570 -80
rect -2550 -100 -2530 -80
rect -2510 -100 -2490 -80
rect -2470 -100 -2450 -80
rect -2430 -100 -2410 -80
rect -2390 -100 -2370 -80
rect -2350 -100 -2330 -80
rect -2310 -100 -2290 -80
rect -2270 -100 -2250 -80
rect -2230 -100 -2210 -80
rect -2190 -100 -2170 -80
rect -2150 -100 -2130 -80
rect -2110 -100 -2090 -80
rect -2070 -100 -2050 -80
rect -2030 -100 -2010 -80
rect -1990 -100 -1970 -80
rect -1950 -100 -1930 -80
rect -1910 -100 -1890 -80
rect -1870 -100 -1850 -80
rect -1830 -100 -1810 -80
rect -1790 -100 -1770 -80
rect -1750 -100 -1730 -80
rect -1710 -100 -1690 -80
rect -1670 -100 -1650 -80
rect -1630 -100 -1610 -80
rect -1590 -100 -1570 -80
rect -1550 -100 -1530 -80
rect -1510 -100 -1490 -80
rect -1470 -100 -1450 -80
rect -1430 -100 -1410 -80
rect -1390 -100 -1370 -80
rect -1350 -100 -1330 -80
rect -1310 -100 -1290 -80
rect -1270 -100 -1250 -80
rect -1230 -100 -1210 -80
rect -1190 -100 -1170 -80
rect -1150 -100 -1130 -80
rect -1110 -100 -1090 -80
rect -1070 -100 -1050 -80
rect -1030 -100 -1005 -80
rect -3470 -630 -3450 -610
rect -3430 -630 -3410 -610
rect -3390 -630 -3370 -610
rect -3350 -630 -3330 -610
rect -3310 -630 -3290 -610
rect -3270 -630 -3250 -610
rect -3230 -630 -3210 -610
rect -3190 -630 -3170 -610
rect -3150 -630 -3130 -610
rect -3110 -630 -3090 -610
rect -3070 -630 -3050 -610
rect -3030 -630 -3010 -610
rect -2990 -630 -2970 -610
rect -2950 -630 -2930 -610
rect -2910 -630 -2890 -610
rect -2870 -630 -2850 -610
rect -2830 -630 -2810 -610
rect -2790 -630 -2770 -610
rect -2750 -630 -2730 -610
rect -2710 -630 -2690 -610
rect -2670 -630 -2650 -610
rect -2630 -630 -2610 -610
rect -2590 -630 -2570 -610
rect -2550 -630 -2530 -610
rect -2510 -630 -2490 -610
rect -2470 -630 -2450 -610
rect -2430 -630 -2410 -610
rect -2390 -630 -2370 -610
rect -2350 -630 -2330 -610
rect -2310 -630 -2290 -610
rect -2270 -630 -2250 -610
rect -2230 -630 -2210 -610
rect -2190 -630 -2170 -610
rect -2150 -630 -2130 -610
rect -2110 -630 -2090 -610
rect -2070 -630 -2050 -610
rect -2030 -630 -2010 -610
rect -1990 -630 -1970 -610
rect -1950 -630 -1930 -610
rect -1910 -630 -1890 -610
rect -1870 -630 -1850 -610
rect -1830 -630 -1810 -610
rect -1790 -630 -1770 -610
rect -1750 -630 -1730 -610
rect -1710 -630 -1690 -610
rect -1670 -630 -1650 -610
rect -1630 -630 -1610 -610
rect -1590 -630 -1570 -610
rect -1550 -630 -1530 -610
rect -1510 -630 -1490 -610
rect -1470 -630 -1450 -610
rect -1430 -630 -1410 -610
rect -1390 -630 -1370 -610
rect -1350 -630 -1330 -610
rect -1310 -630 -1290 -610
rect -1270 -630 -1250 -610
rect -1230 -630 -1210 -610
rect -1190 -630 -1170 -610
rect -1150 -630 -1130 -610
rect -1110 -630 -1090 -610
rect -1070 -630 -1050 -610
rect -1030 -630 -1005 -610
<< nsubdiffcont >>
rect -3470 1415 -3450 1435
rect -3430 1415 -3410 1435
rect -3390 1415 -3370 1435
rect -3350 1415 -3330 1435
rect -3310 1415 -3290 1435
rect -3270 1415 -3250 1435
rect -3230 1415 -3210 1435
rect -3190 1415 -3170 1435
rect -3150 1415 -3130 1435
rect -3110 1415 -3090 1435
rect -3070 1415 -3050 1435
rect -3030 1415 -3010 1435
rect -2990 1415 -2970 1435
rect -2950 1415 -2930 1435
rect -2910 1415 -2890 1435
rect -2870 1415 -2850 1435
rect -2830 1415 -2810 1435
rect -2790 1415 -2770 1435
rect -2750 1415 -2730 1435
rect -2710 1415 -2690 1435
rect -2670 1415 -2650 1435
rect -2630 1415 -2610 1435
rect -2590 1415 -2570 1435
rect -2550 1415 -2530 1435
rect -2510 1415 -2490 1435
rect -2470 1415 -2450 1435
rect -2430 1415 -2410 1435
rect -2390 1415 -2370 1435
rect -2350 1415 -2330 1435
rect -2310 1415 -2290 1435
rect -2270 1415 -2250 1435
rect -2230 1415 -2210 1435
rect -2190 1415 -2170 1435
rect -2150 1415 -2130 1435
rect -2110 1415 -2090 1435
rect -2070 1415 -2050 1435
rect -2030 1415 -2010 1435
rect -1990 1415 -1970 1435
rect -1950 1415 -1930 1435
rect -1910 1415 -1890 1435
rect -1870 1415 -1850 1435
rect -1830 1415 -1810 1435
rect -1790 1415 -1770 1435
rect -1750 1415 -1730 1435
rect -1710 1415 -1690 1435
rect -1670 1415 -1650 1435
rect -1630 1415 -1610 1435
rect -1590 1415 -1570 1435
rect -1550 1415 -1530 1435
rect -1510 1415 -1490 1435
rect -1470 1415 -1450 1435
rect -1430 1415 -1410 1435
rect -1390 1415 -1370 1435
rect -1350 1415 -1330 1435
rect -1310 1415 -1290 1435
rect -1270 1415 -1250 1435
rect -1230 1415 -1210 1435
rect -1190 1415 -1170 1435
rect -1150 1415 -1130 1435
rect -1110 1415 -1090 1435
rect -1070 1415 -1050 1435
rect -1030 1415 -1010 1435
rect -990 1415 -970 1435
rect -950 1415 -930 1435
rect -910 1415 -890 1435
rect -870 1415 -850 1435
rect -830 1415 -810 1435
rect -790 1415 -770 1435
rect -740 1415 -710 1435
rect -3470 -25 -3450 -5
rect -3430 -25 -3410 -5
rect -3390 -25 -3370 -5
rect -3350 -25 -3330 -5
rect -3310 -25 -3290 -5
rect -3270 -25 -3250 -5
rect -3230 -25 -3210 -5
rect -3190 -25 -3170 -5
rect -3150 -25 -3130 -5
rect -3110 -25 -3090 -5
rect -3070 -25 -3050 -5
rect -3030 -25 -3010 -5
rect -2990 -25 -2970 -5
rect -2950 -25 -2930 -5
rect -2910 -25 -2890 -5
rect -2870 -25 -2850 -5
rect -2830 -25 -2810 -5
rect -2790 -25 -2770 -5
rect -2750 -25 -2730 -5
rect -2710 -25 -2690 -5
rect -2670 -25 -2650 -5
rect -2630 -25 -2610 -5
rect -2590 -25 -2570 -5
rect -2550 -25 -2530 -5
rect -2510 -25 -2490 -5
rect -2470 -25 -2450 -5
rect -2430 -25 -2410 -5
rect -2390 -25 -2370 -5
rect -2350 -25 -2330 -5
rect -2310 -25 -2290 -5
rect -2270 -25 -2250 -5
rect -2230 -25 -2210 -5
rect -2190 -25 -2170 -5
rect -2150 -25 -2130 -5
rect -2110 -25 -2090 -5
rect -2070 -25 -2050 -5
rect -2030 -25 -2010 -5
rect -1990 -25 -1970 -5
rect -1950 -25 -1930 -5
rect -1910 -25 -1890 -5
rect -1870 -25 -1850 -5
rect -1830 -25 -1810 -5
rect -1790 -25 -1770 -5
rect -1750 -25 -1730 -5
rect -1710 -25 -1690 -5
rect -1670 -25 -1650 -5
rect -1630 -25 -1610 -5
rect -1590 -25 -1570 -5
rect -1550 -25 -1530 -5
rect -1510 -25 -1490 -5
rect -1470 -25 -1450 -5
rect -1430 -25 -1410 -5
rect -1390 -25 -1370 -5
rect -1350 -25 -1330 -5
rect -1310 -25 -1290 -5
rect -1270 -25 -1250 -5
rect -1230 -25 -1210 -5
rect -1190 -25 -1170 -5
rect -1150 -25 -1130 -5
rect -1110 -25 -1090 -5
rect -1070 -25 -1050 -5
rect -1030 -25 -1010 -5
rect -990 -25 -970 -5
rect -950 -25 -930 -5
rect -910 -25 -890 -5
rect -870 -25 -850 -5
rect -830 -25 -810 -5
rect -790 -25 -770 -5
rect -740 -25 -710 -5
<< poly >>
rect -3665 1360 -3505 1370
rect -3665 1340 -3655 1360
rect -3635 1340 -3615 1360
rect -3595 1340 -3575 1360
rect -3555 1340 -3535 1360
rect -3510 1342 -3485 1360
rect -685 1342 -670 1360
rect -3510 1340 -3505 1342
rect -3665 1330 -3505 1340
rect -3665 1292 -3505 1300
rect -3665 1290 -3485 1292
rect -3665 1270 -3655 1290
rect -3635 1270 -3615 1290
rect -3595 1270 -3575 1290
rect -3555 1270 -3535 1290
rect -3510 1274 -3485 1290
rect -685 1274 -670 1292
rect -3510 1270 -3505 1274
rect -3665 1260 -3505 1270
rect -3665 1225 -3505 1235
rect -3665 1205 -3655 1225
rect -3635 1205 -3615 1225
rect -3595 1205 -3575 1225
rect -3555 1205 -3535 1225
rect -3510 1224 -3505 1225
rect -3510 1206 -3485 1224
rect -685 1206 -670 1224
rect -3510 1205 -3505 1206
rect -3665 1195 -3505 1205
rect -3665 1160 -3505 1170
rect -3665 1140 -3655 1160
rect -3635 1140 -3615 1160
rect -3595 1140 -3575 1160
rect -3555 1140 -3535 1160
rect -3510 1156 -3505 1160
rect -3510 1140 -3485 1156
rect -3665 1138 -3485 1140
rect -685 1138 -670 1156
rect -3665 1130 -3505 1138
rect -3665 1090 -3505 1100
rect -3665 1070 -3655 1090
rect -3635 1070 -3615 1090
rect -3595 1070 -3575 1090
rect -3555 1070 -3535 1090
rect -3510 1088 -3505 1090
rect -3510 1070 -3485 1088
rect -685 1070 -670 1088
rect -3665 1060 -3505 1070
rect -3665 1020 -3505 1030
rect -3665 1000 -3655 1020
rect -3635 1000 -3615 1020
rect -3595 1000 -3575 1020
rect -3555 1000 -3535 1020
rect -3510 1002 -3485 1020
rect -685 1002 -670 1020
rect -3510 1000 -3505 1002
rect -3665 990 -3505 1000
rect -3665 955 -3505 965
rect -3665 935 -3655 955
rect -3635 935 -3615 955
rect -3595 935 -3575 955
rect -3555 935 -3535 955
rect -3510 952 -3505 955
rect -3510 935 -3485 952
rect -3665 934 -3485 935
rect -685 934 -670 952
rect -3665 925 -3505 934
rect -3665 885 -3505 895
rect -3665 865 -3655 885
rect -3635 865 -3615 885
rect -3595 865 -3575 885
rect -3555 865 -3535 885
rect -3510 884 -3505 885
rect -3510 866 -3485 884
rect -685 866 -670 884
rect -3510 865 -3505 866
rect -3665 855 -3505 865
rect -3665 816 -3505 825
rect -3665 815 -3485 816
rect -3665 795 -3655 815
rect -3635 795 -3615 815
rect -3595 795 -3575 815
rect -3555 795 -3535 815
rect -3510 798 -3485 815
rect -685 798 -670 816
rect -3510 795 -3505 798
rect -3665 785 -3505 795
rect -3665 750 -3505 760
rect -3665 730 -3655 750
rect -3635 730 -3615 750
rect -3595 730 -3575 750
rect -3555 730 -3535 750
rect -3510 748 -3505 750
rect -3510 730 -3485 748
rect -685 730 -670 748
rect -3665 720 -3505 730
rect -3665 680 -3505 690
rect -3665 660 -3655 680
rect -3635 660 -3615 680
rect -3595 660 -3575 680
rect -3555 660 -3535 680
rect -3510 662 -3485 680
rect -685 662 -670 680
rect -3510 660 -3505 662
rect -3665 650 -3505 660
rect -3665 615 -3505 625
rect -3665 595 -3655 615
rect -3635 595 -3615 615
rect -3595 595 -3575 615
rect -3555 595 -3535 615
rect -3510 612 -3505 615
rect -3510 595 -3485 612
rect -3665 594 -3485 595
rect -685 594 -670 612
rect -3665 585 -3505 594
rect -3665 545 -3505 555
rect -3665 525 -3655 545
rect -3635 525 -3615 545
rect -3595 525 -3575 545
rect -3555 525 -3535 545
rect -3510 544 -3505 545
rect -3510 526 -3485 544
rect -685 526 -670 544
rect -3510 525 -3505 526
rect -3665 515 -3505 525
rect -3665 476 -3505 485
rect -3665 475 -3485 476
rect -3665 455 -3655 475
rect -3635 455 -3615 475
rect -3595 455 -3575 475
rect -3555 455 -3535 475
rect -3510 458 -3485 475
rect -685 458 -670 476
rect -3510 455 -3505 458
rect -3665 445 -3505 455
rect -3665 408 -3505 415
rect -3665 405 -3485 408
rect -3665 385 -3655 405
rect -3635 385 -3615 405
rect -3595 385 -3575 405
rect -3555 385 -3535 405
rect -3510 390 -3485 405
rect -685 390 -670 408
rect -3510 385 -3505 390
rect -3665 375 -3505 385
rect -3665 340 -3505 350
rect -3665 320 -3655 340
rect -3635 320 -3615 340
rect -3595 320 -3575 340
rect -3555 320 -3535 340
rect -3510 322 -3485 340
rect -685 322 -670 340
rect -3510 320 -3505 322
rect -3665 310 -3505 320
rect -3665 275 -3505 285
rect -3665 255 -3655 275
rect -3635 255 -3615 275
rect -3595 255 -3575 275
rect -3555 255 -3535 275
rect -3510 272 -3505 275
rect -3510 255 -3485 272
rect -3665 254 -3485 255
rect -685 254 -670 272
rect -3665 245 -3505 254
rect -3665 205 -3505 215
rect -3665 185 -3655 205
rect -3635 185 -3615 205
rect -3595 185 -3575 205
rect -3555 185 -3535 205
rect -3510 204 -3505 205
rect -3510 186 -3485 204
rect -685 186 -670 204
rect -3510 185 -3505 186
rect -3665 175 -3505 185
rect -3665 136 -3505 145
rect -3665 135 -3485 136
rect -3665 115 -3655 135
rect -3635 115 -3615 135
rect -3595 115 -3575 135
rect -3555 115 -3535 135
rect -3510 118 -3485 135
rect -685 118 -670 136
rect -3510 115 -3505 118
rect -3665 105 -3505 115
rect -3665 70 -3505 80
rect -3665 50 -3655 70
rect -3635 50 -3615 70
rect -3595 50 -3575 70
rect -3555 50 -3535 70
rect -3510 68 -3505 70
rect -3510 50 -3485 68
rect -685 50 -670 68
rect -3665 40 -3505 50
rect -3660 -180 -3500 -170
rect -3660 -205 -3650 -180
rect -3630 -205 -3610 -180
rect -3590 -205 -3570 -180
rect -3550 -205 -3530 -180
rect -3505 -185 -3500 -180
rect -3505 -200 -3485 -185
rect -985 -200 -970 -185
rect -3505 -205 -3500 -200
rect -3660 -245 -3500 -205
rect -3660 -270 -3650 -245
rect -3630 -270 -3610 -245
rect -3590 -270 -3570 -245
rect -3550 -270 -3530 -245
rect -3505 -250 -3500 -245
rect -3505 -265 -3485 -250
rect -985 -265 -970 -250
rect -3505 -270 -3500 -265
rect -3660 -310 -3500 -270
rect -3660 -335 -3650 -310
rect -3630 -335 -3610 -310
rect -3590 -335 -3570 -310
rect -3550 -335 -3530 -310
rect -3505 -315 -3500 -310
rect -3505 -330 -3485 -315
rect -985 -330 -970 -315
rect -3505 -335 -3500 -330
rect -3660 -375 -3500 -335
rect -3660 -400 -3650 -375
rect -3630 -400 -3610 -375
rect -3590 -400 -3570 -375
rect -3550 -400 -3530 -375
rect -3505 -380 -3500 -375
rect -3505 -395 -3485 -380
rect -985 -395 -970 -380
rect -3505 -400 -3500 -395
rect -3660 -440 -3500 -400
rect -3660 -465 -3650 -440
rect -3630 -465 -3610 -440
rect -3590 -465 -3570 -440
rect -3550 -465 -3530 -440
rect -3505 -445 -3500 -440
rect -3505 -460 -3485 -445
rect -985 -460 -970 -445
rect -3505 -465 -3500 -460
rect -3660 -505 -3500 -465
rect -3660 -530 -3650 -505
rect -3630 -530 -3610 -505
rect -3590 -530 -3570 -505
rect -3550 -530 -3530 -505
rect -3505 -510 -3500 -505
rect -3505 -525 -3485 -510
rect -985 -525 -970 -510
rect -3505 -530 -3500 -525
rect -3660 -540 -3500 -530
<< polycont >>
rect -3655 1340 -3635 1360
rect -3615 1340 -3595 1360
rect -3575 1340 -3555 1360
rect -3535 1340 -3510 1360
rect -3655 1270 -3635 1290
rect -3615 1270 -3595 1290
rect -3575 1270 -3555 1290
rect -3535 1270 -3510 1290
rect -3655 1205 -3635 1225
rect -3615 1205 -3595 1225
rect -3575 1205 -3555 1225
rect -3535 1205 -3510 1225
rect -3655 1140 -3635 1160
rect -3615 1140 -3595 1160
rect -3575 1140 -3555 1160
rect -3535 1140 -3510 1160
rect -3655 1070 -3635 1090
rect -3615 1070 -3595 1090
rect -3575 1070 -3555 1090
rect -3535 1070 -3510 1090
rect -3655 1000 -3635 1020
rect -3615 1000 -3595 1020
rect -3575 1000 -3555 1020
rect -3535 1000 -3510 1020
rect -3655 935 -3635 955
rect -3615 935 -3595 955
rect -3575 935 -3555 955
rect -3535 935 -3510 955
rect -3655 865 -3635 885
rect -3615 865 -3595 885
rect -3575 865 -3555 885
rect -3535 865 -3510 885
rect -3655 795 -3635 815
rect -3615 795 -3595 815
rect -3575 795 -3555 815
rect -3535 795 -3510 815
rect -3655 730 -3635 750
rect -3615 730 -3595 750
rect -3575 730 -3555 750
rect -3535 730 -3510 750
rect -3655 660 -3635 680
rect -3615 660 -3595 680
rect -3575 660 -3555 680
rect -3535 660 -3510 680
rect -3655 595 -3635 615
rect -3615 595 -3595 615
rect -3575 595 -3555 615
rect -3535 595 -3510 615
rect -3655 525 -3635 545
rect -3615 525 -3595 545
rect -3575 525 -3555 545
rect -3535 525 -3510 545
rect -3655 455 -3635 475
rect -3615 455 -3595 475
rect -3575 455 -3555 475
rect -3535 455 -3510 475
rect -3655 385 -3635 405
rect -3615 385 -3595 405
rect -3575 385 -3555 405
rect -3535 385 -3510 405
rect -3655 320 -3635 340
rect -3615 320 -3595 340
rect -3575 320 -3555 340
rect -3535 320 -3510 340
rect -3655 255 -3635 275
rect -3615 255 -3595 275
rect -3575 255 -3555 275
rect -3535 255 -3510 275
rect -3655 185 -3635 205
rect -3615 185 -3595 205
rect -3575 185 -3555 205
rect -3535 185 -3510 205
rect -3655 115 -3635 135
rect -3615 115 -3595 135
rect -3575 115 -3555 135
rect -3535 115 -3510 135
rect -3655 50 -3635 70
rect -3615 50 -3595 70
rect -3575 50 -3555 70
rect -3535 50 -3510 70
rect -3650 -205 -3630 -180
rect -3610 -205 -3590 -180
rect -3570 -205 -3550 -180
rect -3530 -205 -3505 -180
rect -3650 -270 -3630 -245
rect -3610 -270 -3590 -245
rect -3570 -270 -3550 -245
rect -3530 -270 -3505 -245
rect -3650 -335 -3630 -310
rect -3610 -335 -3590 -310
rect -3570 -335 -3550 -310
rect -3530 -335 -3505 -310
rect -3650 -400 -3630 -375
rect -3610 -400 -3590 -375
rect -3570 -400 -3550 -375
rect -3530 -400 -3505 -375
rect -3650 -465 -3630 -440
rect -3610 -465 -3590 -440
rect -3570 -465 -3550 -440
rect -3530 -465 -3505 -440
rect -3650 -530 -3630 -505
rect -3610 -530 -3590 -505
rect -3570 -530 -3550 -505
rect -3530 -530 -3505 -505
<< locali >>
rect -3485 1435 -685 1445
rect -3485 1415 -3470 1435
rect -3450 1415 -3430 1435
rect -3410 1415 -3390 1435
rect -3370 1415 -3350 1435
rect -3330 1415 -3310 1435
rect -3290 1415 -3270 1435
rect -3250 1415 -3230 1435
rect -3210 1415 -3190 1435
rect -3170 1415 -3150 1435
rect -3130 1415 -3110 1435
rect -3090 1415 -3070 1435
rect -3050 1415 -3030 1435
rect -3010 1415 -2990 1435
rect -2970 1415 -2950 1435
rect -2930 1415 -2910 1435
rect -2890 1415 -2870 1435
rect -2850 1415 -2830 1435
rect -2810 1415 -2790 1435
rect -2770 1415 -2750 1435
rect -2730 1415 -2710 1435
rect -2690 1415 -2670 1435
rect -2650 1415 -2630 1435
rect -2610 1415 -2590 1435
rect -2570 1415 -2550 1435
rect -2530 1415 -2510 1435
rect -2490 1415 -2470 1435
rect -2450 1415 -2430 1435
rect -2410 1415 -2390 1435
rect -2370 1415 -2350 1435
rect -2330 1415 -2310 1435
rect -2290 1415 -2270 1435
rect -2250 1415 -2230 1435
rect -2210 1415 -2190 1435
rect -2170 1415 -2150 1435
rect -2130 1415 -2110 1435
rect -2090 1415 -2070 1435
rect -2050 1415 -2030 1435
rect -2010 1415 -1990 1435
rect -1970 1415 -1950 1435
rect -1930 1415 -1910 1435
rect -1890 1415 -1870 1435
rect -1850 1415 -1830 1435
rect -1810 1415 -1790 1435
rect -1770 1415 -1750 1435
rect -1730 1415 -1710 1435
rect -1690 1415 -1670 1435
rect -1650 1415 -1630 1435
rect -1610 1415 -1590 1435
rect -1570 1415 -1550 1435
rect -1530 1415 -1510 1435
rect -1490 1415 -1470 1435
rect -1450 1415 -1430 1435
rect -1410 1415 -1390 1435
rect -1370 1415 -1350 1435
rect -1330 1415 -1310 1435
rect -1290 1415 -1270 1435
rect -1250 1415 -1230 1435
rect -1210 1415 -1190 1435
rect -1170 1415 -1150 1435
rect -1130 1415 -1110 1435
rect -1090 1415 -1070 1435
rect -1050 1415 -1030 1435
rect -1010 1415 -990 1435
rect -970 1415 -950 1435
rect -930 1415 -910 1435
rect -890 1415 -870 1435
rect -850 1415 -830 1435
rect -810 1415 -790 1435
rect -770 1415 -740 1435
rect -710 1415 -685 1435
rect -3485 1395 -685 1415
rect -3485 1375 -3470 1395
rect -3450 1375 -3430 1395
rect -3410 1375 -3390 1395
rect -3370 1375 -3350 1395
rect -3330 1375 -3310 1395
rect -3290 1375 -3270 1395
rect -3250 1375 -3230 1395
rect -3210 1375 -3190 1395
rect -3170 1375 -3150 1395
rect -3130 1375 -3110 1395
rect -3090 1375 -3070 1395
rect -3050 1375 -3030 1395
rect -3010 1375 -2990 1395
rect -2970 1375 -2950 1395
rect -2930 1375 -2910 1395
rect -2890 1375 -2870 1395
rect -2850 1375 -2830 1395
rect -2810 1375 -2790 1395
rect -2770 1375 -2750 1395
rect -2730 1375 -2710 1395
rect -2690 1375 -2670 1395
rect -2650 1375 -2630 1395
rect -2610 1375 -2590 1395
rect -2570 1375 -2550 1395
rect -2530 1375 -2510 1395
rect -2490 1375 -2470 1395
rect -2450 1375 -2430 1395
rect -2410 1375 -2390 1395
rect -2370 1375 -2350 1395
rect -2330 1375 -2310 1395
rect -2290 1375 -2270 1395
rect -2250 1375 -2230 1395
rect -2210 1375 -2190 1395
rect -2170 1375 -2150 1395
rect -2130 1375 -2110 1395
rect -2090 1375 -2070 1395
rect -2050 1375 -2030 1395
rect -2010 1375 -1990 1395
rect -1970 1375 -1950 1395
rect -1930 1375 -1910 1395
rect -1890 1375 -1870 1395
rect -1850 1375 -1830 1395
rect -1810 1375 -1790 1395
rect -1770 1375 -1750 1395
rect -1730 1375 -1710 1395
rect -1690 1375 -1670 1395
rect -1650 1375 -1630 1395
rect -1610 1375 -1590 1395
rect -1570 1375 -1550 1395
rect -1530 1375 -1510 1395
rect -1490 1375 -1470 1395
rect -1450 1375 -1430 1395
rect -1410 1375 -1390 1395
rect -1370 1375 -1350 1395
rect -1330 1375 -1310 1395
rect -1290 1375 -1270 1395
rect -1250 1375 -1230 1395
rect -1210 1375 -1190 1395
rect -1170 1375 -1150 1395
rect -1130 1375 -1110 1395
rect -1090 1375 -1070 1395
rect -1050 1375 -1030 1395
rect -1010 1375 -990 1395
rect -970 1375 -950 1395
rect -930 1375 -910 1395
rect -890 1375 -870 1395
rect -850 1375 -830 1395
rect -810 1375 -790 1395
rect -770 1375 -740 1395
rect -710 1375 -685 1395
rect -3665 1360 -3510 1370
rect -3485 1365 -685 1375
rect -3665 1340 -3655 1360
rect -3635 1340 -3615 1360
rect -3595 1340 -3575 1360
rect -3555 1340 -3535 1360
rect -3665 1330 -3510 1340
rect -3485 1327 -685 1337
rect -3485 1307 -3470 1327
rect -3450 1307 -3430 1327
rect -3410 1307 -3390 1327
rect -3370 1307 -3350 1327
rect -3330 1307 -3310 1327
rect -3290 1307 -3270 1327
rect -3250 1307 -3230 1327
rect -3210 1307 -3190 1327
rect -3170 1307 -3150 1327
rect -3130 1307 -3110 1327
rect -3090 1307 -3070 1327
rect -3050 1307 -3030 1327
rect -3010 1307 -2990 1327
rect -2970 1307 -2950 1327
rect -2930 1307 -2910 1327
rect -2890 1307 -2870 1327
rect -2850 1307 -2830 1327
rect -2810 1307 -2790 1327
rect -2770 1307 -2750 1327
rect -2730 1307 -2710 1327
rect -2690 1307 -2670 1327
rect -2650 1307 -2630 1327
rect -2610 1307 -2590 1327
rect -2570 1307 -2550 1327
rect -2530 1307 -2510 1327
rect -2490 1307 -2470 1327
rect -2450 1307 -2430 1327
rect -2410 1307 -2390 1327
rect -2370 1307 -2350 1327
rect -2330 1307 -2310 1327
rect -2290 1307 -2270 1327
rect -2250 1307 -2230 1327
rect -2210 1307 -2190 1327
rect -2170 1307 -2150 1327
rect -2130 1307 -2110 1327
rect -2090 1307 -2070 1327
rect -2050 1307 -2030 1327
rect -2010 1307 -1990 1327
rect -1970 1307 -1950 1327
rect -1930 1307 -1910 1327
rect -1890 1307 -1870 1327
rect -1850 1307 -1830 1327
rect -1810 1307 -1790 1327
rect -1770 1307 -1750 1327
rect -1730 1307 -1710 1327
rect -1690 1307 -1670 1327
rect -1650 1307 -1630 1327
rect -1610 1307 -1590 1327
rect -1570 1307 -1550 1327
rect -1530 1307 -1510 1327
rect -1490 1307 -1470 1327
rect -1450 1307 -1430 1327
rect -1410 1307 -1390 1327
rect -1370 1307 -1350 1327
rect -1330 1307 -1310 1327
rect -1290 1307 -1270 1327
rect -1250 1307 -1230 1327
rect -1210 1307 -1190 1327
rect -1170 1307 -1150 1327
rect -1130 1307 -1110 1327
rect -1090 1307 -1070 1327
rect -1050 1307 -1030 1327
rect -1010 1307 -990 1327
rect -970 1307 -950 1327
rect -930 1307 -910 1327
rect -890 1307 -870 1327
rect -850 1307 -830 1327
rect -810 1307 -790 1327
rect -770 1307 -740 1327
rect -710 1307 -685 1327
rect -3665 1290 -3510 1300
rect -3485 1297 -685 1307
rect -3665 1270 -3655 1290
rect -3635 1270 -3615 1290
rect -3595 1270 -3575 1290
rect -3555 1270 -3535 1290
rect -3665 1260 -3510 1270
rect -3485 1259 -685 1269
rect -3485 1239 -3470 1259
rect -3450 1239 -3430 1259
rect -3410 1239 -3390 1259
rect -3370 1239 -3350 1259
rect -3330 1239 -3310 1259
rect -3290 1239 -3270 1259
rect -3250 1239 -3230 1259
rect -3210 1239 -3190 1259
rect -3170 1239 -3150 1259
rect -3130 1239 -3110 1259
rect -3090 1239 -3070 1259
rect -3050 1239 -3030 1259
rect -3010 1239 -2990 1259
rect -2970 1239 -2950 1259
rect -2930 1239 -2910 1259
rect -2890 1239 -2870 1259
rect -2850 1239 -2830 1259
rect -2810 1239 -2790 1259
rect -2770 1239 -2750 1259
rect -2730 1239 -2710 1259
rect -2690 1239 -2670 1259
rect -2650 1239 -2630 1259
rect -2610 1239 -2590 1259
rect -2570 1239 -2550 1259
rect -2530 1239 -2510 1259
rect -2490 1239 -2470 1259
rect -2450 1239 -2430 1259
rect -2410 1239 -2390 1259
rect -2370 1239 -2350 1259
rect -2330 1239 -2310 1259
rect -2290 1239 -2270 1259
rect -2250 1239 -2230 1259
rect -2210 1239 -2190 1259
rect -2170 1239 -2150 1259
rect -2130 1239 -2110 1259
rect -2090 1239 -2070 1259
rect -2050 1239 -2030 1259
rect -2010 1239 -1990 1259
rect -1970 1239 -1950 1259
rect -1930 1239 -1910 1259
rect -1890 1239 -1870 1259
rect -1850 1239 -1830 1259
rect -1810 1239 -1790 1259
rect -1770 1239 -1750 1259
rect -1730 1239 -1710 1259
rect -1690 1239 -1670 1259
rect -1650 1239 -1630 1259
rect -1610 1239 -1590 1259
rect -1570 1239 -1550 1259
rect -1530 1239 -1510 1259
rect -1490 1239 -1470 1259
rect -1450 1239 -1430 1259
rect -1410 1239 -1390 1259
rect -1370 1239 -1350 1259
rect -1330 1239 -1310 1259
rect -1290 1239 -1270 1259
rect -1250 1239 -1230 1259
rect -1210 1239 -1190 1259
rect -1170 1239 -1150 1259
rect -1130 1239 -1110 1259
rect -1090 1239 -1070 1259
rect -1050 1239 -1030 1259
rect -1010 1239 -990 1259
rect -970 1239 -950 1259
rect -930 1239 -910 1259
rect -890 1239 -870 1259
rect -850 1239 -830 1259
rect -810 1239 -790 1259
rect -770 1239 -740 1259
rect -710 1239 -685 1259
rect -3665 1225 -3510 1235
rect -3485 1229 -685 1239
rect -3665 1205 -3655 1225
rect -3635 1205 -3615 1225
rect -3595 1205 -3575 1225
rect -3555 1205 -3535 1225
rect -3665 1195 -3510 1205
rect -3485 1191 -685 1201
rect -3485 1171 -3470 1191
rect -3450 1171 -3430 1191
rect -3410 1171 -3390 1191
rect -3370 1171 -3350 1191
rect -3330 1171 -3310 1191
rect -3290 1171 -3270 1191
rect -3250 1171 -3230 1191
rect -3210 1171 -3190 1191
rect -3170 1171 -3150 1191
rect -3130 1171 -3110 1191
rect -3090 1171 -3070 1191
rect -3050 1171 -3030 1191
rect -3010 1171 -2990 1191
rect -2970 1171 -2950 1191
rect -2930 1171 -2910 1191
rect -2890 1171 -2870 1191
rect -2850 1171 -2830 1191
rect -2810 1171 -2790 1191
rect -2770 1171 -2750 1191
rect -2730 1171 -2710 1191
rect -2690 1171 -2670 1191
rect -2650 1171 -2630 1191
rect -2610 1171 -2590 1191
rect -2570 1171 -2550 1191
rect -2530 1171 -2510 1191
rect -2490 1171 -2470 1191
rect -2450 1171 -2430 1191
rect -2410 1171 -2390 1191
rect -2370 1171 -2350 1191
rect -2330 1171 -2310 1191
rect -2290 1171 -2270 1191
rect -2250 1171 -2230 1191
rect -2210 1171 -2190 1191
rect -2170 1171 -2150 1191
rect -2130 1171 -2110 1191
rect -2090 1171 -2070 1191
rect -2050 1171 -2030 1191
rect -2010 1171 -1990 1191
rect -1970 1171 -1950 1191
rect -1930 1171 -1910 1191
rect -1890 1171 -1870 1191
rect -1850 1171 -1830 1191
rect -1810 1171 -1790 1191
rect -1770 1171 -1750 1191
rect -1730 1171 -1710 1191
rect -1690 1171 -1670 1191
rect -1650 1171 -1630 1191
rect -1610 1171 -1590 1191
rect -1570 1171 -1550 1191
rect -1530 1171 -1510 1191
rect -1490 1171 -1470 1191
rect -1450 1171 -1430 1191
rect -1410 1171 -1390 1191
rect -1370 1171 -1350 1191
rect -1330 1171 -1310 1191
rect -1290 1171 -1270 1191
rect -1250 1171 -1230 1191
rect -1210 1171 -1190 1191
rect -1170 1171 -1150 1191
rect -1130 1171 -1110 1191
rect -1090 1171 -1070 1191
rect -1050 1171 -1030 1191
rect -1010 1171 -990 1191
rect -970 1171 -950 1191
rect -930 1171 -910 1191
rect -890 1171 -870 1191
rect -850 1171 -830 1191
rect -810 1171 -790 1191
rect -770 1171 -740 1191
rect -710 1171 -685 1191
rect -3665 1160 -3510 1170
rect -3485 1161 -685 1171
rect -3665 1140 -3655 1160
rect -3635 1140 -3615 1160
rect -3595 1140 -3575 1160
rect -3555 1140 -3535 1160
rect -3665 1130 -3510 1140
rect -3485 1123 -685 1133
rect -3485 1103 -3470 1123
rect -3450 1103 -3430 1123
rect -3410 1103 -3390 1123
rect -3370 1103 -3350 1123
rect -3330 1103 -3310 1123
rect -3290 1103 -3270 1123
rect -3250 1103 -3230 1123
rect -3210 1103 -3190 1123
rect -3170 1103 -3150 1123
rect -3130 1103 -3110 1123
rect -3090 1103 -3070 1123
rect -3050 1103 -3030 1123
rect -3010 1103 -2990 1123
rect -2970 1103 -2950 1123
rect -2930 1103 -2910 1123
rect -2890 1103 -2870 1123
rect -2850 1103 -2830 1123
rect -2810 1103 -2790 1123
rect -2770 1103 -2750 1123
rect -2730 1103 -2710 1123
rect -2690 1103 -2670 1123
rect -2650 1103 -2630 1123
rect -2610 1103 -2590 1123
rect -2570 1103 -2550 1123
rect -2530 1103 -2510 1123
rect -2490 1103 -2470 1123
rect -2450 1103 -2430 1123
rect -2410 1103 -2390 1123
rect -2370 1103 -2350 1123
rect -2330 1103 -2310 1123
rect -2290 1103 -2270 1123
rect -2250 1103 -2230 1123
rect -2210 1103 -2190 1123
rect -2170 1103 -2150 1123
rect -2130 1103 -2110 1123
rect -2090 1103 -2070 1123
rect -2050 1103 -2030 1123
rect -2010 1103 -1990 1123
rect -1970 1103 -1950 1123
rect -1930 1103 -1910 1123
rect -1890 1103 -1870 1123
rect -1850 1103 -1830 1123
rect -1810 1103 -1790 1123
rect -1770 1103 -1750 1123
rect -1730 1103 -1710 1123
rect -1690 1103 -1670 1123
rect -1650 1103 -1630 1123
rect -1610 1103 -1590 1123
rect -1570 1103 -1550 1123
rect -1530 1103 -1510 1123
rect -1490 1103 -1470 1123
rect -1450 1103 -1430 1123
rect -1410 1103 -1390 1123
rect -1370 1103 -1350 1123
rect -1330 1103 -1310 1123
rect -1290 1103 -1270 1123
rect -1250 1103 -1230 1123
rect -1210 1103 -1190 1123
rect -1170 1103 -1150 1123
rect -1130 1103 -1110 1123
rect -1090 1103 -1070 1123
rect -1050 1103 -1030 1123
rect -1010 1103 -990 1123
rect -970 1103 -950 1123
rect -930 1103 -910 1123
rect -890 1103 -870 1123
rect -850 1103 -830 1123
rect -810 1103 -790 1123
rect -770 1103 -740 1123
rect -710 1103 -685 1123
rect -3665 1090 -3510 1100
rect -3485 1093 -685 1103
rect -3665 1070 -3655 1090
rect -3635 1070 -3615 1090
rect -3595 1070 -3575 1090
rect -3555 1070 -3535 1090
rect -3665 1060 -3510 1070
rect -3485 1055 -685 1065
rect -3485 1035 -3470 1055
rect -3450 1035 -3430 1055
rect -3410 1035 -3390 1055
rect -3370 1035 -3350 1055
rect -3330 1035 -3310 1055
rect -3290 1035 -3270 1055
rect -3250 1035 -3230 1055
rect -3210 1035 -3190 1055
rect -3170 1035 -3150 1055
rect -3130 1035 -3110 1055
rect -3090 1035 -3070 1055
rect -3050 1035 -3030 1055
rect -3010 1035 -2990 1055
rect -2970 1035 -2950 1055
rect -2930 1035 -2910 1055
rect -2890 1035 -2870 1055
rect -2850 1035 -2830 1055
rect -2810 1035 -2790 1055
rect -2770 1035 -2750 1055
rect -2730 1035 -2710 1055
rect -2690 1035 -2670 1055
rect -2650 1035 -2630 1055
rect -2610 1035 -2590 1055
rect -2570 1035 -2550 1055
rect -2530 1035 -2510 1055
rect -2490 1035 -2470 1055
rect -2450 1035 -2430 1055
rect -2410 1035 -2390 1055
rect -2370 1035 -2350 1055
rect -2330 1035 -2310 1055
rect -2290 1035 -2270 1055
rect -2250 1035 -2230 1055
rect -2210 1035 -2190 1055
rect -2170 1035 -2150 1055
rect -2130 1035 -2110 1055
rect -2090 1035 -2070 1055
rect -2050 1035 -2030 1055
rect -2010 1035 -1990 1055
rect -1970 1035 -1950 1055
rect -1930 1035 -1910 1055
rect -1890 1035 -1870 1055
rect -1850 1035 -1830 1055
rect -1810 1035 -1790 1055
rect -1770 1035 -1750 1055
rect -1730 1035 -1710 1055
rect -1690 1035 -1670 1055
rect -1650 1035 -1630 1055
rect -1610 1035 -1590 1055
rect -1570 1035 -1550 1055
rect -1530 1035 -1510 1055
rect -1490 1035 -1470 1055
rect -1450 1035 -1430 1055
rect -1410 1035 -1390 1055
rect -1370 1035 -1350 1055
rect -1330 1035 -1310 1055
rect -1290 1035 -1270 1055
rect -1250 1035 -1230 1055
rect -1210 1035 -1190 1055
rect -1170 1035 -1150 1055
rect -1130 1035 -1110 1055
rect -1090 1035 -1070 1055
rect -1050 1035 -1030 1055
rect -1010 1035 -990 1055
rect -970 1035 -950 1055
rect -930 1035 -910 1055
rect -890 1035 -870 1055
rect -850 1035 -830 1055
rect -810 1035 -790 1055
rect -770 1035 -740 1055
rect -710 1035 -685 1055
rect -3665 1020 -3510 1030
rect -3485 1025 -685 1035
rect -3665 1000 -3655 1020
rect -3635 1000 -3615 1020
rect -3595 1000 -3575 1020
rect -3555 1000 -3535 1020
rect -3665 990 -3510 1000
rect -3485 987 -685 997
rect -3485 967 -3470 987
rect -3450 967 -3430 987
rect -3410 967 -3390 987
rect -3370 967 -3350 987
rect -3330 967 -3310 987
rect -3290 967 -3270 987
rect -3250 967 -3230 987
rect -3210 967 -3190 987
rect -3170 967 -3150 987
rect -3130 967 -3110 987
rect -3090 967 -3070 987
rect -3050 967 -3030 987
rect -3010 967 -2990 987
rect -2970 967 -2950 987
rect -2930 967 -2910 987
rect -2890 967 -2870 987
rect -2850 967 -2830 987
rect -2810 967 -2790 987
rect -2770 967 -2750 987
rect -2730 967 -2710 987
rect -2690 967 -2670 987
rect -2650 967 -2630 987
rect -2610 967 -2590 987
rect -2570 967 -2550 987
rect -2530 967 -2510 987
rect -2490 967 -2470 987
rect -2450 967 -2430 987
rect -2410 967 -2390 987
rect -2370 967 -2350 987
rect -2330 967 -2310 987
rect -2290 967 -2270 987
rect -2250 967 -2230 987
rect -2210 967 -2190 987
rect -2170 967 -2150 987
rect -2130 967 -2110 987
rect -2090 967 -2070 987
rect -2050 967 -2030 987
rect -2010 967 -1990 987
rect -1970 967 -1950 987
rect -1930 967 -1910 987
rect -1890 967 -1870 987
rect -1850 967 -1830 987
rect -1810 967 -1790 987
rect -1770 967 -1750 987
rect -1730 967 -1710 987
rect -1690 967 -1670 987
rect -1650 967 -1630 987
rect -1610 967 -1590 987
rect -1570 967 -1550 987
rect -1530 967 -1510 987
rect -1490 967 -1470 987
rect -1450 967 -1430 987
rect -1410 967 -1390 987
rect -1370 967 -1350 987
rect -1330 967 -1310 987
rect -1290 967 -1270 987
rect -1250 967 -1230 987
rect -1210 967 -1190 987
rect -1170 967 -1150 987
rect -1130 967 -1110 987
rect -1090 967 -1070 987
rect -1050 967 -1030 987
rect -1010 967 -990 987
rect -970 967 -950 987
rect -930 967 -910 987
rect -890 967 -870 987
rect -850 967 -830 987
rect -810 967 -790 987
rect -770 967 -740 987
rect -710 967 -685 987
rect -3665 955 -3510 965
rect -3485 957 -685 967
rect -3665 935 -3655 955
rect -3635 935 -3615 955
rect -3595 935 -3575 955
rect -3555 935 -3535 955
rect -3665 925 -3510 935
rect -3485 919 -685 929
rect -3485 899 -3470 919
rect -3450 899 -3430 919
rect -3410 899 -3390 919
rect -3370 899 -3350 919
rect -3330 899 -3310 919
rect -3290 899 -3270 919
rect -3250 899 -3230 919
rect -3210 899 -3190 919
rect -3170 899 -3150 919
rect -3130 899 -3110 919
rect -3090 899 -3070 919
rect -3050 899 -3030 919
rect -3010 899 -2990 919
rect -2970 899 -2950 919
rect -2930 899 -2910 919
rect -2890 899 -2870 919
rect -2850 899 -2830 919
rect -2810 899 -2790 919
rect -2770 899 -2750 919
rect -2730 899 -2710 919
rect -2690 899 -2670 919
rect -2650 899 -2630 919
rect -2610 899 -2590 919
rect -2570 899 -2550 919
rect -2530 899 -2510 919
rect -2490 899 -2470 919
rect -2450 899 -2430 919
rect -2410 899 -2390 919
rect -2370 899 -2350 919
rect -2330 899 -2310 919
rect -2290 899 -2270 919
rect -2250 899 -2230 919
rect -2210 899 -2190 919
rect -2170 899 -2150 919
rect -2130 899 -2110 919
rect -2090 899 -2070 919
rect -2050 899 -2030 919
rect -2010 899 -1990 919
rect -1970 899 -1950 919
rect -1930 899 -1910 919
rect -1890 899 -1870 919
rect -1850 899 -1830 919
rect -1810 899 -1790 919
rect -1770 899 -1750 919
rect -1730 899 -1710 919
rect -1690 899 -1670 919
rect -1650 899 -1630 919
rect -1610 899 -1590 919
rect -1570 899 -1550 919
rect -1530 899 -1510 919
rect -1490 899 -1470 919
rect -1450 899 -1430 919
rect -1410 899 -1390 919
rect -1370 899 -1350 919
rect -1330 899 -1310 919
rect -1290 899 -1270 919
rect -1250 899 -1230 919
rect -1210 899 -1190 919
rect -1170 899 -1150 919
rect -1130 899 -1110 919
rect -1090 899 -1070 919
rect -1050 899 -1030 919
rect -1010 899 -990 919
rect -970 899 -950 919
rect -930 899 -910 919
rect -890 899 -870 919
rect -850 899 -830 919
rect -810 899 -790 919
rect -770 899 -740 919
rect -710 899 -685 919
rect -3665 885 -3510 895
rect -3485 889 -685 899
rect -3665 865 -3655 885
rect -3635 865 -3615 885
rect -3595 865 -3575 885
rect -3555 865 -3535 885
rect -3665 855 -3510 865
rect -3485 851 -685 861
rect -3485 831 -3470 851
rect -3450 831 -3430 851
rect -3410 831 -3390 851
rect -3370 831 -3350 851
rect -3330 831 -3310 851
rect -3290 831 -3270 851
rect -3250 831 -3230 851
rect -3210 831 -3190 851
rect -3170 831 -3150 851
rect -3130 831 -3110 851
rect -3090 831 -3070 851
rect -3050 831 -3030 851
rect -3010 831 -2990 851
rect -2970 831 -2950 851
rect -2930 831 -2910 851
rect -2890 831 -2870 851
rect -2850 831 -2830 851
rect -2810 831 -2790 851
rect -2770 831 -2750 851
rect -2730 831 -2710 851
rect -2690 831 -2670 851
rect -2650 831 -2630 851
rect -2610 831 -2590 851
rect -2570 831 -2550 851
rect -2530 831 -2510 851
rect -2490 831 -2470 851
rect -2450 831 -2430 851
rect -2410 831 -2390 851
rect -2370 831 -2350 851
rect -2330 831 -2310 851
rect -2290 831 -2270 851
rect -2250 831 -2230 851
rect -2210 831 -2190 851
rect -2170 831 -2150 851
rect -2130 831 -2110 851
rect -2090 831 -2070 851
rect -2050 831 -2030 851
rect -2010 831 -1990 851
rect -1970 831 -1950 851
rect -1930 831 -1910 851
rect -1890 831 -1870 851
rect -1850 831 -1830 851
rect -1810 831 -1790 851
rect -1770 831 -1750 851
rect -1730 831 -1710 851
rect -1690 831 -1670 851
rect -1650 831 -1630 851
rect -1610 831 -1590 851
rect -1570 831 -1550 851
rect -1530 831 -1510 851
rect -1490 831 -1470 851
rect -1450 831 -1430 851
rect -1410 831 -1390 851
rect -1370 831 -1350 851
rect -1330 831 -1310 851
rect -1290 831 -1270 851
rect -1250 831 -1230 851
rect -1210 831 -1190 851
rect -1170 831 -1150 851
rect -1130 831 -1110 851
rect -1090 831 -1070 851
rect -1050 831 -1030 851
rect -1010 831 -990 851
rect -970 831 -950 851
rect -930 831 -910 851
rect -890 831 -870 851
rect -850 831 -830 851
rect -810 831 -790 851
rect -770 831 -740 851
rect -710 831 -685 851
rect -3665 815 -3510 825
rect -3485 821 -685 831
rect -3665 795 -3655 815
rect -3635 795 -3615 815
rect -3595 795 -3575 815
rect -3555 795 -3535 815
rect -3665 785 -3510 795
rect -3485 783 -685 793
rect -3485 763 -3470 783
rect -3450 763 -3430 783
rect -3410 763 -3390 783
rect -3370 763 -3350 783
rect -3330 763 -3310 783
rect -3290 763 -3270 783
rect -3250 763 -3230 783
rect -3210 763 -3190 783
rect -3170 763 -3150 783
rect -3130 763 -3110 783
rect -3090 763 -3070 783
rect -3050 763 -3030 783
rect -3010 763 -2990 783
rect -2970 763 -2950 783
rect -2930 763 -2910 783
rect -2890 763 -2870 783
rect -2850 763 -2830 783
rect -2810 763 -2790 783
rect -2770 763 -2750 783
rect -2730 763 -2710 783
rect -2690 763 -2670 783
rect -2650 763 -2630 783
rect -2610 763 -2590 783
rect -2570 763 -2550 783
rect -2530 763 -2510 783
rect -2490 763 -2470 783
rect -2450 763 -2430 783
rect -2410 763 -2390 783
rect -2370 763 -2350 783
rect -2330 763 -2310 783
rect -2290 763 -2270 783
rect -2250 763 -2230 783
rect -2210 763 -2190 783
rect -2170 763 -2150 783
rect -2130 763 -2110 783
rect -2090 763 -2070 783
rect -2050 763 -2030 783
rect -2010 763 -1990 783
rect -1970 763 -1950 783
rect -1930 763 -1910 783
rect -1890 763 -1870 783
rect -1850 763 -1830 783
rect -1810 763 -1790 783
rect -1770 763 -1750 783
rect -1730 763 -1710 783
rect -1690 763 -1670 783
rect -1650 763 -1630 783
rect -1610 763 -1590 783
rect -1570 763 -1550 783
rect -1530 763 -1510 783
rect -1490 763 -1470 783
rect -1450 763 -1430 783
rect -1410 763 -1390 783
rect -1370 763 -1350 783
rect -1330 763 -1310 783
rect -1290 763 -1270 783
rect -1250 763 -1230 783
rect -1210 763 -1190 783
rect -1170 763 -1150 783
rect -1130 763 -1110 783
rect -1090 763 -1070 783
rect -1050 763 -1030 783
rect -1010 763 -990 783
rect -970 763 -950 783
rect -930 763 -910 783
rect -890 763 -870 783
rect -850 763 -830 783
rect -810 763 -790 783
rect -770 763 -740 783
rect -710 763 -685 783
rect -3665 750 -3510 760
rect -3485 753 -685 763
rect -3665 730 -3655 750
rect -3635 730 -3615 750
rect -3595 730 -3575 750
rect -3555 730 -3535 750
rect -3665 720 -3510 730
rect -3485 715 -685 725
rect -3485 695 -3470 715
rect -3450 695 -3430 715
rect -3410 695 -3390 715
rect -3370 695 -3350 715
rect -3330 695 -3310 715
rect -3290 695 -3270 715
rect -3250 695 -3230 715
rect -3210 695 -3190 715
rect -3170 695 -3150 715
rect -3130 695 -3110 715
rect -3090 695 -3070 715
rect -3050 695 -3030 715
rect -3010 695 -2990 715
rect -2970 695 -2950 715
rect -2930 695 -2910 715
rect -2890 695 -2870 715
rect -2850 695 -2830 715
rect -2810 695 -2790 715
rect -2770 695 -2750 715
rect -2730 695 -2710 715
rect -2690 695 -2670 715
rect -2650 695 -2630 715
rect -2610 695 -2590 715
rect -2570 695 -2550 715
rect -2530 695 -2510 715
rect -2490 695 -2470 715
rect -2450 695 -2430 715
rect -2410 695 -2390 715
rect -2370 695 -2350 715
rect -2330 695 -2310 715
rect -2290 695 -2270 715
rect -2250 695 -2230 715
rect -2210 695 -2190 715
rect -2170 695 -2150 715
rect -2130 695 -2110 715
rect -2090 695 -2070 715
rect -2050 695 -2030 715
rect -2010 695 -1990 715
rect -1970 695 -1950 715
rect -1930 695 -1910 715
rect -1890 695 -1870 715
rect -1850 695 -1830 715
rect -1810 695 -1790 715
rect -1770 695 -1750 715
rect -1730 695 -1710 715
rect -1690 695 -1670 715
rect -1650 695 -1630 715
rect -1610 695 -1590 715
rect -1570 695 -1550 715
rect -1530 695 -1510 715
rect -1490 695 -1470 715
rect -1450 695 -1430 715
rect -1410 695 -1390 715
rect -1370 695 -1350 715
rect -1330 695 -1310 715
rect -1290 695 -1270 715
rect -1250 695 -1230 715
rect -1210 695 -1190 715
rect -1170 695 -1150 715
rect -1130 695 -1110 715
rect -1090 695 -1070 715
rect -1050 695 -1030 715
rect -1010 695 -990 715
rect -970 695 -950 715
rect -930 695 -910 715
rect -890 695 -870 715
rect -850 695 -830 715
rect -810 695 -790 715
rect -770 695 -740 715
rect -710 695 -685 715
rect -3665 680 -3510 690
rect -3485 685 -685 695
rect -3665 660 -3655 680
rect -3635 660 -3615 680
rect -3595 660 -3575 680
rect -3555 660 -3535 680
rect -3665 650 -3510 660
rect -3485 647 -685 657
rect -3485 627 -3470 647
rect -3450 627 -3430 647
rect -3410 627 -3390 647
rect -3370 627 -3350 647
rect -3330 627 -3310 647
rect -3290 627 -3270 647
rect -3250 627 -3230 647
rect -3210 627 -3190 647
rect -3170 627 -3150 647
rect -3130 627 -3110 647
rect -3090 627 -3070 647
rect -3050 627 -3030 647
rect -3010 627 -2990 647
rect -2970 627 -2950 647
rect -2930 627 -2910 647
rect -2890 627 -2870 647
rect -2850 627 -2830 647
rect -2810 627 -2790 647
rect -2770 627 -2750 647
rect -2730 627 -2710 647
rect -2690 627 -2670 647
rect -2650 627 -2630 647
rect -2610 627 -2590 647
rect -2570 627 -2550 647
rect -2530 627 -2510 647
rect -2490 627 -2470 647
rect -2450 627 -2430 647
rect -2410 627 -2390 647
rect -2370 627 -2350 647
rect -2330 627 -2310 647
rect -2290 627 -2270 647
rect -2250 627 -2230 647
rect -2210 627 -2190 647
rect -2170 627 -2150 647
rect -2130 627 -2110 647
rect -2090 627 -2070 647
rect -2050 627 -2030 647
rect -2010 627 -1990 647
rect -1970 627 -1950 647
rect -1930 627 -1910 647
rect -1890 627 -1870 647
rect -1850 627 -1830 647
rect -1810 627 -1790 647
rect -1770 627 -1750 647
rect -1730 627 -1710 647
rect -1690 627 -1670 647
rect -1650 627 -1630 647
rect -1610 627 -1590 647
rect -1570 627 -1550 647
rect -1530 627 -1510 647
rect -1490 627 -1470 647
rect -1450 627 -1430 647
rect -1410 627 -1390 647
rect -1370 627 -1350 647
rect -1330 627 -1310 647
rect -1290 627 -1270 647
rect -1250 627 -1230 647
rect -1210 627 -1190 647
rect -1170 627 -1150 647
rect -1130 627 -1110 647
rect -1090 627 -1070 647
rect -1050 627 -1030 647
rect -1010 627 -990 647
rect -970 627 -950 647
rect -930 627 -910 647
rect -890 627 -870 647
rect -850 627 -830 647
rect -810 627 -790 647
rect -770 627 -740 647
rect -710 627 -685 647
rect -3665 615 -3510 625
rect -3485 617 -685 627
rect -3665 595 -3655 615
rect -3635 595 -3615 615
rect -3595 595 -3575 615
rect -3555 595 -3535 615
rect -3665 585 -3510 595
rect -3485 579 -685 589
rect -3485 559 -3470 579
rect -3450 559 -3430 579
rect -3410 559 -3390 579
rect -3370 559 -3350 579
rect -3330 559 -3310 579
rect -3290 559 -3270 579
rect -3250 559 -3230 579
rect -3210 559 -3190 579
rect -3170 559 -3150 579
rect -3130 559 -3110 579
rect -3090 559 -3070 579
rect -3050 559 -3030 579
rect -3010 559 -2990 579
rect -2970 559 -2950 579
rect -2930 559 -2910 579
rect -2890 559 -2870 579
rect -2850 559 -2830 579
rect -2810 559 -2790 579
rect -2770 559 -2750 579
rect -2730 559 -2710 579
rect -2690 559 -2670 579
rect -2650 559 -2630 579
rect -2610 559 -2590 579
rect -2570 559 -2550 579
rect -2530 559 -2510 579
rect -2490 559 -2470 579
rect -2450 559 -2430 579
rect -2410 559 -2390 579
rect -2370 559 -2350 579
rect -2330 559 -2310 579
rect -2290 559 -2270 579
rect -2250 559 -2230 579
rect -2210 559 -2190 579
rect -2170 559 -2150 579
rect -2130 559 -2110 579
rect -2090 559 -2070 579
rect -2050 559 -2030 579
rect -2010 559 -1990 579
rect -1970 559 -1950 579
rect -1930 559 -1910 579
rect -1890 559 -1870 579
rect -1850 559 -1830 579
rect -1810 559 -1790 579
rect -1770 559 -1750 579
rect -1730 559 -1710 579
rect -1690 559 -1670 579
rect -1650 559 -1630 579
rect -1610 559 -1590 579
rect -1570 559 -1550 579
rect -1530 559 -1510 579
rect -1490 559 -1470 579
rect -1450 559 -1430 579
rect -1410 559 -1390 579
rect -1370 559 -1350 579
rect -1330 559 -1310 579
rect -1290 559 -1270 579
rect -1250 559 -1230 579
rect -1210 559 -1190 579
rect -1170 559 -1150 579
rect -1130 559 -1110 579
rect -1090 559 -1070 579
rect -1050 559 -1030 579
rect -1010 559 -990 579
rect -970 559 -950 579
rect -930 559 -910 579
rect -890 559 -870 579
rect -850 559 -830 579
rect -810 559 -790 579
rect -770 559 -740 579
rect -710 559 -685 579
rect -3665 545 -3510 555
rect -3485 549 -685 559
rect -3665 525 -3655 545
rect -3635 525 -3615 545
rect -3595 525 -3575 545
rect -3555 525 -3535 545
rect -3665 515 -3510 525
rect -3485 511 -685 521
rect -3485 491 -3470 511
rect -3450 491 -3430 511
rect -3410 491 -3390 511
rect -3370 491 -3350 511
rect -3330 491 -3310 511
rect -3290 491 -3270 511
rect -3250 491 -3230 511
rect -3210 491 -3190 511
rect -3170 491 -3150 511
rect -3130 491 -3110 511
rect -3090 491 -3070 511
rect -3050 491 -3030 511
rect -3010 491 -2990 511
rect -2970 491 -2950 511
rect -2930 491 -2910 511
rect -2890 491 -2870 511
rect -2850 491 -2830 511
rect -2810 491 -2790 511
rect -2770 491 -2750 511
rect -2730 491 -2710 511
rect -2690 491 -2670 511
rect -2650 491 -2630 511
rect -2610 491 -2590 511
rect -2570 491 -2550 511
rect -2530 491 -2510 511
rect -2490 491 -2470 511
rect -2450 491 -2430 511
rect -2410 491 -2390 511
rect -2370 491 -2350 511
rect -2330 491 -2310 511
rect -2290 491 -2270 511
rect -2250 491 -2230 511
rect -2210 491 -2190 511
rect -2170 491 -2150 511
rect -2130 491 -2110 511
rect -2090 491 -2070 511
rect -2050 491 -2030 511
rect -2010 491 -1990 511
rect -1970 491 -1950 511
rect -1930 491 -1910 511
rect -1890 491 -1870 511
rect -1850 491 -1830 511
rect -1810 491 -1790 511
rect -1770 491 -1750 511
rect -1730 491 -1710 511
rect -1690 491 -1670 511
rect -1650 491 -1630 511
rect -1610 491 -1590 511
rect -1570 491 -1550 511
rect -1530 491 -1510 511
rect -1490 491 -1470 511
rect -1450 491 -1430 511
rect -1410 491 -1390 511
rect -1370 491 -1350 511
rect -1330 491 -1310 511
rect -1290 491 -1270 511
rect -1250 491 -1230 511
rect -1210 491 -1190 511
rect -1170 491 -1150 511
rect -1130 491 -1110 511
rect -1090 491 -1070 511
rect -1050 491 -1030 511
rect -1010 491 -990 511
rect -970 491 -950 511
rect -930 491 -910 511
rect -890 491 -870 511
rect -850 491 -830 511
rect -810 491 -790 511
rect -770 491 -740 511
rect -710 491 -685 511
rect -3665 475 -3510 485
rect -3485 481 -685 491
rect -3665 455 -3655 475
rect -3635 455 -3615 475
rect -3595 455 -3575 475
rect -3555 455 -3535 475
rect -3665 445 -3510 455
rect -3485 443 -685 453
rect -3485 423 -3470 443
rect -3450 423 -3430 443
rect -3410 423 -3390 443
rect -3370 423 -3350 443
rect -3330 423 -3310 443
rect -3290 423 -3270 443
rect -3250 423 -3230 443
rect -3210 423 -3190 443
rect -3170 423 -3150 443
rect -3130 423 -3110 443
rect -3090 423 -3070 443
rect -3050 423 -3030 443
rect -3010 423 -2990 443
rect -2970 423 -2950 443
rect -2930 423 -2910 443
rect -2890 423 -2870 443
rect -2850 423 -2830 443
rect -2810 423 -2790 443
rect -2770 423 -2750 443
rect -2730 423 -2710 443
rect -2690 423 -2670 443
rect -2650 423 -2630 443
rect -2610 423 -2590 443
rect -2570 423 -2550 443
rect -2530 423 -2510 443
rect -2490 423 -2470 443
rect -2450 423 -2430 443
rect -2410 423 -2390 443
rect -2370 423 -2350 443
rect -2330 423 -2310 443
rect -2290 423 -2270 443
rect -2250 423 -2230 443
rect -2210 423 -2190 443
rect -2170 423 -2150 443
rect -2130 423 -2110 443
rect -2090 423 -2070 443
rect -2050 423 -2030 443
rect -2010 423 -1990 443
rect -1970 423 -1950 443
rect -1930 423 -1910 443
rect -1890 423 -1870 443
rect -1850 423 -1830 443
rect -1810 423 -1790 443
rect -1770 423 -1750 443
rect -1730 423 -1710 443
rect -1690 423 -1670 443
rect -1650 423 -1630 443
rect -1610 423 -1590 443
rect -1570 423 -1550 443
rect -1530 423 -1510 443
rect -1490 423 -1470 443
rect -1450 423 -1430 443
rect -1410 423 -1390 443
rect -1370 423 -1350 443
rect -1330 423 -1310 443
rect -1290 423 -1270 443
rect -1250 423 -1230 443
rect -1210 423 -1190 443
rect -1170 423 -1150 443
rect -1130 423 -1110 443
rect -1090 423 -1070 443
rect -1050 423 -1030 443
rect -1010 423 -990 443
rect -970 423 -950 443
rect -930 423 -910 443
rect -890 423 -870 443
rect -850 423 -830 443
rect -810 423 -790 443
rect -770 423 -740 443
rect -710 423 -685 443
rect -3665 405 -3510 415
rect -3485 413 -685 423
rect -3665 385 -3655 405
rect -3635 385 -3615 405
rect -3595 385 -3575 405
rect -3555 385 -3535 405
rect -3665 375 -3510 385
rect -3485 375 -685 385
rect -3485 355 -3470 375
rect -3450 355 -3430 375
rect -3410 355 -3390 375
rect -3370 355 -3350 375
rect -3330 355 -3310 375
rect -3290 355 -3270 375
rect -3250 355 -3230 375
rect -3210 355 -3190 375
rect -3170 355 -3150 375
rect -3130 355 -3110 375
rect -3090 355 -3070 375
rect -3050 355 -3030 375
rect -3010 355 -2990 375
rect -2970 355 -2950 375
rect -2930 355 -2910 375
rect -2890 355 -2870 375
rect -2850 355 -2830 375
rect -2810 355 -2790 375
rect -2770 355 -2750 375
rect -2730 355 -2710 375
rect -2690 355 -2670 375
rect -2650 355 -2630 375
rect -2610 355 -2590 375
rect -2570 355 -2550 375
rect -2530 355 -2510 375
rect -2490 355 -2470 375
rect -2450 355 -2430 375
rect -2410 355 -2390 375
rect -2370 355 -2350 375
rect -2330 355 -2310 375
rect -2290 355 -2270 375
rect -2250 355 -2230 375
rect -2210 355 -2190 375
rect -2170 355 -2150 375
rect -2130 355 -2110 375
rect -2090 355 -2070 375
rect -2050 355 -2030 375
rect -2010 355 -1990 375
rect -1970 355 -1950 375
rect -1930 355 -1910 375
rect -1890 355 -1870 375
rect -1850 355 -1830 375
rect -1810 355 -1790 375
rect -1770 355 -1750 375
rect -1730 355 -1710 375
rect -1690 355 -1670 375
rect -1650 355 -1630 375
rect -1610 355 -1590 375
rect -1570 355 -1550 375
rect -1530 355 -1510 375
rect -1490 355 -1470 375
rect -1450 355 -1430 375
rect -1410 355 -1390 375
rect -1370 355 -1350 375
rect -1330 355 -1310 375
rect -1290 355 -1270 375
rect -1250 355 -1230 375
rect -1210 355 -1190 375
rect -1170 355 -1150 375
rect -1130 355 -1110 375
rect -1090 355 -1070 375
rect -1050 355 -1030 375
rect -1010 355 -990 375
rect -970 355 -950 375
rect -930 355 -910 375
rect -890 355 -870 375
rect -850 355 -830 375
rect -810 355 -790 375
rect -770 355 -740 375
rect -710 355 -685 375
rect -3665 340 -3510 350
rect -3485 345 -685 355
rect -3665 320 -3655 340
rect -3635 320 -3615 340
rect -3595 320 -3575 340
rect -3555 320 -3535 340
rect -3665 310 -3510 320
rect -3485 307 -685 317
rect -3485 287 -3470 307
rect -3450 287 -3430 307
rect -3410 287 -3390 307
rect -3370 287 -3350 307
rect -3330 287 -3310 307
rect -3290 287 -3270 307
rect -3250 287 -3230 307
rect -3210 287 -3190 307
rect -3170 287 -3150 307
rect -3130 287 -3110 307
rect -3090 287 -3070 307
rect -3050 287 -3030 307
rect -3010 287 -2990 307
rect -2970 287 -2950 307
rect -2930 287 -2910 307
rect -2890 287 -2870 307
rect -2850 287 -2830 307
rect -2810 287 -2790 307
rect -2770 287 -2750 307
rect -2730 287 -2710 307
rect -2690 287 -2670 307
rect -2650 287 -2630 307
rect -2610 287 -2590 307
rect -2570 287 -2550 307
rect -2530 287 -2510 307
rect -2490 287 -2470 307
rect -2450 287 -2430 307
rect -2410 287 -2390 307
rect -2370 287 -2350 307
rect -2330 287 -2310 307
rect -2290 287 -2270 307
rect -2250 287 -2230 307
rect -2210 287 -2190 307
rect -2170 287 -2150 307
rect -2130 287 -2110 307
rect -2090 287 -2070 307
rect -2050 287 -2030 307
rect -2010 287 -1990 307
rect -1970 287 -1950 307
rect -1930 287 -1910 307
rect -1890 287 -1870 307
rect -1850 287 -1830 307
rect -1810 287 -1790 307
rect -1770 287 -1750 307
rect -1730 287 -1710 307
rect -1690 287 -1670 307
rect -1650 287 -1630 307
rect -1610 287 -1590 307
rect -1570 287 -1550 307
rect -1530 287 -1510 307
rect -1490 287 -1470 307
rect -1450 287 -1430 307
rect -1410 287 -1390 307
rect -1370 287 -1350 307
rect -1330 287 -1310 307
rect -1290 287 -1270 307
rect -1250 287 -1230 307
rect -1210 287 -1190 307
rect -1170 287 -1150 307
rect -1130 287 -1110 307
rect -1090 287 -1070 307
rect -1050 287 -1030 307
rect -1010 287 -990 307
rect -970 287 -950 307
rect -930 287 -910 307
rect -890 287 -870 307
rect -850 287 -830 307
rect -810 287 -790 307
rect -770 287 -740 307
rect -710 287 -685 307
rect -3665 275 -3510 285
rect -3485 277 -685 287
rect -3665 255 -3655 275
rect -3635 255 -3615 275
rect -3595 255 -3575 275
rect -3555 255 -3535 275
rect -3665 245 -3510 255
rect -3485 239 -685 249
rect -3485 219 -3470 239
rect -3450 219 -3430 239
rect -3410 219 -3390 239
rect -3370 219 -3350 239
rect -3330 219 -3310 239
rect -3290 219 -3270 239
rect -3250 219 -3230 239
rect -3210 219 -3190 239
rect -3170 219 -3150 239
rect -3130 219 -3110 239
rect -3090 219 -3070 239
rect -3050 219 -3030 239
rect -3010 219 -2990 239
rect -2970 219 -2950 239
rect -2930 219 -2910 239
rect -2890 219 -2870 239
rect -2850 219 -2830 239
rect -2810 219 -2790 239
rect -2770 219 -2750 239
rect -2730 219 -2710 239
rect -2690 219 -2670 239
rect -2650 219 -2630 239
rect -2610 219 -2590 239
rect -2570 219 -2550 239
rect -2530 219 -2510 239
rect -2490 219 -2470 239
rect -2450 219 -2430 239
rect -2410 219 -2390 239
rect -2370 219 -2350 239
rect -2330 219 -2310 239
rect -2290 219 -2270 239
rect -2250 219 -2230 239
rect -2210 219 -2190 239
rect -2170 219 -2150 239
rect -2130 219 -2110 239
rect -2090 219 -2070 239
rect -2050 219 -2030 239
rect -2010 219 -1990 239
rect -1970 219 -1950 239
rect -1930 219 -1910 239
rect -1890 219 -1870 239
rect -1850 219 -1830 239
rect -1810 219 -1790 239
rect -1770 219 -1750 239
rect -1730 219 -1710 239
rect -1690 219 -1670 239
rect -1650 219 -1630 239
rect -1610 219 -1590 239
rect -1570 219 -1550 239
rect -1530 219 -1510 239
rect -1490 219 -1470 239
rect -1450 219 -1430 239
rect -1410 219 -1390 239
rect -1370 219 -1350 239
rect -1330 219 -1310 239
rect -1290 219 -1270 239
rect -1250 219 -1230 239
rect -1210 219 -1190 239
rect -1170 219 -1150 239
rect -1130 219 -1110 239
rect -1090 219 -1070 239
rect -1050 219 -1030 239
rect -1010 219 -990 239
rect -970 219 -950 239
rect -930 219 -910 239
rect -890 219 -870 239
rect -850 219 -830 239
rect -810 219 -790 239
rect -770 219 -740 239
rect -710 219 -685 239
rect -3665 205 -3510 215
rect -3485 209 -685 219
rect -3665 185 -3655 205
rect -3635 185 -3615 205
rect -3595 185 -3575 205
rect -3555 185 -3535 205
rect -3665 175 -3510 185
rect -3485 171 -685 181
rect -3485 151 -3470 171
rect -3450 151 -3430 171
rect -3410 151 -3390 171
rect -3370 151 -3350 171
rect -3330 151 -3310 171
rect -3290 151 -3270 171
rect -3250 151 -3230 171
rect -3210 151 -3190 171
rect -3170 151 -3150 171
rect -3130 151 -3110 171
rect -3090 151 -3070 171
rect -3050 151 -3030 171
rect -3010 151 -2990 171
rect -2970 151 -2950 171
rect -2930 151 -2910 171
rect -2890 151 -2870 171
rect -2850 151 -2830 171
rect -2810 151 -2790 171
rect -2770 151 -2750 171
rect -2730 151 -2710 171
rect -2690 151 -2670 171
rect -2650 151 -2630 171
rect -2610 151 -2590 171
rect -2570 151 -2550 171
rect -2530 151 -2510 171
rect -2490 151 -2470 171
rect -2450 151 -2430 171
rect -2410 151 -2390 171
rect -2370 151 -2350 171
rect -2330 151 -2310 171
rect -2290 151 -2270 171
rect -2250 151 -2230 171
rect -2210 151 -2190 171
rect -2170 151 -2150 171
rect -2130 151 -2110 171
rect -2090 151 -2070 171
rect -2050 151 -2030 171
rect -2010 151 -1990 171
rect -1970 151 -1950 171
rect -1930 151 -1910 171
rect -1890 151 -1870 171
rect -1850 151 -1830 171
rect -1810 151 -1790 171
rect -1770 151 -1750 171
rect -1730 151 -1710 171
rect -1690 151 -1670 171
rect -1650 151 -1630 171
rect -1610 151 -1590 171
rect -1570 151 -1550 171
rect -1530 151 -1510 171
rect -1490 151 -1470 171
rect -1450 151 -1430 171
rect -1410 151 -1390 171
rect -1370 151 -1350 171
rect -1330 151 -1310 171
rect -1290 151 -1270 171
rect -1250 151 -1230 171
rect -1210 151 -1190 171
rect -1170 151 -1150 171
rect -1130 151 -1110 171
rect -1090 151 -1070 171
rect -1050 151 -1030 171
rect -1010 151 -990 171
rect -970 151 -950 171
rect -930 151 -910 171
rect -890 151 -870 171
rect -850 151 -830 171
rect -810 151 -790 171
rect -770 151 -740 171
rect -710 151 -685 171
rect -3665 135 -3510 145
rect -3485 141 -685 151
rect -3665 115 -3655 135
rect -3635 115 -3615 135
rect -3595 115 -3575 135
rect -3555 115 -3535 135
rect -3665 105 -3510 115
rect -3485 103 -685 113
rect -3485 83 -3470 103
rect -3450 83 -3430 103
rect -3410 83 -3390 103
rect -3370 83 -3350 103
rect -3330 83 -3310 103
rect -3290 83 -3270 103
rect -3250 83 -3230 103
rect -3210 83 -3190 103
rect -3170 83 -3150 103
rect -3130 83 -3110 103
rect -3090 83 -3070 103
rect -3050 83 -3030 103
rect -3010 83 -2990 103
rect -2970 83 -2950 103
rect -2930 83 -2910 103
rect -2890 83 -2870 103
rect -2850 83 -2830 103
rect -2810 83 -2790 103
rect -2770 83 -2750 103
rect -2730 83 -2710 103
rect -2690 83 -2670 103
rect -2650 83 -2630 103
rect -2610 83 -2590 103
rect -2570 83 -2550 103
rect -2530 83 -2510 103
rect -2490 83 -2470 103
rect -2450 83 -2430 103
rect -2410 83 -2390 103
rect -2370 83 -2350 103
rect -2330 83 -2310 103
rect -2290 83 -2270 103
rect -2250 83 -2230 103
rect -2210 83 -2190 103
rect -2170 83 -2150 103
rect -2130 83 -2110 103
rect -2090 83 -2070 103
rect -2050 83 -2030 103
rect -2010 83 -1990 103
rect -1970 83 -1950 103
rect -1930 83 -1910 103
rect -1890 83 -1870 103
rect -1850 83 -1830 103
rect -1810 83 -1790 103
rect -1770 83 -1750 103
rect -1730 83 -1710 103
rect -1690 83 -1670 103
rect -1650 83 -1630 103
rect -1610 83 -1590 103
rect -1570 83 -1550 103
rect -1530 83 -1510 103
rect -1490 83 -1470 103
rect -1450 83 -1430 103
rect -1410 83 -1390 103
rect -1370 83 -1350 103
rect -1330 83 -1310 103
rect -1290 83 -1270 103
rect -1250 83 -1230 103
rect -1210 83 -1190 103
rect -1170 83 -1150 103
rect -1130 83 -1110 103
rect -1090 83 -1070 103
rect -1050 83 -1030 103
rect -1010 83 -990 103
rect -970 83 -950 103
rect -930 83 -910 103
rect -890 83 -870 103
rect -850 83 -830 103
rect -810 83 -790 103
rect -770 83 -740 103
rect -710 83 -685 103
rect -3665 70 -3510 80
rect -3485 73 -685 83
rect -3665 50 -3655 70
rect -3635 50 -3615 70
rect -3595 50 -3575 70
rect -3555 50 -3535 70
rect -3665 40 -3510 50
rect -3485 35 -685 45
rect -3485 15 -3470 35
rect -3450 15 -3430 35
rect -3410 15 -3390 35
rect -3370 15 -3350 35
rect -3330 15 -3310 35
rect -3290 15 -3270 35
rect -3250 15 -3230 35
rect -3210 15 -3190 35
rect -3170 15 -3150 35
rect -3130 15 -3110 35
rect -3090 15 -3070 35
rect -3050 15 -3030 35
rect -3010 15 -2990 35
rect -2970 15 -2950 35
rect -2930 15 -2910 35
rect -2890 15 -2870 35
rect -2850 15 -2830 35
rect -2810 15 -2790 35
rect -2770 15 -2750 35
rect -2730 15 -2710 35
rect -2690 15 -2670 35
rect -2650 15 -2630 35
rect -2610 15 -2590 35
rect -2570 15 -2550 35
rect -2530 15 -2510 35
rect -2490 15 -2470 35
rect -2450 15 -2430 35
rect -2410 15 -2390 35
rect -2370 15 -2350 35
rect -2330 15 -2310 35
rect -2290 15 -2270 35
rect -2250 15 -2230 35
rect -2210 15 -2190 35
rect -2170 15 -2150 35
rect -2130 15 -2110 35
rect -2090 15 -2070 35
rect -2050 15 -2030 35
rect -2010 15 -1990 35
rect -1970 15 -1950 35
rect -1930 15 -1910 35
rect -1890 15 -1870 35
rect -1850 15 -1830 35
rect -1810 15 -1790 35
rect -1770 15 -1750 35
rect -1730 15 -1710 35
rect -1690 15 -1670 35
rect -1650 15 -1630 35
rect -1610 15 -1590 35
rect -1570 15 -1550 35
rect -1530 15 -1510 35
rect -1490 15 -1470 35
rect -1450 15 -1430 35
rect -1410 15 -1390 35
rect -1370 15 -1350 35
rect -1330 15 -1310 35
rect -1290 15 -1270 35
rect -1250 15 -1230 35
rect -1210 15 -1190 35
rect -1170 15 -1150 35
rect -1130 15 -1110 35
rect -1090 15 -1070 35
rect -1050 15 -1030 35
rect -1010 15 -990 35
rect -970 15 -950 35
rect -930 15 -910 35
rect -890 15 -870 35
rect -850 15 -830 35
rect -810 15 -790 35
rect -770 15 -740 35
rect -710 15 -685 35
rect -3485 -5 -685 15
rect -3485 -25 -3470 -5
rect -3450 -25 -3430 -5
rect -3410 -25 -3390 -5
rect -3370 -25 -3350 -5
rect -3330 -25 -3310 -5
rect -3290 -25 -3270 -5
rect -3250 -25 -3230 -5
rect -3210 -25 -3190 -5
rect -3170 -25 -3150 -5
rect -3130 -25 -3110 -5
rect -3090 -25 -3070 -5
rect -3050 -25 -3030 -5
rect -3010 -25 -2990 -5
rect -2970 -25 -2950 -5
rect -2930 -25 -2910 -5
rect -2890 -25 -2870 -5
rect -2850 -25 -2830 -5
rect -2810 -25 -2790 -5
rect -2770 -25 -2750 -5
rect -2730 -25 -2710 -5
rect -2690 -25 -2670 -5
rect -2650 -25 -2630 -5
rect -2610 -25 -2590 -5
rect -2570 -25 -2550 -5
rect -2530 -25 -2510 -5
rect -2490 -25 -2470 -5
rect -2450 -25 -2430 -5
rect -2410 -25 -2390 -5
rect -2370 -25 -2350 -5
rect -2330 -25 -2310 -5
rect -2290 -25 -2270 -5
rect -2250 -25 -2230 -5
rect -2210 -25 -2190 -5
rect -2170 -25 -2150 -5
rect -2130 -25 -2110 -5
rect -2090 -25 -2070 -5
rect -2050 -25 -2030 -5
rect -2010 -25 -1990 -5
rect -1970 -25 -1950 -5
rect -1930 -25 -1910 -5
rect -1890 -25 -1870 -5
rect -1850 -25 -1830 -5
rect -1810 -25 -1790 -5
rect -1770 -25 -1750 -5
rect -1730 -25 -1710 -5
rect -1690 -25 -1670 -5
rect -1650 -25 -1630 -5
rect -1610 -25 -1590 -5
rect -1570 -25 -1550 -5
rect -1530 -25 -1510 -5
rect -1490 -25 -1470 -5
rect -1450 -25 -1430 -5
rect -1410 -25 -1390 -5
rect -1370 -25 -1350 -5
rect -1330 -25 -1310 -5
rect -1290 -25 -1270 -5
rect -1250 -25 -1230 -5
rect -1210 -25 -1190 -5
rect -1170 -25 -1150 -5
rect -1130 -25 -1110 -5
rect -1090 -25 -1070 -5
rect -1050 -25 -1030 -5
rect -1010 -25 -990 -5
rect -970 -25 -950 -5
rect -930 -25 -910 -5
rect -890 -25 -870 -5
rect -850 -25 -830 -5
rect -810 -25 -790 -5
rect -770 -25 -740 -5
rect -710 -25 -685 -5
rect -3485 -35 -685 -25
rect -3485 -80 -985 -70
rect -3485 -100 -3470 -80
rect -3450 -100 -3430 -80
rect -3410 -100 -3390 -80
rect -3370 -100 -3350 -80
rect -3330 -100 -3310 -80
rect -3290 -100 -3270 -80
rect -3250 -100 -3230 -80
rect -3210 -100 -3190 -80
rect -3170 -100 -3150 -80
rect -3130 -100 -3110 -80
rect -3090 -100 -3070 -80
rect -3050 -100 -3030 -80
rect -3010 -100 -2990 -80
rect -2970 -100 -2950 -80
rect -2930 -100 -2910 -80
rect -2890 -100 -2870 -80
rect -2850 -100 -2830 -80
rect -2810 -100 -2790 -80
rect -2770 -100 -2750 -80
rect -2730 -100 -2710 -80
rect -2690 -100 -2670 -80
rect -2650 -100 -2630 -80
rect -2610 -100 -2590 -80
rect -2570 -100 -2550 -80
rect -2530 -100 -2510 -80
rect -2490 -100 -2470 -80
rect -2450 -100 -2430 -80
rect -2410 -100 -2390 -80
rect -2370 -100 -2350 -80
rect -2330 -100 -2310 -80
rect -2290 -100 -2270 -80
rect -2250 -100 -2230 -80
rect -2210 -100 -2190 -80
rect -2170 -100 -2150 -80
rect -2130 -100 -2110 -80
rect -2090 -100 -2070 -80
rect -2050 -100 -2030 -80
rect -2010 -100 -1990 -80
rect -1970 -100 -1950 -80
rect -1930 -100 -1910 -80
rect -1890 -100 -1870 -80
rect -1850 -100 -1830 -80
rect -1810 -100 -1790 -80
rect -1770 -100 -1750 -80
rect -1730 -100 -1710 -80
rect -1690 -100 -1670 -80
rect -1650 -100 -1630 -80
rect -1610 -100 -1590 -80
rect -1570 -100 -1550 -80
rect -1530 -100 -1510 -80
rect -1490 -100 -1470 -80
rect -1450 -100 -1430 -80
rect -1410 -100 -1390 -80
rect -1370 -100 -1350 -80
rect -1330 -100 -1310 -80
rect -1290 -100 -1270 -80
rect -1250 -100 -1230 -80
rect -1210 -100 -1190 -80
rect -1170 -100 -1150 -80
rect -1130 -100 -1110 -80
rect -1090 -100 -1070 -80
rect -1050 -100 -1030 -80
rect -1005 -100 -985 -80
rect -3485 -110 -985 -100
rect -3485 -150 -985 -140
rect -3485 -170 -3470 -150
rect -3450 -170 -3430 -150
rect -3410 -170 -3390 -150
rect -3370 -170 -3350 -150
rect -3330 -170 -3310 -150
rect -3290 -170 -3270 -150
rect -3250 -170 -3230 -150
rect -3210 -170 -3190 -150
rect -3170 -170 -3150 -150
rect -3130 -170 -3110 -150
rect -3090 -170 -3070 -150
rect -3050 -170 -3030 -150
rect -3010 -170 -2990 -150
rect -2970 -170 -2950 -150
rect -2930 -170 -2910 -150
rect -2890 -170 -2870 -150
rect -2850 -170 -2830 -150
rect -2810 -170 -2790 -150
rect -2770 -170 -2750 -150
rect -2730 -170 -2710 -150
rect -2690 -170 -2670 -150
rect -2650 -170 -2630 -150
rect -2610 -170 -2590 -150
rect -2570 -170 -2550 -150
rect -2530 -170 -2510 -150
rect -2490 -170 -2470 -150
rect -2450 -170 -2430 -150
rect -2410 -170 -2390 -150
rect -2370 -170 -2350 -150
rect -2330 -170 -2310 -150
rect -2290 -170 -2270 -150
rect -2250 -170 -2230 -150
rect -2210 -170 -2190 -150
rect -2170 -170 -2150 -150
rect -2130 -170 -2110 -150
rect -2090 -170 -2070 -150
rect -2050 -170 -2030 -150
rect -2010 -170 -1990 -150
rect -1970 -170 -1950 -150
rect -1930 -170 -1910 -150
rect -1890 -170 -1870 -150
rect -1850 -170 -1830 -150
rect -1810 -170 -1790 -150
rect -1770 -170 -1750 -150
rect -1730 -170 -1710 -150
rect -1690 -170 -1670 -150
rect -1650 -170 -1630 -150
rect -1610 -170 -1590 -150
rect -1570 -170 -1550 -150
rect -1530 -170 -1510 -150
rect -1490 -170 -1470 -150
rect -1450 -170 -1430 -150
rect -1410 -170 -1390 -150
rect -1370 -170 -1350 -150
rect -1330 -170 -1310 -150
rect -1290 -170 -1270 -150
rect -1250 -170 -1230 -150
rect -1210 -170 -1190 -150
rect -1170 -170 -1150 -150
rect -1130 -170 -1110 -150
rect -1090 -170 -1070 -150
rect -1050 -170 -1030 -150
rect -1005 -170 -985 -150
rect -3660 -180 -3505 -170
rect -3485 -180 -985 -170
rect -3660 -205 -3650 -180
rect -3630 -205 -3610 -180
rect -3590 -205 -3570 -180
rect -3550 -205 -3530 -180
rect -3660 -215 -3505 -205
rect -3485 -215 -985 -205
rect -3485 -235 -3470 -215
rect -3450 -235 -3430 -215
rect -3410 -235 -3390 -215
rect -3370 -235 -3350 -215
rect -3330 -235 -3310 -215
rect -3290 -235 -3270 -215
rect -3250 -235 -3230 -215
rect -3210 -235 -3190 -215
rect -3170 -235 -3150 -215
rect -3130 -235 -3110 -215
rect -3090 -235 -3070 -215
rect -3050 -235 -3030 -215
rect -3010 -235 -2990 -215
rect -2970 -235 -2950 -215
rect -2930 -235 -2910 -215
rect -2890 -235 -2870 -215
rect -2850 -235 -2830 -215
rect -2810 -235 -2790 -215
rect -2770 -235 -2750 -215
rect -2730 -235 -2710 -215
rect -2690 -235 -2670 -215
rect -2650 -235 -2630 -215
rect -2610 -235 -2590 -215
rect -2570 -235 -2550 -215
rect -2530 -235 -2510 -215
rect -2490 -235 -2470 -215
rect -2450 -235 -2430 -215
rect -2410 -235 -2390 -215
rect -2370 -235 -2350 -215
rect -2330 -235 -2310 -215
rect -2290 -235 -2270 -215
rect -2250 -235 -2230 -215
rect -2210 -235 -2190 -215
rect -2170 -235 -2150 -215
rect -2130 -235 -2110 -215
rect -2090 -235 -2070 -215
rect -2050 -235 -2030 -215
rect -2010 -235 -1990 -215
rect -1970 -235 -1950 -215
rect -1930 -235 -1910 -215
rect -1890 -235 -1870 -215
rect -1850 -235 -1830 -215
rect -1810 -235 -1790 -215
rect -1770 -235 -1750 -215
rect -1730 -235 -1710 -215
rect -1690 -235 -1670 -215
rect -1650 -235 -1630 -215
rect -1610 -235 -1590 -215
rect -1570 -235 -1550 -215
rect -1530 -235 -1510 -215
rect -1490 -235 -1470 -215
rect -1450 -235 -1430 -215
rect -1410 -235 -1390 -215
rect -1370 -235 -1350 -215
rect -1330 -235 -1310 -215
rect -1290 -235 -1270 -215
rect -1250 -235 -1230 -215
rect -1210 -235 -1190 -215
rect -1170 -235 -1150 -215
rect -1130 -235 -1110 -215
rect -1090 -235 -1070 -215
rect -1050 -235 -1030 -215
rect -1005 -235 -985 -215
rect -3660 -245 -3505 -235
rect -3485 -245 -985 -235
rect -3660 -270 -3650 -245
rect -3630 -270 -3610 -245
rect -3590 -270 -3570 -245
rect -3550 -270 -3530 -245
rect -3660 -280 -3505 -270
rect -3485 -280 -985 -270
rect -3485 -300 -3470 -280
rect -3450 -300 -3430 -280
rect -3410 -300 -3390 -280
rect -3370 -300 -3350 -280
rect -3330 -300 -3310 -280
rect -3290 -300 -3270 -280
rect -3250 -300 -3230 -280
rect -3210 -300 -3190 -280
rect -3170 -300 -3150 -280
rect -3130 -300 -3110 -280
rect -3090 -300 -3070 -280
rect -3050 -300 -3030 -280
rect -3010 -300 -2990 -280
rect -2970 -300 -2950 -280
rect -2930 -300 -2910 -280
rect -2890 -300 -2870 -280
rect -2850 -300 -2830 -280
rect -2810 -300 -2790 -280
rect -2770 -300 -2750 -280
rect -2730 -300 -2710 -280
rect -2690 -300 -2670 -280
rect -2650 -300 -2630 -280
rect -2610 -300 -2590 -280
rect -2570 -300 -2550 -280
rect -2530 -300 -2510 -280
rect -2490 -300 -2470 -280
rect -2450 -300 -2430 -280
rect -2410 -300 -2390 -280
rect -2370 -300 -2350 -280
rect -2330 -300 -2310 -280
rect -2290 -300 -2270 -280
rect -2250 -300 -2230 -280
rect -2210 -300 -2190 -280
rect -2170 -300 -2150 -280
rect -2130 -300 -2110 -280
rect -2090 -300 -2070 -280
rect -2050 -300 -2030 -280
rect -2010 -300 -1990 -280
rect -1970 -300 -1950 -280
rect -1930 -300 -1910 -280
rect -1890 -300 -1870 -280
rect -1850 -300 -1830 -280
rect -1810 -300 -1790 -280
rect -1770 -300 -1750 -280
rect -1730 -300 -1710 -280
rect -1690 -300 -1670 -280
rect -1650 -300 -1630 -280
rect -1610 -300 -1590 -280
rect -1570 -300 -1550 -280
rect -1530 -300 -1510 -280
rect -1490 -300 -1470 -280
rect -1450 -300 -1430 -280
rect -1410 -300 -1390 -280
rect -1370 -300 -1350 -280
rect -1330 -300 -1310 -280
rect -1290 -300 -1270 -280
rect -1250 -300 -1230 -280
rect -1210 -300 -1190 -280
rect -1170 -300 -1150 -280
rect -1130 -300 -1110 -280
rect -1090 -300 -1070 -280
rect -1050 -300 -1030 -280
rect -1005 -300 -985 -280
rect -3660 -310 -3505 -300
rect -3485 -310 -985 -300
rect -3660 -335 -3650 -310
rect -3630 -335 -3610 -310
rect -3590 -335 -3570 -310
rect -3550 -335 -3530 -310
rect -3660 -345 -3505 -335
rect -3485 -345 -985 -335
rect -3485 -365 -3470 -345
rect -3450 -365 -3430 -345
rect -3410 -365 -3390 -345
rect -3370 -365 -3350 -345
rect -3330 -365 -3310 -345
rect -3290 -365 -3270 -345
rect -3250 -365 -3230 -345
rect -3210 -365 -3190 -345
rect -3170 -365 -3150 -345
rect -3130 -365 -3110 -345
rect -3090 -365 -3070 -345
rect -3050 -365 -3030 -345
rect -3010 -365 -2990 -345
rect -2970 -365 -2950 -345
rect -2930 -365 -2910 -345
rect -2890 -365 -2870 -345
rect -2850 -365 -2830 -345
rect -2810 -365 -2790 -345
rect -2770 -365 -2750 -345
rect -2730 -365 -2710 -345
rect -2690 -365 -2670 -345
rect -2650 -365 -2630 -345
rect -2610 -365 -2590 -345
rect -2570 -365 -2550 -345
rect -2530 -365 -2510 -345
rect -2490 -365 -2470 -345
rect -2450 -365 -2430 -345
rect -2410 -365 -2390 -345
rect -2370 -365 -2350 -345
rect -2330 -365 -2310 -345
rect -2290 -365 -2270 -345
rect -2250 -365 -2230 -345
rect -2210 -365 -2190 -345
rect -2170 -365 -2150 -345
rect -2130 -365 -2110 -345
rect -2090 -365 -2070 -345
rect -2050 -365 -2030 -345
rect -2010 -365 -1990 -345
rect -1970 -365 -1950 -345
rect -1930 -365 -1910 -345
rect -1890 -365 -1870 -345
rect -1850 -365 -1830 -345
rect -1810 -365 -1790 -345
rect -1770 -365 -1750 -345
rect -1730 -365 -1710 -345
rect -1690 -365 -1670 -345
rect -1650 -365 -1630 -345
rect -1610 -365 -1590 -345
rect -1570 -365 -1550 -345
rect -1530 -365 -1510 -345
rect -1490 -365 -1470 -345
rect -1450 -365 -1430 -345
rect -1410 -365 -1390 -345
rect -1370 -365 -1350 -345
rect -1330 -365 -1310 -345
rect -1290 -365 -1270 -345
rect -1250 -365 -1230 -345
rect -1210 -365 -1190 -345
rect -1170 -365 -1150 -345
rect -1130 -365 -1110 -345
rect -1090 -365 -1070 -345
rect -1050 -365 -1030 -345
rect -1005 -365 -985 -345
rect -3660 -375 -3505 -365
rect -3485 -375 -985 -365
rect -3660 -400 -3650 -375
rect -3630 -400 -3610 -375
rect -3590 -400 -3570 -375
rect -3550 -400 -3530 -375
rect -3660 -410 -3505 -400
rect -3485 -410 -985 -400
rect -3485 -430 -3470 -410
rect -3450 -430 -3430 -410
rect -3410 -430 -3390 -410
rect -3370 -430 -3350 -410
rect -3330 -430 -3310 -410
rect -3290 -430 -3270 -410
rect -3250 -430 -3230 -410
rect -3210 -430 -3190 -410
rect -3170 -430 -3150 -410
rect -3130 -430 -3110 -410
rect -3090 -430 -3070 -410
rect -3050 -430 -3030 -410
rect -3010 -430 -2990 -410
rect -2970 -430 -2950 -410
rect -2930 -430 -2910 -410
rect -2890 -430 -2870 -410
rect -2850 -430 -2830 -410
rect -2810 -430 -2790 -410
rect -2770 -430 -2750 -410
rect -2730 -430 -2710 -410
rect -2690 -430 -2670 -410
rect -2650 -430 -2630 -410
rect -2610 -430 -2590 -410
rect -2570 -430 -2550 -410
rect -2530 -430 -2510 -410
rect -2490 -430 -2470 -410
rect -2450 -430 -2430 -410
rect -2410 -430 -2390 -410
rect -2370 -430 -2350 -410
rect -2330 -430 -2310 -410
rect -2290 -430 -2270 -410
rect -2250 -430 -2230 -410
rect -2210 -430 -2190 -410
rect -2170 -430 -2150 -410
rect -2130 -430 -2110 -410
rect -2090 -430 -2070 -410
rect -2050 -430 -2030 -410
rect -2010 -430 -1990 -410
rect -1970 -430 -1950 -410
rect -1930 -430 -1910 -410
rect -1890 -430 -1870 -410
rect -1850 -430 -1830 -410
rect -1810 -430 -1790 -410
rect -1770 -430 -1750 -410
rect -1730 -430 -1710 -410
rect -1690 -430 -1670 -410
rect -1650 -430 -1630 -410
rect -1610 -430 -1590 -410
rect -1570 -430 -1550 -410
rect -1530 -430 -1510 -410
rect -1490 -430 -1470 -410
rect -1450 -430 -1430 -410
rect -1410 -430 -1390 -410
rect -1370 -430 -1350 -410
rect -1330 -430 -1310 -410
rect -1290 -430 -1270 -410
rect -1250 -430 -1230 -410
rect -1210 -430 -1190 -410
rect -1170 -430 -1150 -410
rect -1130 -430 -1110 -410
rect -1090 -430 -1070 -410
rect -1050 -430 -1030 -410
rect -1005 -430 -985 -410
rect -3660 -440 -3505 -430
rect -3485 -440 -985 -430
rect -3660 -465 -3650 -440
rect -3630 -465 -3610 -440
rect -3590 -465 -3570 -440
rect -3550 -465 -3530 -440
rect -3660 -475 -3505 -465
rect -3485 -475 -985 -465
rect -3485 -495 -3470 -475
rect -3450 -495 -3430 -475
rect -3410 -495 -3390 -475
rect -3370 -495 -3350 -475
rect -3330 -495 -3310 -475
rect -3290 -495 -3270 -475
rect -3250 -495 -3230 -475
rect -3210 -495 -3190 -475
rect -3170 -495 -3150 -475
rect -3130 -495 -3110 -475
rect -3090 -495 -3070 -475
rect -3050 -495 -3030 -475
rect -3010 -495 -2990 -475
rect -2970 -495 -2950 -475
rect -2930 -495 -2910 -475
rect -2890 -495 -2870 -475
rect -2850 -495 -2830 -475
rect -2810 -495 -2790 -475
rect -2770 -495 -2750 -475
rect -2730 -495 -2710 -475
rect -2690 -495 -2670 -475
rect -2650 -495 -2630 -475
rect -2610 -495 -2590 -475
rect -2570 -495 -2550 -475
rect -2530 -495 -2510 -475
rect -2490 -495 -2470 -475
rect -2450 -495 -2430 -475
rect -2410 -495 -2390 -475
rect -2370 -495 -2350 -475
rect -2330 -495 -2310 -475
rect -2290 -495 -2270 -475
rect -2250 -495 -2230 -475
rect -2210 -495 -2190 -475
rect -2170 -495 -2150 -475
rect -2130 -495 -2110 -475
rect -2090 -495 -2070 -475
rect -2050 -495 -2030 -475
rect -2010 -495 -1990 -475
rect -1970 -495 -1950 -475
rect -1930 -495 -1910 -475
rect -1890 -495 -1870 -475
rect -1850 -495 -1830 -475
rect -1810 -495 -1790 -475
rect -1770 -495 -1750 -475
rect -1730 -495 -1710 -475
rect -1690 -495 -1670 -475
rect -1650 -495 -1630 -475
rect -1610 -495 -1590 -475
rect -1570 -495 -1550 -475
rect -1530 -495 -1510 -475
rect -1490 -495 -1470 -475
rect -1450 -495 -1430 -475
rect -1410 -495 -1390 -475
rect -1370 -495 -1350 -475
rect -1330 -495 -1310 -475
rect -1290 -495 -1270 -475
rect -1250 -495 -1230 -475
rect -1210 -495 -1190 -475
rect -1170 -495 -1150 -475
rect -1130 -495 -1110 -475
rect -1090 -495 -1070 -475
rect -1050 -495 -1030 -475
rect -1005 -495 -985 -475
rect -3660 -505 -3505 -495
rect -3485 -505 -985 -495
rect -3660 -530 -3650 -505
rect -3630 -530 -3610 -505
rect -3590 -530 -3570 -505
rect -3550 -530 -3530 -505
rect -3660 -540 -3505 -530
rect -3485 -540 -985 -530
rect -3485 -560 -3470 -540
rect -3450 -560 -3430 -540
rect -3410 -560 -3390 -540
rect -3370 -560 -3350 -540
rect -3330 -560 -3310 -540
rect -3290 -560 -3270 -540
rect -3250 -560 -3230 -540
rect -3210 -560 -3190 -540
rect -3170 -560 -3150 -540
rect -3130 -560 -3110 -540
rect -3090 -560 -3070 -540
rect -3050 -560 -3030 -540
rect -3010 -560 -2990 -540
rect -2970 -560 -2950 -540
rect -2930 -560 -2910 -540
rect -2890 -560 -2870 -540
rect -2850 -560 -2830 -540
rect -2810 -560 -2790 -540
rect -2770 -560 -2750 -540
rect -2730 -560 -2710 -540
rect -2690 -560 -2670 -540
rect -2650 -560 -2630 -540
rect -2610 -560 -2590 -540
rect -2570 -560 -2550 -540
rect -2530 -560 -2510 -540
rect -2490 -560 -2470 -540
rect -2450 -560 -2430 -540
rect -2410 -560 -2390 -540
rect -2370 -560 -2350 -540
rect -2330 -560 -2310 -540
rect -2290 -560 -2270 -540
rect -2250 -560 -2230 -540
rect -2210 -560 -2190 -540
rect -2170 -560 -2150 -540
rect -2130 -560 -2110 -540
rect -2090 -560 -2070 -540
rect -2050 -560 -2030 -540
rect -2010 -560 -1990 -540
rect -1970 -560 -1950 -540
rect -1930 -560 -1910 -540
rect -1890 -560 -1870 -540
rect -1850 -560 -1830 -540
rect -1810 -560 -1790 -540
rect -1770 -560 -1750 -540
rect -1730 -560 -1710 -540
rect -1690 -560 -1670 -540
rect -1650 -560 -1630 -540
rect -1610 -560 -1590 -540
rect -1570 -560 -1550 -540
rect -1530 -560 -1510 -540
rect -1490 -560 -1470 -540
rect -1450 -560 -1430 -540
rect -1410 -560 -1390 -540
rect -1370 -560 -1350 -540
rect -1330 -560 -1310 -540
rect -1290 -560 -1270 -540
rect -1250 -560 -1230 -540
rect -1210 -560 -1190 -540
rect -1170 -560 -1150 -540
rect -1130 -560 -1110 -540
rect -1090 -560 -1070 -540
rect -1050 -560 -1030 -540
rect -1005 -560 -985 -540
rect -3485 -570 -985 -560
rect -3485 -610 -985 -600
rect -3485 -630 -3470 -610
rect -3450 -630 -3430 -610
rect -3410 -630 -3390 -610
rect -3370 -630 -3350 -610
rect -3330 -630 -3310 -610
rect -3290 -630 -3270 -610
rect -3250 -630 -3230 -610
rect -3210 -630 -3190 -610
rect -3170 -630 -3150 -610
rect -3130 -630 -3110 -610
rect -3090 -630 -3070 -610
rect -3050 -630 -3030 -610
rect -3010 -630 -2990 -610
rect -2970 -630 -2950 -610
rect -2930 -630 -2910 -610
rect -2890 -630 -2870 -610
rect -2850 -630 -2830 -610
rect -2810 -630 -2790 -610
rect -2770 -630 -2750 -610
rect -2730 -630 -2710 -610
rect -2690 -630 -2670 -610
rect -2650 -630 -2630 -610
rect -2610 -630 -2590 -610
rect -2570 -630 -2550 -610
rect -2530 -630 -2510 -610
rect -2490 -630 -2470 -610
rect -2450 -630 -2430 -610
rect -2410 -630 -2390 -610
rect -2370 -630 -2350 -610
rect -2330 -630 -2310 -610
rect -2290 -630 -2270 -610
rect -2250 -630 -2230 -610
rect -2210 -630 -2190 -610
rect -2170 -630 -2150 -610
rect -2130 -630 -2110 -610
rect -2090 -630 -2070 -610
rect -2050 -630 -2030 -610
rect -2010 -630 -1990 -610
rect -1970 -630 -1950 -610
rect -1930 -630 -1910 -610
rect -1890 -630 -1870 -610
rect -1850 -630 -1830 -610
rect -1810 -630 -1790 -610
rect -1770 -630 -1750 -610
rect -1730 -630 -1710 -610
rect -1690 -630 -1670 -610
rect -1650 -630 -1630 -610
rect -1610 -630 -1590 -610
rect -1570 -630 -1550 -610
rect -1530 -630 -1510 -610
rect -1490 -630 -1470 -610
rect -1450 -630 -1430 -610
rect -1410 -630 -1390 -610
rect -1370 -630 -1350 -610
rect -1330 -630 -1310 -610
rect -1290 -630 -1270 -610
rect -1250 -630 -1230 -610
rect -1210 -630 -1190 -610
rect -1170 -630 -1150 -610
rect -1130 -630 -1110 -610
rect -1090 -630 -1070 -610
rect -1050 -630 -1030 -610
rect -1005 -630 -985 -610
rect -3485 -640 -985 -630
<< viali >>
rect -1550 1415 -1530 1435
rect -1510 1415 -1490 1435
rect -1470 1415 -1450 1435
rect -1430 1415 -1410 1435
rect -1390 1415 -1370 1435
rect -1350 1415 -1330 1435
rect -1310 1415 -1290 1435
rect -1270 1415 -1250 1435
rect -1230 1415 -1210 1435
rect -1190 1415 -1170 1435
rect -1150 1415 -1130 1435
rect -1110 1415 -1090 1435
rect -1070 1415 -1050 1435
rect -1030 1415 -1010 1435
rect -990 1415 -970 1435
rect -950 1415 -930 1435
rect -910 1415 -890 1435
rect -870 1415 -850 1435
rect -830 1415 -810 1435
rect -790 1415 -770 1435
rect -1550 1375 -1530 1395
rect -1510 1375 -1490 1395
rect -1470 1375 -1450 1395
rect -1430 1375 -1410 1395
rect -1390 1375 -1370 1395
rect -1350 1375 -1330 1395
rect -1310 1375 -1290 1395
rect -1270 1375 -1250 1395
rect -1230 1375 -1210 1395
rect -1190 1375 -1170 1395
rect -1150 1375 -1130 1395
rect -1110 1375 -1090 1395
rect -1070 1375 -1050 1395
rect -1030 1375 -1010 1395
rect -990 1375 -970 1395
rect -950 1375 -930 1395
rect -910 1375 -890 1395
rect -870 1375 -850 1395
rect -830 1375 -810 1395
rect -790 1375 -770 1395
rect -3655 1340 -3635 1360
rect -3615 1340 -3595 1360
rect -3575 1340 -3555 1360
rect -3535 1340 -3515 1360
rect -2510 1307 -2490 1327
rect -2470 1307 -2450 1327
rect -2430 1307 -2410 1327
rect -2390 1307 -2370 1327
rect -2350 1307 -2330 1327
rect -2310 1307 -2290 1327
rect -2270 1307 -2250 1327
rect -2230 1307 -2210 1327
rect -2190 1307 -2170 1327
rect -2150 1307 -2130 1327
rect -2110 1307 -2090 1327
rect -2070 1307 -2050 1327
rect -2030 1307 -2010 1327
rect -1990 1307 -1970 1327
rect -1950 1307 -1930 1327
rect -1910 1307 -1890 1327
rect -1870 1307 -1850 1327
rect -1830 1307 -1810 1327
rect -1790 1307 -1770 1327
rect -1750 1307 -1730 1327
rect -3655 1270 -3635 1290
rect -3615 1270 -3595 1290
rect -3575 1270 -3555 1290
rect -3535 1270 -3515 1290
rect -1550 1239 -1530 1259
rect -1510 1239 -1490 1259
rect -1470 1239 -1450 1259
rect -1430 1239 -1410 1259
rect -1390 1239 -1370 1259
rect -1350 1239 -1330 1259
rect -1310 1239 -1290 1259
rect -1270 1239 -1250 1259
rect -1230 1239 -1210 1259
rect -1190 1239 -1170 1259
rect -1150 1239 -1130 1259
rect -1110 1239 -1090 1259
rect -1070 1239 -1050 1259
rect -1030 1239 -1010 1259
rect -990 1239 -970 1259
rect -950 1239 -930 1259
rect -910 1239 -890 1259
rect -870 1239 -850 1259
rect -830 1239 -810 1259
rect -790 1239 -770 1259
rect -3655 1205 -3635 1225
rect -3615 1205 -3595 1225
rect -3575 1205 -3555 1225
rect -3535 1205 -3515 1225
rect -2510 1171 -2490 1191
rect -2470 1171 -2450 1191
rect -2430 1171 -2410 1191
rect -2390 1171 -2370 1191
rect -2350 1171 -2330 1191
rect -2310 1171 -2290 1191
rect -2270 1171 -2250 1191
rect -2230 1171 -2210 1191
rect -2190 1171 -2170 1191
rect -2150 1171 -2130 1191
rect -2110 1171 -2090 1191
rect -2070 1171 -2050 1191
rect -2030 1171 -2010 1191
rect -1990 1171 -1970 1191
rect -1950 1171 -1930 1191
rect -1910 1171 -1890 1191
rect -1870 1171 -1850 1191
rect -1830 1171 -1810 1191
rect -1790 1171 -1770 1191
rect -1750 1171 -1730 1191
rect -3655 1140 -3635 1160
rect -3615 1140 -3595 1160
rect -3575 1140 -3555 1160
rect -3535 1140 -3515 1160
rect -1550 1103 -1530 1123
rect -1510 1103 -1490 1123
rect -1470 1103 -1450 1123
rect -1430 1103 -1410 1123
rect -1390 1103 -1370 1123
rect -1350 1103 -1330 1123
rect -1310 1103 -1290 1123
rect -1270 1103 -1250 1123
rect -1230 1103 -1210 1123
rect -1190 1103 -1170 1123
rect -1150 1103 -1130 1123
rect -1110 1103 -1090 1123
rect -1070 1103 -1050 1123
rect -1030 1103 -1010 1123
rect -990 1103 -970 1123
rect -950 1103 -930 1123
rect -910 1103 -890 1123
rect -870 1103 -850 1123
rect -830 1103 -810 1123
rect -790 1103 -770 1123
rect -3655 1070 -3635 1090
rect -3615 1070 -3595 1090
rect -3575 1070 -3555 1090
rect -3535 1070 -3515 1090
rect -2510 1035 -2490 1055
rect -2470 1035 -2450 1055
rect -2430 1035 -2410 1055
rect -2390 1035 -2370 1055
rect -2350 1035 -2330 1055
rect -2310 1035 -2290 1055
rect -2270 1035 -2250 1055
rect -2230 1035 -2210 1055
rect -2190 1035 -2170 1055
rect -2150 1035 -2130 1055
rect -2110 1035 -2090 1055
rect -2070 1035 -2050 1055
rect -2030 1035 -2010 1055
rect -1990 1035 -1970 1055
rect -1950 1035 -1930 1055
rect -1910 1035 -1890 1055
rect -1870 1035 -1850 1055
rect -1830 1035 -1810 1055
rect -1790 1035 -1770 1055
rect -1750 1035 -1730 1055
rect -3655 1000 -3635 1020
rect -3615 1000 -3595 1020
rect -3575 1000 -3555 1020
rect -3535 1000 -3515 1020
rect -1550 967 -1530 987
rect -1510 967 -1490 987
rect -1470 967 -1450 987
rect -1430 967 -1410 987
rect -1390 967 -1370 987
rect -1350 967 -1330 987
rect -1310 967 -1290 987
rect -1270 967 -1250 987
rect -1230 967 -1210 987
rect -1190 967 -1170 987
rect -1150 967 -1130 987
rect -1110 967 -1090 987
rect -1070 967 -1050 987
rect -1030 967 -1010 987
rect -990 967 -970 987
rect -950 967 -930 987
rect -910 967 -890 987
rect -870 967 -850 987
rect -830 967 -810 987
rect -790 967 -770 987
rect -3655 935 -3635 955
rect -3615 935 -3595 955
rect -3575 935 -3555 955
rect -3535 935 -3515 955
rect -2510 899 -2490 919
rect -2470 899 -2450 919
rect -2430 899 -2410 919
rect -2390 899 -2370 919
rect -2350 899 -2330 919
rect -2310 899 -2290 919
rect -2270 899 -2250 919
rect -2230 899 -2210 919
rect -2190 899 -2170 919
rect -2150 899 -2130 919
rect -2110 899 -2090 919
rect -2070 899 -2050 919
rect -2030 899 -2010 919
rect -1990 899 -1970 919
rect -1950 899 -1930 919
rect -1910 899 -1890 919
rect -1870 899 -1850 919
rect -1830 899 -1810 919
rect -1790 899 -1770 919
rect -1750 899 -1730 919
rect -3655 865 -3635 885
rect -3615 865 -3595 885
rect -3575 865 -3555 885
rect -3535 865 -3515 885
rect -1550 831 -1530 851
rect -1510 831 -1490 851
rect -1470 831 -1450 851
rect -1430 831 -1410 851
rect -1390 831 -1370 851
rect -1350 831 -1330 851
rect -1310 831 -1290 851
rect -1270 831 -1250 851
rect -1230 831 -1210 851
rect -1190 831 -1170 851
rect -1150 831 -1130 851
rect -1110 831 -1090 851
rect -1070 831 -1050 851
rect -1030 831 -1010 851
rect -990 831 -970 851
rect -950 831 -930 851
rect -910 831 -890 851
rect -870 831 -850 851
rect -830 831 -810 851
rect -790 831 -770 851
rect -3655 795 -3635 815
rect -3615 795 -3595 815
rect -3575 795 -3555 815
rect -3535 795 -3515 815
rect -2510 763 -2490 783
rect -2470 763 -2450 783
rect -2430 763 -2410 783
rect -2390 763 -2370 783
rect -2350 763 -2330 783
rect -2310 763 -2290 783
rect -2270 763 -2250 783
rect -2230 763 -2210 783
rect -2190 763 -2170 783
rect -2150 763 -2130 783
rect -2110 763 -2090 783
rect -2070 763 -2050 783
rect -2030 763 -2010 783
rect -1990 763 -1970 783
rect -1950 763 -1930 783
rect -1910 763 -1890 783
rect -1870 763 -1850 783
rect -1830 763 -1810 783
rect -1790 763 -1770 783
rect -1750 763 -1730 783
rect -3655 730 -3635 750
rect -3615 730 -3595 750
rect -3575 730 -3555 750
rect -3535 730 -3515 750
rect -1550 695 -1530 715
rect -1510 695 -1490 715
rect -1470 695 -1450 715
rect -1430 695 -1410 715
rect -1390 695 -1370 715
rect -1350 695 -1330 715
rect -1310 695 -1290 715
rect -1270 695 -1250 715
rect -1230 695 -1210 715
rect -1190 695 -1170 715
rect -1150 695 -1130 715
rect -1110 695 -1090 715
rect -1070 695 -1050 715
rect -1030 695 -1010 715
rect -990 695 -970 715
rect -950 695 -930 715
rect -910 695 -890 715
rect -870 695 -850 715
rect -830 695 -810 715
rect -790 695 -770 715
rect -3655 660 -3635 680
rect -3615 660 -3595 680
rect -3575 660 -3555 680
rect -3535 660 -3515 680
rect -2510 627 -2490 647
rect -2470 627 -2450 647
rect -2430 627 -2410 647
rect -2390 627 -2370 647
rect -2350 627 -2330 647
rect -2310 627 -2290 647
rect -2270 627 -2250 647
rect -2230 627 -2210 647
rect -2190 627 -2170 647
rect -2150 627 -2130 647
rect -2110 627 -2090 647
rect -2070 627 -2050 647
rect -2030 627 -2010 647
rect -1990 627 -1970 647
rect -1950 627 -1930 647
rect -1910 627 -1890 647
rect -1870 627 -1850 647
rect -1830 627 -1810 647
rect -1790 627 -1770 647
rect -1750 627 -1730 647
rect -3655 595 -3635 615
rect -3615 595 -3595 615
rect -3575 595 -3555 615
rect -3535 595 -3515 615
rect -1550 559 -1530 579
rect -1510 559 -1490 579
rect -1470 559 -1450 579
rect -1430 559 -1410 579
rect -1390 559 -1370 579
rect -1350 559 -1330 579
rect -1310 559 -1290 579
rect -1270 559 -1250 579
rect -1230 559 -1210 579
rect -1190 559 -1170 579
rect -1150 559 -1130 579
rect -1110 559 -1090 579
rect -1070 559 -1050 579
rect -1030 559 -1010 579
rect -990 559 -970 579
rect -950 559 -930 579
rect -910 559 -890 579
rect -870 559 -850 579
rect -830 559 -810 579
rect -790 559 -770 579
rect -3655 525 -3635 545
rect -3615 525 -3595 545
rect -3575 525 -3555 545
rect -3535 525 -3515 545
rect -2510 491 -2490 511
rect -2470 491 -2450 511
rect -2430 491 -2410 511
rect -2390 491 -2370 511
rect -2350 491 -2330 511
rect -2310 491 -2290 511
rect -2270 491 -2250 511
rect -2230 491 -2210 511
rect -2190 491 -2170 511
rect -2150 491 -2130 511
rect -2110 491 -2090 511
rect -2070 491 -2050 511
rect -2030 491 -2010 511
rect -1990 491 -1970 511
rect -1950 491 -1930 511
rect -1910 491 -1890 511
rect -1870 491 -1850 511
rect -1830 491 -1810 511
rect -1790 491 -1770 511
rect -1750 491 -1730 511
rect -3655 455 -3635 475
rect -3615 455 -3595 475
rect -3575 455 -3555 475
rect -3535 455 -3515 475
rect -1550 423 -1530 443
rect -1510 423 -1490 443
rect -1470 423 -1450 443
rect -1430 423 -1410 443
rect -1390 423 -1370 443
rect -1350 423 -1330 443
rect -1310 423 -1290 443
rect -1270 423 -1250 443
rect -1230 423 -1210 443
rect -1190 423 -1170 443
rect -1150 423 -1130 443
rect -1110 423 -1090 443
rect -1070 423 -1050 443
rect -1030 423 -1010 443
rect -990 423 -970 443
rect -950 423 -930 443
rect -910 423 -890 443
rect -870 423 -850 443
rect -830 423 -810 443
rect -790 423 -770 443
rect -3655 385 -3635 405
rect -3615 385 -3595 405
rect -3575 385 -3555 405
rect -3535 385 -3515 405
rect -2510 355 -2490 375
rect -2470 355 -2450 375
rect -2430 355 -2410 375
rect -2390 355 -2370 375
rect -2350 355 -2330 375
rect -2310 355 -2290 375
rect -2270 355 -2250 375
rect -2230 355 -2210 375
rect -2190 355 -2170 375
rect -2150 355 -2130 375
rect -2110 355 -2090 375
rect -2070 355 -2050 375
rect -2030 355 -2010 375
rect -1990 355 -1970 375
rect -1950 355 -1930 375
rect -1910 355 -1890 375
rect -1870 355 -1850 375
rect -1830 355 -1810 375
rect -1790 355 -1770 375
rect -1750 355 -1730 375
rect -3655 320 -3635 340
rect -3615 320 -3595 340
rect -3575 320 -3555 340
rect -3535 320 -3515 340
rect -1550 287 -1530 307
rect -1510 287 -1490 307
rect -1470 287 -1450 307
rect -1430 287 -1410 307
rect -1390 287 -1370 307
rect -1350 287 -1330 307
rect -1310 287 -1290 307
rect -1270 287 -1250 307
rect -1230 287 -1210 307
rect -1190 287 -1170 307
rect -1150 287 -1130 307
rect -1110 287 -1090 307
rect -1070 287 -1050 307
rect -1030 287 -1010 307
rect -990 287 -970 307
rect -950 287 -930 307
rect -910 287 -890 307
rect -870 287 -850 307
rect -830 287 -810 307
rect -790 287 -770 307
rect -3655 255 -3635 275
rect -3615 255 -3595 275
rect -3575 255 -3555 275
rect -3535 255 -3515 275
rect -2510 219 -2490 239
rect -2470 219 -2450 239
rect -2430 219 -2410 239
rect -2390 219 -2370 239
rect -2350 219 -2330 239
rect -2310 219 -2290 239
rect -2270 219 -2250 239
rect -2230 219 -2210 239
rect -2190 219 -2170 239
rect -2150 219 -2130 239
rect -2110 219 -2090 239
rect -2070 219 -2050 239
rect -2030 219 -2010 239
rect -1990 219 -1970 239
rect -1950 219 -1930 239
rect -1910 219 -1890 239
rect -1870 219 -1850 239
rect -1830 219 -1810 239
rect -1790 219 -1770 239
rect -1750 219 -1730 239
rect -3655 185 -3635 205
rect -3615 185 -3595 205
rect -3575 185 -3555 205
rect -3535 185 -3515 205
rect -1550 151 -1530 171
rect -1510 151 -1490 171
rect -1470 151 -1450 171
rect -1430 151 -1410 171
rect -1390 151 -1370 171
rect -1350 151 -1330 171
rect -1310 151 -1290 171
rect -1270 151 -1250 171
rect -1230 151 -1210 171
rect -1190 151 -1170 171
rect -1150 151 -1130 171
rect -1110 151 -1090 171
rect -1070 151 -1050 171
rect -1030 151 -1010 171
rect -990 151 -970 171
rect -950 151 -930 171
rect -910 151 -890 171
rect -870 151 -850 171
rect -830 151 -810 171
rect -790 151 -770 171
rect -3655 115 -3635 135
rect -3615 115 -3595 135
rect -3575 115 -3555 135
rect -3535 115 -3515 135
rect -2510 83 -2490 103
rect -2470 83 -2450 103
rect -2430 83 -2410 103
rect -2390 83 -2370 103
rect -2350 83 -2330 103
rect -2310 83 -2290 103
rect -2270 83 -2250 103
rect -2230 83 -2210 103
rect -2190 83 -2170 103
rect -2150 83 -2130 103
rect -2110 83 -2090 103
rect -2070 83 -2050 103
rect -2030 83 -2010 103
rect -1990 83 -1970 103
rect -1950 83 -1930 103
rect -1910 83 -1890 103
rect -1870 83 -1850 103
rect -1830 83 -1810 103
rect -1790 83 -1770 103
rect -1750 83 -1730 103
rect -3655 50 -3635 70
rect -3615 50 -3595 70
rect -3575 50 -3555 70
rect -3535 50 -3515 70
rect -1550 15 -1530 35
rect -1510 15 -1490 35
rect -1470 15 -1450 35
rect -1430 15 -1410 35
rect -1390 15 -1370 35
rect -1350 15 -1330 35
rect -1310 15 -1290 35
rect -1270 15 -1250 35
rect -1230 15 -1210 35
rect -1190 15 -1170 35
rect -1150 15 -1130 35
rect -1110 15 -1090 35
rect -1070 15 -1050 35
rect -1030 15 -1010 35
rect -990 15 -970 35
rect -950 15 -930 35
rect -910 15 -890 35
rect -870 15 -850 35
rect -830 15 -810 35
rect -790 15 -770 35
rect -1550 -25 -1530 -5
rect -1510 -25 -1490 -5
rect -1470 -25 -1450 -5
rect -1430 -25 -1410 -5
rect -1390 -25 -1370 -5
rect -1350 -25 -1330 -5
rect -1310 -25 -1290 -5
rect -1270 -25 -1250 -5
rect -1230 -25 -1210 -5
rect -1190 -25 -1170 -5
rect -1150 -25 -1130 -5
rect -1110 -25 -1090 -5
rect -1070 -25 -1050 -5
rect -1030 -25 -1010 -5
rect -990 -25 -970 -5
rect -950 -25 -930 -5
rect -910 -25 -890 -5
rect -870 -25 -850 -5
rect -830 -25 -810 -5
rect -790 -25 -770 -5
rect -1270 -100 -1250 -80
rect -1230 -100 -1210 -80
rect -1190 -100 -1170 -80
rect -3390 -170 -3370 -150
rect -3350 -170 -3330 -150
rect -3310 -170 -3290 -150
rect -3270 -170 -3250 -150
rect -3230 -170 -3210 -150
rect -3190 -170 -3170 -150
rect -3150 -170 -3130 -150
rect -3110 -170 -3090 -150
rect -3070 -170 -3050 -150
rect -3030 -170 -3010 -150
rect -2990 -170 -2970 -150
rect -2950 -170 -2930 -150
rect -2910 -170 -2890 -150
rect -2870 -170 -2850 -150
rect -2830 -170 -2810 -150
rect -2790 -170 -2770 -150
rect -2750 -170 -2730 -150
rect -2710 -170 -2690 -150
rect -2670 -170 -2650 -150
rect -2630 -170 -2610 -150
rect -3650 -205 -3630 -180
rect -3610 -205 -3590 -180
rect -3570 -205 -3550 -180
rect -3530 -205 -3510 -180
rect -2510 -235 -2490 -215
rect -2470 -235 -2450 -215
rect -2430 -235 -2410 -215
rect -2390 -235 -2370 -215
rect -2350 -235 -2330 -215
rect -2310 -235 -2290 -215
rect -2270 -235 -2250 -215
rect -2230 -235 -2210 -215
rect -2190 -235 -2170 -215
rect -2150 -235 -2130 -215
rect -2110 -235 -2090 -215
rect -2070 -235 -2050 -215
rect -2030 -235 -2010 -215
rect -1990 -235 -1970 -215
rect -1950 -235 -1930 -215
rect -1910 -235 -1890 -215
rect -1870 -235 -1850 -215
rect -1830 -235 -1810 -215
rect -1790 -235 -1770 -215
rect -1750 -235 -1730 -215
rect -3650 -270 -3630 -245
rect -3610 -270 -3590 -245
rect -3570 -270 -3550 -245
rect -3530 -270 -3510 -245
rect -3390 -300 -3370 -280
rect -3350 -300 -3330 -280
rect -3310 -300 -3290 -280
rect -3270 -300 -3250 -280
rect -3230 -300 -3210 -280
rect -3190 -300 -3170 -280
rect -3150 -300 -3130 -280
rect -3110 -300 -3090 -280
rect -3070 -300 -3050 -280
rect -3030 -300 -3010 -280
rect -2990 -300 -2970 -280
rect -2950 -300 -2930 -280
rect -2910 -300 -2890 -280
rect -2870 -300 -2850 -280
rect -2830 -300 -2810 -280
rect -2790 -300 -2770 -280
rect -2750 -300 -2730 -280
rect -2710 -300 -2690 -280
rect -2670 -300 -2650 -280
rect -2630 -300 -2610 -280
rect -3650 -335 -3630 -310
rect -3610 -335 -3590 -310
rect -3570 -335 -3550 -310
rect -3530 -335 -3510 -310
rect -2510 -365 -2490 -345
rect -2470 -365 -2450 -345
rect -2430 -365 -2410 -345
rect -2390 -365 -2370 -345
rect -2350 -365 -2330 -345
rect -2310 -365 -2290 -345
rect -2270 -365 -2250 -345
rect -2230 -365 -2210 -345
rect -2190 -365 -2170 -345
rect -2150 -365 -2130 -345
rect -2110 -365 -2090 -345
rect -2070 -365 -2050 -345
rect -2030 -365 -2010 -345
rect -1990 -365 -1970 -345
rect -1950 -365 -1930 -345
rect -1910 -365 -1890 -345
rect -1870 -365 -1850 -345
rect -1830 -365 -1810 -345
rect -1790 -365 -1770 -345
rect -1750 -365 -1730 -345
rect -3650 -400 -3630 -375
rect -3610 -400 -3590 -375
rect -3570 -400 -3550 -375
rect -3530 -400 -3510 -375
rect -3390 -430 -3370 -410
rect -3350 -430 -3330 -410
rect -3310 -430 -3290 -410
rect -3270 -430 -3250 -410
rect -3230 -430 -3210 -410
rect -3190 -430 -3170 -410
rect -3150 -430 -3130 -410
rect -3110 -430 -3090 -410
rect -3070 -430 -3050 -410
rect -3030 -430 -3010 -410
rect -2990 -430 -2970 -410
rect -2950 -430 -2930 -410
rect -2910 -430 -2890 -410
rect -2870 -430 -2850 -410
rect -2830 -430 -2810 -410
rect -2790 -430 -2770 -410
rect -2750 -430 -2730 -410
rect -2710 -430 -2690 -410
rect -2670 -430 -2650 -410
rect -2630 -430 -2610 -410
rect -3650 -465 -3630 -440
rect -3610 -465 -3590 -440
rect -3570 -465 -3550 -440
rect -3530 -465 -3510 -440
rect -2510 -495 -2490 -475
rect -2470 -495 -2450 -475
rect -2430 -495 -2410 -475
rect -2390 -495 -2370 -475
rect -2350 -495 -2330 -475
rect -2310 -495 -2290 -475
rect -2270 -495 -2250 -475
rect -2230 -495 -2210 -475
rect -2190 -495 -2170 -475
rect -2150 -495 -2130 -475
rect -2110 -495 -2090 -475
rect -2070 -495 -2050 -475
rect -2030 -495 -2010 -475
rect -1990 -495 -1970 -475
rect -1950 -495 -1930 -475
rect -1910 -495 -1890 -475
rect -1870 -495 -1850 -475
rect -1830 -495 -1810 -475
rect -1790 -495 -1770 -475
rect -1750 -495 -1730 -475
rect -3650 -530 -3630 -505
rect -3610 -530 -3590 -505
rect -3570 -530 -3550 -505
rect -3530 -530 -3510 -505
rect -3390 -560 -3370 -540
rect -3350 -560 -3330 -540
rect -3310 -560 -3290 -540
rect -3270 -560 -3250 -540
rect -3230 -560 -3210 -540
rect -3190 -560 -3170 -540
rect -3150 -560 -3130 -540
rect -3110 -560 -3090 -540
rect -3070 -560 -3050 -540
rect -3030 -560 -3010 -540
rect -2990 -560 -2970 -540
rect -2950 -560 -2930 -540
rect -2910 -560 -2890 -540
rect -2870 -560 -2850 -540
rect -2830 -560 -2810 -540
rect -2790 -560 -2770 -540
rect -2750 -560 -2730 -540
rect -2710 -560 -2690 -540
rect -2670 -560 -2650 -540
rect -2630 -560 -2610 -540
rect -1270 -630 -1250 -610
rect -1230 -630 -1210 -610
rect -1190 -630 -1170 -610
<< metal1 >>
rect -1560 1435 -760 1460
rect -1560 1415 -1550 1435
rect -1530 1415 -1510 1435
rect -1490 1415 -1470 1435
rect -1450 1415 -1430 1435
rect -1410 1415 -1390 1435
rect -1370 1415 -1350 1435
rect -1330 1415 -1310 1435
rect -1290 1415 -1270 1435
rect -1250 1415 -1230 1435
rect -1210 1415 -1190 1435
rect -1170 1415 -1150 1435
rect -1130 1415 -1110 1435
rect -1090 1415 -1070 1435
rect -1050 1415 -1030 1435
rect -1010 1415 -990 1435
rect -970 1415 -950 1435
rect -930 1415 -910 1435
rect -890 1415 -870 1435
rect -850 1415 -830 1435
rect -810 1415 -790 1435
rect -770 1415 -760 1435
rect -1560 1395 -760 1415
rect -1560 1375 -1550 1395
rect -1530 1375 -1510 1395
rect -1490 1375 -1470 1395
rect -1450 1375 -1430 1395
rect -1410 1375 -1390 1395
rect -1370 1375 -1350 1395
rect -1330 1375 -1310 1395
rect -1290 1375 -1270 1395
rect -1250 1375 -1230 1395
rect -1210 1375 -1190 1395
rect -1170 1375 -1150 1395
rect -1130 1375 -1110 1395
rect -1090 1375 -1070 1395
rect -1050 1375 -1030 1395
rect -1010 1375 -990 1395
rect -970 1375 -950 1395
rect -930 1375 -910 1395
rect -890 1375 -870 1395
rect -850 1375 -830 1395
rect -810 1375 -790 1395
rect -770 1375 -760 1395
rect -3665 1360 -3510 1370
rect -3665 1340 -3655 1360
rect -3635 1340 -3615 1360
rect -3595 1340 -3575 1360
rect -3555 1340 -3535 1360
rect -3515 1340 -3510 1360
rect -3665 1290 -3510 1340
rect -3665 1270 -3655 1290
rect -3635 1270 -3615 1290
rect -3595 1270 -3575 1290
rect -3555 1270 -3535 1290
rect -3515 1270 -3510 1290
rect -3665 1225 -3510 1270
rect -3665 1205 -3655 1225
rect -3635 1205 -3615 1225
rect -3595 1205 -3575 1225
rect -3555 1205 -3535 1225
rect -3515 1205 -3510 1225
rect -3665 1160 -3510 1205
rect -3665 1140 -3655 1160
rect -3635 1140 -3615 1160
rect -3595 1140 -3575 1160
rect -3555 1140 -3535 1160
rect -3515 1140 -3510 1160
rect -3665 1130 -3510 1140
rect -2520 1327 -1720 1337
rect -2520 1307 -2510 1327
rect -2490 1307 -2470 1327
rect -2450 1307 -2430 1327
rect -2410 1307 -2390 1327
rect -2370 1307 -2350 1327
rect -2330 1307 -2310 1327
rect -2290 1307 -2270 1327
rect -2250 1307 -2230 1327
rect -2210 1307 -2190 1327
rect -2170 1307 -2150 1327
rect -2130 1307 -2110 1327
rect -2090 1307 -2070 1327
rect -2050 1307 -2030 1327
rect -2010 1307 -1990 1327
rect -1970 1307 -1950 1327
rect -1930 1307 -1910 1327
rect -1890 1307 -1870 1327
rect -1850 1307 -1830 1327
rect -1810 1307 -1790 1327
rect -1770 1307 -1750 1327
rect -1730 1307 -1720 1327
rect -2520 1191 -1720 1307
rect -2520 1171 -2510 1191
rect -2490 1171 -2470 1191
rect -2450 1171 -2430 1191
rect -2410 1171 -2390 1191
rect -2370 1171 -2350 1191
rect -2330 1171 -2310 1191
rect -2290 1171 -2270 1191
rect -2250 1171 -2230 1191
rect -2210 1171 -2190 1191
rect -2170 1171 -2150 1191
rect -2130 1171 -2110 1191
rect -2090 1171 -2070 1191
rect -2050 1171 -2030 1191
rect -2010 1171 -1990 1191
rect -1970 1171 -1950 1191
rect -1930 1171 -1910 1191
rect -1890 1171 -1870 1191
rect -1850 1171 -1830 1191
rect -1810 1171 -1790 1191
rect -1770 1171 -1750 1191
rect -1730 1171 -1720 1191
rect -3665 1090 -3510 1100
rect -3665 1070 -3655 1090
rect -3635 1070 -3615 1090
rect -3595 1070 -3575 1090
rect -3555 1070 -3535 1090
rect -3515 1070 -3510 1090
rect -3665 1020 -3510 1070
rect -3665 1000 -3655 1020
rect -3635 1000 -3615 1020
rect -3595 1000 -3575 1020
rect -3555 1000 -3535 1020
rect -3515 1000 -3510 1020
rect -3665 955 -3510 1000
rect -3665 935 -3655 955
rect -3635 935 -3615 955
rect -3595 935 -3575 955
rect -3555 935 -3535 955
rect -3515 935 -3510 955
rect -3665 885 -3510 935
rect -3665 865 -3655 885
rect -3635 865 -3615 885
rect -3595 865 -3575 885
rect -3555 865 -3535 885
rect -3515 865 -3510 885
rect -3665 815 -3510 865
rect -3665 795 -3655 815
rect -3635 795 -3615 815
rect -3595 795 -3575 815
rect -3555 795 -3535 815
rect -3515 795 -3510 815
rect -3665 750 -3510 795
rect -3665 730 -3655 750
rect -3635 730 -3615 750
rect -3595 730 -3575 750
rect -3555 730 -3535 750
rect -3515 730 -3510 750
rect -3665 680 -3510 730
rect -3665 660 -3655 680
rect -3635 660 -3615 680
rect -3595 660 -3575 680
rect -3555 660 -3535 680
rect -3515 660 -3510 680
rect -3665 615 -3510 660
rect -3665 595 -3655 615
rect -3635 595 -3615 615
rect -3595 595 -3575 615
rect -3555 595 -3535 615
rect -3515 595 -3510 615
rect -3665 545 -3510 595
rect -3665 525 -3655 545
rect -3635 525 -3615 545
rect -3595 525 -3575 545
rect -3555 525 -3535 545
rect -3515 525 -3510 545
rect -3665 475 -3510 525
rect -3665 455 -3655 475
rect -3635 455 -3615 475
rect -3595 455 -3575 475
rect -3555 455 -3535 475
rect -3515 455 -3510 475
rect -3665 405 -3510 455
rect -3665 385 -3655 405
rect -3635 385 -3615 405
rect -3595 385 -3575 405
rect -3555 385 -3535 405
rect -3515 385 -3510 405
rect -3665 340 -3510 385
rect -3665 320 -3655 340
rect -3635 320 -3615 340
rect -3595 320 -3575 340
rect -3555 320 -3535 340
rect -3515 320 -3510 340
rect -3665 275 -3510 320
rect -3665 255 -3655 275
rect -3635 255 -3615 275
rect -3595 255 -3575 275
rect -3555 255 -3535 275
rect -3515 255 -3510 275
rect -3665 205 -3510 255
rect -3665 185 -3655 205
rect -3635 185 -3615 205
rect -3595 185 -3575 205
rect -3555 185 -3535 205
rect -3515 185 -3510 205
rect -3665 135 -3510 185
rect -3665 115 -3655 135
rect -3635 115 -3615 135
rect -3595 115 -3575 135
rect -3555 115 -3535 135
rect -3515 115 -3510 135
rect -3665 70 -3510 115
rect -3665 50 -3655 70
rect -3635 50 -3615 70
rect -3595 50 -3575 70
rect -3555 50 -3535 70
rect -3515 50 -3510 70
rect -3665 40 -3510 50
rect -2520 1055 -1720 1171
rect -2520 1035 -2510 1055
rect -2490 1035 -2470 1055
rect -2450 1035 -2430 1055
rect -2410 1035 -2390 1055
rect -2370 1035 -2350 1055
rect -2330 1035 -2310 1055
rect -2290 1035 -2270 1055
rect -2250 1035 -2230 1055
rect -2210 1035 -2190 1055
rect -2170 1035 -2150 1055
rect -2130 1035 -2110 1055
rect -2090 1035 -2070 1055
rect -2050 1035 -2030 1055
rect -2010 1035 -1990 1055
rect -1970 1035 -1950 1055
rect -1930 1035 -1910 1055
rect -1890 1035 -1870 1055
rect -1850 1035 -1830 1055
rect -1810 1035 -1790 1055
rect -1770 1035 -1750 1055
rect -1730 1035 -1720 1055
rect -2520 919 -1720 1035
rect -2520 899 -2510 919
rect -2490 899 -2470 919
rect -2450 899 -2430 919
rect -2410 899 -2390 919
rect -2370 899 -2350 919
rect -2330 899 -2310 919
rect -2290 899 -2270 919
rect -2250 899 -2230 919
rect -2210 899 -2190 919
rect -2170 899 -2150 919
rect -2130 899 -2110 919
rect -2090 899 -2070 919
rect -2050 899 -2030 919
rect -2010 899 -1990 919
rect -1970 899 -1950 919
rect -1930 899 -1910 919
rect -1890 899 -1870 919
rect -1850 899 -1830 919
rect -1810 899 -1790 919
rect -1770 899 -1750 919
rect -1730 899 -1720 919
rect -2520 783 -1720 899
rect -2520 763 -2510 783
rect -2490 763 -2470 783
rect -2450 763 -2430 783
rect -2410 763 -2390 783
rect -2370 763 -2350 783
rect -2330 763 -2310 783
rect -2290 763 -2270 783
rect -2250 763 -2230 783
rect -2210 763 -2190 783
rect -2170 763 -2150 783
rect -2130 763 -2110 783
rect -2090 763 -2070 783
rect -2050 763 -2030 783
rect -2010 763 -1990 783
rect -1970 763 -1950 783
rect -1930 763 -1910 783
rect -1890 763 -1870 783
rect -1850 763 -1830 783
rect -1810 763 -1790 783
rect -1770 763 -1750 783
rect -1730 763 -1720 783
rect -2520 647 -1720 763
rect -2520 627 -2510 647
rect -2490 627 -2470 647
rect -2450 627 -2430 647
rect -2410 627 -2390 647
rect -2370 627 -2350 647
rect -2330 627 -2310 647
rect -2290 627 -2270 647
rect -2250 627 -2230 647
rect -2210 627 -2190 647
rect -2170 627 -2150 647
rect -2130 627 -2110 647
rect -2090 627 -2070 647
rect -2050 627 -2030 647
rect -2010 627 -1990 647
rect -1970 627 -1950 647
rect -1930 627 -1910 647
rect -1890 627 -1870 647
rect -1850 627 -1830 647
rect -1810 627 -1790 647
rect -1770 627 -1750 647
rect -1730 627 -1720 647
rect -2520 511 -1720 627
rect -2520 491 -2510 511
rect -2490 491 -2470 511
rect -2450 491 -2430 511
rect -2410 491 -2390 511
rect -2370 491 -2350 511
rect -2330 491 -2310 511
rect -2290 491 -2270 511
rect -2250 491 -2230 511
rect -2210 491 -2190 511
rect -2170 491 -2150 511
rect -2130 491 -2110 511
rect -2090 491 -2070 511
rect -2050 491 -2030 511
rect -2010 491 -1990 511
rect -1970 491 -1950 511
rect -1930 491 -1910 511
rect -1890 491 -1870 511
rect -1850 491 -1830 511
rect -1810 491 -1790 511
rect -1770 491 -1750 511
rect -1730 491 -1720 511
rect -2520 375 -1720 491
rect -2520 355 -2510 375
rect -2490 355 -2470 375
rect -2450 355 -2430 375
rect -2410 355 -2390 375
rect -2370 355 -2350 375
rect -2330 355 -2310 375
rect -2290 355 -2270 375
rect -2250 355 -2230 375
rect -2210 355 -2190 375
rect -2170 355 -2150 375
rect -2130 355 -2110 375
rect -2090 355 -2070 375
rect -2050 355 -2030 375
rect -2010 355 -1990 375
rect -1970 355 -1950 375
rect -1930 355 -1910 375
rect -1890 355 -1870 375
rect -1850 355 -1830 375
rect -1810 355 -1790 375
rect -1770 355 -1750 375
rect -1730 355 -1720 375
rect -2520 239 -1720 355
rect -2520 219 -2510 239
rect -2490 219 -2470 239
rect -2450 219 -2430 239
rect -2410 219 -2390 239
rect -2370 219 -2350 239
rect -2330 219 -2310 239
rect -2290 219 -2270 239
rect -2250 219 -2230 239
rect -2210 219 -2190 239
rect -2170 219 -2150 239
rect -2130 219 -2110 239
rect -2090 219 -2070 239
rect -2050 219 -2030 239
rect -2010 219 -1990 239
rect -1970 219 -1950 239
rect -1930 219 -1910 239
rect -1890 219 -1870 239
rect -1850 219 -1830 239
rect -1810 219 -1790 239
rect -1770 219 -1750 239
rect -1730 219 -1720 239
rect -2520 103 -1720 219
rect -2520 83 -2510 103
rect -2490 83 -2470 103
rect -2450 83 -2430 103
rect -2410 83 -2390 103
rect -2370 83 -2350 103
rect -2330 83 -2310 103
rect -2290 83 -2270 103
rect -2250 83 -2230 103
rect -2210 83 -2190 103
rect -2170 83 -2150 103
rect -2130 83 -2110 103
rect -2090 83 -2070 103
rect -2050 83 -2030 103
rect -2010 83 -1990 103
rect -1970 83 -1950 103
rect -1930 83 -1910 103
rect -1890 83 -1870 103
rect -1850 83 -1830 103
rect -1810 83 -1790 103
rect -1770 83 -1750 103
rect -1730 83 -1720 103
rect -3400 -150 -2600 -140
rect -3400 -170 -3390 -150
rect -3370 -170 -3350 -150
rect -3330 -170 -3310 -150
rect -3290 -170 -3270 -150
rect -3250 -170 -3230 -150
rect -3210 -170 -3190 -150
rect -3170 -170 -3150 -150
rect -3130 -170 -3110 -150
rect -3090 -170 -3070 -150
rect -3050 -170 -3030 -150
rect -3010 -170 -2990 -150
rect -2970 -170 -2950 -150
rect -2930 -170 -2910 -150
rect -2890 -170 -2870 -150
rect -2850 -170 -2830 -150
rect -2810 -170 -2790 -150
rect -2770 -170 -2750 -150
rect -2730 -170 -2710 -150
rect -2690 -170 -2670 -150
rect -2650 -170 -2630 -150
rect -2610 -170 -2600 -150
rect -3660 -180 -3505 -170
rect -3660 -205 -3650 -180
rect -3630 -205 -3610 -180
rect -3590 -205 -3570 -180
rect -3550 -205 -3530 -180
rect -3510 -205 -3505 -180
rect -3660 -245 -3505 -205
rect -3660 -270 -3650 -245
rect -3630 -270 -3610 -245
rect -3590 -270 -3570 -245
rect -3550 -270 -3530 -245
rect -3510 -270 -3505 -245
rect -3660 -310 -3505 -270
rect -3660 -335 -3650 -310
rect -3630 -335 -3610 -310
rect -3590 -335 -3570 -310
rect -3550 -335 -3530 -310
rect -3510 -335 -3505 -310
rect -3660 -375 -3505 -335
rect -3660 -400 -3650 -375
rect -3630 -400 -3610 -375
rect -3590 -400 -3570 -375
rect -3550 -400 -3530 -375
rect -3510 -400 -3505 -375
rect -3660 -440 -3505 -400
rect -3660 -465 -3650 -440
rect -3630 -465 -3610 -440
rect -3590 -465 -3570 -440
rect -3550 -465 -3530 -440
rect -3510 -465 -3505 -440
rect -3660 -505 -3505 -465
rect -3660 -530 -3650 -505
rect -3630 -530 -3610 -505
rect -3590 -530 -3570 -505
rect -3550 -530 -3530 -505
rect -3510 -530 -3505 -505
rect -3660 -540 -3505 -530
rect -3400 -280 -2600 -170
rect -3400 -300 -3390 -280
rect -3370 -300 -3350 -280
rect -3330 -300 -3310 -280
rect -3290 -300 -3270 -280
rect -3250 -300 -3230 -280
rect -3210 -300 -3190 -280
rect -3170 -300 -3150 -280
rect -3130 -300 -3110 -280
rect -3090 -300 -3070 -280
rect -3050 -300 -3030 -280
rect -3010 -300 -2990 -280
rect -2970 -300 -2950 -280
rect -2930 -300 -2910 -280
rect -2890 -300 -2870 -280
rect -2850 -300 -2830 -280
rect -2810 -300 -2790 -280
rect -2770 -300 -2750 -280
rect -2730 -300 -2710 -280
rect -2690 -300 -2670 -280
rect -2650 -300 -2630 -280
rect -2610 -300 -2600 -280
rect -3400 -410 -2600 -300
rect -3400 -430 -3390 -410
rect -3370 -430 -3350 -410
rect -3330 -430 -3310 -410
rect -3290 -430 -3270 -410
rect -3250 -430 -3230 -410
rect -3210 -430 -3190 -410
rect -3170 -430 -3150 -410
rect -3130 -430 -3110 -410
rect -3090 -430 -3070 -410
rect -3050 -430 -3030 -410
rect -3010 -430 -2990 -410
rect -2970 -430 -2950 -410
rect -2930 -430 -2910 -410
rect -2890 -430 -2870 -410
rect -2850 -430 -2830 -410
rect -2810 -430 -2790 -410
rect -2770 -430 -2750 -410
rect -2730 -430 -2710 -410
rect -2690 -430 -2670 -410
rect -2650 -430 -2630 -410
rect -2610 -430 -2600 -410
rect -3400 -540 -2600 -430
rect -2520 -215 -1720 83
rect -1560 1259 -760 1375
rect -1560 1239 -1550 1259
rect -1530 1239 -1510 1259
rect -1490 1239 -1470 1259
rect -1450 1239 -1430 1259
rect -1410 1239 -1390 1259
rect -1370 1239 -1350 1259
rect -1330 1239 -1310 1259
rect -1290 1239 -1270 1259
rect -1250 1239 -1230 1259
rect -1210 1239 -1190 1259
rect -1170 1239 -1150 1259
rect -1130 1239 -1110 1259
rect -1090 1239 -1070 1259
rect -1050 1239 -1030 1259
rect -1010 1239 -990 1259
rect -970 1239 -950 1259
rect -930 1239 -910 1259
rect -890 1239 -870 1259
rect -850 1239 -830 1259
rect -810 1239 -790 1259
rect -770 1239 -760 1259
rect -1560 1123 -760 1239
rect -1560 1103 -1550 1123
rect -1530 1103 -1510 1123
rect -1490 1103 -1470 1123
rect -1450 1103 -1430 1123
rect -1410 1103 -1390 1123
rect -1370 1103 -1350 1123
rect -1330 1103 -1310 1123
rect -1290 1103 -1270 1123
rect -1250 1103 -1230 1123
rect -1210 1103 -1190 1123
rect -1170 1103 -1150 1123
rect -1130 1103 -1110 1123
rect -1090 1103 -1070 1123
rect -1050 1103 -1030 1123
rect -1010 1103 -990 1123
rect -970 1103 -950 1123
rect -930 1103 -910 1123
rect -890 1103 -870 1123
rect -850 1103 -830 1123
rect -810 1103 -790 1123
rect -770 1103 -760 1123
rect -1560 987 -760 1103
rect -1560 967 -1550 987
rect -1530 967 -1510 987
rect -1490 967 -1470 987
rect -1450 967 -1430 987
rect -1410 967 -1390 987
rect -1370 967 -1350 987
rect -1330 967 -1310 987
rect -1290 967 -1270 987
rect -1250 967 -1230 987
rect -1210 967 -1190 987
rect -1170 967 -1150 987
rect -1130 967 -1110 987
rect -1090 967 -1070 987
rect -1050 967 -1030 987
rect -1010 967 -990 987
rect -970 967 -950 987
rect -930 967 -910 987
rect -890 967 -870 987
rect -850 967 -830 987
rect -810 967 -790 987
rect -770 967 -760 987
rect -1560 851 -760 967
rect -1560 831 -1550 851
rect -1530 831 -1510 851
rect -1490 831 -1470 851
rect -1450 831 -1430 851
rect -1410 831 -1390 851
rect -1370 831 -1350 851
rect -1330 831 -1310 851
rect -1290 831 -1270 851
rect -1250 831 -1230 851
rect -1210 831 -1190 851
rect -1170 831 -1150 851
rect -1130 831 -1110 851
rect -1090 831 -1070 851
rect -1050 831 -1030 851
rect -1010 831 -990 851
rect -970 831 -950 851
rect -930 831 -910 851
rect -890 831 -870 851
rect -850 831 -830 851
rect -810 831 -790 851
rect -770 831 -760 851
rect -1560 715 -760 831
rect -1560 695 -1550 715
rect -1530 695 -1510 715
rect -1490 695 -1470 715
rect -1450 695 -1430 715
rect -1410 695 -1390 715
rect -1370 695 -1350 715
rect -1330 695 -1310 715
rect -1290 695 -1270 715
rect -1250 695 -1230 715
rect -1210 695 -1190 715
rect -1170 695 -1150 715
rect -1130 695 -1110 715
rect -1090 695 -1070 715
rect -1050 695 -1030 715
rect -1010 695 -990 715
rect -970 695 -950 715
rect -930 695 -910 715
rect -890 695 -870 715
rect -850 695 -830 715
rect -810 695 -790 715
rect -770 695 -760 715
rect -1560 579 -760 695
rect -1560 559 -1550 579
rect -1530 559 -1510 579
rect -1490 559 -1470 579
rect -1450 559 -1430 579
rect -1410 559 -1390 579
rect -1370 559 -1350 579
rect -1330 559 -1310 579
rect -1290 559 -1270 579
rect -1250 559 -1230 579
rect -1210 559 -1190 579
rect -1170 559 -1150 579
rect -1130 559 -1110 579
rect -1090 559 -1070 579
rect -1050 559 -1030 579
rect -1010 559 -990 579
rect -970 559 -950 579
rect -930 559 -910 579
rect -890 559 -870 579
rect -850 559 -830 579
rect -810 559 -790 579
rect -770 559 -760 579
rect -1560 443 -760 559
rect -1560 423 -1550 443
rect -1530 423 -1510 443
rect -1490 423 -1470 443
rect -1450 423 -1430 443
rect -1410 423 -1390 443
rect -1370 423 -1350 443
rect -1330 423 -1310 443
rect -1290 423 -1270 443
rect -1250 423 -1230 443
rect -1210 423 -1190 443
rect -1170 423 -1150 443
rect -1130 423 -1110 443
rect -1090 423 -1070 443
rect -1050 423 -1030 443
rect -1010 423 -990 443
rect -970 423 -950 443
rect -930 423 -910 443
rect -890 423 -870 443
rect -850 423 -830 443
rect -810 423 -790 443
rect -770 423 -760 443
rect -1560 307 -760 423
rect -1560 287 -1550 307
rect -1530 287 -1510 307
rect -1490 287 -1470 307
rect -1450 287 -1430 307
rect -1410 287 -1390 307
rect -1370 287 -1350 307
rect -1330 287 -1310 307
rect -1290 287 -1270 307
rect -1250 287 -1230 307
rect -1210 287 -1190 307
rect -1170 287 -1150 307
rect -1130 287 -1110 307
rect -1090 287 -1070 307
rect -1050 287 -1030 307
rect -1010 287 -990 307
rect -970 287 -950 307
rect -930 287 -910 307
rect -890 287 -870 307
rect -850 287 -830 307
rect -810 287 -790 307
rect -770 287 -760 307
rect -1560 171 -760 287
rect -1560 151 -1550 171
rect -1530 151 -1510 171
rect -1490 151 -1470 171
rect -1450 151 -1430 171
rect -1410 151 -1390 171
rect -1370 151 -1350 171
rect -1330 151 -1310 171
rect -1290 151 -1270 171
rect -1250 151 -1230 171
rect -1210 151 -1190 171
rect -1170 151 -1150 171
rect -1130 151 -1110 171
rect -1090 151 -1070 171
rect -1050 151 -1030 171
rect -1010 151 -990 171
rect -970 151 -950 171
rect -930 151 -910 171
rect -890 151 -870 171
rect -850 151 -830 171
rect -810 151 -790 171
rect -770 151 -760 171
rect -1560 35 -760 151
rect -1560 15 -1550 35
rect -1530 15 -1510 35
rect -1490 15 -1470 35
rect -1450 15 -1430 35
rect -1410 15 -1390 35
rect -1370 15 -1350 35
rect -1330 15 -1310 35
rect -1290 15 -1270 35
rect -1250 15 -1230 35
rect -1210 15 -1190 35
rect -1170 15 -1150 35
rect -1130 15 -1110 35
rect -1090 15 -1070 35
rect -1050 15 -1030 35
rect -1010 15 -990 35
rect -970 15 -950 35
rect -930 15 -910 35
rect -890 15 -870 35
rect -850 15 -830 35
rect -810 15 -790 35
rect -770 15 -760 35
rect -1560 -5 -760 15
rect -1560 -25 -1550 -5
rect -1530 -25 -1510 -5
rect -1490 -25 -1470 -5
rect -1450 -25 -1430 -5
rect -1410 -25 -1390 -5
rect -1370 -25 -1350 -5
rect -1330 -25 -1310 -5
rect -1290 -25 -1270 -5
rect -1250 -25 -1230 -5
rect -1210 -25 -1190 -5
rect -1170 -25 -1150 -5
rect -1130 -25 -1110 -5
rect -1090 -25 -1070 -5
rect -1050 -25 -1030 -5
rect -1010 -25 -990 -5
rect -970 -25 -950 -5
rect -930 -25 -910 -5
rect -890 -25 -870 -5
rect -850 -25 -830 -5
rect -810 -25 -790 -5
rect -770 -25 -760 -5
rect -1560 -35 -760 -25
rect -2520 -235 -2510 -215
rect -2490 -235 -2470 -215
rect -2450 -235 -2430 -215
rect -2410 -235 -2390 -215
rect -2370 -235 -2350 -215
rect -2330 -235 -2310 -215
rect -2290 -235 -2270 -215
rect -2250 -235 -2230 -215
rect -2210 -235 -2190 -215
rect -2170 -235 -2150 -215
rect -2130 -235 -2110 -215
rect -2090 -235 -2070 -215
rect -2050 -235 -2030 -215
rect -2010 -235 -1990 -215
rect -1970 -235 -1950 -215
rect -1930 -235 -1910 -215
rect -1890 -235 -1870 -215
rect -1850 -235 -1830 -215
rect -1810 -235 -1790 -215
rect -1770 -235 -1750 -215
rect -1730 -235 -1720 -215
rect -2520 -345 -1720 -235
rect -2520 -365 -2510 -345
rect -2490 -365 -2470 -345
rect -2450 -365 -2430 -345
rect -2410 -365 -2390 -345
rect -2370 -365 -2350 -345
rect -2330 -365 -2310 -345
rect -2290 -365 -2270 -345
rect -2250 -365 -2230 -345
rect -2210 -365 -2190 -345
rect -2170 -365 -2150 -345
rect -2130 -365 -2110 -345
rect -2090 -365 -2070 -345
rect -2050 -365 -2030 -345
rect -2010 -365 -1990 -345
rect -1970 -365 -1950 -345
rect -1930 -365 -1910 -345
rect -1890 -365 -1870 -345
rect -1850 -365 -1830 -345
rect -1810 -365 -1790 -345
rect -1770 -365 -1750 -345
rect -1730 -365 -1720 -345
rect -2520 -475 -1720 -365
rect -2520 -495 -2510 -475
rect -2490 -495 -2470 -475
rect -2450 -495 -2430 -475
rect -2410 -495 -2390 -475
rect -2370 -495 -2350 -475
rect -2330 -495 -2310 -475
rect -2290 -495 -2270 -475
rect -2250 -495 -2230 -475
rect -2210 -495 -2190 -475
rect -2170 -495 -2150 -475
rect -2130 -495 -2110 -475
rect -2090 -495 -2070 -475
rect -2050 -495 -2030 -475
rect -2010 -495 -1990 -475
rect -1970 -495 -1950 -475
rect -1930 -495 -1910 -475
rect -1890 -495 -1870 -475
rect -1850 -495 -1830 -475
rect -1810 -495 -1790 -475
rect -1770 -495 -1750 -475
rect -1730 -495 -1720 -475
rect -2520 -505 -1720 -495
rect -1280 -80 -1160 -70
rect -1280 -100 -1270 -80
rect -1250 -100 -1230 -80
rect -1210 -100 -1190 -80
rect -1170 -100 -1160 -80
rect -3400 -560 -3390 -540
rect -3370 -560 -3350 -540
rect -3330 -560 -3310 -540
rect -3290 -560 -3270 -540
rect -3250 -560 -3230 -540
rect -3210 -560 -3190 -540
rect -3170 -560 -3150 -540
rect -3130 -560 -3110 -540
rect -3090 -560 -3070 -540
rect -3050 -560 -3030 -540
rect -3010 -560 -2990 -540
rect -2970 -560 -2950 -540
rect -2930 -560 -2910 -540
rect -2890 -560 -2870 -540
rect -2850 -560 -2830 -540
rect -2810 -560 -2790 -540
rect -2770 -560 -2750 -540
rect -2730 -560 -2710 -540
rect -2690 -560 -2670 -540
rect -2650 -560 -2630 -540
rect -2610 -560 -2600 -540
rect -3400 -655 -2600 -560
rect -1280 -610 -1160 -100
rect -1280 -630 -1270 -610
rect -1250 -630 -1230 -610
rect -1210 -630 -1190 -610
rect -1170 -630 -1160 -610
rect -1280 -655 -1160 -630
<< labels >>
rlabel metal1 -2160 -65 -2160 -65 1 Vout
port 1 n
rlabel metal1 -1165 1455 -1165 1455 1 VDD
port 5 n
rlabel metal1 -3650 -310 -3650 -310 1 Vin
port 2 n
rlabel metal1 -3655 1250 -3655 1250 1 Vcmfb
port 7 n
rlabel metal1 -3655 705 -3655 705 1 Vb2
port 8 n
rlabel metal1 -1220 -650 -1220 -650 1 GND
port 11 n
rlabel metal1 -3000 -650 -3000 -650 1 s
port 3 n
rlabel pdiff -2935 1360 -2935 1360 1 S$
rlabel pdiff -2935 1342 -2935 1342 1 D$
rlabel pdiff -2935 1224 -2935 1224 1 S$
rlabel pdiff -2935 1206 -2935 1206 1 D$
rlabel pdiff -2935 1088 -2935 1088 1 S$
rlabel pdiff -2935 1070 -2935 1070 1 D$
rlabel pdiff -2935 952 -2935 952 1 S$
rlabel pdiff -2935 934 -2935 934 1 D$
rlabel pdiff -2935 816 -2935 816 1 S$
rlabel pdiff -2935 798 -2935 798 1 D$
rlabel pdiff -2935 680 -2935 680 1 S$
rlabel pdiff -2935 662 -2935 662 1 D$
rlabel pdiff -2935 544 -2935 544 1 S$
rlabel pdiff -2935 526 -2935 526 1 D$
rlabel pdiff -2935 408 -2935 408 1 S$
rlabel pdiff -2935 390 -2935 390 1 D$
rlabel pdiff -2935 272 -2935 272 1 S$
rlabel pdiff -2935 254 -2935 254 1 D$
rlabel pdiff -2935 136 -2935 136 1 S$
rlabel pdiff -2935 118 -2935 118 1 D$
rlabel pdiff -2955 68 -2955 68 1 D$
rlabel pdiff -2955 50 -2955 50 1 S$
rlabel pdiff -2955 204 -2955 204 1 D$
rlabel pdiff -2955 186 -2955 186 1 S$
rlabel pdiff -2955 340 -2955 340 1 D$
rlabel pdiff -2955 322 -2955 322 1 S$
rlabel pdiff -2955 476 -2955 476 1 D$
rlabel pdiff -2955 458 -2955 458 1 S$
rlabel pdiff -2955 612 -2955 612 1 D$
rlabel pdiff -2955 594 -2955 594 1 S$
rlabel pdiff -2955 748 -2955 748 1 D$
rlabel pdiff -2955 730 -2955 730 1 S$
rlabel pdiff -2955 884 -2955 884 1 D$
rlabel pdiff -2955 866 -2955 866 1 S$
rlabel pdiff -2955 1020 -2955 1020 1 D$
rlabel pdiff -2955 1002 -2955 1002 1 S$
rlabel pdiff -2955 1156 -2955 1156 1 D$
rlabel pdiff -2955 1138 -2955 1138 1 S$
rlabel pdiff -2955 1292 -2955 1292 1 D$
rlabel pdiff -2955 1274 -2955 1274 1 S$
rlabel ndiff -2565 -525 -2565 -525 1 S$
rlabel ndiff -2565 -510 -2565 -510 1 D$
rlabel ndiff -2565 -395 -2565 -395 1 S$
rlabel ndiff -2565 -380 -2565 -380 1 D$
rlabel ndiff -2565 -265 -2565 -265 1 S$
rlabel ndiff -2565 -250 -2565 -250 1 D$
rlabel ndiff -2565 -185 -2565 -185 1 S$
rlabel ndiff -2565 -200 -2565 -200 1 D$
rlabel ndiff -2565 -315 -2565 -315 1 S$
rlabel ndiff -2565 -330 -2565 -330 1 D$
rlabel ndiff -2565 -445 -2565 -445 1 S$
rlabel ndiff -2565 -460 -2565 -460 1 D$
<< end >>
