magic
tech sky130A
magscale 1 2
timestamp 1636480389
<< nwell >>
rect 1508 2690 7002 4058
<< pmoslvt >>
rect 1704 2910 1904 3910
rect 1962 2910 2162 3910
rect 2220 2910 2420 3910
rect 2478 2910 2678 3910
rect 2736 2910 2936 3910
rect 2994 2910 3194 3910
rect 3252 2910 3452 3910
rect 3510 2910 3710 3910
rect 3768 2910 3968 3910
rect 4026 2910 4226 3910
rect 4284 2910 4484 3910
rect 4542 2910 4742 3910
rect 4800 2910 5000 3910
rect 5058 2910 5258 3910
rect 5316 2910 5516 3910
rect 5574 2910 5774 3910
rect 5832 2910 6032 3910
rect 6090 2910 6290 3910
rect 6348 2910 6548 3910
rect 6606 2910 6806 3910
<< pdiff >>
rect 1646 3898 1704 3910
rect 1646 2922 1658 3898
rect 1692 2922 1704 3898
rect 1646 2910 1704 2922
rect 1904 3898 1962 3910
rect 1904 2922 1916 3898
rect 1950 2922 1962 3898
rect 1904 2910 1962 2922
rect 2162 3898 2220 3910
rect 2162 2922 2174 3898
rect 2208 2922 2220 3898
rect 2162 2910 2220 2922
rect 2420 3898 2478 3910
rect 2420 2922 2432 3898
rect 2466 2922 2478 3898
rect 2420 2910 2478 2922
rect 2678 3898 2736 3910
rect 2678 2922 2690 3898
rect 2724 2922 2736 3898
rect 2678 2910 2736 2922
rect 2936 3898 2994 3910
rect 2936 2922 2948 3898
rect 2982 2922 2994 3898
rect 2936 2910 2994 2922
rect 3194 3898 3252 3910
rect 3194 2922 3206 3898
rect 3240 2922 3252 3898
rect 3194 2910 3252 2922
rect 3452 3898 3510 3910
rect 3452 2922 3464 3898
rect 3498 2922 3510 3898
rect 3452 2910 3510 2922
rect 3710 3898 3768 3910
rect 3710 2922 3722 3898
rect 3756 2922 3768 3898
rect 3710 2910 3768 2922
rect 3968 3898 4026 3910
rect 3968 2922 3980 3898
rect 4014 2922 4026 3898
rect 3968 2910 4026 2922
rect 4226 3898 4284 3910
rect 4226 2922 4238 3898
rect 4272 2922 4284 3898
rect 4226 2910 4284 2922
rect 4484 3898 4542 3910
rect 4484 2922 4496 3898
rect 4530 2922 4542 3898
rect 4484 2910 4542 2922
rect 4742 3898 4800 3910
rect 4742 2922 4754 3898
rect 4788 2922 4800 3898
rect 4742 2910 4800 2922
rect 5000 3898 5058 3910
rect 5000 2922 5012 3898
rect 5046 2922 5058 3898
rect 5000 2910 5058 2922
rect 5258 3898 5316 3910
rect 5258 2922 5270 3898
rect 5304 2922 5316 3898
rect 5258 2910 5316 2922
rect 5516 3898 5574 3910
rect 5516 2922 5528 3898
rect 5562 2922 5574 3898
rect 5516 2910 5574 2922
rect 5774 3898 5832 3910
rect 5774 2922 5786 3898
rect 5820 2922 5832 3898
rect 5774 2910 5832 2922
rect 6032 3898 6090 3910
rect 6032 2922 6044 3898
rect 6078 2922 6090 3898
rect 6032 2910 6090 2922
rect 6290 3898 6348 3910
rect 6290 2922 6302 3898
rect 6336 2922 6348 3898
rect 6290 2910 6348 2922
rect 6548 3898 6606 3910
rect 6548 2922 6560 3898
rect 6594 2922 6606 3898
rect 6548 2910 6606 2922
rect 6806 3898 6864 3910
rect 6806 2922 6818 3898
rect 6852 2922 6864 3898
rect 6806 2910 6864 2922
<< pdiffc >>
rect 1658 2922 1692 3898
rect 1916 2922 1950 3898
rect 2174 2922 2208 3898
rect 2432 2922 2466 3898
rect 2690 2922 2724 3898
rect 2948 2922 2982 3898
rect 3206 2922 3240 3898
rect 3464 2922 3498 3898
rect 3722 2922 3756 3898
rect 3980 2922 4014 3898
rect 4238 2922 4272 3898
rect 4496 2922 4530 3898
rect 4754 2922 4788 3898
rect 5012 2922 5046 3898
rect 5270 2922 5304 3898
rect 5528 2922 5562 3898
rect 5786 2922 5820 3898
rect 6044 2922 6078 3898
rect 6302 2922 6336 3898
rect 6560 2922 6594 3898
rect 6818 2922 6852 3898
<< nsubdiff >>
rect 1544 3988 1640 4022
rect 6870 3988 6966 4022
rect 1544 3925 1578 3988
rect 6932 3925 6966 3988
rect 1544 2760 1578 2823
rect 6932 2760 6966 2823
rect 1544 2726 1640 2760
rect 6870 2726 6966 2760
<< nsubdiffcont >>
rect 1640 3988 6870 4022
rect 1544 2823 1578 3925
rect 6932 2823 6966 3925
rect 1640 2726 6870 2760
<< poly >>
rect 1704 3910 1904 3936
rect 1962 3910 2162 3936
rect 2220 3910 2420 3936
rect 2478 3910 2678 3936
rect 2736 3910 2936 3936
rect 2994 3910 3194 3936
rect 3252 3910 3452 3936
rect 3510 3910 3710 3936
rect 3768 3910 3968 3936
rect 4026 3910 4226 3936
rect 4284 3910 4484 3936
rect 4542 3910 4742 3936
rect 4800 3910 5000 3936
rect 5058 3910 5258 3936
rect 5316 3910 5516 3936
rect 5574 3910 5774 3936
rect 5832 3910 6032 3936
rect 6090 3910 6290 3936
rect 6348 3910 6548 3936
rect 6606 3910 6806 3936
rect 1704 2863 1904 2910
rect 1704 2829 1720 2863
rect 1888 2829 1904 2863
rect 1704 2813 1904 2829
rect 1962 2863 2162 2910
rect 1962 2829 1978 2863
rect 2146 2829 2162 2863
rect 1962 2813 2162 2829
rect 2220 2863 2420 2910
rect 2220 2829 2236 2863
rect 2404 2829 2420 2863
rect 2220 2813 2420 2829
rect 2478 2863 2678 2910
rect 2478 2829 2494 2863
rect 2662 2829 2678 2863
rect 2478 2813 2678 2829
rect 2736 2863 2936 2910
rect 2736 2829 2752 2863
rect 2920 2829 2936 2863
rect 2736 2813 2936 2829
rect 2994 2863 3194 2910
rect 2994 2829 3010 2863
rect 3178 2829 3194 2863
rect 2994 2813 3194 2829
rect 3252 2863 3452 2910
rect 3252 2829 3268 2863
rect 3436 2829 3452 2863
rect 3252 2813 3452 2829
rect 3510 2863 3710 2910
rect 3510 2829 3526 2863
rect 3694 2829 3710 2863
rect 3510 2813 3710 2829
rect 3768 2863 3968 2910
rect 3768 2829 3784 2863
rect 3952 2829 3968 2863
rect 3768 2813 3968 2829
rect 4026 2863 4226 2910
rect 4026 2829 4042 2863
rect 4210 2829 4226 2863
rect 4026 2813 4226 2829
rect 4284 2863 4484 2910
rect 4284 2829 4300 2863
rect 4468 2829 4484 2863
rect 4284 2813 4484 2829
rect 4542 2863 4742 2910
rect 4542 2829 4558 2863
rect 4726 2829 4742 2863
rect 4542 2813 4742 2829
rect 4800 2863 5000 2910
rect 4800 2829 4816 2863
rect 4984 2829 5000 2863
rect 4800 2813 5000 2829
rect 5058 2863 5258 2910
rect 5058 2829 5074 2863
rect 5242 2829 5258 2863
rect 5058 2813 5258 2829
rect 5316 2863 5516 2910
rect 5316 2829 5332 2863
rect 5500 2829 5516 2863
rect 5316 2813 5516 2829
rect 5574 2863 5774 2910
rect 5574 2829 5590 2863
rect 5758 2829 5774 2863
rect 5574 2813 5774 2829
rect 5832 2863 6032 2910
rect 5832 2829 5848 2863
rect 6016 2829 6032 2863
rect 5832 2813 6032 2829
rect 6090 2863 6290 2910
rect 6090 2829 6106 2863
rect 6274 2829 6290 2863
rect 6090 2813 6290 2829
rect 6348 2863 6548 2910
rect 6348 2829 6364 2863
rect 6532 2829 6548 2863
rect 6348 2813 6548 2829
rect 6606 2863 6806 2910
rect 6606 2829 6622 2863
rect 6790 2829 6806 2863
rect 6606 2813 6806 2829
<< polycont >>
rect 1720 2829 1888 2863
rect 1978 2829 2146 2863
rect 2236 2829 2404 2863
rect 2494 2829 2662 2863
rect 2752 2829 2920 2863
rect 3010 2829 3178 2863
rect 3268 2829 3436 2863
rect 3526 2829 3694 2863
rect 3784 2829 3952 2863
rect 4042 2829 4210 2863
rect 4300 2829 4468 2863
rect 4558 2829 4726 2863
rect 4816 2829 4984 2863
rect 5074 2829 5242 2863
rect 5332 2829 5500 2863
rect 5590 2829 5758 2863
rect 5848 2829 6016 2863
rect 6106 2829 6274 2863
rect 6364 2829 6532 2863
rect 6622 2829 6790 2863
<< locali >>
rect 1544 3925 1578 4022
rect 6932 3925 6966 4022
rect 1658 3898 1692 3914
rect 1658 2906 1692 2922
rect 1916 3898 1950 3914
rect 1916 2863 1950 2922
rect 2174 3898 2208 3914
rect 2174 2906 2208 2922
rect 2432 3898 2466 3914
rect 2432 2863 2466 2922
rect 2690 3898 2724 3914
rect 2690 2906 2724 2922
rect 2948 3898 2982 3914
rect 2948 2863 2982 2922
rect 3206 3898 3240 3914
rect 3206 2906 3240 2922
rect 3464 3898 3498 3914
rect 3464 2863 3498 2922
rect 3722 3898 3756 3914
rect 3722 2906 3756 2922
rect 3980 3898 4014 3914
rect 3980 2863 4014 2922
rect 4238 3898 4272 3914
rect 4238 2906 4272 2922
rect 4496 3898 4530 3914
rect 4496 2863 4530 2922
rect 4754 3898 4788 3914
rect 4754 2906 4788 2922
rect 5012 3898 5046 3914
rect 5012 2863 5046 2922
rect 5270 3898 5304 3914
rect 5270 2906 5304 2922
rect 5528 3898 5562 3914
rect 5528 2863 5562 2922
rect 5786 3898 5820 3914
rect 5786 2906 5820 2922
rect 6044 3898 6078 3914
rect 6044 2863 6078 2922
rect 6302 3898 6336 3914
rect 6302 2906 6336 2922
rect 6560 3898 6594 3914
rect 6560 2863 6594 2922
rect 6818 3898 6852 3914
rect 6818 2906 6852 2922
rect 1658 2829 1720 2863
rect 1888 2829 1978 2863
rect 2146 2829 2236 2863
rect 2404 2829 2494 2863
rect 2662 2829 2752 2863
rect 2920 2829 3010 2863
rect 3178 2829 3268 2863
rect 3436 2829 3526 2863
rect 3694 2829 3784 2863
rect 3952 2829 4042 2863
rect 4210 2829 4300 2863
rect 4468 2829 4558 2863
rect 4726 2829 4816 2863
rect 4984 2829 5074 2863
rect 5242 2829 5332 2863
rect 5500 2829 5590 2863
rect 5758 2829 5848 2863
rect 6016 2829 6106 2863
rect 6274 2829 6364 2863
rect 6532 2829 6622 2863
rect 6790 2829 6852 2863
rect 1544 2760 1578 2823
rect 6932 2760 6966 2823
rect 1544 2726 1640 2760
rect 6870 2726 6966 2760
<< viali >>
rect 1578 3988 1640 4022
rect 1640 3988 6870 4022
rect 6870 3988 6932 4022
rect 1544 2883 1578 3865
rect 1658 2922 1692 3898
rect 1916 2922 1950 3898
rect 2174 2922 2208 3898
rect 2432 2922 2466 3898
rect 2690 2922 2724 3898
rect 2948 2922 2982 3898
rect 3206 2922 3240 3898
rect 3464 2922 3498 3898
rect 3722 2922 3756 3898
rect 3980 2922 4014 3898
rect 4238 2922 4272 3898
rect 4496 2922 4530 3898
rect 4754 2922 4788 3898
rect 5012 2922 5046 3898
rect 5270 2922 5304 3898
rect 5528 2922 5562 3898
rect 5786 2922 5820 3898
rect 6044 2922 6078 3898
rect 6302 2922 6336 3898
rect 6560 2922 6594 3898
rect 6818 2922 6852 3898
rect 6932 2883 6966 3865
rect 1762 2829 1846 2863
rect 2020 2829 2104 2863
rect 2278 2829 2362 2863
rect 2536 2829 2620 2863
rect 2794 2829 2878 2863
rect 3052 2829 3136 2863
rect 3310 2829 3394 2863
rect 3568 2829 3652 2863
rect 3826 2829 3910 2863
rect 4084 2829 4168 2863
rect 4342 2829 4426 2863
rect 4600 2829 4684 2863
rect 4858 2829 4942 2863
rect 5116 2829 5200 2863
rect 5374 2829 5458 2863
rect 5632 2829 5716 2863
rect 5890 2829 5974 2863
rect 6148 2829 6232 2863
rect 6406 2829 6490 2863
rect 6664 2829 6748 2863
<< metal1 >>
rect 1538 4250 6972 4283
rect 1538 4170 1868 4250
rect 1948 4170 2028 4250
rect 2108 4170 2188 4250
rect 2268 4170 2348 4250
rect 2428 4170 2508 4250
rect 2588 4170 2668 4250
rect 2748 4170 2828 4250
rect 2908 4170 2988 4250
rect 3068 4170 3148 4250
rect 3228 4170 3308 4250
rect 3388 4170 3468 4250
rect 3548 4170 3628 4250
rect 3708 4170 3788 4250
rect 3868 4170 3948 4250
rect 4028 4170 4108 4250
rect 4188 4170 4268 4250
rect 4348 4170 4428 4250
rect 4508 4170 4588 4250
rect 4668 4170 4748 4250
rect 4828 4170 4908 4250
rect 4988 4170 5068 4250
rect 5148 4170 5228 4250
rect 5308 4170 5388 4250
rect 5468 4170 5548 4250
rect 5628 4170 5708 4250
rect 5788 4170 5868 4250
rect 5948 4170 6028 4250
rect 6108 4170 6188 4250
rect 6268 4170 6348 4250
rect 6428 4170 6508 4250
rect 6588 4170 6668 4250
rect 6748 4170 6972 4250
rect 1538 4090 6972 4170
rect 1538 4022 1868 4090
rect 1948 4022 2028 4090
rect 2108 4022 2188 4090
rect 2268 4022 2348 4090
rect 2428 4022 2508 4090
rect 2588 4022 2668 4090
rect 2748 4022 2828 4090
rect 2908 4022 2988 4090
rect 3068 4022 3148 4090
rect 3228 4022 3308 4090
rect 3388 4022 3468 4090
rect 3548 4022 3628 4090
rect 3708 4022 3788 4090
rect 3868 4022 3948 4090
rect 4028 4022 4108 4090
rect 4188 4022 4268 4090
rect 4348 4022 4428 4090
rect 4508 4022 4588 4090
rect 4668 4022 4748 4090
rect 4828 4022 4908 4090
rect 4988 4022 5068 4090
rect 5148 4022 5228 4090
rect 5308 4022 5388 4090
rect 5468 4022 5548 4090
rect 5628 4022 5708 4090
rect 5788 4022 5868 4090
rect 5948 4022 6028 4090
rect 6108 4022 6188 4090
rect 6268 4022 6348 4090
rect 6428 4022 6508 4090
rect 6588 4022 6668 4090
rect 6748 4022 6972 4090
rect 1538 3988 1578 4022
rect 6932 3988 6972 4022
rect 1538 3982 6972 3988
rect 1538 3865 1584 3982
rect 1538 2883 1544 3865
rect 1578 2883 1584 3865
rect 1538 2871 1584 2883
rect 1652 3898 1698 3910
rect 1652 2922 1658 3898
rect 1692 2922 1698 3898
rect 1652 2785 1698 2922
rect 1910 3898 1956 3982
rect 1910 2922 1916 3898
rect 1950 2922 1956 3898
rect 1910 2910 1956 2922
rect 2168 3898 2214 3910
rect 2168 2922 2174 3898
rect 2208 2922 2214 3898
rect 1750 2863 1858 2869
rect 1750 2829 1762 2863
rect 1846 2829 1858 2863
rect 1750 2823 1858 2829
rect 2008 2863 2116 2869
rect 2008 2829 2020 2863
rect 2104 2829 2116 2863
rect 2008 2823 2116 2829
rect 2168 2785 2214 2922
rect 2426 3898 2472 3982
rect 2426 2922 2432 3898
rect 2466 2922 2472 3898
rect 2426 2910 2472 2922
rect 2684 3898 2730 3910
rect 2684 2922 2690 3898
rect 2724 2922 2730 3898
rect 2266 2863 2374 2869
rect 2266 2829 2278 2863
rect 2362 2829 2374 2863
rect 2266 2823 2374 2829
rect 2524 2863 2632 2869
rect 2524 2829 2536 2863
rect 2620 2829 2632 2863
rect 2524 2823 2632 2829
rect 2684 2785 2730 2922
rect 2942 3898 2988 3982
rect 2942 2922 2948 3898
rect 2982 2922 2988 3898
rect 2942 2910 2988 2922
rect 3200 3898 3246 3910
rect 3200 2922 3206 3898
rect 3240 2922 3246 3898
rect 2782 2863 2890 2869
rect 2782 2829 2794 2863
rect 2878 2829 2890 2863
rect 2782 2823 2890 2829
rect 3040 2863 3148 2869
rect 3040 2829 3052 2863
rect 3136 2829 3148 2863
rect 3040 2823 3148 2829
rect 3200 2785 3246 2922
rect 3458 3898 3504 3982
rect 3458 2922 3464 3898
rect 3498 2922 3504 3898
rect 3458 2910 3504 2922
rect 3716 3898 3762 3910
rect 3716 2922 3722 3898
rect 3756 2922 3762 3898
rect 3298 2863 3406 2869
rect 3298 2829 3310 2863
rect 3394 2829 3406 2863
rect 3298 2823 3406 2829
rect 3556 2863 3664 2869
rect 3556 2829 3568 2863
rect 3652 2829 3664 2863
rect 3556 2823 3664 2829
rect 3716 2785 3762 2922
rect 3974 3898 4020 3982
rect 3974 2922 3980 3898
rect 4014 2922 4020 3898
rect 3974 2910 4020 2922
rect 4232 3898 4278 3910
rect 4232 2922 4238 3898
rect 4272 2922 4278 3898
rect 3814 2863 3922 2869
rect 3814 2829 3826 2863
rect 3910 2829 3922 2863
rect 3814 2823 3922 2829
rect 4072 2863 4180 2869
rect 4072 2829 4084 2863
rect 4168 2829 4180 2863
rect 4072 2823 4180 2829
rect 4232 2785 4278 2922
rect 4490 3898 4536 3982
rect 4490 2922 4496 3898
rect 4530 2922 4536 3898
rect 4490 2910 4536 2922
rect 4748 3898 4794 3910
rect 4748 2922 4754 3898
rect 4788 2922 4794 3898
rect 4330 2863 4438 2869
rect 4330 2829 4342 2863
rect 4426 2829 4438 2863
rect 4330 2823 4438 2829
rect 4588 2863 4696 2869
rect 4588 2829 4600 2863
rect 4684 2829 4696 2863
rect 4588 2823 4696 2829
rect 4748 2785 4794 2922
rect 5006 3898 5052 3982
rect 5006 2922 5012 3898
rect 5046 2922 5052 3898
rect 5006 2910 5052 2922
rect 5264 3898 5310 3910
rect 5264 2922 5270 3898
rect 5304 2922 5310 3898
rect 4846 2863 4954 2869
rect 4846 2829 4858 2863
rect 4942 2829 4954 2863
rect 4846 2823 4954 2829
rect 5104 2863 5212 2869
rect 5104 2829 5116 2863
rect 5200 2829 5212 2863
rect 5104 2823 5212 2829
rect 5264 2785 5310 2922
rect 5522 3898 5568 3982
rect 5522 2922 5528 3898
rect 5562 2922 5568 3898
rect 5522 2910 5568 2922
rect 5780 3898 5826 3910
rect 5780 2922 5786 3898
rect 5820 2922 5826 3898
rect 5362 2863 5470 2869
rect 5362 2829 5374 2863
rect 5458 2829 5470 2863
rect 5362 2823 5470 2829
rect 5620 2863 5728 2869
rect 5620 2829 5632 2863
rect 5716 2829 5728 2863
rect 5620 2823 5728 2829
rect 5780 2785 5826 2922
rect 6038 3898 6084 3982
rect 6038 2922 6044 3898
rect 6078 2922 6084 3898
rect 6038 2910 6084 2922
rect 6296 3898 6342 3910
rect 6296 2922 6302 3898
rect 6336 2922 6342 3898
rect 5878 2863 5986 2869
rect 5878 2829 5890 2863
rect 5974 2829 5986 2863
rect 5878 2823 5986 2829
rect 6136 2863 6244 2869
rect 6136 2829 6148 2863
rect 6232 2829 6244 2863
rect 6136 2823 6244 2829
rect 6296 2785 6342 2922
rect 6554 3898 6600 3982
rect 6554 2922 6560 3898
rect 6594 2922 6600 3898
rect 6554 2910 6600 2922
rect 6812 3898 6858 3910
rect 6812 2922 6818 3898
rect 6852 2922 6858 3898
rect 6394 2863 6502 2869
rect 6394 2829 6406 2863
rect 6490 2829 6502 2863
rect 6394 2823 6502 2829
rect 6652 2863 6760 2869
rect 6652 2829 6664 2863
rect 6748 2829 6760 2863
rect 6652 2823 6760 2829
rect 6812 2785 6858 2922
rect 6926 3865 6972 3982
rect 6926 2883 6932 3865
rect 6966 2883 6972 3865
rect 6926 2871 6972 2883
rect 1508 2729 7002 2785
rect 1508 2669 1610 2729
rect 1670 2669 1730 2729
rect 1790 2669 1850 2729
rect 1910 2669 1970 2729
rect 2030 2669 2090 2729
rect 2150 2669 2210 2729
rect 2270 2669 2330 2729
rect 2390 2669 2450 2729
rect 2510 2669 2570 2729
rect 2630 2669 2690 2729
rect 2750 2669 2810 2729
rect 2870 2669 2930 2729
rect 2990 2669 3050 2729
rect 3110 2669 3170 2729
rect 3230 2669 3290 2729
rect 3350 2669 3410 2729
rect 3470 2669 3530 2729
rect 3590 2669 3650 2729
rect 3710 2669 3770 2729
rect 3830 2669 3890 2729
rect 3950 2669 4010 2729
rect 4070 2669 4130 2729
rect 4190 2669 4250 2729
rect 4310 2669 4370 2729
rect 4430 2669 4490 2729
rect 4550 2669 4610 2729
rect 4670 2669 4730 2729
rect 4790 2669 4850 2729
rect 4910 2669 4970 2729
rect 5030 2669 5090 2729
rect 5150 2669 5210 2729
rect 5270 2669 5330 2729
rect 5390 2669 5450 2729
rect 5510 2669 5570 2729
rect 5630 2669 5690 2729
rect 5750 2669 5810 2729
rect 5870 2669 5930 2729
rect 5990 2669 6050 2729
rect 6110 2669 6170 2729
rect 6230 2669 6290 2729
rect 6350 2669 6410 2729
rect 6470 2669 6530 2729
rect 6590 2669 6650 2729
rect 6710 2669 6770 2729
rect 6830 2669 6890 2729
rect 6950 2669 7002 2729
rect 1508 2609 7002 2669
rect 1508 2549 1610 2609
rect 1670 2549 1730 2609
rect 1790 2549 1850 2609
rect 1910 2549 1970 2609
rect 2030 2549 2090 2609
rect 2150 2549 2210 2609
rect 2270 2549 2330 2609
rect 2390 2549 2450 2609
rect 2510 2549 2570 2609
rect 2630 2549 2690 2609
rect 2750 2549 2810 2609
rect 2870 2549 2930 2609
rect 2990 2549 3050 2609
rect 3110 2549 3170 2609
rect 3230 2549 3290 2609
rect 3350 2549 3410 2609
rect 3470 2549 3530 2609
rect 3590 2549 3650 2609
rect 3710 2549 3770 2609
rect 3830 2549 3890 2609
rect 3950 2549 4010 2609
rect 4070 2549 4130 2609
rect 4190 2549 4250 2609
rect 4310 2549 4370 2609
rect 4430 2549 4490 2609
rect 4550 2549 4610 2609
rect 4670 2549 4730 2609
rect 4790 2549 4850 2609
rect 4910 2549 4970 2609
rect 5030 2549 5090 2609
rect 5150 2549 5210 2609
rect 5270 2549 5330 2609
rect 5390 2549 5450 2609
rect 5510 2549 5570 2609
rect 5630 2549 5690 2609
rect 5750 2549 5810 2609
rect 5870 2549 5930 2609
rect 5990 2549 6050 2609
rect 6110 2549 6170 2609
rect 6230 2549 6290 2609
rect 6350 2549 6410 2609
rect 6470 2549 6530 2609
rect 6590 2549 6650 2609
rect 6710 2549 6770 2609
rect 6830 2549 6890 2609
rect 6950 2549 7002 2609
rect 1508 2510 7002 2549
<< via1 >>
rect 1868 4170 1948 4250
rect 2028 4170 2108 4250
rect 2188 4170 2268 4250
rect 2348 4170 2428 4250
rect 2508 4170 2588 4250
rect 2668 4170 2748 4250
rect 2828 4170 2908 4250
rect 2988 4170 3068 4250
rect 3148 4170 3228 4250
rect 3308 4170 3388 4250
rect 3468 4170 3548 4250
rect 3628 4170 3708 4250
rect 3788 4170 3868 4250
rect 3948 4170 4028 4250
rect 4108 4170 4188 4250
rect 4268 4170 4348 4250
rect 4428 4170 4508 4250
rect 4588 4170 4668 4250
rect 4748 4170 4828 4250
rect 4908 4170 4988 4250
rect 5068 4170 5148 4250
rect 5228 4170 5308 4250
rect 5388 4170 5468 4250
rect 5548 4170 5628 4250
rect 5708 4170 5788 4250
rect 5868 4170 5948 4250
rect 6028 4170 6108 4250
rect 6188 4170 6268 4250
rect 6348 4170 6428 4250
rect 6508 4170 6588 4250
rect 6668 4170 6748 4250
rect 1868 4022 1948 4090
rect 2028 4022 2108 4090
rect 2188 4022 2268 4090
rect 2348 4022 2428 4090
rect 2508 4022 2588 4090
rect 2668 4022 2748 4090
rect 2828 4022 2908 4090
rect 2988 4022 3068 4090
rect 3148 4022 3228 4090
rect 3308 4022 3388 4090
rect 3468 4022 3548 4090
rect 3628 4022 3708 4090
rect 3788 4022 3868 4090
rect 3948 4022 4028 4090
rect 4108 4022 4188 4090
rect 4268 4022 4348 4090
rect 4428 4022 4508 4090
rect 4588 4022 4668 4090
rect 4748 4022 4828 4090
rect 4908 4022 4988 4090
rect 5068 4022 5148 4090
rect 5228 4022 5308 4090
rect 5388 4022 5468 4090
rect 5548 4022 5628 4090
rect 5708 4022 5788 4090
rect 5868 4022 5948 4090
rect 6028 4022 6108 4090
rect 6188 4022 6268 4090
rect 6348 4022 6428 4090
rect 6508 4022 6588 4090
rect 6668 4022 6748 4090
rect 1868 4010 1948 4022
rect 2028 4010 2108 4022
rect 2188 4010 2268 4022
rect 2348 4010 2428 4022
rect 2508 4010 2588 4022
rect 2668 4010 2748 4022
rect 2828 4010 2908 4022
rect 2988 4010 3068 4022
rect 3148 4010 3228 4022
rect 3308 4010 3388 4022
rect 3468 4010 3548 4022
rect 3628 4010 3708 4022
rect 3788 4010 3868 4022
rect 3948 4010 4028 4022
rect 4108 4010 4188 4022
rect 4268 4010 4348 4022
rect 4428 4010 4508 4022
rect 4588 4010 4668 4022
rect 4748 4010 4828 4022
rect 4908 4010 4988 4022
rect 5068 4010 5148 4022
rect 5228 4010 5308 4022
rect 5388 4010 5468 4022
rect 5548 4010 5628 4022
rect 5708 4010 5788 4022
rect 5868 4010 5948 4022
rect 6028 4010 6108 4022
rect 6188 4010 6268 4022
rect 6348 4010 6428 4022
rect 6508 4010 6588 4022
rect 6668 4010 6748 4022
rect 1610 2669 1670 2729
rect 1730 2669 1790 2729
rect 1850 2669 1910 2729
rect 1970 2669 2030 2729
rect 2090 2669 2150 2729
rect 2210 2669 2270 2729
rect 2330 2669 2390 2729
rect 2450 2669 2510 2729
rect 2570 2669 2630 2729
rect 2690 2669 2750 2729
rect 2810 2669 2870 2729
rect 2930 2669 2990 2729
rect 3050 2669 3110 2729
rect 3170 2669 3230 2729
rect 3290 2669 3350 2729
rect 3410 2669 3470 2729
rect 3530 2669 3590 2729
rect 3650 2669 3710 2729
rect 3770 2669 3830 2729
rect 3890 2669 3950 2729
rect 4010 2669 4070 2729
rect 4130 2669 4190 2729
rect 4250 2669 4310 2729
rect 4370 2669 4430 2729
rect 4490 2669 4550 2729
rect 4610 2669 4670 2729
rect 4730 2669 4790 2729
rect 4850 2669 4910 2729
rect 4970 2669 5030 2729
rect 5090 2669 5150 2729
rect 5210 2669 5270 2729
rect 5330 2669 5390 2729
rect 5450 2669 5510 2729
rect 5570 2669 5630 2729
rect 5690 2669 5750 2729
rect 5810 2669 5870 2729
rect 5930 2669 5990 2729
rect 6050 2669 6110 2729
rect 6170 2669 6230 2729
rect 6290 2669 6350 2729
rect 6410 2669 6470 2729
rect 6530 2669 6590 2729
rect 6650 2669 6710 2729
rect 6770 2669 6830 2729
rect 6890 2669 6950 2729
rect 1610 2549 1670 2609
rect 1730 2549 1790 2609
rect 1850 2549 1910 2609
rect 1970 2549 2030 2609
rect 2090 2549 2150 2609
rect 2210 2549 2270 2609
rect 2330 2549 2390 2609
rect 2450 2549 2510 2609
rect 2570 2549 2630 2609
rect 2690 2549 2750 2609
rect 2810 2549 2870 2609
rect 2930 2549 2990 2609
rect 3050 2549 3110 2609
rect 3170 2549 3230 2609
rect 3290 2549 3350 2609
rect 3410 2549 3470 2609
rect 3530 2549 3590 2609
rect 3650 2549 3710 2609
rect 3770 2549 3830 2609
rect 3890 2549 3950 2609
rect 4010 2549 4070 2609
rect 4130 2549 4190 2609
rect 4250 2549 4310 2609
rect 4370 2549 4430 2609
rect 4490 2549 4550 2609
rect 4610 2549 4670 2609
rect 4730 2549 4790 2609
rect 4850 2549 4910 2609
rect 4970 2549 5030 2609
rect 5090 2549 5150 2609
rect 5210 2549 5270 2609
rect 5330 2549 5390 2609
rect 5450 2549 5510 2609
rect 5570 2549 5630 2609
rect 5690 2549 5750 2609
rect 5810 2549 5870 2609
rect 5930 2549 5990 2609
rect 6050 2549 6110 2609
rect 6170 2549 6230 2609
rect 6290 2549 6350 2609
rect 6410 2549 6470 2609
rect 6530 2549 6590 2609
rect 6650 2549 6710 2609
rect 6770 2549 6830 2609
rect 6890 2549 6950 2609
<< metal2 >>
rect 1768 4250 6868 4330
rect 1768 4170 1868 4250
rect 1948 4170 2028 4250
rect 2108 4170 2188 4250
rect 2268 4170 2348 4250
rect 2428 4170 2508 4250
rect 2588 4170 2668 4250
rect 2748 4170 2828 4250
rect 2908 4170 2988 4250
rect 3068 4170 3148 4250
rect 3228 4170 3308 4250
rect 3388 4170 3468 4250
rect 3548 4170 3628 4250
rect 3708 4170 3788 4250
rect 3868 4170 3948 4250
rect 4028 4170 4108 4250
rect 4188 4170 4268 4250
rect 4348 4170 4428 4250
rect 4508 4170 4588 4250
rect 4668 4170 4748 4250
rect 4828 4170 4908 4250
rect 4988 4170 5068 4250
rect 5148 4170 5228 4250
rect 5308 4170 5388 4250
rect 5468 4170 5548 4250
rect 5628 4170 5708 4250
rect 5788 4170 5868 4250
rect 5948 4170 6028 4250
rect 6108 4170 6188 4250
rect 6268 4170 6348 4250
rect 6428 4170 6508 4250
rect 6588 4170 6668 4250
rect 6748 4170 6868 4250
rect 1768 4090 6868 4170
rect 1768 4010 1868 4090
rect 1948 4010 2028 4090
rect 2108 4010 2188 4090
rect 2268 4010 2348 4090
rect 2428 4010 2508 4090
rect 2588 4010 2668 4090
rect 2748 4010 2828 4090
rect 2908 4010 2988 4090
rect 3068 4010 3148 4090
rect 3228 4010 3308 4090
rect 3388 4010 3468 4090
rect 3548 4010 3628 4090
rect 3708 4010 3788 4090
rect 3868 4010 3948 4090
rect 4028 4010 4108 4090
rect 4188 4010 4268 4090
rect 4348 4010 4428 4090
rect 4508 4010 4588 4090
rect 4668 4010 4748 4090
rect 4828 4010 4908 4090
rect 4988 4010 5068 4090
rect 5148 4010 5228 4090
rect 5308 4010 5388 4090
rect 5468 4010 5548 4090
rect 5628 4010 5708 4090
rect 5788 4010 5868 4090
rect 5948 4010 6028 4090
rect 6108 4010 6188 4090
rect 6268 4010 6348 4090
rect 6428 4010 6508 4090
rect 6588 4010 6668 4090
rect 6748 4010 6868 4090
rect 1768 3970 6868 4010
rect 1490 2729 7010 2789
rect 1490 2669 1610 2729
rect 1670 2669 1730 2729
rect 1790 2669 1850 2729
rect 1910 2669 1970 2729
rect 2030 2669 2090 2729
rect 2150 2669 2210 2729
rect 2270 2669 2330 2729
rect 2390 2669 2450 2729
rect 2510 2669 2570 2729
rect 2630 2669 2690 2729
rect 2750 2669 2810 2729
rect 2870 2669 2930 2729
rect 2990 2669 3050 2729
rect 3110 2669 3170 2729
rect 3230 2669 3290 2729
rect 3350 2669 3410 2729
rect 3470 2669 3530 2729
rect 3590 2669 3650 2729
rect 3710 2669 3770 2729
rect 3830 2669 3890 2729
rect 3950 2669 4010 2729
rect 4070 2669 4130 2729
rect 4190 2669 4250 2729
rect 4310 2669 4370 2729
rect 4430 2669 4490 2729
rect 4550 2669 4610 2729
rect 4670 2669 4730 2729
rect 4790 2669 4850 2729
rect 4910 2669 4970 2729
rect 5030 2669 5090 2729
rect 5150 2669 5210 2729
rect 5270 2669 5330 2729
rect 5390 2669 5450 2729
rect 5510 2669 5570 2729
rect 5630 2669 5690 2729
rect 5750 2669 5810 2729
rect 5870 2669 5930 2729
rect 5990 2669 6050 2729
rect 6110 2669 6170 2729
rect 6230 2669 6290 2729
rect 6350 2669 6410 2729
rect 6470 2669 6530 2729
rect 6590 2669 6650 2729
rect 6710 2669 6770 2729
rect 6830 2669 6890 2729
rect 6950 2669 7010 2729
rect 1490 2609 7010 2669
rect 1490 2549 1610 2609
rect 1670 2549 1730 2609
rect 1790 2549 1850 2609
rect 1910 2549 1970 2609
rect 2030 2549 2090 2609
rect 2150 2549 2210 2609
rect 2270 2549 2330 2609
rect 2390 2549 2450 2609
rect 2510 2549 2570 2609
rect 2630 2549 2690 2609
rect 2750 2549 2810 2609
rect 2870 2549 2930 2609
rect 2990 2549 3050 2609
rect 3110 2549 3170 2609
rect 3230 2549 3290 2609
rect 3350 2549 3410 2609
rect 3470 2549 3530 2609
rect 3590 2549 3650 2609
rect 3710 2549 3770 2609
rect 3830 2549 3890 2609
rect 3950 2549 4010 2609
rect 4070 2549 4130 2609
rect 4190 2549 4250 2609
rect 4310 2549 4370 2609
rect 4430 2549 4490 2609
rect 4550 2549 4610 2609
rect 4670 2549 4730 2609
rect 4790 2549 4850 2609
rect 4910 2549 4970 2609
rect 5030 2549 5090 2609
rect 5150 2549 5210 2609
rect 5270 2549 5330 2609
rect 5390 2549 5450 2609
rect 5510 2549 5570 2609
rect 5630 2549 5690 2609
rect 5750 2549 5810 2609
rect 5870 2549 5930 2609
rect 5990 2549 6050 2609
rect 6110 2549 6170 2609
rect 6230 2549 6290 2609
rect 6350 2549 6410 2609
rect 6470 2549 6530 2609
rect 6590 2549 6650 2609
rect 6710 2549 6770 2609
rect 6830 2549 6890 2609
rect 6950 2549 7010 2609
rect 1490 2489 7010 2549
<< via2 >>
rect 1868 4170 1948 4250
rect 2028 4170 2108 4250
rect 2188 4170 2268 4250
rect 2348 4170 2428 4250
rect 2508 4170 2588 4250
rect 2668 4170 2748 4250
rect 2828 4170 2908 4250
rect 2988 4170 3068 4250
rect 3148 4170 3228 4250
rect 3308 4170 3388 4250
rect 3468 4170 3548 4250
rect 3628 4170 3708 4250
rect 3788 4170 3868 4250
rect 3948 4170 4028 4250
rect 4108 4170 4188 4250
rect 4268 4170 4348 4250
rect 4428 4170 4508 4250
rect 4588 4170 4668 4250
rect 4748 4170 4828 4250
rect 4908 4170 4988 4250
rect 5068 4170 5148 4250
rect 5228 4170 5308 4250
rect 5388 4170 5468 4250
rect 5548 4170 5628 4250
rect 5708 4170 5788 4250
rect 5868 4170 5948 4250
rect 6028 4170 6108 4250
rect 6188 4170 6268 4250
rect 6348 4170 6428 4250
rect 6508 4170 6588 4250
rect 6668 4170 6748 4250
rect 1868 4010 1948 4090
rect 2028 4010 2108 4090
rect 2188 4010 2268 4090
rect 2348 4010 2428 4090
rect 2508 4010 2588 4090
rect 2668 4010 2748 4090
rect 2828 4010 2908 4090
rect 2988 4010 3068 4090
rect 3148 4010 3228 4090
rect 3308 4010 3388 4090
rect 3468 4010 3548 4090
rect 3628 4010 3708 4090
rect 3788 4010 3868 4090
rect 3948 4010 4028 4090
rect 4108 4010 4188 4090
rect 4268 4010 4348 4090
rect 4428 4010 4508 4090
rect 4588 4010 4668 4090
rect 4748 4010 4828 4090
rect 4908 4010 4988 4090
rect 5068 4010 5148 4090
rect 5228 4010 5308 4090
rect 5388 4010 5468 4090
rect 5548 4010 5628 4090
rect 5708 4010 5788 4090
rect 5868 4010 5948 4090
rect 6028 4010 6108 4090
rect 6188 4010 6268 4090
rect 6348 4010 6428 4090
rect 6508 4010 6588 4090
rect 6668 4010 6748 4090
rect 1610 2669 1670 2729
rect 1730 2669 1790 2729
rect 1850 2669 1910 2729
rect 1970 2669 2030 2729
rect 2090 2669 2150 2729
rect 2210 2669 2270 2729
rect 2330 2669 2390 2729
rect 2450 2669 2510 2729
rect 2570 2669 2630 2729
rect 2690 2669 2750 2729
rect 2810 2669 2870 2729
rect 2930 2669 2990 2729
rect 3050 2669 3110 2729
rect 3170 2669 3230 2729
rect 3290 2669 3350 2729
rect 3410 2669 3470 2729
rect 3530 2669 3590 2729
rect 3650 2669 3710 2729
rect 3770 2669 3830 2729
rect 3890 2669 3950 2729
rect 4010 2669 4070 2729
rect 4130 2669 4190 2729
rect 4250 2669 4310 2729
rect 4370 2669 4430 2729
rect 4490 2669 4550 2729
rect 4610 2669 4670 2729
rect 4730 2669 4790 2729
rect 4850 2669 4910 2729
rect 4970 2669 5030 2729
rect 5090 2669 5150 2729
rect 5210 2669 5270 2729
rect 5330 2669 5390 2729
rect 5450 2669 5510 2729
rect 5570 2669 5630 2729
rect 5690 2669 5750 2729
rect 5810 2669 5870 2729
rect 5930 2669 5990 2729
rect 6050 2669 6110 2729
rect 6170 2669 6230 2729
rect 6290 2669 6350 2729
rect 6410 2669 6470 2729
rect 6530 2669 6590 2729
rect 6650 2669 6710 2729
rect 6770 2669 6830 2729
rect 6890 2669 6950 2729
rect 1610 2549 1670 2609
rect 1730 2549 1790 2609
rect 1850 2549 1910 2609
rect 1970 2549 2030 2609
rect 2090 2549 2150 2609
rect 2210 2549 2270 2609
rect 2330 2549 2390 2609
rect 2450 2549 2510 2609
rect 2570 2549 2630 2609
rect 2690 2549 2750 2609
rect 2810 2549 2870 2609
rect 2930 2549 2990 2609
rect 3050 2549 3110 2609
rect 3170 2549 3230 2609
rect 3290 2549 3350 2609
rect 3410 2549 3470 2609
rect 3530 2549 3590 2609
rect 3650 2549 3710 2609
rect 3770 2549 3830 2609
rect 3890 2549 3950 2609
rect 4010 2549 4070 2609
rect 4130 2549 4190 2609
rect 4250 2549 4310 2609
rect 4370 2549 4430 2609
rect 4490 2549 4550 2609
rect 4610 2549 4670 2609
rect 4730 2549 4790 2609
rect 4850 2549 4910 2609
rect 4970 2549 5030 2609
rect 5090 2549 5150 2609
rect 5210 2549 5270 2609
rect 5330 2549 5390 2609
rect 5450 2549 5510 2609
rect 5570 2549 5630 2609
rect 5690 2549 5750 2609
rect 5810 2549 5870 2609
rect 5930 2549 5990 2609
rect 6050 2549 6110 2609
rect 6170 2549 6230 2609
rect 6290 2549 6350 2609
rect 6410 2549 6470 2609
rect 6530 2549 6590 2609
rect 6650 2549 6710 2609
rect 6770 2549 6830 2609
rect 6890 2549 6950 2609
<< metal3 >>
rect 1768 4250 6868 4330
rect 1768 4170 1868 4250
rect 1948 4170 2028 4250
rect 2108 4170 2188 4250
rect 2268 4170 2348 4250
rect 2428 4170 2508 4250
rect 2588 4170 2668 4250
rect 2748 4170 2828 4250
rect 2908 4170 2988 4250
rect 3068 4170 3148 4250
rect 3228 4170 3308 4250
rect 3388 4170 3468 4250
rect 3548 4170 3628 4250
rect 3708 4170 3788 4250
rect 3868 4170 3948 4250
rect 4028 4170 4108 4250
rect 4188 4170 4268 4250
rect 4348 4170 4428 4250
rect 4508 4170 4588 4250
rect 4668 4170 4748 4250
rect 4828 4170 4908 4250
rect 4988 4170 5068 4250
rect 5148 4170 5228 4250
rect 5308 4170 5388 4250
rect 5468 4170 5548 4250
rect 5628 4170 5708 4250
rect 5788 4170 5868 4250
rect 5948 4170 6028 4250
rect 6108 4170 6188 4250
rect 6268 4170 6348 4250
rect 6428 4170 6508 4250
rect 6588 4170 6668 4250
rect 6748 4170 6868 4250
rect 1768 4090 6868 4170
rect 1768 4010 1868 4090
rect 1948 4010 2028 4090
rect 2108 4010 2188 4090
rect 2268 4010 2348 4090
rect 2428 4010 2508 4090
rect 2588 4010 2668 4090
rect 2748 4010 2828 4090
rect 2908 4010 2988 4090
rect 3068 4010 3148 4090
rect 3228 4010 3308 4090
rect 3388 4010 3468 4090
rect 3548 4010 3628 4090
rect 3708 4010 3788 4090
rect 3868 4010 3948 4090
rect 4028 4010 4108 4090
rect 4188 4010 4268 4090
rect 4348 4010 4428 4090
rect 4508 4010 4588 4090
rect 4668 4010 4748 4090
rect 4828 4010 4908 4090
rect 4988 4010 5068 4090
rect 5148 4010 5228 4090
rect 5308 4010 5388 4090
rect 5468 4010 5548 4090
rect 5628 4010 5708 4090
rect 5788 4010 5868 4090
rect 5948 4010 6028 4090
rect 6108 4010 6188 4090
rect 6268 4010 6348 4090
rect 6428 4010 6508 4090
rect 6588 4010 6668 4090
rect 6748 4010 6868 4090
rect 1768 3970 6868 4010
rect 0 2729 8084 2966
rect 0 2669 1610 2729
rect 1670 2669 1730 2729
rect 1790 2669 1850 2729
rect 1910 2669 1970 2729
rect 2030 2669 2090 2729
rect 2150 2669 2210 2729
rect 2270 2669 2330 2729
rect 2390 2669 2450 2729
rect 2510 2669 2570 2729
rect 2630 2669 2690 2729
rect 2750 2669 2810 2729
rect 2870 2669 2930 2729
rect 2990 2669 3050 2729
rect 3110 2669 3170 2729
rect 3230 2669 3290 2729
rect 3350 2669 3410 2729
rect 3470 2669 3530 2729
rect 3590 2669 3650 2729
rect 3710 2669 3770 2729
rect 3830 2669 3890 2729
rect 3950 2669 4010 2729
rect 4070 2669 4130 2729
rect 4190 2669 4250 2729
rect 4310 2669 4370 2729
rect 4430 2669 4490 2729
rect 4550 2669 4610 2729
rect 4670 2669 4730 2729
rect 4790 2669 4850 2729
rect 4910 2669 4970 2729
rect 5030 2669 5090 2729
rect 5150 2669 5210 2729
rect 5270 2669 5330 2729
rect 5390 2669 5450 2729
rect 5510 2669 5570 2729
rect 5630 2669 5690 2729
rect 5750 2669 5810 2729
rect 5870 2669 5930 2729
rect 5990 2669 6050 2729
rect 6110 2669 6170 2729
rect 6230 2669 6290 2729
rect 6350 2669 6410 2729
rect 6470 2669 6530 2729
rect 6590 2669 6650 2729
rect 6710 2669 6770 2729
rect 6830 2669 6890 2729
rect 6950 2669 8084 2729
rect 0 2609 8084 2669
rect 0 2549 1610 2609
rect 1670 2549 1730 2609
rect 1790 2549 1850 2609
rect 1910 2549 1970 2609
rect 2030 2549 2090 2609
rect 2150 2549 2210 2609
rect 2270 2549 2330 2609
rect 2390 2549 2450 2609
rect 2510 2549 2570 2609
rect 2630 2549 2690 2609
rect 2750 2549 2810 2609
rect 2870 2549 2930 2609
rect 2990 2549 3050 2609
rect 3110 2549 3170 2609
rect 3230 2549 3290 2609
rect 3350 2549 3410 2609
rect 3470 2549 3530 2609
rect 3590 2549 3650 2609
rect 3710 2549 3770 2609
rect 3830 2549 3890 2609
rect 3950 2549 4010 2609
rect 4070 2549 4130 2609
rect 4190 2549 4250 2609
rect 4310 2549 4370 2609
rect 4430 2549 4490 2609
rect 4550 2549 4610 2609
rect 4670 2549 4730 2609
rect 4790 2549 4850 2609
rect 4910 2549 4970 2609
rect 5030 2549 5090 2609
rect 5150 2549 5210 2609
rect 5270 2549 5330 2609
rect 5390 2549 5450 2609
rect 5510 2549 5570 2609
rect 5630 2549 5690 2609
rect 5750 2549 5810 2609
rect 5870 2549 5930 2609
rect 5990 2549 6050 2609
rect 6110 2549 6170 2609
rect 6230 2549 6290 2609
rect 6350 2549 6410 2609
rect 6470 2549 6530 2609
rect 6590 2549 6650 2609
rect 6710 2549 6770 2609
rect 6830 2549 6890 2609
rect 6950 2549 8084 2609
rect 0 0 8084 2549
<< via3 >>
rect 1868 4170 1948 4250
rect 2028 4170 2108 4250
rect 2188 4170 2268 4250
rect 2348 4170 2428 4250
rect 2508 4170 2588 4250
rect 2668 4170 2748 4250
rect 2828 4170 2908 4250
rect 2988 4170 3068 4250
rect 3148 4170 3228 4250
rect 3308 4170 3388 4250
rect 3468 4170 3548 4250
rect 3628 4170 3708 4250
rect 3788 4170 3868 4250
rect 3948 4170 4028 4250
rect 4108 4170 4188 4250
rect 4268 4170 4348 4250
rect 4428 4170 4508 4250
rect 4588 4170 4668 4250
rect 4748 4170 4828 4250
rect 4908 4170 4988 4250
rect 5068 4170 5148 4250
rect 5228 4170 5308 4250
rect 5388 4170 5468 4250
rect 5548 4170 5628 4250
rect 5708 4170 5788 4250
rect 5868 4170 5948 4250
rect 6028 4170 6108 4250
rect 6188 4170 6268 4250
rect 6348 4170 6428 4250
rect 6508 4170 6588 4250
rect 6668 4170 6748 4250
rect 1868 4010 1948 4090
rect 2028 4010 2108 4090
rect 2188 4010 2268 4090
rect 2348 4010 2428 4090
rect 2508 4010 2588 4090
rect 2668 4010 2748 4090
rect 2828 4010 2908 4090
rect 2988 4010 3068 4090
rect 3148 4010 3228 4090
rect 3308 4010 3388 4090
rect 3468 4010 3548 4090
rect 3628 4010 3708 4090
rect 3788 4010 3868 4090
rect 3948 4010 4028 4090
rect 4108 4010 4188 4090
rect 4268 4010 4348 4090
rect 4428 4010 4508 4090
rect 4588 4010 4668 4090
rect 4748 4010 4828 4090
rect 4908 4010 4988 4090
rect 5068 4010 5148 4090
rect 5228 4010 5308 4090
rect 5388 4010 5468 4090
rect 5548 4010 5628 4090
rect 5708 4010 5788 4090
rect 5868 4010 5948 4090
rect 6028 4010 6108 4090
rect 6188 4010 6268 4090
rect 6348 4010 6428 4090
rect 6508 4010 6588 4090
rect 6668 4010 6748 4090
<< metal4 >>
rect 1768 4290 6868 4330
rect 1768 4250 2012 4290
rect 2248 4250 2484 4290
rect 2720 4250 2956 4290
rect 3192 4250 3428 4290
rect 3664 4250 3900 4290
rect 4136 4250 4372 4290
rect 4608 4250 4844 4290
rect 5080 4250 5316 4290
rect 5552 4250 5788 4290
rect 6024 4250 6260 4290
rect 6496 4250 6868 4290
rect 1768 4170 1868 4250
rect 1948 4170 2012 4250
rect 2268 4170 2348 4250
rect 2428 4170 2484 4250
rect 2748 4170 2828 4250
rect 2908 4170 2956 4250
rect 3228 4170 3308 4250
rect 3388 4170 3428 4250
rect 3708 4170 3788 4250
rect 3868 4170 3900 4250
rect 4188 4170 4268 4250
rect 4348 4170 4372 4250
rect 4668 4170 4748 4250
rect 4828 4170 4844 4250
rect 5148 4170 5228 4250
rect 5308 4170 5316 4250
rect 5628 4170 5708 4250
rect 6024 4170 6028 4250
rect 6108 4170 6188 4250
rect 6496 4170 6508 4250
rect 6588 4170 6668 4250
rect 6748 4170 6868 4250
rect 1768 4090 2012 4170
rect 2248 4090 2484 4170
rect 2720 4090 2956 4170
rect 3192 4090 3428 4170
rect 3664 4090 3900 4170
rect 4136 4090 4372 4170
rect 4608 4090 4844 4170
rect 5080 4090 5316 4170
rect 5552 4090 5788 4170
rect 6024 4090 6260 4170
rect 6496 4090 6868 4170
rect 1768 4010 1868 4090
rect 1948 4054 2012 4090
rect 1948 4010 2028 4054
rect 2108 4010 2188 4054
rect 2268 4010 2348 4090
rect 2428 4054 2484 4090
rect 2428 4010 2508 4054
rect 2588 4010 2668 4054
rect 2748 4010 2828 4090
rect 2908 4054 2956 4090
rect 2908 4010 2988 4054
rect 3068 4010 3148 4054
rect 3228 4010 3308 4090
rect 3388 4054 3428 4090
rect 3388 4010 3468 4054
rect 3548 4010 3628 4054
rect 3708 4010 3788 4090
rect 3868 4054 3900 4090
rect 3868 4010 3948 4054
rect 4028 4010 4108 4054
rect 4188 4010 4268 4090
rect 4348 4054 4372 4090
rect 4348 4010 4428 4054
rect 4508 4010 4588 4054
rect 4668 4010 4748 4090
rect 4828 4054 4844 4090
rect 4828 4010 4908 4054
rect 4988 4010 5068 4054
rect 5148 4010 5228 4090
rect 5308 4054 5316 4090
rect 5308 4010 5388 4054
rect 5468 4010 5548 4054
rect 5628 4010 5708 4090
rect 6024 4054 6028 4090
rect 5788 4010 5868 4054
rect 5948 4010 6028 4054
rect 6108 4010 6188 4090
rect 6496 4054 6508 4090
rect 6268 4010 6348 4054
rect 6428 4010 6508 4054
rect 6588 4010 6668 4090
rect 6748 4010 6868 4090
rect 1768 3970 6868 4010
<< via4 >>
rect 2012 4250 2248 4290
rect 2484 4250 2720 4290
rect 2956 4250 3192 4290
rect 3428 4250 3664 4290
rect 3900 4250 4136 4290
rect 4372 4250 4608 4290
rect 4844 4250 5080 4290
rect 5316 4250 5552 4290
rect 5788 4250 6024 4290
rect 6260 4250 6496 4290
rect 2012 4170 2028 4250
rect 2028 4170 2108 4250
rect 2108 4170 2188 4250
rect 2188 4170 2248 4250
rect 2484 4170 2508 4250
rect 2508 4170 2588 4250
rect 2588 4170 2668 4250
rect 2668 4170 2720 4250
rect 2956 4170 2988 4250
rect 2988 4170 3068 4250
rect 3068 4170 3148 4250
rect 3148 4170 3192 4250
rect 3428 4170 3468 4250
rect 3468 4170 3548 4250
rect 3548 4170 3628 4250
rect 3628 4170 3664 4250
rect 3900 4170 3948 4250
rect 3948 4170 4028 4250
rect 4028 4170 4108 4250
rect 4108 4170 4136 4250
rect 4372 4170 4428 4250
rect 4428 4170 4508 4250
rect 4508 4170 4588 4250
rect 4588 4170 4608 4250
rect 4844 4170 4908 4250
rect 4908 4170 4988 4250
rect 4988 4170 5068 4250
rect 5068 4170 5080 4250
rect 5316 4170 5388 4250
rect 5388 4170 5468 4250
rect 5468 4170 5548 4250
rect 5548 4170 5552 4250
rect 5788 4170 5868 4250
rect 5868 4170 5948 4250
rect 5948 4170 6024 4250
rect 6260 4170 6268 4250
rect 6268 4170 6348 4250
rect 6348 4170 6428 4250
rect 6428 4170 6496 4250
rect 2012 4090 2248 4170
rect 2484 4090 2720 4170
rect 2956 4090 3192 4170
rect 3428 4090 3664 4170
rect 3900 4090 4136 4170
rect 4372 4090 4608 4170
rect 4844 4090 5080 4170
rect 5316 4090 5552 4170
rect 5788 4090 6024 4170
rect 6260 4090 6496 4170
rect 2012 4054 2028 4090
rect 2028 4054 2108 4090
rect 2108 4054 2188 4090
rect 2188 4054 2248 4090
rect 2484 4054 2508 4090
rect 2508 4054 2588 4090
rect 2588 4054 2668 4090
rect 2668 4054 2720 4090
rect 2956 4054 2988 4090
rect 2988 4054 3068 4090
rect 3068 4054 3148 4090
rect 3148 4054 3192 4090
rect 3428 4054 3468 4090
rect 3468 4054 3548 4090
rect 3548 4054 3628 4090
rect 3628 4054 3664 4090
rect 3900 4054 3948 4090
rect 3948 4054 4028 4090
rect 4028 4054 4108 4090
rect 4108 4054 4136 4090
rect 4372 4054 4428 4090
rect 4428 4054 4508 4090
rect 4508 4054 4588 4090
rect 4588 4054 4608 4090
rect 4844 4054 4908 4090
rect 4908 4054 4988 4090
rect 4988 4054 5068 4090
rect 5068 4054 5080 4090
rect 5316 4054 5388 4090
rect 5388 4054 5468 4090
rect 5468 4054 5548 4090
rect 5548 4054 5552 4090
rect 5788 4054 5868 4090
rect 5868 4054 5948 4090
rect 5948 4054 6024 4090
rect 6260 4054 6268 4090
rect 6268 4054 6348 4090
rect 6348 4054 6428 4090
rect 6428 4054 6496 4090
<< metal5 >>
rect 1844 4290 6812 6390
rect 1844 4054 2012 4290
rect 2248 4054 2484 4290
rect 2720 4054 2956 4290
rect 3192 4054 3428 4290
rect 3664 4054 3900 4290
rect 4136 4054 4372 4290
rect 4608 4054 4844 4290
rect 5080 4054 5316 4290
rect 5552 4054 5788 4290
rect 6024 4054 6260 4290
rect 6496 4054 6812 4290
rect 1844 0 6812 4054
<< end >>
