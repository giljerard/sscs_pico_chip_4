magic
tech sky130A
magscale 1 2
timestamp 1636532148
<< nwell >>
rect 227356 690078 232850 691446
<< pwell >>
rect 165334 690070 170828 691426
rect 165334 690068 170520 690070
rect 170590 690068 170828 690070
<< pmoslvt >>
rect 227552 690226 227752 691226
rect 227810 690226 228010 691226
rect 228068 690226 228268 691226
rect 228326 690226 228526 691226
rect 228584 690226 228784 691226
rect 228842 690226 229042 691226
rect 229100 690226 229300 691226
rect 229358 690226 229558 691226
rect 229616 690226 229816 691226
rect 229874 690226 230074 691226
rect 230132 690226 230332 691226
rect 230390 690226 230590 691226
rect 230648 690226 230848 691226
rect 230906 690226 231106 691226
rect 231164 690226 231364 691226
rect 231422 690226 231622 691226
rect 231680 690226 231880 691226
rect 231938 690226 232138 691226
rect 232196 690226 232396 691226
rect 232454 690226 232654 691226
<< nmoslvt >>
rect 165530 690216 165730 691216
rect 165788 690216 165988 691216
rect 166046 690216 166246 691216
rect 166304 690216 166504 691216
rect 166562 690216 166762 691216
rect 166820 690216 167020 691216
rect 167078 690216 167278 691216
rect 167336 690216 167536 691216
rect 167594 690216 167794 691216
rect 167852 690216 168052 691216
rect 168110 690216 168310 691216
rect 168368 690216 168568 691216
rect 168626 690216 168826 691216
rect 168884 690216 169084 691216
rect 169142 690216 169342 691216
rect 169400 690216 169600 691216
rect 169658 690216 169858 691216
rect 169916 690216 170116 691216
rect 170174 690216 170374 691216
rect 170432 690216 170632 691216
<< ndiff >>
rect 165472 691204 165530 691216
rect 165472 690228 165484 691204
rect 165518 690228 165530 691204
rect 165472 690216 165530 690228
rect 165730 691204 165788 691216
rect 165730 690228 165742 691204
rect 165776 690228 165788 691204
rect 165730 690216 165788 690228
rect 165988 691204 166046 691216
rect 165988 690228 166000 691204
rect 166034 690228 166046 691204
rect 165988 690216 166046 690228
rect 166246 691204 166304 691216
rect 166246 690228 166258 691204
rect 166292 690228 166304 691204
rect 166246 690216 166304 690228
rect 166504 691204 166562 691216
rect 166504 690228 166516 691204
rect 166550 690228 166562 691204
rect 166504 690216 166562 690228
rect 166762 691204 166820 691216
rect 166762 690228 166774 691204
rect 166808 690228 166820 691204
rect 166762 690216 166820 690228
rect 167020 691204 167078 691216
rect 167020 690228 167032 691204
rect 167066 690228 167078 691204
rect 167020 690216 167078 690228
rect 167278 691204 167336 691216
rect 167278 690228 167290 691204
rect 167324 690228 167336 691204
rect 167278 690216 167336 690228
rect 167536 691204 167594 691216
rect 167536 690228 167548 691204
rect 167582 690228 167594 691204
rect 167536 690216 167594 690228
rect 167794 691204 167852 691216
rect 167794 690228 167806 691204
rect 167840 690228 167852 691204
rect 167794 690216 167852 690228
rect 168052 691204 168110 691216
rect 168052 690228 168064 691204
rect 168098 690228 168110 691204
rect 168052 690216 168110 690228
rect 168310 691204 168368 691216
rect 168310 690228 168322 691204
rect 168356 690228 168368 691204
rect 168310 690216 168368 690228
rect 168568 691204 168626 691216
rect 168568 690228 168580 691204
rect 168614 690228 168626 691204
rect 168568 690216 168626 690228
rect 168826 691204 168884 691216
rect 168826 690228 168838 691204
rect 168872 690228 168884 691204
rect 168826 690216 168884 690228
rect 169084 691204 169142 691216
rect 169084 690228 169096 691204
rect 169130 690228 169142 691204
rect 169084 690216 169142 690228
rect 169342 691204 169400 691216
rect 169342 690228 169354 691204
rect 169388 690228 169400 691204
rect 169342 690216 169400 690228
rect 169600 691204 169658 691216
rect 169600 690228 169612 691204
rect 169646 690228 169658 691204
rect 169600 690216 169658 690228
rect 169858 691204 169916 691216
rect 169858 690228 169870 691204
rect 169904 690228 169916 691204
rect 169858 690216 169916 690228
rect 170116 691204 170174 691216
rect 170116 690228 170128 691204
rect 170162 690228 170174 691204
rect 170116 690216 170174 690228
rect 170374 691204 170432 691216
rect 170374 690228 170386 691204
rect 170420 690228 170432 691204
rect 170374 690216 170432 690228
rect 170632 691204 170690 691216
rect 170632 690228 170644 691204
rect 170678 690228 170690 691204
rect 170632 690216 170690 690228
<< pdiff >>
rect 227494 691214 227552 691226
rect 227494 690238 227506 691214
rect 227540 690238 227552 691214
rect 227494 690226 227552 690238
rect 227752 691214 227810 691226
rect 227752 690238 227764 691214
rect 227798 690238 227810 691214
rect 227752 690226 227810 690238
rect 228010 691214 228068 691226
rect 228010 690238 228022 691214
rect 228056 690238 228068 691214
rect 228010 690226 228068 690238
rect 228268 691214 228326 691226
rect 228268 690238 228280 691214
rect 228314 690238 228326 691214
rect 228268 690226 228326 690238
rect 228526 691214 228584 691226
rect 228526 690238 228538 691214
rect 228572 690238 228584 691214
rect 228526 690226 228584 690238
rect 228784 691214 228842 691226
rect 228784 690238 228796 691214
rect 228830 690238 228842 691214
rect 228784 690226 228842 690238
rect 229042 691214 229100 691226
rect 229042 690238 229054 691214
rect 229088 690238 229100 691214
rect 229042 690226 229100 690238
rect 229300 691214 229358 691226
rect 229300 690238 229312 691214
rect 229346 690238 229358 691214
rect 229300 690226 229358 690238
rect 229558 691214 229616 691226
rect 229558 690238 229570 691214
rect 229604 690238 229616 691214
rect 229558 690226 229616 690238
rect 229816 691214 229874 691226
rect 229816 690238 229828 691214
rect 229862 690238 229874 691214
rect 229816 690226 229874 690238
rect 230074 691214 230132 691226
rect 230074 690238 230086 691214
rect 230120 690238 230132 691214
rect 230074 690226 230132 690238
rect 230332 691214 230390 691226
rect 230332 690238 230344 691214
rect 230378 690238 230390 691214
rect 230332 690226 230390 690238
rect 230590 691214 230648 691226
rect 230590 690238 230602 691214
rect 230636 690238 230648 691214
rect 230590 690226 230648 690238
rect 230848 691214 230906 691226
rect 230848 690238 230860 691214
rect 230894 690238 230906 691214
rect 230848 690226 230906 690238
rect 231106 691214 231164 691226
rect 231106 690238 231118 691214
rect 231152 690238 231164 691214
rect 231106 690226 231164 690238
rect 231364 691214 231422 691226
rect 231364 690238 231376 691214
rect 231410 690238 231422 691214
rect 231364 690226 231422 690238
rect 231622 691214 231680 691226
rect 231622 690238 231634 691214
rect 231668 690238 231680 691214
rect 231622 690226 231680 690238
rect 231880 691214 231938 691226
rect 231880 690238 231892 691214
rect 231926 690238 231938 691214
rect 231880 690226 231938 690238
rect 232138 691214 232196 691226
rect 232138 690238 232150 691214
rect 232184 690238 232196 691214
rect 232138 690226 232196 690238
rect 232396 691214 232454 691226
rect 232396 690238 232408 691214
rect 232442 690238 232454 691214
rect 232396 690226 232454 690238
rect 232654 691214 232712 691226
rect 232654 690238 232666 691214
rect 232700 690238 232712 691214
rect 232654 690226 232712 690238
<< ndiffc >>
rect 165484 690228 165518 691204
rect 165742 690228 165776 691204
rect 166000 690228 166034 691204
rect 166258 690228 166292 691204
rect 166516 690228 166550 691204
rect 166774 690228 166808 691204
rect 167032 690228 167066 691204
rect 167290 690228 167324 691204
rect 167548 690228 167582 691204
rect 167806 690228 167840 691204
rect 168064 690228 168098 691204
rect 168322 690228 168356 691204
rect 168580 690228 168614 691204
rect 168838 690228 168872 691204
rect 169096 690228 169130 691204
rect 169354 690228 169388 691204
rect 169612 690228 169646 691204
rect 169870 690228 169904 691204
rect 170128 690228 170162 691204
rect 170386 690228 170420 691204
rect 170644 690228 170678 691204
<< pdiffc >>
rect 227506 690238 227540 691214
rect 227764 690238 227798 691214
rect 228022 690238 228056 691214
rect 228280 690238 228314 691214
rect 228538 690238 228572 691214
rect 228796 690238 228830 691214
rect 229054 690238 229088 691214
rect 229312 690238 229346 691214
rect 229570 690238 229604 691214
rect 229828 690238 229862 691214
rect 230086 690238 230120 691214
rect 230344 690238 230378 691214
rect 230602 690238 230636 691214
rect 230860 690238 230894 691214
rect 231118 690238 231152 691214
rect 231376 690238 231410 691214
rect 231634 690238 231668 691214
rect 231892 690238 231926 691214
rect 232150 690238 232184 691214
rect 232408 690238 232442 691214
rect 232666 690238 232700 691214
<< psubdiff >>
rect 165370 691356 165466 691390
rect 170696 691356 170792 691390
rect 165370 691294 165404 691356
rect 170758 691294 170792 691356
rect 165370 690138 165404 690200
rect 170758 690138 170792 690200
rect 165370 690104 165466 690138
rect 170696 690104 170792 690138
<< nsubdiff >>
rect 227392 691376 227488 691410
rect 232718 691376 232814 691410
rect 227392 691313 227426 691376
rect 232780 691313 232814 691376
rect 227392 690148 227426 690211
rect 232780 690148 232814 690211
rect 227392 690114 227488 690148
rect 232718 690114 232814 690148
<< psubdiffcont >>
rect 165466 691356 170696 691390
rect 165370 690200 165404 691294
rect 170758 690200 170792 691294
rect 165466 690104 170696 690138
<< nsubdiffcont >>
rect 227488 691376 232718 691410
rect 227392 690211 227426 691313
rect 232780 690211 232814 691313
rect 227488 690114 232718 690148
<< poly >>
rect 165530 691288 165730 691304
rect 165530 691254 165546 691288
rect 165714 691254 165730 691288
rect 165530 691216 165730 691254
rect 165788 691288 165988 691304
rect 165788 691254 165804 691288
rect 165972 691254 165988 691288
rect 165788 691216 165988 691254
rect 166046 691288 166246 691304
rect 166046 691254 166062 691288
rect 166230 691254 166246 691288
rect 166046 691216 166246 691254
rect 166304 691288 166504 691304
rect 166304 691254 166320 691288
rect 166488 691254 166504 691288
rect 166304 691216 166504 691254
rect 166562 691288 166762 691304
rect 166562 691254 166578 691288
rect 166746 691254 166762 691288
rect 166562 691216 166762 691254
rect 166820 691288 167020 691304
rect 166820 691254 166836 691288
rect 167004 691254 167020 691288
rect 166820 691216 167020 691254
rect 167078 691288 167278 691304
rect 167078 691254 167094 691288
rect 167262 691254 167278 691288
rect 167078 691216 167278 691254
rect 167336 691288 167536 691304
rect 167336 691254 167352 691288
rect 167520 691254 167536 691288
rect 167336 691216 167536 691254
rect 167594 691288 167794 691304
rect 167594 691254 167610 691288
rect 167778 691254 167794 691288
rect 167594 691216 167794 691254
rect 167852 691288 168052 691304
rect 167852 691254 167868 691288
rect 168036 691254 168052 691288
rect 167852 691216 168052 691254
rect 168110 691288 168310 691304
rect 168110 691254 168126 691288
rect 168294 691254 168310 691288
rect 168110 691216 168310 691254
rect 168368 691288 168568 691304
rect 168368 691254 168384 691288
rect 168552 691254 168568 691288
rect 168368 691216 168568 691254
rect 168626 691288 168826 691304
rect 168626 691254 168642 691288
rect 168810 691254 168826 691288
rect 168626 691216 168826 691254
rect 168884 691288 169084 691304
rect 168884 691254 168900 691288
rect 169068 691254 169084 691288
rect 168884 691216 169084 691254
rect 169142 691288 169342 691304
rect 169142 691254 169158 691288
rect 169326 691254 169342 691288
rect 169142 691216 169342 691254
rect 169400 691288 169600 691304
rect 169400 691254 169416 691288
rect 169584 691254 169600 691288
rect 169400 691216 169600 691254
rect 169658 691288 169858 691304
rect 169658 691254 169674 691288
rect 169842 691254 169858 691288
rect 169658 691216 169858 691254
rect 169916 691288 170116 691304
rect 169916 691254 169932 691288
rect 170100 691254 170116 691288
rect 169916 691216 170116 691254
rect 170174 691288 170374 691304
rect 170174 691254 170190 691288
rect 170358 691254 170374 691288
rect 170174 691216 170374 691254
rect 170432 691288 170632 691304
rect 170432 691254 170448 691288
rect 170616 691254 170632 691288
rect 170432 691216 170632 691254
rect 165530 690190 165730 690216
rect 165788 690190 165988 690216
rect 166046 690190 166246 690216
rect 166304 690190 166504 690216
rect 166562 690190 166762 690216
rect 166820 690190 167020 690216
rect 167078 690190 167278 690216
rect 167336 690190 167536 690216
rect 167594 690190 167794 690216
rect 167852 690190 168052 690216
rect 168110 690190 168310 690216
rect 168368 690190 168568 690216
rect 168626 690190 168826 690216
rect 168884 690190 169084 690216
rect 169142 690190 169342 690216
rect 169400 690190 169600 690216
rect 169658 690190 169858 690216
rect 169916 690190 170116 690216
rect 170174 690190 170374 690216
rect 170432 690190 170632 690216
rect 227552 691307 227752 691323
rect 227552 691273 227568 691307
rect 227736 691273 227752 691307
rect 227552 691226 227752 691273
rect 227810 691307 228010 691323
rect 227810 691273 227826 691307
rect 227994 691273 228010 691307
rect 227810 691226 228010 691273
rect 228068 691307 228268 691323
rect 228068 691273 228084 691307
rect 228252 691273 228268 691307
rect 228068 691226 228268 691273
rect 228326 691307 228526 691323
rect 228326 691273 228342 691307
rect 228510 691273 228526 691307
rect 228326 691226 228526 691273
rect 228584 691307 228784 691323
rect 228584 691273 228600 691307
rect 228768 691273 228784 691307
rect 228584 691226 228784 691273
rect 228842 691307 229042 691323
rect 228842 691273 228858 691307
rect 229026 691273 229042 691307
rect 228842 691226 229042 691273
rect 229100 691307 229300 691323
rect 229100 691273 229116 691307
rect 229284 691273 229300 691307
rect 229100 691226 229300 691273
rect 229358 691307 229558 691323
rect 229358 691273 229374 691307
rect 229542 691273 229558 691307
rect 229358 691226 229558 691273
rect 229616 691307 229816 691323
rect 229616 691273 229632 691307
rect 229800 691273 229816 691307
rect 229616 691226 229816 691273
rect 229874 691307 230074 691323
rect 229874 691273 229890 691307
rect 230058 691273 230074 691307
rect 229874 691226 230074 691273
rect 230132 691307 230332 691323
rect 230132 691273 230148 691307
rect 230316 691273 230332 691307
rect 230132 691226 230332 691273
rect 230390 691307 230590 691323
rect 230390 691273 230406 691307
rect 230574 691273 230590 691307
rect 230390 691226 230590 691273
rect 230648 691307 230848 691323
rect 230648 691273 230664 691307
rect 230832 691273 230848 691307
rect 230648 691226 230848 691273
rect 230906 691307 231106 691323
rect 230906 691273 230922 691307
rect 231090 691273 231106 691307
rect 230906 691226 231106 691273
rect 231164 691307 231364 691323
rect 231164 691273 231180 691307
rect 231348 691273 231364 691307
rect 231164 691226 231364 691273
rect 231422 691307 231622 691323
rect 231422 691273 231438 691307
rect 231606 691273 231622 691307
rect 231422 691226 231622 691273
rect 231680 691307 231880 691323
rect 231680 691273 231696 691307
rect 231864 691273 231880 691307
rect 231680 691226 231880 691273
rect 231938 691307 232138 691323
rect 231938 691273 231954 691307
rect 232122 691273 232138 691307
rect 231938 691226 232138 691273
rect 232196 691307 232396 691323
rect 232196 691273 232212 691307
rect 232380 691273 232396 691307
rect 232196 691226 232396 691273
rect 232454 691307 232654 691323
rect 232454 691273 232470 691307
rect 232638 691273 232654 691307
rect 232454 691226 232654 691273
rect 227552 690200 227752 690226
rect 227810 690200 228010 690226
rect 228068 690200 228268 690226
rect 228326 690200 228526 690226
rect 228584 690200 228784 690226
rect 228842 690200 229042 690226
rect 229100 690200 229300 690226
rect 229358 690200 229558 690226
rect 229616 690200 229816 690226
rect 229874 690200 230074 690226
rect 230132 690200 230332 690226
rect 230390 690200 230590 690226
rect 230648 690200 230848 690226
rect 230906 690200 231106 690226
rect 231164 690200 231364 690226
rect 231422 690200 231622 690226
rect 231680 690200 231880 690226
rect 231938 690200 232138 690226
rect 232196 690200 232396 690226
rect 232454 690200 232654 690226
<< polycont >>
rect 165546 691254 165714 691288
rect 165804 691254 165972 691288
rect 166062 691254 166230 691288
rect 166320 691254 166488 691288
rect 166578 691254 166746 691288
rect 166836 691254 167004 691288
rect 167094 691254 167262 691288
rect 167352 691254 167520 691288
rect 167610 691254 167778 691288
rect 167868 691254 168036 691288
rect 168126 691254 168294 691288
rect 168384 691254 168552 691288
rect 168642 691254 168810 691288
rect 168900 691254 169068 691288
rect 169158 691254 169326 691288
rect 169416 691254 169584 691288
rect 169674 691254 169842 691288
rect 169932 691254 170100 691288
rect 170190 691254 170358 691288
rect 170448 691254 170616 691288
rect 227568 691273 227736 691307
rect 227826 691273 227994 691307
rect 228084 691273 228252 691307
rect 228342 691273 228510 691307
rect 228600 691273 228768 691307
rect 228858 691273 229026 691307
rect 229116 691273 229284 691307
rect 229374 691273 229542 691307
rect 229632 691273 229800 691307
rect 229890 691273 230058 691307
rect 230148 691273 230316 691307
rect 230406 691273 230574 691307
rect 230664 691273 230832 691307
rect 230922 691273 231090 691307
rect 231180 691273 231348 691307
rect 231438 691273 231606 691307
rect 231696 691273 231864 691307
rect 231954 691273 232122 691307
rect 232212 691273 232380 691307
rect 232470 691273 232638 691307
<< locali >>
rect 165370 691356 165466 691390
rect 170696 691356 170792 691390
rect 165370 691294 165404 691356
rect 170758 691294 170792 691356
rect 165482 691254 165546 691288
rect 165714 691254 165804 691288
rect 165972 691254 166062 691288
rect 166230 691254 166320 691288
rect 166488 691254 166578 691288
rect 166746 691254 166836 691288
rect 167004 691254 167094 691288
rect 167262 691254 167352 691288
rect 167520 691254 167610 691288
rect 167778 691254 167868 691288
rect 168036 691254 168126 691288
rect 168294 691254 168384 691288
rect 168552 691254 168642 691288
rect 168810 691254 168900 691288
rect 169068 691254 169158 691288
rect 169326 691254 169416 691288
rect 169584 691254 169674 691288
rect 169842 691254 169932 691288
rect 170100 691254 170190 691288
rect 170358 691254 170448 691288
rect 170616 691254 170679 691288
rect 165484 691204 165518 691220
rect 165484 690212 165518 690228
rect 165742 691204 165776 691254
rect 165742 690212 165776 690228
rect 166000 691204 166034 691220
rect 166000 690212 166034 690228
rect 166258 691204 166292 691254
rect 166258 690212 166292 690228
rect 166516 691204 166550 691220
rect 166516 690212 166550 690228
rect 166774 691204 166808 691254
rect 166774 690212 166808 690228
rect 167032 691204 167066 691220
rect 167032 690212 167066 690228
rect 167290 691204 167324 691254
rect 167290 690212 167324 690228
rect 167548 691204 167582 691220
rect 167548 690212 167582 690228
rect 167806 691204 167840 691254
rect 167806 690212 167840 690228
rect 168064 691204 168098 691220
rect 168064 690212 168098 690228
rect 168322 691204 168356 691254
rect 168322 690212 168356 690228
rect 168580 691204 168614 691220
rect 168580 690212 168614 690228
rect 168838 691204 168872 691254
rect 168838 690212 168872 690228
rect 169096 691204 169130 691220
rect 169096 690212 169130 690228
rect 169354 691204 169388 691254
rect 169354 690212 169388 690228
rect 169612 691204 169646 691220
rect 169612 690212 169646 690228
rect 169870 691204 169904 691254
rect 169870 690212 169904 690228
rect 170128 691204 170162 691220
rect 170128 690212 170162 690228
rect 170386 691204 170420 691254
rect 170386 690212 170420 690228
rect 170644 691204 170678 691220
rect 170644 690212 170678 690228
rect 165370 690104 165404 690200
rect 170758 690104 170792 690200
rect 227392 691376 227488 691410
rect 232718 691376 232814 691410
rect 227392 691313 227426 691376
rect 232780 691313 232814 691376
rect 227506 691273 227568 691307
rect 227736 691273 227826 691307
rect 227994 691273 228084 691307
rect 228252 691273 228342 691307
rect 228510 691273 228600 691307
rect 228768 691273 228858 691307
rect 229026 691273 229116 691307
rect 229284 691273 229374 691307
rect 229542 691273 229632 691307
rect 229800 691273 229890 691307
rect 230058 691273 230148 691307
rect 230316 691273 230406 691307
rect 230574 691273 230664 691307
rect 230832 691273 230922 691307
rect 231090 691273 231180 691307
rect 231348 691273 231438 691307
rect 231606 691273 231696 691307
rect 231864 691273 231954 691307
rect 232122 691273 232212 691307
rect 232380 691273 232470 691307
rect 232638 691273 232700 691307
rect 227506 691214 227540 691230
rect 227506 690222 227540 690238
rect 227764 691214 227798 691273
rect 227764 690222 227798 690238
rect 228022 691214 228056 691230
rect 228022 690222 228056 690238
rect 228280 691214 228314 691273
rect 228280 690222 228314 690238
rect 228538 691214 228572 691230
rect 228538 690222 228572 690238
rect 228796 691214 228830 691273
rect 228796 690222 228830 690238
rect 229054 691214 229088 691230
rect 229054 690222 229088 690238
rect 229312 691214 229346 691273
rect 229312 690222 229346 690238
rect 229570 691214 229604 691230
rect 229570 690222 229604 690238
rect 229828 691214 229862 691273
rect 229828 690222 229862 690238
rect 230086 691214 230120 691230
rect 230086 690222 230120 690238
rect 230344 691214 230378 691273
rect 230344 690222 230378 690238
rect 230602 691214 230636 691230
rect 230602 690222 230636 690238
rect 230860 691214 230894 691273
rect 230860 690222 230894 690238
rect 231118 691214 231152 691230
rect 231118 690222 231152 690238
rect 231376 691214 231410 691273
rect 231376 690222 231410 690238
rect 231634 691214 231668 691230
rect 231634 690222 231668 690238
rect 231892 691214 231926 691273
rect 231892 690222 231926 690238
rect 232150 691214 232184 691230
rect 232150 690222 232184 690238
rect 232408 691214 232442 691273
rect 232408 690222 232442 690238
rect 232666 691214 232700 691230
rect 232666 690222 232700 690238
rect 227392 690114 227426 690211
rect 232780 690114 232814 690211
<< viali >>
rect 165588 691254 165672 691288
rect 165846 691254 165930 691288
rect 166104 691254 166188 691288
rect 166362 691254 166446 691288
rect 166620 691254 166704 691288
rect 166878 691254 166962 691288
rect 167136 691254 167220 691288
rect 167394 691254 167478 691288
rect 167652 691254 167736 691288
rect 167910 691254 167994 691288
rect 168168 691254 168252 691288
rect 168426 691254 168510 691288
rect 168684 691254 168768 691288
rect 168942 691254 169026 691288
rect 169200 691254 169284 691288
rect 169458 691254 169542 691288
rect 169716 691254 169800 691288
rect 169974 691254 170058 691288
rect 170232 691254 170316 691288
rect 170490 691254 170574 691288
rect 165370 690260 165404 691234
rect 165484 690228 165518 691204
rect 165742 690228 165776 691204
rect 166000 690228 166034 691204
rect 166258 690228 166292 691204
rect 166516 690228 166550 691204
rect 166774 690228 166808 691204
rect 167032 690228 167066 691204
rect 167290 690228 167324 691204
rect 167548 690228 167582 691204
rect 167806 690228 167840 691204
rect 168064 690228 168098 691204
rect 168322 690228 168356 691204
rect 168580 690228 168614 691204
rect 168838 690228 168872 691204
rect 169096 690228 169130 691204
rect 169354 690228 169388 691204
rect 169612 690228 169646 691204
rect 169870 690228 169904 691204
rect 170128 690228 170162 691204
rect 170386 690228 170420 691204
rect 170644 690228 170678 691204
rect 170758 690260 170792 691234
rect 165404 690104 165466 690138
rect 165466 690104 170696 690138
rect 170696 690104 170758 690138
rect 227610 691273 227694 691307
rect 227868 691273 227952 691307
rect 228126 691273 228210 691307
rect 228384 691273 228468 691307
rect 228642 691273 228726 691307
rect 228900 691273 228984 691307
rect 229158 691273 229242 691307
rect 229416 691273 229500 691307
rect 229674 691273 229758 691307
rect 229932 691273 230016 691307
rect 230190 691273 230274 691307
rect 230448 691273 230532 691307
rect 230706 691273 230790 691307
rect 230964 691273 231048 691307
rect 231222 691273 231306 691307
rect 231480 691273 231564 691307
rect 231738 691273 231822 691307
rect 231996 691273 232080 691307
rect 232254 691273 232338 691307
rect 232512 691273 232596 691307
rect 227392 690271 227426 691253
rect 227506 690238 227540 691214
rect 227764 690238 227798 691214
rect 228022 690238 228056 691214
rect 228280 690238 228314 691214
rect 228538 690238 228572 691214
rect 228796 690238 228830 691214
rect 229054 690238 229088 691214
rect 229312 690238 229346 691214
rect 229570 690238 229604 691214
rect 229828 690238 229862 691214
rect 230086 690238 230120 691214
rect 230344 690238 230378 691214
rect 230602 690238 230636 691214
rect 230860 690238 230894 691214
rect 231118 690238 231152 691214
rect 231376 690238 231410 691214
rect 231634 690238 231668 691214
rect 231892 690238 231926 691214
rect 232150 690238 232184 691214
rect 232408 690238 232442 691214
rect 232666 690238 232700 691214
rect 232780 690271 232814 691253
rect 227426 690114 227488 690148
rect 227488 690114 232718 690148
rect 232718 690114 232780 690148
<< metal1 >>
rect 165334 691580 170828 691635
rect 165334 691510 165360 691580
rect 165430 691510 165460 691580
rect 165530 691510 165560 691580
rect 165630 691510 165660 691580
rect 165730 691510 165760 691580
rect 165830 691510 165860 691580
rect 165930 691510 165960 691580
rect 166030 691510 166060 691580
rect 166130 691510 166160 691580
rect 166230 691510 166260 691580
rect 166330 691510 166360 691580
rect 166430 691510 166460 691580
rect 166530 691510 166560 691580
rect 166630 691510 166660 691580
rect 166730 691510 166760 691580
rect 166830 691510 166860 691580
rect 166930 691510 166960 691580
rect 167030 691510 167060 691580
rect 167130 691510 167160 691580
rect 167230 691510 167260 691580
rect 167330 691510 167360 691580
rect 167430 691510 167460 691580
rect 167530 691510 167560 691580
rect 167630 691510 167660 691580
rect 167730 691510 167760 691580
rect 167830 691510 167860 691580
rect 167930 691510 167960 691580
rect 168030 691510 168060 691580
rect 168130 691510 168160 691580
rect 168230 691510 168260 691580
rect 168330 691510 168360 691580
rect 168430 691510 168460 691580
rect 168530 691510 168560 691580
rect 168630 691510 168660 691580
rect 168730 691510 168760 691580
rect 168830 691510 168860 691580
rect 168930 691510 168960 691580
rect 169030 691510 169060 691580
rect 169130 691510 169160 691580
rect 169230 691510 169260 691580
rect 169330 691510 169360 691580
rect 169430 691510 169460 691580
rect 169530 691510 169560 691580
rect 169630 691510 169660 691580
rect 169730 691510 169760 691580
rect 169830 691510 169860 691580
rect 169930 691510 169960 691580
rect 170030 691510 170060 691580
rect 170130 691510 170160 691580
rect 170230 691510 170260 691580
rect 170330 691510 170360 691580
rect 170430 691510 170460 691580
rect 170530 691510 170828 691580
rect 165334 691470 170828 691510
rect 165334 691400 165360 691470
rect 165430 691400 165460 691470
rect 165530 691400 165560 691470
rect 165630 691400 165660 691470
rect 165730 691400 165760 691470
rect 165830 691400 165860 691470
rect 165930 691400 165960 691470
rect 166030 691400 166060 691470
rect 166130 691400 166160 691470
rect 166230 691400 166260 691470
rect 166330 691400 166360 691470
rect 166430 691400 166460 691470
rect 166530 691400 166560 691470
rect 166630 691400 166660 691470
rect 166730 691400 166760 691470
rect 166830 691400 166860 691470
rect 166930 691400 166960 691470
rect 167030 691400 167060 691470
rect 167130 691400 167160 691470
rect 167230 691400 167260 691470
rect 167330 691400 167360 691470
rect 167430 691400 167460 691470
rect 167530 691400 167560 691470
rect 167630 691400 167660 691470
rect 167730 691400 167760 691470
rect 167830 691400 167860 691470
rect 167930 691400 167960 691470
rect 168030 691400 168060 691470
rect 168130 691400 168160 691470
rect 168230 691400 168260 691470
rect 168330 691400 168360 691470
rect 168430 691400 168460 691470
rect 168530 691400 168560 691470
rect 168630 691400 168660 691470
rect 168730 691400 168760 691470
rect 168830 691400 168860 691470
rect 168930 691400 168960 691470
rect 169030 691400 169060 691470
rect 169130 691400 169160 691470
rect 169230 691400 169260 691470
rect 169330 691400 169360 691470
rect 169430 691400 169460 691470
rect 169530 691400 169560 691470
rect 169630 691400 169660 691470
rect 169730 691400 169760 691470
rect 169830 691400 169860 691470
rect 169930 691400 169960 691470
rect 170030 691400 170060 691470
rect 170130 691400 170160 691470
rect 170230 691400 170260 691470
rect 170330 691400 170360 691470
rect 170430 691400 170460 691470
rect 170530 691400 170828 691470
rect 165334 691360 170828 691400
rect 227356 691600 232850 691626
rect 227356 691540 227370 691600
rect 227430 691540 227460 691600
rect 227520 691540 227550 691600
rect 227610 691540 227640 691600
rect 227700 691540 227730 691600
rect 227790 691540 227820 691600
rect 227880 691540 227910 691600
rect 227970 691540 228000 691600
rect 228060 691540 228090 691600
rect 228150 691540 228180 691600
rect 228240 691540 228270 691600
rect 228330 691540 228360 691600
rect 228420 691540 228450 691600
rect 228510 691540 228540 691600
rect 228600 691540 228630 691600
rect 228690 691540 228720 691600
rect 228780 691540 228810 691600
rect 228870 691540 228900 691600
rect 228960 691540 228990 691600
rect 229050 691540 229080 691600
rect 229140 691540 229170 691600
rect 229230 691540 229260 691600
rect 229320 691540 229350 691600
rect 229410 691540 229440 691600
rect 229500 691540 229530 691600
rect 229590 691540 229620 691600
rect 229680 691540 229710 691600
rect 229770 691540 229800 691600
rect 229860 691540 229890 691600
rect 229950 691540 229980 691600
rect 230040 691540 230070 691600
rect 230130 691540 230160 691600
rect 230220 691540 230250 691600
rect 230310 691540 230340 691600
rect 230400 691540 230430 691600
rect 230490 691540 230520 691600
rect 230580 691540 230610 691600
rect 230670 691540 230700 691600
rect 230760 691540 230790 691600
rect 230850 691540 230880 691600
rect 230940 691540 230970 691600
rect 231030 691540 231060 691600
rect 231120 691540 231150 691600
rect 231210 691540 231240 691600
rect 231300 691540 231330 691600
rect 231390 691540 231420 691600
rect 231480 691540 231510 691600
rect 231570 691540 231600 691600
rect 231660 691540 231690 691600
rect 231750 691540 231780 691600
rect 231840 691540 231870 691600
rect 231930 691540 231960 691600
rect 232020 691540 232050 691600
rect 232110 691540 232140 691600
rect 232200 691540 232230 691600
rect 232290 691540 232320 691600
rect 232380 691540 232410 691600
rect 232470 691540 232500 691600
rect 232560 691540 232590 691600
rect 232650 691540 232680 691600
rect 232740 691540 232770 691600
rect 232830 691540 232850 691600
rect 227356 691510 232850 691540
rect 227356 691450 227370 691510
rect 227430 691450 227460 691510
rect 227520 691450 227550 691510
rect 227610 691450 227640 691510
rect 227700 691450 227730 691510
rect 227790 691450 227820 691510
rect 227880 691450 227910 691510
rect 227970 691450 228000 691510
rect 228060 691450 228090 691510
rect 228150 691450 228180 691510
rect 228240 691450 228270 691510
rect 228330 691450 228360 691510
rect 228420 691450 228450 691510
rect 228510 691450 228540 691510
rect 228600 691450 228630 691510
rect 228690 691450 228720 691510
rect 228780 691450 228810 691510
rect 228870 691450 228900 691510
rect 228960 691450 228990 691510
rect 229050 691450 229080 691510
rect 229140 691450 229170 691510
rect 229230 691450 229260 691510
rect 229320 691450 229350 691510
rect 229410 691450 229440 691510
rect 229500 691450 229530 691510
rect 229590 691450 229620 691510
rect 229680 691450 229710 691510
rect 229770 691450 229800 691510
rect 229860 691450 229890 691510
rect 229950 691450 229980 691510
rect 230040 691450 230070 691510
rect 230130 691450 230160 691510
rect 230220 691450 230250 691510
rect 230310 691450 230340 691510
rect 230400 691450 230430 691510
rect 230490 691450 230520 691510
rect 230580 691450 230610 691510
rect 230670 691450 230700 691510
rect 230760 691450 230790 691510
rect 230850 691450 230880 691510
rect 230940 691450 230970 691510
rect 231030 691450 231060 691510
rect 231120 691450 231150 691510
rect 231210 691450 231240 691510
rect 231300 691450 231330 691510
rect 231390 691450 231420 691510
rect 231480 691450 231510 691510
rect 231570 691450 231600 691510
rect 231660 691450 231690 691510
rect 231750 691450 231780 691510
rect 231840 691450 231870 691510
rect 231930 691450 231960 691510
rect 232020 691450 232050 691510
rect 232110 691450 232140 691510
rect 232200 691450 232230 691510
rect 232290 691450 232320 691510
rect 232380 691450 232410 691510
rect 232470 691450 232500 691510
rect 232560 691450 232590 691510
rect 232650 691450 232680 691510
rect 232740 691450 232770 691510
rect 232830 691450 232850 691510
rect 227356 691420 232850 691450
rect 227356 691360 227370 691420
rect 227430 691360 227460 691420
rect 227520 691360 227550 691420
rect 227610 691360 227640 691420
rect 227700 691360 227730 691420
rect 227790 691360 227820 691420
rect 227880 691360 227910 691420
rect 227970 691360 228000 691420
rect 228060 691360 228090 691420
rect 228150 691360 228180 691420
rect 228240 691360 228270 691420
rect 228330 691360 228360 691420
rect 228420 691360 228450 691420
rect 228510 691360 228540 691420
rect 228600 691360 228630 691420
rect 228690 691360 228720 691420
rect 228780 691360 228810 691420
rect 228870 691360 228900 691420
rect 228960 691360 228990 691420
rect 229050 691360 229080 691420
rect 229140 691360 229170 691420
rect 229230 691360 229260 691420
rect 229320 691360 229350 691420
rect 229410 691360 229440 691420
rect 229500 691360 229530 691420
rect 229590 691360 229620 691420
rect 229680 691360 229710 691420
rect 229770 691360 229800 691420
rect 229860 691360 229890 691420
rect 229950 691360 229980 691420
rect 230040 691360 230070 691420
rect 230130 691360 230160 691420
rect 230220 691360 230250 691420
rect 230310 691360 230340 691420
rect 230400 691360 230430 691420
rect 230490 691360 230520 691420
rect 230580 691360 230610 691420
rect 230670 691360 230700 691420
rect 230760 691360 230790 691420
rect 230850 691360 230880 691420
rect 230940 691360 230970 691420
rect 231030 691360 231060 691420
rect 231120 691360 231150 691420
rect 231210 691360 231240 691420
rect 231300 691360 231330 691420
rect 231390 691360 231420 691420
rect 231480 691360 231510 691420
rect 231570 691360 231600 691420
rect 231660 691360 231690 691420
rect 231750 691360 231780 691420
rect 231840 691360 231870 691420
rect 231930 691360 231960 691420
rect 232020 691360 232050 691420
rect 232110 691360 232140 691420
rect 232200 691360 232230 691420
rect 232290 691360 232320 691420
rect 232380 691360 232410 691420
rect 232470 691360 232500 691420
rect 232560 691360 232590 691420
rect 232650 691360 232680 691420
rect 232740 691360 232770 691420
rect 232830 691360 232850 691420
rect 165364 691234 165410 691246
rect 165364 690260 165370 691234
rect 165404 690260 165410 691234
rect 165364 690178 165410 690260
rect 165478 691204 165524 691360
rect 165576 691288 165684 691294
rect 165576 691254 165588 691288
rect 165672 691254 165684 691288
rect 165576 691248 165684 691254
rect 165834 691288 165942 691294
rect 165834 691254 165846 691288
rect 165930 691254 165942 691288
rect 165834 691248 165942 691254
rect 165478 690228 165484 691204
rect 165518 690228 165524 691204
rect 165478 690216 165524 690228
rect 165736 691204 165782 691216
rect 165736 690228 165742 691204
rect 165776 690228 165782 691204
rect 165736 690216 165782 690228
rect 165994 691204 166040 691360
rect 166092 691288 166200 691294
rect 166092 691254 166104 691288
rect 166188 691254 166200 691288
rect 166092 691248 166200 691254
rect 166350 691288 166458 691294
rect 166350 691254 166362 691288
rect 166446 691254 166458 691288
rect 166350 691248 166458 691254
rect 165994 690228 166000 691204
rect 166034 690228 166040 691204
rect 165994 690216 166040 690228
rect 166252 691204 166298 691216
rect 166252 690228 166258 691204
rect 166292 690228 166298 691204
rect 166252 690216 166298 690228
rect 166510 691204 166556 691360
rect 166608 691288 166716 691294
rect 166608 691254 166620 691288
rect 166704 691254 166716 691288
rect 166608 691248 166716 691254
rect 166866 691288 166974 691294
rect 166866 691254 166878 691288
rect 166962 691254 166974 691288
rect 166866 691248 166974 691254
rect 166510 690228 166516 691204
rect 166550 690228 166556 691204
rect 166510 690216 166556 690228
rect 166768 691204 166814 691216
rect 166768 690228 166774 691204
rect 166808 690228 166814 691204
rect 166768 690216 166814 690228
rect 167026 691204 167072 691360
rect 167124 691288 167232 691294
rect 167124 691254 167136 691288
rect 167220 691254 167232 691288
rect 167124 691248 167232 691254
rect 167382 691288 167490 691294
rect 167382 691254 167394 691288
rect 167478 691254 167490 691288
rect 167382 691248 167490 691254
rect 167026 690228 167032 691204
rect 167066 690228 167072 691204
rect 167026 690216 167072 690228
rect 167284 691204 167330 691216
rect 167284 690228 167290 691204
rect 167324 690228 167330 691204
rect 167284 690216 167330 690228
rect 167542 691204 167588 691360
rect 167640 691288 167748 691294
rect 167640 691254 167652 691288
rect 167736 691254 167748 691288
rect 167640 691248 167748 691254
rect 167898 691288 168006 691294
rect 167898 691254 167910 691288
rect 167994 691254 168006 691288
rect 167898 691248 168006 691254
rect 167542 690228 167548 691204
rect 167582 690228 167588 691204
rect 167542 690216 167588 690228
rect 167800 691204 167846 691216
rect 167800 690228 167806 691204
rect 167840 690228 167846 691204
rect 167800 690216 167846 690228
rect 168058 691204 168104 691360
rect 168156 691288 168264 691294
rect 168156 691254 168168 691288
rect 168252 691254 168264 691288
rect 168156 691248 168264 691254
rect 168414 691288 168522 691294
rect 168414 691254 168426 691288
rect 168510 691254 168522 691288
rect 168414 691248 168522 691254
rect 168058 690228 168064 691204
rect 168098 690228 168104 691204
rect 168058 690216 168104 690228
rect 168316 691204 168362 691216
rect 168316 690228 168322 691204
rect 168356 690228 168362 691204
rect 168316 690216 168362 690228
rect 168574 691204 168620 691360
rect 168672 691288 168780 691294
rect 168672 691254 168684 691288
rect 168768 691254 168780 691288
rect 168672 691248 168780 691254
rect 168930 691288 169038 691294
rect 168930 691254 168942 691288
rect 169026 691254 169038 691288
rect 168930 691248 169038 691254
rect 168574 690228 168580 691204
rect 168614 690228 168620 691204
rect 168574 690216 168620 690228
rect 168832 691204 168878 691216
rect 168832 690228 168838 691204
rect 168872 690228 168878 691204
rect 168832 690216 168878 690228
rect 169090 691204 169136 691360
rect 169188 691288 169296 691294
rect 169188 691254 169200 691288
rect 169284 691254 169296 691288
rect 169188 691248 169296 691254
rect 169446 691288 169554 691294
rect 169446 691254 169458 691288
rect 169542 691254 169554 691288
rect 169446 691248 169554 691254
rect 169090 690228 169096 691204
rect 169130 690228 169136 691204
rect 169090 690216 169136 690228
rect 169348 691204 169394 691216
rect 169348 690228 169354 691204
rect 169388 690228 169394 691204
rect 169348 690216 169394 690228
rect 169606 691204 169652 691360
rect 169704 691288 169812 691294
rect 169704 691254 169716 691288
rect 169800 691254 169812 691288
rect 169704 691248 169812 691254
rect 169962 691288 170070 691294
rect 169962 691254 169974 691288
rect 170058 691254 170070 691288
rect 169962 691248 170070 691254
rect 169606 690228 169612 691204
rect 169646 690228 169652 691204
rect 169606 690216 169652 690228
rect 169864 691204 169910 691216
rect 169864 690228 169870 691204
rect 169904 690228 169910 691204
rect 169864 690216 169910 690228
rect 170122 691204 170168 691360
rect 170220 691288 170328 691294
rect 170220 691254 170232 691288
rect 170316 691254 170328 691288
rect 170220 691248 170328 691254
rect 170478 691288 170586 691294
rect 170478 691254 170490 691288
rect 170574 691254 170586 691288
rect 170478 691248 170586 691254
rect 170122 690228 170128 691204
rect 170162 690228 170168 691204
rect 170122 690216 170168 690228
rect 170380 691204 170426 691216
rect 170380 690228 170386 691204
rect 170420 690228 170426 691204
rect 170380 690216 170426 690228
rect 170638 691204 170684 691360
rect 227356 691351 232850 691360
rect 227386 691253 227432 691265
rect 170638 690228 170644 691204
rect 170678 690228 170684 691204
rect 170638 690216 170684 690228
rect 170752 691234 170798 691246
rect 170752 690260 170758 691234
rect 170792 690260 170798 691234
rect 165742 690178 165776 690216
rect 166258 690178 166292 690216
rect 166774 690178 166808 690216
rect 167290 690178 167324 690216
rect 167806 690178 167840 690216
rect 168322 690178 168356 690216
rect 168838 690178 168872 690216
rect 169354 690178 169388 690216
rect 169870 690178 169904 690216
rect 170386 690178 170420 690216
rect 170752 690178 170798 690260
rect 165364 690138 170798 690178
rect 165364 690104 165404 690138
rect 170758 690104 170798 690138
rect 165364 690070 170798 690104
rect 165364 690000 165620 690070
rect 165690 690000 165720 690070
rect 165790 690000 165820 690070
rect 165890 690000 165920 690070
rect 165990 690000 166020 690070
rect 166090 690000 166120 690070
rect 166190 690000 166220 690070
rect 166290 690000 166320 690070
rect 166390 690000 166420 690070
rect 166490 690000 166520 690070
rect 166590 690000 166620 690070
rect 166690 690000 166720 690070
rect 166790 690000 166820 690070
rect 166890 690000 166920 690070
rect 166990 690000 167020 690070
rect 167090 690000 167120 690070
rect 167190 690000 167220 690070
rect 167290 690000 167320 690070
rect 167390 690000 167420 690070
rect 167490 690000 167520 690070
rect 167590 690000 167620 690070
rect 167690 690000 167720 690070
rect 167790 690000 167820 690070
rect 167890 690000 167920 690070
rect 167990 690000 168020 690070
rect 168090 690000 168120 690070
rect 168190 690000 168220 690070
rect 168290 690000 168320 690070
rect 168390 690000 168420 690070
rect 168490 690000 168520 690070
rect 168590 690000 168620 690070
rect 168690 690000 168720 690070
rect 168790 690000 168820 690070
rect 168890 690000 168920 690070
rect 168990 690000 169020 690070
rect 169090 690000 169120 690070
rect 169190 690000 169220 690070
rect 169290 690000 169320 690070
rect 169390 690000 169420 690070
rect 169490 690000 169520 690070
rect 169590 690000 169620 690070
rect 169690 690000 169720 690070
rect 169790 690000 169820 690070
rect 169890 690000 169920 690070
rect 169990 690000 170020 690070
rect 170090 690000 170120 690070
rect 170190 690000 170220 690070
rect 170290 690000 170320 690070
rect 170390 690000 170420 690070
rect 170490 690000 170798 690070
rect 165364 689970 170798 690000
rect 165364 689900 165620 689970
rect 165690 689900 165720 689970
rect 165790 689900 165820 689970
rect 165890 689900 165920 689970
rect 165990 689900 166020 689970
rect 166090 689900 166120 689970
rect 166190 689900 166220 689970
rect 166290 689900 166320 689970
rect 166390 689900 166420 689970
rect 166490 689900 166520 689970
rect 166590 689900 166620 689970
rect 166690 689900 166720 689970
rect 166790 689900 166820 689970
rect 166890 689900 166920 689970
rect 166990 689900 167020 689970
rect 167090 689900 167120 689970
rect 167190 689900 167220 689970
rect 167290 689900 167320 689970
rect 167390 689900 167420 689970
rect 167490 689900 167520 689970
rect 167590 689900 167620 689970
rect 167690 689900 167720 689970
rect 167790 689900 167820 689970
rect 167890 689900 167920 689970
rect 167990 689900 168020 689970
rect 168090 689900 168120 689970
rect 168190 689900 168220 689970
rect 168290 689900 168320 689970
rect 168390 689900 168420 689970
rect 168490 689900 168520 689970
rect 168590 689900 168620 689970
rect 168690 689900 168720 689970
rect 168790 689900 168820 689970
rect 168890 689900 168920 689970
rect 168990 689900 169020 689970
rect 169090 689900 169120 689970
rect 169190 689900 169220 689970
rect 169290 689900 169320 689970
rect 169390 689900 169420 689970
rect 169490 689900 169520 689970
rect 169590 689900 169620 689970
rect 169690 689900 169720 689970
rect 169790 689900 169820 689970
rect 169890 689900 169920 689970
rect 169990 689900 170020 689970
rect 170090 689900 170120 689970
rect 170190 689900 170220 689970
rect 170290 689900 170320 689970
rect 170390 689900 170420 689970
rect 170490 689900 170798 689970
rect 165364 689877 170798 689900
rect 227386 690271 227392 691253
rect 227426 690271 227432 691253
rect 227386 690154 227432 690271
rect 227500 691214 227546 691351
rect 227598 691307 227706 691313
rect 227598 691273 227610 691307
rect 227694 691273 227706 691307
rect 227598 691267 227706 691273
rect 227856 691307 227964 691313
rect 227856 691273 227868 691307
rect 227952 691273 227964 691307
rect 227856 691267 227964 691273
rect 227500 690238 227506 691214
rect 227540 690238 227546 691214
rect 227500 690226 227546 690238
rect 227758 691214 227804 691226
rect 227758 690238 227764 691214
rect 227798 690238 227804 691214
rect 227758 690154 227804 690238
rect 228016 691214 228062 691351
rect 228114 691307 228222 691313
rect 228114 691273 228126 691307
rect 228210 691273 228222 691307
rect 228114 691267 228222 691273
rect 228372 691307 228480 691313
rect 228372 691273 228384 691307
rect 228468 691273 228480 691307
rect 228372 691267 228480 691273
rect 228016 690238 228022 691214
rect 228056 690238 228062 691214
rect 228016 690226 228062 690238
rect 228274 691214 228320 691226
rect 228274 690238 228280 691214
rect 228314 690238 228320 691214
rect 228274 690154 228320 690238
rect 228532 691214 228578 691351
rect 228630 691307 228738 691313
rect 228630 691273 228642 691307
rect 228726 691273 228738 691307
rect 228630 691267 228738 691273
rect 228888 691307 228996 691313
rect 228888 691273 228900 691307
rect 228984 691273 228996 691307
rect 228888 691267 228996 691273
rect 228532 690238 228538 691214
rect 228572 690238 228578 691214
rect 228532 690226 228578 690238
rect 228790 691214 228836 691226
rect 228790 690238 228796 691214
rect 228830 690238 228836 691214
rect 228790 690154 228836 690238
rect 229048 691214 229094 691351
rect 229146 691307 229254 691313
rect 229146 691273 229158 691307
rect 229242 691273 229254 691307
rect 229146 691267 229254 691273
rect 229404 691307 229512 691313
rect 229404 691273 229416 691307
rect 229500 691273 229512 691307
rect 229404 691267 229512 691273
rect 229048 690238 229054 691214
rect 229088 690238 229094 691214
rect 229048 690226 229094 690238
rect 229306 691214 229352 691226
rect 229306 690238 229312 691214
rect 229346 690238 229352 691214
rect 229306 690154 229352 690238
rect 229564 691214 229610 691351
rect 229662 691307 229770 691313
rect 229662 691273 229674 691307
rect 229758 691273 229770 691307
rect 229662 691267 229770 691273
rect 229920 691307 230028 691313
rect 229920 691273 229932 691307
rect 230016 691273 230028 691307
rect 229920 691267 230028 691273
rect 229564 690238 229570 691214
rect 229604 690238 229610 691214
rect 229564 690226 229610 690238
rect 229822 691214 229868 691226
rect 229822 690238 229828 691214
rect 229862 690238 229868 691214
rect 229822 690154 229868 690238
rect 230080 691214 230126 691351
rect 230178 691307 230286 691313
rect 230178 691273 230190 691307
rect 230274 691273 230286 691307
rect 230178 691267 230286 691273
rect 230436 691307 230544 691313
rect 230436 691273 230448 691307
rect 230532 691273 230544 691307
rect 230436 691267 230544 691273
rect 230080 690238 230086 691214
rect 230120 690238 230126 691214
rect 230080 690226 230126 690238
rect 230338 691214 230384 691226
rect 230338 690238 230344 691214
rect 230378 690238 230384 691214
rect 230338 690154 230384 690238
rect 230596 691214 230642 691351
rect 230694 691307 230802 691313
rect 230694 691273 230706 691307
rect 230790 691273 230802 691307
rect 230694 691267 230802 691273
rect 230952 691307 231060 691313
rect 230952 691273 230964 691307
rect 231048 691273 231060 691307
rect 230952 691267 231060 691273
rect 230596 690238 230602 691214
rect 230636 690238 230642 691214
rect 230596 690226 230642 690238
rect 230854 691214 230900 691226
rect 230854 690238 230860 691214
rect 230894 690238 230900 691214
rect 230854 690154 230900 690238
rect 231112 691214 231158 691351
rect 231210 691307 231318 691313
rect 231210 691273 231222 691307
rect 231306 691273 231318 691307
rect 231210 691267 231318 691273
rect 231468 691307 231576 691313
rect 231468 691273 231480 691307
rect 231564 691273 231576 691307
rect 231468 691267 231576 691273
rect 231112 690238 231118 691214
rect 231152 690238 231158 691214
rect 231112 690226 231158 690238
rect 231370 691214 231416 691226
rect 231370 690238 231376 691214
rect 231410 690238 231416 691214
rect 231370 690154 231416 690238
rect 231628 691214 231674 691351
rect 231726 691307 231834 691313
rect 231726 691273 231738 691307
rect 231822 691273 231834 691307
rect 231726 691267 231834 691273
rect 231984 691307 232092 691313
rect 231984 691273 231996 691307
rect 232080 691273 232092 691307
rect 231984 691267 232092 691273
rect 231628 690238 231634 691214
rect 231668 690238 231674 691214
rect 231628 690226 231674 690238
rect 231886 691214 231932 691226
rect 231886 690238 231892 691214
rect 231926 690238 231932 691214
rect 231886 690154 231932 690238
rect 232144 691214 232190 691351
rect 232242 691307 232350 691313
rect 232242 691273 232254 691307
rect 232338 691273 232350 691307
rect 232242 691267 232350 691273
rect 232500 691307 232608 691313
rect 232500 691273 232512 691307
rect 232596 691273 232608 691307
rect 232500 691267 232608 691273
rect 232144 690238 232150 691214
rect 232184 690238 232190 691214
rect 232144 690226 232190 690238
rect 232402 691214 232448 691226
rect 232402 690238 232408 691214
rect 232442 690238 232448 691214
rect 232402 690154 232448 690238
rect 232660 691214 232706 691351
rect 232660 690238 232666 691214
rect 232700 690238 232706 691214
rect 232660 690226 232706 690238
rect 232774 691253 232820 691265
rect 232774 690271 232780 691253
rect 232814 690271 232820 691253
rect 232774 690154 232820 690271
rect 227386 690148 232820 690154
rect 227386 690114 227426 690148
rect 232780 690114 232820 690148
rect 227386 690060 232820 690114
rect 227386 689990 227640 690060
rect 227710 689990 227740 690060
rect 227810 689990 227840 690060
rect 227910 689990 227940 690060
rect 228010 689990 228040 690060
rect 228110 689990 228140 690060
rect 228210 689990 228240 690060
rect 228310 689990 228340 690060
rect 228410 689990 228440 690060
rect 228510 689990 228540 690060
rect 228610 689990 228640 690060
rect 228710 689990 228740 690060
rect 228810 689990 228840 690060
rect 228910 689990 228940 690060
rect 229010 689990 229040 690060
rect 229110 689990 229140 690060
rect 229210 689990 229240 690060
rect 229310 689990 229340 690060
rect 229410 689990 229440 690060
rect 229510 689990 229540 690060
rect 229610 689990 229640 690060
rect 229710 689990 229740 690060
rect 229810 689990 229840 690060
rect 229910 689990 229940 690060
rect 230010 689990 230040 690060
rect 230110 689990 230140 690060
rect 230210 689990 230240 690060
rect 230310 689990 230340 690060
rect 230410 689990 230440 690060
rect 230510 689990 230540 690060
rect 230610 689990 230640 690060
rect 230710 689990 230740 690060
rect 230810 689990 230840 690060
rect 230910 689990 230940 690060
rect 231010 689990 231040 690060
rect 231110 689990 231140 690060
rect 231210 689990 231240 690060
rect 231310 689990 231340 690060
rect 231410 689990 231440 690060
rect 231510 689990 231540 690060
rect 231610 689990 231640 690060
rect 231710 689990 231740 690060
rect 231810 689990 231840 690060
rect 231910 689990 231940 690060
rect 232010 689990 232040 690060
rect 232110 689990 232140 690060
rect 232210 689990 232240 690060
rect 232310 689990 232340 690060
rect 232410 689990 232440 690060
rect 232510 689990 232820 690060
rect 227386 689960 232820 689990
rect 227386 689890 227640 689960
rect 227710 689890 227740 689960
rect 227810 689890 227840 689960
rect 227910 689890 227940 689960
rect 228010 689890 228040 689960
rect 228110 689890 228140 689960
rect 228210 689890 228240 689960
rect 228310 689890 228340 689960
rect 228410 689890 228440 689960
rect 228510 689890 228540 689960
rect 228610 689890 228640 689960
rect 228710 689890 228740 689960
rect 228810 689890 228840 689960
rect 228910 689890 228940 689960
rect 229010 689890 229040 689960
rect 229110 689890 229140 689960
rect 229210 689890 229240 689960
rect 229310 689890 229340 689960
rect 229410 689890 229440 689960
rect 229510 689890 229540 689960
rect 229610 689890 229640 689960
rect 229710 689890 229740 689960
rect 229810 689890 229840 689960
rect 229910 689890 229940 689960
rect 230010 689890 230040 689960
rect 230110 689890 230140 689960
rect 230210 689890 230240 689960
rect 230310 689890 230340 689960
rect 230410 689890 230440 689960
rect 230510 689890 230540 689960
rect 230610 689890 230640 689960
rect 230710 689890 230740 689960
rect 230810 689890 230840 689960
rect 230910 689890 230940 689960
rect 231010 689890 231040 689960
rect 231110 689890 231140 689960
rect 231210 689890 231240 689960
rect 231310 689890 231340 689960
rect 231410 689890 231440 689960
rect 231510 689890 231540 689960
rect 231610 689890 231640 689960
rect 231710 689890 231740 689960
rect 231810 689890 231840 689960
rect 231910 689890 231940 689960
rect 232010 689890 232040 689960
rect 232110 689890 232140 689960
rect 232210 689890 232240 689960
rect 232310 689890 232340 689960
rect 232410 689890 232440 689960
rect 232510 689890 232820 689960
rect 227386 689853 232820 689890
<< via1 >>
rect 165360 691510 165430 691580
rect 165460 691510 165530 691580
rect 165560 691510 165630 691580
rect 165660 691510 165730 691580
rect 165760 691510 165830 691580
rect 165860 691510 165930 691580
rect 165960 691510 166030 691580
rect 166060 691510 166130 691580
rect 166160 691510 166230 691580
rect 166260 691510 166330 691580
rect 166360 691510 166430 691580
rect 166460 691510 166530 691580
rect 166560 691510 166630 691580
rect 166660 691510 166730 691580
rect 166760 691510 166830 691580
rect 166860 691510 166930 691580
rect 166960 691510 167030 691580
rect 167060 691510 167130 691580
rect 167160 691510 167230 691580
rect 167260 691510 167330 691580
rect 167360 691510 167430 691580
rect 167460 691510 167530 691580
rect 167560 691510 167630 691580
rect 167660 691510 167730 691580
rect 167760 691510 167830 691580
rect 167860 691510 167930 691580
rect 167960 691510 168030 691580
rect 168060 691510 168130 691580
rect 168160 691510 168230 691580
rect 168260 691510 168330 691580
rect 168360 691510 168430 691580
rect 168460 691510 168530 691580
rect 168560 691510 168630 691580
rect 168660 691510 168730 691580
rect 168760 691510 168830 691580
rect 168860 691510 168930 691580
rect 168960 691510 169030 691580
rect 169060 691510 169130 691580
rect 169160 691510 169230 691580
rect 169260 691510 169330 691580
rect 169360 691510 169430 691580
rect 169460 691510 169530 691580
rect 169560 691510 169630 691580
rect 169660 691510 169730 691580
rect 169760 691510 169830 691580
rect 169860 691510 169930 691580
rect 169960 691510 170030 691580
rect 170060 691510 170130 691580
rect 170160 691510 170230 691580
rect 170260 691510 170330 691580
rect 170360 691510 170430 691580
rect 170460 691510 170530 691580
rect 165360 691400 165430 691470
rect 165460 691400 165530 691470
rect 165560 691400 165630 691470
rect 165660 691400 165730 691470
rect 165760 691400 165830 691470
rect 165860 691400 165930 691470
rect 165960 691400 166030 691470
rect 166060 691400 166130 691470
rect 166160 691400 166230 691470
rect 166260 691400 166330 691470
rect 166360 691400 166430 691470
rect 166460 691400 166530 691470
rect 166560 691400 166630 691470
rect 166660 691400 166730 691470
rect 166760 691400 166830 691470
rect 166860 691400 166930 691470
rect 166960 691400 167030 691470
rect 167060 691400 167130 691470
rect 167160 691400 167230 691470
rect 167260 691400 167330 691470
rect 167360 691400 167430 691470
rect 167460 691400 167530 691470
rect 167560 691400 167630 691470
rect 167660 691400 167730 691470
rect 167760 691400 167830 691470
rect 167860 691400 167930 691470
rect 167960 691400 168030 691470
rect 168060 691400 168130 691470
rect 168160 691400 168230 691470
rect 168260 691400 168330 691470
rect 168360 691400 168430 691470
rect 168460 691400 168530 691470
rect 168560 691400 168630 691470
rect 168660 691400 168730 691470
rect 168760 691400 168830 691470
rect 168860 691400 168930 691470
rect 168960 691400 169030 691470
rect 169060 691400 169130 691470
rect 169160 691400 169230 691470
rect 169260 691400 169330 691470
rect 169360 691400 169430 691470
rect 169460 691400 169530 691470
rect 169560 691400 169630 691470
rect 169660 691400 169730 691470
rect 169760 691400 169830 691470
rect 169860 691400 169930 691470
rect 169960 691400 170030 691470
rect 170060 691400 170130 691470
rect 170160 691400 170230 691470
rect 170260 691400 170330 691470
rect 170360 691400 170430 691470
rect 170460 691400 170530 691470
rect 227370 691540 227430 691600
rect 227460 691540 227520 691600
rect 227550 691540 227610 691600
rect 227640 691540 227700 691600
rect 227730 691540 227790 691600
rect 227820 691540 227880 691600
rect 227910 691540 227970 691600
rect 228000 691540 228060 691600
rect 228090 691540 228150 691600
rect 228180 691540 228240 691600
rect 228270 691540 228330 691600
rect 228360 691540 228420 691600
rect 228450 691540 228510 691600
rect 228540 691540 228600 691600
rect 228630 691540 228690 691600
rect 228720 691540 228780 691600
rect 228810 691540 228870 691600
rect 228900 691540 228960 691600
rect 228990 691540 229050 691600
rect 229080 691540 229140 691600
rect 229170 691540 229230 691600
rect 229260 691540 229320 691600
rect 229350 691540 229410 691600
rect 229440 691540 229500 691600
rect 229530 691540 229590 691600
rect 229620 691540 229680 691600
rect 229710 691540 229770 691600
rect 229800 691540 229860 691600
rect 229890 691540 229950 691600
rect 229980 691540 230040 691600
rect 230070 691540 230130 691600
rect 230160 691540 230220 691600
rect 230250 691540 230310 691600
rect 230340 691540 230400 691600
rect 230430 691540 230490 691600
rect 230520 691540 230580 691600
rect 230610 691540 230670 691600
rect 230700 691540 230760 691600
rect 230790 691540 230850 691600
rect 230880 691540 230940 691600
rect 230970 691540 231030 691600
rect 231060 691540 231120 691600
rect 231150 691540 231210 691600
rect 231240 691540 231300 691600
rect 231330 691540 231390 691600
rect 231420 691540 231480 691600
rect 231510 691540 231570 691600
rect 231600 691540 231660 691600
rect 231690 691540 231750 691600
rect 231780 691540 231840 691600
rect 231870 691540 231930 691600
rect 231960 691540 232020 691600
rect 232050 691540 232110 691600
rect 232140 691540 232200 691600
rect 232230 691540 232290 691600
rect 232320 691540 232380 691600
rect 232410 691540 232470 691600
rect 232500 691540 232560 691600
rect 232590 691540 232650 691600
rect 232680 691540 232740 691600
rect 232770 691540 232830 691600
rect 227370 691450 227430 691510
rect 227460 691450 227520 691510
rect 227550 691450 227610 691510
rect 227640 691450 227700 691510
rect 227730 691450 227790 691510
rect 227820 691450 227880 691510
rect 227910 691450 227970 691510
rect 228000 691450 228060 691510
rect 228090 691450 228150 691510
rect 228180 691450 228240 691510
rect 228270 691450 228330 691510
rect 228360 691450 228420 691510
rect 228450 691450 228510 691510
rect 228540 691450 228600 691510
rect 228630 691450 228690 691510
rect 228720 691450 228780 691510
rect 228810 691450 228870 691510
rect 228900 691450 228960 691510
rect 228990 691450 229050 691510
rect 229080 691450 229140 691510
rect 229170 691450 229230 691510
rect 229260 691450 229320 691510
rect 229350 691450 229410 691510
rect 229440 691450 229500 691510
rect 229530 691450 229590 691510
rect 229620 691450 229680 691510
rect 229710 691450 229770 691510
rect 229800 691450 229860 691510
rect 229890 691450 229950 691510
rect 229980 691450 230040 691510
rect 230070 691450 230130 691510
rect 230160 691450 230220 691510
rect 230250 691450 230310 691510
rect 230340 691450 230400 691510
rect 230430 691450 230490 691510
rect 230520 691450 230580 691510
rect 230610 691450 230670 691510
rect 230700 691450 230760 691510
rect 230790 691450 230850 691510
rect 230880 691450 230940 691510
rect 230970 691450 231030 691510
rect 231060 691450 231120 691510
rect 231150 691450 231210 691510
rect 231240 691450 231300 691510
rect 231330 691450 231390 691510
rect 231420 691450 231480 691510
rect 231510 691450 231570 691510
rect 231600 691450 231660 691510
rect 231690 691450 231750 691510
rect 231780 691450 231840 691510
rect 231870 691450 231930 691510
rect 231960 691450 232020 691510
rect 232050 691450 232110 691510
rect 232140 691450 232200 691510
rect 232230 691450 232290 691510
rect 232320 691450 232380 691510
rect 232410 691450 232470 691510
rect 232500 691450 232560 691510
rect 232590 691450 232650 691510
rect 232680 691450 232740 691510
rect 232770 691450 232830 691510
rect 227370 691360 227430 691420
rect 227460 691360 227520 691420
rect 227550 691360 227610 691420
rect 227640 691360 227700 691420
rect 227730 691360 227790 691420
rect 227820 691360 227880 691420
rect 227910 691360 227970 691420
rect 228000 691360 228060 691420
rect 228090 691360 228150 691420
rect 228180 691360 228240 691420
rect 228270 691360 228330 691420
rect 228360 691360 228420 691420
rect 228450 691360 228510 691420
rect 228540 691360 228600 691420
rect 228630 691360 228690 691420
rect 228720 691360 228780 691420
rect 228810 691360 228870 691420
rect 228900 691360 228960 691420
rect 228990 691360 229050 691420
rect 229080 691360 229140 691420
rect 229170 691360 229230 691420
rect 229260 691360 229320 691420
rect 229350 691360 229410 691420
rect 229440 691360 229500 691420
rect 229530 691360 229590 691420
rect 229620 691360 229680 691420
rect 229710 691360 229770 691420
rect 229800 691360 229860 691420
rect 229890 691360 229950 691420
rect 229980 691360 230040 691420
rect 230070 691360 230130 691420
rect 230160 691360 230220 691420
rect 230250 691360 230310 691420
rect 230340 691360 230400 691420
rect 230430 691360 230490 691420
rect 230520 691360 230580 691420
rect 230610 691360 230670 691420
rect 230700 691360 230760 691420
rect 230790 691360 230850 691420
rect 230880 691360 230940 691420
rect 230970 691360 231030 691420
rect 231060 691360 231120 691420
rect 231150 691360 231210 691420
rect 231240 691360 231300 691420
rect 231330 691360 231390 691420
rect 231420 691360 231480 691420
rect 231510 691360 231570 691420
rect 231600 691360 231660 691420
rect 231690 691360 231750 691420
rect 231780 691360 231840 691420
rect 231870 691360 231930 691420
rect 231960 691360 232020 691420
rect 232050 691360 232110 691420
rect 232140 691360 232200 691420
rect 232230 691360 232290 691420
rect 232320 691360 232380 691420
rect 232410 691360 232470 691420
rect 232500 691360 232560 691420
rect 232590 691360 232650 691420
rect 232680 691360 232740 691420
rect 232770 691360 232830 691420
rect 165620 690000 165690 690070
rect 165720 690000 165790 690070
rect 165820 690000 165890 690070
rect 165920 690000 165990 690070
rect 166020 690000 166090 690070
rect 166120 690000 166190 690070
rect 166220 690000 166290 690070
rect 166320 690000 166390 690070
rect 166420 690000 166490 690070
rect 166520 690000 166590 690070
rect 166620 690000 166690 690070
rect 166720 690000 166790 690070
rect 166820 690000 166890 690070
rect 166920 690000 166990 690070
rect 167020 690000 167090 690070
rect 167120 690000 167190 690070
rect 167220 690000 167290 690070
rect 167320 690000 167390 690070
rect 167420 690000 167490 690070
rect 167520 690000 167590 690070
rect 167620 690000 167690 690070
rect 167720 690000 167790 690070
rect 167820 690000 167890 690070
rect 167920 690000 167990 690070
rect 168020 690000 168090 690070
rect 168120 690000 168190 690070
rect 168220 690000 168290 690070
rect 168320 690000 168390 690070
rect 168420 690000 168490 690070
rect 168520 690000 168590 690070
rect 168620 690000 168690 690070
rect 168720 690000 168790 690070
rect 168820 690000 168890 690070
rect 168920 690000 168990 690070
rect 169020 690000 169090 690070
rect 169120 690000 169190 690070
rect 169220 690000 169290 690070
rect 169320 690000 169390 690070
rect 169420 690000 169490 690070
rect 169520 690000 169590 690070
rect 169620 690000 169690 690070
rect 169720 690000 169790 690070
rect 169820 690000 169890 690070
rect 169920 690000 169990 690070
rect 170020 690000 170090 690070
rect 170120 690000 170190 690070
rect 170220 690000 170290 690070
rect 170320 690000 170390 690070
rect 170420 690000 170490 690070
rect 165620 689900 165690 689970
rect 165720 689900 165790 689970
rect 165820 689900 165890 689970
rect 165920 689900 165990 689970
rect 166020 689900 166090 689970
rect 166120 689900 166190 689970
rect 166220 689900 166290 689970
rect 166320 689900 166390 689970
rect 166420 689900 166490 689970
rect 166520 689900 166590 689970
rect 166620 689900 166690 689970
rect 166720 689900 166790 689970
rect 166820 689900 166890 689970
rect 166920 689900 166990 689970
rect 167020 689900 167090 689970
rect 167120 689900 167190 689970
rect 167220 689900 167290 689970
rect 167320 689900 167390 689970
rect 167420 689900 167490 689970
rect 167520 689900 167590 689970
rect 167620 689900 167690 689970
rect 167720 689900 167790 689970
rect 167820 689900 167890 689970
rect 167920 689900 167990 689970
rect 168020 689900 168090 689970
rect 168120 689900 168190 689970
rect 168220 689900 168290 689970
rect 168320 689900 168390 689970
rect 168420 689900 168490 689970
rect 168520 689900 168590 689970
rect 168620 689900 168690 689970
rect 168720 689900 168790 689970
rect 168820 689900 168890 689970
rect 168920 689900 168990 689970
rect 169020 689900 169090 689970
rect 169120 689900 169190 689970
rect 169220 689900 169290 689970
rect 169320 689900 169390 689970
rect 169420 689900 169490 689970
rect 169520 689900 169590 689970
rect 169620 689900 169690 689970
rect 169720 689900 169790 689970
rect 169820 689900 169890 689970
rect 169920 689900 169990 689970
rect 170020 689900 170090 689970
rect 170120 689900 170190 689970
rect 170220 689900 170290 689970
rect 170320 689900 170390 689970
rect 170420 689900 170490 689970
rect 227640 689990 227710 690060
rect 227740 689990 227810 690060
rect 227840 689990 227910 690060
rect 227940 689990 228010 690060
rect 228040 689990 228110 690060
rect 228140 689990 228210 690060
rect 228240 689990 228310 690060
rect 228340 689990 228410 690060
rect 228440 689990 228510 690060
rect 228540 689990 228610 690060
rect 228640 689990 228710 690060
rect 228740 689990 228810 690060
rect 228840 689990 228910 690060
rect 228940 689990 229010 690060
rect 229040 689990 229110 690060
rect 229140 689990 229210 690060
rect 229240 689990 229310 690060
rect 229340 689990 229410 690060
rect 229440 689990 229510 690060
rect 229540 689990 229610 690060
rect 229640 689990 229710 690060
rect 229740 689990 229810 690060
rect 229840 689990 229910 690060
rect 229940 689990 230010 690060
rect 230040 689990 230110 690060
rect 230140 689990 230210 690060
rect 230240 689990 230310 690060
rect 230340 689990 230410 690060
rect 230440 689990 230510 690060
rect 230540 689990 230610 690060
rect 230640 689990 230710 690060
rect 230740 689990 230810 690060
rect 230840 689990 230910 690060
rect 230940 689990 231010 690060
rect 231040 689990 231110 690060
rect 231140 689990 231210 690060
rect 231240 689990 231310 690060
rect 231340 689990 231410 690060
rect 231440 689990 231510 690060
rect 231540 689990 231610 690060
rect 231640 689990 231710 690060
rect 231740 689990 231810 690060
rect 231840 689990 231910 690060
rect 231940 689990 232010 690060
rect 232040 689990 232110 690060
rect 232140 689990 232210 690060
rect 232240 689990 232310 690060
rect 232340 689990 232410 690060
rect 232440 689990 232510 690060
rect 227640 689890 227710 689960
rect 227740 689890 227810 689960
rect 227840 689890 227910 689960
rect 227940 689890 228010 689960
rect 228040 689890 228110 689960
rect 228140 689890 228210 689960
rect 228240 689890 228310 689960
rect 228340 689890 228410 689960
rect 228440 689890 228510 689960
rect 228540 689890 228610 689960
rect 228640 689890 228710 689960
rect 228740 689890 228810 689960
rect 228840 689890 228910 689960
rect 228940 689890 229010 689960
rect 229040 689890 229110 689960
rect 229140 689890 229210 689960
rect 229240 689890 229310 689960
rect 229340 689890 229410 689960
rect 229440 689890 229510 689960
rect 229540 689890 229610 689960
rect 229640 689890 229710 689960
rect 229740 689890 229810 689960
rect 229840 689890 229910 689960
rect 229940 689890 230010 689960
rect 230040 689890 230110 689960
rect 230140 689890 230210 689960
rect 230240 689890 230310 689960
rect 230340 689890 230410 689960
rect 230440 689890 230510 689960
rect 230540 689890 230610 689960
rect 230640 689890 230710 689960
rect 230740 689890 230810 689960
rect 230840 689890 230910 689960
rect 230940 689890 231010 689960
rect 231040 689890 231110 689960
rect 231140 689890 231210 689960
rect 231240 689890 231310 689960
rect 231340 689890 231410 689960
rect 231440 689890 231510 689960
rect 231540 689890 231610 689960
rect 231640 689890 231710 689960
rect 231740 689890 231810 689960
rect 231840 689890 231910 689960
rect 231940 689890 232010 689960
rect 232040 689890 232110 689960
rect 232140 689890 232210 689960
rect 232240 689890 232310 689960
rect 232340 689890 232410 689960
rect 232440 689890 232510 689960
<< metal2 >>
rect 165334 691580 170828 691635
rect 165334 691510 165360 691580
rect 165430 691510 165460 691580
rect 165530 691510 165560 691580
rect 165630 691510 165660 691580
rect 165730 691510 165760 691580
rect 165830 691510 165860 691580
rect 165930 691510 165960 691580
rect 166030 691510 166060 691580
rect 166130 691510 166160 691580
rect 166230 691510 166260 691580
rect 166330 691510 166360 691580
rect 166430 691510 166460 691580
rect 166530 691510 166560 691580
rect 166630 691510 166660 691580
rect 166730 691510 166760 691580
rect 166830 691510 166860 691580
rect 166930 691510 166960 691580
rect 167030 691510 167060 691580
rect 167130 691510 167160 691580
rect 167230 691510 167260 691580
rect 167330 691510 167360 691580
rect 167430 691510 167460 691580
rect 167530 691510 167560 691580
rect 167630 691510 167660 691580
rect 167730 691510 167760 691580
rect 167830 691510 167860 691580
rect 167930 691510 167960 691580
rect 168030 691510 168060 691580
rect 168130 691510 168160 691580
rect 168230 691510 168260 691580
rect 168330 691510 168360 691580
rect 168430 691510 168460 691580
rect 168530 691510 168560 691580
rect 168630 691510 168660 691580
rect 168730 691510 168760 691580
rect 168830 691510 168860 691580
rect 168930 691510 168960 691580
rect 169030 691510 169060 691580
rect 169130 691510 169160 691580
rect 169230 691510 169260 691580
rect 169330 691510 169360 691580
rect 169430 691510 169460 691580
rect 169530 691510 169560 691580
rect 169630 691510 169660 691580
rect 169730 691510 169760 691580
rect 169830 691510 169860 691580
rect 169930 691510 169960 691580
rect 170030 691510 170060 691580
rect 170130 691510 170160 691580
rect 170230 691510 170260 691580
rect 170330 691510 170360 691580
rect 170430 691510 170460 691580
rect 170530 691510 170828 691580
rect 165334 691470 170828 691510
rect 165334 691400 165360 691470
rect 165430 691400 165460 691470
rect 165530 691400 165560 691470
rect 165630 691400 165660 691470
rect 165730 691400 165760 691470
rect 165830 691400 165860 691470
rect 165930 691400 165960 691470
rect 166030 691400 166060 691470
rect 166130 691400 166160 691470
rect 166230 691400 166260 691470
rect 166330 691400 166360 691470
rect 166430 691400 166460 691470
rect 166530 691400 166560 691470
rect 166630 691400 166660 691470
rect 166730 691400 166760 691470
rect 166830 691400 166860 691470
rect 166930 691400 166960 691470
rect 167030 691400 167060 691470
rect 167130 691400 167160 691470
rect 167230 691400 167260 691470
rect 167330 691400 167360 691470
rect 167430 691400 167460 691470
rect 167530 691400 167560 691470
rect 167630 691400 167660 691470
rect 167730 691400 167760 691470
rect 167830 691400 167860 691470
rect 167930 691400 167960 691470
rect 168030 691400 168060 691470
rect 168130 691400 168160 691470
rect 168230 691400 168260 691470
rect 168330 691400 168360 691470
rect 168430 691400 168460 691470
rect 168530 691400 168560 691470
rect 168630 691400 168660 691470
rect 168730 691400 168760 691470
rect 168830 691400 168860 691470
rect 168930 691400 168960 691470
rect 169030 691400 169060 691470
rect 169130 691400 169160 691470
rect 169230 691400 169260 691470
rect 169330 691400 169360 691470
rect 169430 691400 169460 691470
rect 169530 691400 169560 691470
rect 169630 691400 169660 691470
rect 169730 691400 169760 691470
rect 169830 691400 169860 691470
rect 169930 691400 169960 691470
rect 170030 691400 170060 691470
rect 170130 691400 170160 691470
rect 170230 691400 170260 691470
rect 170330 691400 170360 691470
rect 170430 691400 170460 691470
rect 170530 691400 170828 691470
rect 165334 691360 170828 691400
rect 227356 691600 232850 691626
rect 227356 691540 227370 691600
rect 227430 691540 227460 691600
rect 227520 691540 227550 691600
rect 227610 691540 227640 691600
rect 227700 691540 227730 691600
rect 227790 691540 227820 691600
rect 227880 691540 227910 691600
rect 227970 691540 228000 691600
rect 228060 691540 228090 691600
rect 228150 691540 228180 691600
rect 228240 691540 228270 691600
rect 228330 691540 228360 691600
rect 228420 691540 228450 691600
rect 228510 691540 228540 691600
rect 228600 691540 228630 691600
rect 228690 691540 228720 691600
rect 228780 691540 228810 691600
rect 228870 691540 228900 691600
rect 228960 691540 228990 691600
rect 229050 691540 229080 691600
rect 229140 691540 229170 691600
rect 229230 691540 229260 691600
rect 229320 691540 229350 691600
rect 229410 691540 229440 691600
rect 229500 691540 229530 691600
rect 229590 691540 229620 691600
rect 229680 691540 229710 691600
rect 229770 691540 229800 691600
rect 229860 691540 229890 691600
rect 229950 691540 229980 691600
rect 230040 691540 230070 691600
rect 230130 691540 230160 691600
rect 230220 691540 230250 691600
rect 230310 691540 230340 691600
rect 230400 691540 230430 691600
rect 230490 691540 230520 691600
rect 230580 691540 230610 691600
rect 230670 691540 230700 691600
rect 230760 691540 230790 691600
rect 230850 691540 230880 691600
rect 230940 691540 230970 691600
rect 231030 691540 231060 691600
rect 231120 691540 231150 691600
rect 231210 691540 231240 691600
rect 231300 691540 231330 691600
rect 231390 691540 231420 691600
rect 231480 691540 231510 691600
rect 231570 691540 231600 691600
rect 231660 691540 231690 691600
rect 231750 691540 231780 691600
rect 231840 691540 231870 691600
rect 231930 691540 231960 691600
rect 232020 691540 232050 691600
rect 232110 691540 232140 691600
rect 232200 691540 232230 691600
rect 232290 691540 232320 691600
rect 232380 691540 232410 691600
rect 232470 691540 232500 691600
rect 232560 691540 232590 691600
rect 232650 691540 232680 691600
rect 232740 691540 232770 691600
rect 232830 691540 232850 691600
rect 227356 691510 232850 691540
rect 227356 691450 227370 691510
rect 227430 691450 227460 691510
rect 227520 691450 227550 691510
rect 227610 691450 227640 691510
rect 227700 691450 227730 691510
rect 227790 691450 227820 691510
rect 227880 691450 227910 691510
rect 227970 691450 228000 691510
rect 228060 691450 228090 691510
rect 228150 691450 228180 691510
rect 228240 691450 228270 691510
rect 228330 691450 228360 691510
rect 228420 691450 228450 691510
rect 228510 691450 228540 691510
rect 228600 691450 228630 691510
rect 228690 691450 228720 691510
rect 228780 691450 228810 691510
rect 228870 691450 228900 691510
rect 228960 691450 228990 691510
rect 229050 691450 229080 691510
rect 229140 691450 229170 691510
rect 229230 691450 229260 691510
rect 229320 691450 229350 691510
rect 229410 691450 229440 691510
rect 229500 691450 229530 691510
rect 229590 691450 229620 691510
rect 229680 691450 229710 691510
rect 229770 691450 229800 691510
rect 229860 691450 229890 691510
rect 229950 691450 229980 691510
rect 230040 691450 230070 691510
rect 230130 691450 230160 691510
rect 230220 691450 230250 691510
rect 230310 691450 230340 691510
rect 230400 691450 230430 691510
rect 230490 691450 230520 691510
rect 230580 691450 230610 691510
rect 230670 691450 230700 691510
rect 230760 691450 230790 691510
rect 230850 691450 230880 691510
rect 230940 691450 230970 691510
rect 231030 691450 231060 691510
rect 231120 691450 231150 691510
rect 231210 691450 231240 691510
rect 231300 691450 231330 691510
rect 231390 691450 231420 691510
rect 231480 691450 231510 691510
rect 231570 691450 231600 691510
rect 231660 691450 231690 691510
rect 231750 691450 231780 691510
rect 231840 691450 231870 691510
rect 231930 691450 231960 691510
rect 232020 691450 232050 691510
rect 232110 691450 232140 691510
rect 232200 691450 232230 691510
rect 232290 691450 232320 691510
rect 232380 691450 232410 691510
rect 232470 691450 232500 691510
rect 232560 691450 232590 691510
rect 232650 691450 232680 691510
rect 232740 691450 232770 691510
rect 232830 691450 232850 691510
rect 227356 691420 232850 691450
rect 227356 691360 227370 691420
rect 227430 691360 227460 691420
rect 227520 691360 227550 691420
rect 227610 691360 227640 691420
rect 227700 691360 227730 691420
rect 227790 691360 227820 691420
rect 227880 691360 227910 691420
rect 227970 691360 228000 691420
rect 228060 691360 228090 691420
rect 228150 691360 228180 691420
rect 228240 691360 228270 691420
rect 228330 691360 228360 691420
rect 228420 691360 228450 691420
rect 228510 691360 228540 691420
rect 228600 691360 228630 691420
rect 228690 691360 228720 691420
rect 228780 691360 228810 691420
rect 228870 691360 228900 691420
rect 228960 691360 228990 691420
rect 229050 691360 229080 691420
rect 229140 691360 229170 691420
rect 229230 691360 229260 691420
rect 229320 691360 229350 691420
rect 229410 691360 229440 691420
rect 229500 691360 229530 691420
rect 229590 691360 229620 691420
rect 229680 691360 229710 691420
rect 229770 691360 229800 691420
rect 229860 691360 229890 691420
rect 229950 691360 229980 691420
rect 230040 691360 230070 691420
rect 230130 691360 230160 691420
rect 230220 691360 230250 691420
rect 230310 691360 230340 691420
rect 230400 691360 230430 691420
rect 230490 691360 230520 691420
rect 230580 691360 230610 691420
rect 230670 691360 230700 691420
rect 230760 691360 230790 691420
rect 230850 691360 230880 691420
rect 230940 691360 230970 691420
rect 231030 691360 231060 691420
rect 231120 691360 231150 691420
rect 231210 691360 231240 691420
rect 231300 691360 231330 691420
rect 231390 691360 231420 691420
rect 231480 691360 231510 691420
rect 231570 691360 231600 691420
rect 231660 691360 231690 691420
rect 231750 691360 231780 691420
rect 231840 691360 231870 691420
rect 231930 691360 231960 691420
rect 232020 691360 232050 691420
rect 232110 691360 232140 691420
rect 232200 691360 232230 691420
rect 232290 691360 232320 691420
rect 232380 691360 232410 691420
rect 232470 691360 232500 691420
rect 232560 691360 232590 691420
rect 232650 691360 232680 691420
rect 232740 691360 232770 691420
rect 232830 691360 232850 691420
rect 227356 691351 232850 691360
rect 165364 690070 170798 690104
rect 165364 690000 165620 690070
rect 165690 690000 165720 690070
rect 165790 690000 165820 690070
rect 165890 690000 165920 690070
rect 165990 690000 166020 690070
rect 166090 690000 166120 690070
rect 166190 690000 166220 690070
rect 166290 690000 166320 690070
rect 166390 690000 166420 690070
rect 166490 690000 166520 690070
rect 166590 690000 166620 690070
rect 166690 690000 166720 690070
rect 166790 690000 166820 690070
rect 166890 690000 166920 690070
rect 166990 690000 167020 690070
rect 167090 690000 167120 690070
rect 167190 690000 167220 690070
rect 167290 690000 167320 690070
rect 167390 690000 167420 690070
rect 167490 690000 167520 690070
rect 167590 690000 167620 690070
rect 167690 690000 167720 690070
rect 167790 690000 167820 690070
rect 167890 690000 167920 690070
rect 167990 690000 168020 690070
rect 168090 690000 168120 690070
rect 168190 690000 168220 690070
rect 168290 690000 168320 690070
rect 168390 690000 168420 690070
rect 168490 690000 168520 690070
rect 168590 690000 168620 690070
rect 168690 690000 168720 690070
rect 168790 690000 168820 690070
rect 168890 690000 168920 690070
rect 168990 690000 169020 690070
rect 169090 690000 169120 690070
rect 169190 690000 169220 690070
rect 169290 690000 169320 690070
rect 169390 690000 169420 690070
rect 169490 690000 169520 690070
rect 169590 690000 169620 690070
rect 169690 690000 169720 690070
rect 169790 690000 169820 690070
rect 169890 690000 169920 690070
rect 169990 690000 170020 690070
rect 170090 690000 170120 690070
rect 170190 690000 170220 690070
rect 170290 690000 170320 690070
rect 170390 690000 170420 690070
rect 170490 690000 170798 690070
rect 165364 689970 170798 690000
rect 165364 689900 165620 689970
rect 165690 689900 165720 689970
rect 165790 689900 165820 689970
rect 165890 689900 165920 689970
rect 165990 689900 166020 689970
rect 166090 689900 166120 689970
rect 166190 689900 166220 689970
rect 166290 689900 166320 689970
rect 166390 689900 166420 689970
rect 166490 689900 166520 689970
rect 166590 689900 166620 689970
rect 166690 689900 166720 689970
rect 166790 689900 166820 689970
rect 166890 689900 166920 689970
rect 166990 689900 167020 689970
rect 167090 689900 167120 689970
rect 167190 689900 167220 689970
rect 167290 689900 167320 689970
rect 167390 689900 167420 689970
rect 167490 689900 167520 689970
rect 167590 689900 167620 689970
rect 167690 689900 167720 689970
rect 167790 689900 167820 689970
rect 167890 689900 167920 689970
rect 167990 689900 168020 689970
rect 168090 689900 168120 689970
rect 168190 689900 168220 689970
rect 168290 689900 168320 689970
rect 168390 689900 168420 689970
rect 168490 689900 168520 689970
rect 168590 689900 168620 689970
rect 168690 689900 168720 689970
rect 168790 689900 168820 689970
rect 168890 689900 168920 689970
rect 168990 689900 169020 689970
rect 169090 689900 169120 689970
rect 169190 689900 169220 689970
rect 169290 689900 169320 689970
rect 169390 689900 169420 689970
rect 169490 689900 169520 689970
rect 169590 689900 169620 689970
rect 169690 689900 169720 689970
rect 169790 689900 169820 689970
rect 169890 689900 169920 689970
rect 169990 689900 170020 689970
rect 170090 689900 170120 689970
rect 170190 689900 170220 689970
rect 170290 689900 170320 689970
rect 170390 689900 170420 689970
rect 170490 689900 170798 689970
rect 165364 689877 170798 689900
rect 227386 690060 232820 690114
rect 227386 689990 227640 690060
rect 227710 689990 227740 690060
rect 227810 689990 227840 690060
rect 227910 689990 227940 690060
rect 228010 689990 228040 690060
rect 228110 689990 228140 690060
rect 228210 689990 228240 690060
rect 228310 689990 228340 690060
rect 228410 689990 228440 690060
rect 228510 689990 228540 690060
rect 228610 689990 228640 690060
rect 228710 689990 228740 690060
rect 228810 689990 228840 690060
rect 228910 689990 228940 690060
rect 229010 689990 229040 690060
rect 229110 689990 229140 690060
rect 229210 689990 229240 690060
rect 229310 689990 229340 690060
rect 229410 689990 229440 690060
rect 229510 689990 229540 690060
rect 229610 689990 229640 690060
rect 229710 689990 229740 690060
rect 229810 689990 229840 690060
rect 229910 689990 229940 690060
rect 230010 689990 230040 690060
rect 230110 689990 230140 690060
rect 230210 689990 230240 690060
rect 230310 689990 230340 690060
rect 230410 689990 230440 690060
rect 230510 689990 230540 690060
rect 230610 689990 230640 690060
rect 230710 689990 230740 690060
rect 230810 689990 230840 690060
rect 230910 689990 230940 690060
rect 231010 689990 231040 690060
rect 231110 689990 231140 690060
rect 231210 689990 231240 690060
rect 231310 689990 231340 690060
rect 231410 689990 231440 690060
rect 231510 689990 231540 690060
rect 231610 689990 231640 690060
rect 231710 689990 231740 690060
rect 231810 689990 231840 690060
rect 231910 689990 231940 690060
rect 232010 689990 232040 690060
rect 232110 689990 232140 690060
rect 232210 689990 232240 690060
rect 232310 689990 232340 690060
rect 232410 689990 232440 690060
rect 232510 689990 232820 690060
rect 227386 689960 232820 689990
rect 227386 689890 227640 689960
rect 227710 689890 227740 689960
rect 227810 689890 227840 689960
rect 227910 689890 227940 689960
rect 228010 689890 228040 689960
rect 228110 689890 228140 689960
rect 228210 689890 228240 689960
rect 228310 689890 228340 689960
rect 228410 689890 228440 689960
rect 228510 689890 228540 689960
rect 228610 689890 228640 689960
rect 228710 689890 228740 689960
rect 228810 689890 228840 689960
rect 228910 689890 228940 689960
rect 229010 689890 229040 689960
rect 229110 689890 229140 689960
rect 229210 689890 229240 689960
rect 229310 689890 229340 689960
rect 229410 689890 229440 689960
rect 229510 689890 229540 689960
rect 229610 689890 229640 689960
rect 229710 689890 229740 689960
rect 229810 689890 229840 689960
rect 229910 689890 229940 689960
rect 230010 689890 230040 689960
rect 230110 689890 230140 689960
rect 230210 689890 230240 689960
rect 230310 689890 230340 689960
rect 230410 689890 230440 689960
rect 230510 689890 230540 689960
rect 230610 689890 230640 689960
rect 230710 689890 230740 689960
rect 230810 689890 230840 689960
rect 230910 689890 230940 689960
rect 231010 689890 231040 689960
rect 231110 689890 231140 689960
rect 231210 689890 231240 689960
rect 231310 689890 231340 689960
rect 231410 689890 231440 689960
rect 231510 689890 231540 689960
rect 231610 689890 231640 689960
rect 231710 689890 231740 689960
rect 231810 689890 231840 689960
rect 231910 689890 231940 689960
rect 232010 689890 232040 689960
rect 232110 689890 232140 689960
rect 232210 689890 232240 689960
rect 232310 689890 232340 689960
rect 232410 689890 232440 689960
rect 232510 689890 232820 689960
rect 227386 689853 232820 689890
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 165360 691510 165430 691580
rect 165460 691510 165530 691580
rect 165560 691510 165630 691580
rect 165660 691510 165730 691580
rect 165760 691510 165830 691580
rect 165860 691510 165930 691580
rect 165960 691510 166030 691580
rect 166060 691510 166130 691580
rect 166160 691510 166230 691580
rect 166260 691510 166330 691580
rect 166360 691510 166430 691580
rect 166460 691510 166530 691580
rect 166560 691510 166630 691580
rect 166660 691510 166730 691580
rect 166760 691510 166830 691580
rect 166860 691510 166930 691580
rect 166960 691510 167030 691580
rect 167060 691510 167130 691580
rect 167160 691510 167230 691580
rect 167260 691510 167330 691580
rect 167360 691510 167430 691580
rect 167460 691510 167530 691580
rect 167560 691510 167630 691580
rect 167660 691510 167730 691580
rect 167760 691510 167830 691580
rect 167860 691510 167930 691580
rect 167960 691510 168030 691580
rect 168060 691510 168130 691580
rect 168160 691510 168230 691580
rect 168260 691510 168330 691580
rect 168360 691510 168430 691580
rect 168460 691510 168530 691580
rect 168560 691510 168630 691580
rect 168660 691510 168730 691580
rect 168760 691510 168830 691580
rect 168860 691510 168930 691580
rect 168960 691510 169030 691580
rect 169060 691510 169130 691580
rect 169160 691510 169230 691580
rect 169260 691510 169330 691580
rect 169360 691510 169430 691580
rect 169460 691510 169530 691580
rect 169560 691510 169630 691580
rect 169660 691510 169730 691580
rect 169760 691510 169830 691580
rect 169860 691510 169930 691580
rect 169960 691510 170030 691580
rect 170060 691510 170130 691580
rect 170160 691510 170230 691580
rect 170260 691510 170330 691580
rect 170360 691510 170430 691580
rect 170460 691510 170530 691580
rect 165360 691400 165430 691470
rect 165460 691400 165530 691470
rect 165560 691400 165630 691470
rect 165660 691400 165730 691470
rect 165760 691400 165830 691470
rect 165860 691400 165930 691470
rect 165960 691400 166030 691470
rect 166060 691400 166130 691470
rect 166160 691400 166230 691470
rect 166260 691400 166330 691470
rect 166360 691400 166430 691470
rect 166460 691400 166530 691470
rect 166560 691400 166630 691470
rect 166660 691400 166730 691470
rect 166760 691400 166830 691470
rect 166860 691400 166930 691470
rect 166960 691400 167030 691470
rect 167060 691400 167130 691470
rect 167160 691400 167230 691470
rect 167260 691400 167330 691470
rect 167360 691400 167430 691470
rect 167460 691400 167530 691470
rect 167560 691400 167630 691470
rect 167660 691400 167730 691470
rect 167760 691400 167830 691470
rect 167860 691400 167930 691470
rect 167960 691400 168030 691470
rect 168060 691400 168130 691470
rect 168160 691400 168230 691470
rect 168260 691400 168330 691470
rect 168360 691400 168430 691470
rect 168460 691400 168530 691470
rect 168560 691400 168630 691470
rect 168660 691400 168730 691470
rect 168760 691400 168830 691470
rect 168860 691400 168930 691470
rect 168960 691400 169030 691470
rect 169060 691400 169130 691470
rect 169160 691400 169230 691470
rect 169260 691400 169330 691470
rect 169360 691400 169430 691470
rect 169460 691400 169530 691470
rect 169560 691400 169630 691470
rect 169660 691400 169730 691470
rect 169760 691400 169830 691470
rect 169860 691400 169930 691470
rect 169960 691400 170030 691470
rect 170060 691400 170130 691470
rect 170160 691400 170230 691470
rect 170260 691400 170330 691470
rect 170360 691400 170430 691470
rect 170460 691400 170530 691470
rect 227370 691540 227430 691600
rect 227460 691540 227520 691600
rect 227550 691540 227610 691600
rect 227640 691540 227700 691600
rect 227730 691540 227790 691600
rect 227820 691540 227880 691600
rect 227910 691540 227970 691600
rect 228000 691540 228060 691600
rect 228090 691540 228150 691600
rect 228180 691540 228240 691600
rect 228270 691540 228330 691600
rect 228360 691540 228420 691600
rect 228450 691540 228510 691600
rect 228540 691540 228600 691600
rect 228630 691540 228690 691600
rect 228720 691540 228780 691600
rect 228810 691540 228870 691600
rect 228900 691540 228960 691600
rect 228990 691540 229050 691600
rect 229080 691540 229140 691600
rect 229170 691540 229230 691600
rect 229260 691540 229320 691600
rect 229350 691540 229410 691600
rect 229440 691540 229500 691600
rect 229530 691540 229590 691600
rect 229620 691540 229680 691600
rect 229710 691540 229770 691600
rect 229800 691540 229860 691600
rect 229890 691540 229950 691600
rect 229980 691540 230040 691600
rect 230070 691540 230130 691600
rect 230160 691540 230220 691600
rect 230250 691540 230310 691600
rect 230340 691540 230400 691600
rect 230430 691540 230490 691600
rect 230520 691540 230580 691600
rect 230610 691540 230670 691600
rect 230700 691540 230760 691600
rect 230790 691540 230850 691600
rect 230880 691540 230940 691600
rect 230970 691540 231030 691600
rect 231060 691540 231120 691600
rect 231150 691540 231210 691600
rect 231240 691540 231300 691600
rect 231330 691540 231390 691600
rect 231420 691540 231480 691600
rect 231510 691540 231570 691600
rect 231600 691540 231660 691600
rect 231690 691540 231750 691600
rect 231780 691540 231840 691600
rect 231870 691540 231930 691600
rect 231960 691540 232020 691600
rect 232050 691540 232110 691600
rect 232140 691540 232200 691600
rect 232230 691540 232290 691600
rect 232320 691540 232380 691600
rect 232410 691540 232470 691600
rect 232500 691540 232560 691600
rect 232590 691540 232650 691600
rect 232680 691540 232740 691600
rect 232770 691540 232830 691600
rect 227370 691450 227430 691510
rect 227460 691450 227520 691510
rect 227550 691450 227610 691510
rect 227640 691450 227700 691510
rect 227730 691450 227790 691510
rect 227820 691450 227880 691510
rect 227910 691450 227970 691510
rect 228000 691450 228060 691510
rect 228090 691450 228150 691510
rect 228180 691450 228240 691510
rect 228270 691450 228330 691510
rect 228360 691450 228420 691510
rect 228450 691450 228510 691510
rect 228540 691450 228600 691510
rect 228630 691450 228690 691510
rect 228720 691450 228780 691510
rect 228810 691450 228870 691510
rect 228900 691450 228960 691510
rect 228990 691450 229050 691510
rect 229080 691450 229140 691510
rect 229170 691450 229230 691510
rect 229260 691450 229320 691510
rect 229350 691450 229410 691510
rect 229440 691450 229500 691510
rect 229530 691450 229590 691510
rect 229620 691450 229680 691510
rect 229710 691450 229770 691510
rect 229800 691450 229860 691510
rect 229890 691450 229950 691510
rect 229980 691450 230040 691510
rect 230070 691450 230130 691510
rect 230160 691450 230220 691510
rect 230250 691450 230310 691510
rect 230340 691450 230400 691510
rect 230430 691450 230490 691510
rect 230520 691450 230580 691510
rect 230610 691450 230670 691510
rect 230700 691450 230760 691510
rect 230790 691450 230850 691510
rect 230880 691450 230940 691510
rect 230970 691450 231030 691510
rect 231060 691450 231120 691510
rect 231150 691450 231210 691510
rect 231240 691450 231300 691510
rect 231330 691450 231390 691510
rect 231420 691450 231480 691510
rect 231510 691450 231570 691510
rect 231600 691450 231660 691510
rect 231690 691450 231750 691510
rect 231780 691450 231840 691510
rect 231870 691450 231930 691510
rect 231960 691450 232020 691510
rect 232050 691450 232110 691510
rect 232140 691450 232200 691510
rect 232230 691450 232290 691510
rect 232320 691450 232380 691510
rect 232410 691450 232470 691510
rect 232500 691450 232560 691510
rect 232590 691450 232650 691510
rect 232680 691450 232740 691510
rect 232770 691450 232830 691510
rect 227370 691360 227430 691420
rect 227460 691360 227520 691420
rect 227550 691360 227610 691420
rect 227640 691360 227700 691420
rect 227730 691360 227790 691420
rect 227820 691360 227880 691420
rect 227910 691360 227970 691420
rect 228000 691360 228060 691420
rect 228090 691360 228150 691420
rect 228180 691360 228240 691420
rect 228270 691360 228330 691420
rect 228360 691360 228420 691420
rect 228450 691360 228510 691420
rect 228540 691360 228600 691420
rect 228630 691360 228690 691420
rect 228720 691360 228780 691420
rect 228810 691360 228870 691420
rect 228900 691360 228960 691420
rect 228990 691360 229050 691420
rect 229080 691360 229140 691420
rect 229170 691360 229230 691420
rect 229260 691360 229320 691420
rect 229350 691360 229410 691420
rect 229440 691360 229500 691420
rect 229530 691360 229590 691420
rect 229620 691360 229680 691420
rect 229710 691360 229770 691420
rect 229800 691360 229860 691420
rect 229890 691360 229950 691420
rect 229980 691360 230040 691420
rect 230070 691360 230130 691420
rect 230160 691360 230220 691420
rect 230250 691360 230310 691420
rect 230340 691360 230400 691420
rect 230430 691360 230490 691420
rect 230520 691360 230580 691420
rect 230610 691360 230670 691420
rect 230700 691360 230760 691420
rect 230790 691360 230850 691420
rect 230880 691360 230940 691420
rect 230970 691360 231030 691420
rect 231060 691360 231120 691420
rect 231150 691360 231210 691420
rect 231240 691360 231300 691420
rect 231330 691360 231390 691420
rect 231420 691360 231480 691420
rect 231510 691360 231570 691420
rect 231600 691360 231660 691420
rect 231690 691360 231750 691420
rect 231780 691360 231840 691420
rect 231870 691360 231930 691420
rect 231960 691360 232020 691420
rect 232050 691360 232110 691420
rect 232140 691360 232200 691420
rect 232230 691360 232290 691420
rect 232320 691360 232380 691420
rect 232410 691360 232470 691420
rect 232500 691360 232560 691420
rect 232590 691360 232650 691420
rect 232680 691360 232740 691420
rect 232770 691360 232830 691420
rect 165620 690000 165690 690070
rect 165720 690000 165790 690070
rect 165820 690000 165890 690070
rect 165920 690000 165990 690070
rect 166020 690000 166090 690070
rect 166120 690000 166190 690070
rect 166220 690000 166290 690070
rect 166320 690000 166390 690070
rect 166420 690000 166490 690070
rect 166520 690000 166590 690070
rect 166620 690000 166690 690070
rect 166720 690000 166790 690070
rect 166820 690000 166890 690070
rect 166920 690000 166990 690070
rect 167020 690000 167090 690070
rect 167120 690000 167190 690070
rect 167220 690000 167290 690070
rect 167320 690000 167390 690070
rect 167420 690000 167490 690070
rect 167520 690000 167590 690070
rect 167620 690000 167690 690070
rect 167720 690000 167790 690070
rect 167820 690000 167890 690070
rect 167920 690000 167990 690070
rect 168020 690000 168090 690070
rect 168120 690000 168190 690070
rect 168220 690000 168290 690070
rect 168320 690000 168390 690070
rect 168420 690000 168490 690070
rect 168520 690000 168590 690070
rect 168620 690000 168690 690070
rect 168720 690000 168790 690070
rect 168820 690000 168890 690070
rect 168920 690000 168990 690070
rect 169020 690000 169090 690070
rect 169120 690000 169190 690070
rect 169220 690000 169290 690070
rect 169320 690000 169390 690070
rect 169420 690000 169490 690070
rect 169520 690000 169590 690070
rect 169620 690000 169690 690070
rect 169720 690000 169790 690070
rect 169820 690000 169890 690070
rect 169920 690000 169990 690070
rect 170020 690000 170090 690070
rect 170120 690000 170190 690070
rect 170220 690000 170290 690070
rect 170320 690000 170390 690070
rect 170420 690000 170490 690070
rect 165620 689900 165690 689970
rect 165720 689900 165790 689970
rect 165820 689900 165890 689970
rect 165920 689900 165990 689970
rect 166020 689900 166090 689970
rect 166120 689900 166190 689970
rect 166220 689900 166290 689970
rect 166320 689900 166390 689970
rect 166420 689900 166490 689970
rect 166520 689900 166590 689970
rect 166620 689900 166690 689970
rect 166720 689900 166790 689970
rect 166820 689900 166890 689970
rect 166920 689900 166990 689970
rect 167020 689900 167090 689970
rect 167120 689900 167190 689970
rect 167220 689900 167290 689970
rect 167320 689900 167390 689970
rect 167420 689900 167490 689970
rect 167520 689900 167590 689970
rect 167620 689900 167690 689970
rect 167720 689900 167790 689970
rect 167820 689900 167890 689970
rect 167920 689900 167990 689970
rect 168020 689900 168090 689970
rect 168120 689900 168190 689970
rect 168220 689900 168290 689970
rect 168320 689900 168390 689970
rect 168420 689900 168490 689970
rect 168520 689900 168590 689970
rect 168620 689900 168690 689970
rect 168720 689900 168790 689970
rect 168820 689900 168890 689970
rect 168920 689900 168990 689970
rect 169020 689900 169090 689970
rect 169120 689900 169190 689970
rect 169220 689900 169290 689970
rect 169320 689900 169390 689970
rect 169420 689900 169490 689970
rect 169520 689900 169590 689970
rect 169620 689900 169690 689970
rect 169720 689900 169790 689970
rect 169820 689900 169890 689970
rect 169920 689900 169990 689970
rect 170020 689900 170090 689970
rect 170120 689900 170190 689970
rect 170220 689900 170290 689970
rect 170320 689900 170390 689970
rect 170420 689900 170490 689970
rect 227640 689990 227710 690060
rect 227740 689990 227810 690060
rect 227840 689990 227910 690060
rect 227940 689990 228010 690060
rect 228040 689990 228110 690060
rect 228140 689990 228210 690060
rect 228240 689990 228310 690060
rect 228340 689990 228410 690060
rect 228440 689990 228510 690060
rect 228540 689990 228610 690060
rect 228640 689990 228710 690060
rect 228740 689990 228810 690060
rect 228840 689990 228910 690060
rect 228940 689990 229010 690060
rect 229040 689990 229110 690060
rect 229140 689990 229210 690060
rect 229240 689990 229310 690060
rect 229340 689990 229410 690060
rect 229440 689990 229510 690060
rect 229540 689990 229610 690060
rect 229640 689990 229710 690060
rect 229740 689990 229810 690060
rect 229840 689990 229910 690060
rect 229940 689990 230010 690060
rect 230040 689990 230110 690060
rect 230140 689990 230210 690060
rect 230240 689990 230310 690060
rect 230340 689990 230410 690060
rect 230440 689990 230510 690060
rect 230540 689990 230610 690060
rect 230640 689990 230710 690060
rect 230740 689990 230810 690060
rect 230840 689990 230910 690060
rect 230940 689990 231010 690060
rect 231040 689990 231110 690060
rect 231140 689990 231210 690060
rect 231240 689990 231310 690060
rect 231340 689990 231410 690060
rect 231440 689990 231510 690060
rect 231540 689990 231610 690060
rect 231640 689990 231710 690060
rect 231740 689990 231810 690060
rect 231840 689990 231910 690060
rect 231940 689990 232010 690060
rect 232040 689990 232110 690060
rect 232140 689990 232210 690060
rect 232240 689990 232310 690060
rect 232340 689990 232410 690060
rect 232440 689990 232510 690060
rect 227640 689890 227710 689960
rect 227740 689890 227810 689960
rect 227840 689890 227910 689960
rect 227940 689890 228010 689960
rect 228040 689890 228110 689960
rect 228140 689890 228210 689960
rect 228240 689890 228310 689960
rect 228340 689890 228410 689960
rect 228440 689890 228510 689960
rect 228540 689890 228610 689960
rect 228640 689890 228710 689960
rect 228740 689890 228810 689960
rect 228840 689890 228910 689960
rect 228940 689890 229010 689960
rect 229040 689890 229110 689960
rect 229140 689890 229210 689960
rect 229240 689890 229310 689960
rect 229340 689890 229410 689960
rect 229440 689890 229510 689960
rect 229540 689890 229610 689960
rect 229640 689890 229710 689960
rect 229740 689890 229810 689960
rect 229840 689890 229910 689960
rect 229940 689890 230010 689960
rect 230040 689890 230110 689960
rect 230140 689890 230210 689960
rect 230240 689890 230310 689960
rect 230340 689890 230410 689960
rect 230440 689890 230510 689960
rect 230540 689890 230610 689960
rect 230640 689890 230710 689960
rect 230740 689890 230810 689960
rect 230840 689890 230910 689960
rect 230940 689890 231010 689960
rect 231040 689890 231110 689960
rect 231140 689890 231210 689960
rect 231240 689890 231310 689960
rect 231340 689890 231410 689960
rect 231440 689890 231510 689960
rect 231540 689890 231610 689960
rect 231640 689890 231710 689960
rect 231740 689890 231810 689960
rect 231840 689890 231910 689960
rect 231940 689890 232010 689960
rect 232040 689890 232110 689960
rect 232140 689890 232210 689960
rect 232240 689890 232310 689960
rect 232340 689890 232410 689960
rect 232440 689890 232510 689960
<< metal3 >>
rect 16194 703650 21194 704800
rect 16194 703580 17270 703650
rect 17340 703580 17360 703650
rect 17430 703580 17450 703650
rect 17520 703580 17540 703650
rect 17610 703580 17630 703650
rect 17700 703580 17720 703650
rect 17790 703580 17810 703650
rect 17880 703580 17900 703650
rect 17970 703580 17990 703650
rect 18060 703580 18080 703650
rect 18150 703580 18170 703650
rect 18240 703580 18260 703650
rect 18330 703580 18350 703650
rect 18420 703580 18440 703650
rect 18510 703580 18530 703650
rect 18600 703580 18620 703650
rect 18690 703580 18710 703650
rect 18780 703580 18800 703650
rect 18870 703580 18890 703650
rect 18960 703580 18980 703650
rect 19050 703580 19070 703650
rect 19140 703580 19160 703650
rect 19230 703580 21194 703650
rect 16194 703560 21194 703580
rect 16194 703490 17270 703560
rect 17340 703490 17360 703560
rect 17430 703490 17450 703560
rect 17520 703490 17540 703560
rect 17610 703490 17630 703560
rect 17700 703490 17720 703560
rect 17790 703490 17810 703560
rect 17880 703490 17900 703560
rect 17970 703490 17990 703560
rect 18060 703490 18080 703560
rect 18150 703490 18170 703560
rect 18240 703490 18260 703560
rect 18330 703490 18350 703560
rect 18420 703490 18440 703560
rect 18510 703490 18530 703560
rect 18600 703490 18620 703560
rect 18690 703490 18710 703560
rect 18780 703490 18800 703560
rect 18870 703490 18890 703560
rect 18960 703490 18980 703560
rect 19050 703490 19070 703560
rect 19140 703490 19160 703560
rect 19230 703490 21194 703560
rect 16194 703470 21194 703490
rect 16194 703400 17270 703470
rect 17340 703400 17360 703470
rect 17430 703400 17450 703470
rect 17520 703400 17540 703470
rect 17610 703400 17630 703470
rect 17700 703400 17720 703470
rect 17790 703400 17810 703470
rect 17880 703400 17900 703470
rect 17970 703400 17990 703470
rect 18060 703400 18080 703470
rect 18150 703400 18170 703470
rect 18240 703400 18260 703470
rect 18330 703400 18350 703470
rect 18420 703400 18440 703470
rect 18510 703400 18530 703470
rect 18600 703400 18620 703470
rect 18690 703400 18710 703470
rect 18780 703400 18800 703470
rect 18870 703400 18890 703470
rect 18960 703400 18980 703470
rect 19050 703400 19070 703470
rect 19140 703400 19160 703470
rect 19230 703400 21194 703470
rect 16194 703380 21194 703400
rect 16194 703310 17270 703380
rect 17340 703310 17360 703380
rect 17430 703310 17450 703380
rect 17520 703310 17540 703380
rect 17610 703310 17630 703380
rect 17700 703310 17720 703380
rect 17790 703310 17810 703380
rect 17880 703310 17900 703380
rect 17970 703310 17990 703380
rect 18060 703310 18080 703380
rect 18150 703310 18170 703380
rect 18240 703310 18260 703380
rect 18330 703310 18350 703380
rect 18420 703310 18440 703380
rect 18510 703310 18530 703380
rect 18600 703310 18620 703380
rect 18690 703310 18710 703380
rect 18780 703310 18800 703380
rect 18870 703310 18890 703380
rect 18960 703310 18980 703380
rect 19050 703310 19070 703380
rect 19140 703310 19160 703380
rect 19230 703310 21194 703380
rect 16194 703290 21194 703310
rect 16194 703220 17270 703290
rect 17340 703220 17360 703290
rect 17430 703220 17450 703290
rect 17520 703220 17540 703290
rect 17610 703220 17630 703290
rect 17700 703220 17720 703290
rect 17790 703220 17810 703290
rect 17880 703220 17900 703290
rect 17970 703220 17990 703290
rect 18060 703220 18080 703290
rect 18150 703220 18170 703290
rect 18240 703220 18260 703290
rect 18330 703220 18350 703290
rect 18420 703220 18440 703290
rect 18510 703220 18530 703290
rect 18600 703220 18620 703290
rect 18690 703220 18710 703290
rect 18780 703220 18800 703290
rect 18870 703220 18890 703290
rect 18960 703220 18980 703290
rect 19050 703220 19070 703290
rect 19140 703220 19160 703290
rect 19230 703220 21194 703290
rect 16194 703200 21194 703220
rect 16194 703130 17270 703200
rect 17340 703130 17360 703200
rect 17430 703130 17450 703200
rect 17520 703130 17540 703200
rect 17610 703130 17630 703200
rect 17700 703130 17720 703200
rect 17790 703130 17810 703200
rect 17880 703130 17900 703200
rect 17970 703130 17990 703200
rect 18060 703130 18080 703200
rect 18150 703130 18170 703200
rect 18240 703130 18260 703200
rect 18330 703130 18350 703200
rect 18420 703130 18440 703200
rect 18510 703130 18530 703200
rect 18600 703130 18620 703200
rect 18690 703130 18710 703200
rect 18780 703130 18800 703200
rect 18870 703130 18890 703200
rect 18960 703130 18980 703200
rect 19050 703130 19070 703200
rect 19140 703130 19160 703200
rect 19230 703130 21194 703200
rect 16194 703110 21194 703130
rect 16194 703040 17270 703110
rect 17340 703040 17360 703110
rect 17430 703040 17450 703110
rect 17520 703040 17540 703110
rect 17610 703040 17630 703110
rect 17700 703040 17720 703110
rect 17790 703040 17810 703110
rect 17880 703040 17900 703110
rect 17970 703040 17990 703110
rect 18060 703040 18080 703110
rect 18150 703040 18170 703110
rect 18240 703040 18260 703110
rect 18330 703040 18350 703110
rect 18420 703040 18440 703110
rect 18510 703040 18530 703110
rect 18600 703040 18620 703110
rect 18690 703040 18710 703110
rect 18780 703040 18800 703110
rect 18870 703040 18890 703110
rect 18960 703040 18980 703110
rect 19050 703040 19070 703110
rect 19140 703040 19160 703110
rect 19230 703040 21194 703110
rect 16194 703020 21194 703040
rect 16194 702950 17270 703020
rect 17340 702950 17360 703020
rect 17430 702950 17450 703020
rect 17520 702950 17540 703020
rect 17610 702950 17630 703020
rect 17700 702950 17720 703020
rect 17790 702950 17810 703020
rect 17880 702950 17900 703020
rect 17970 702950 17990 703020
rect 18060 702950 18080 703020
rect 18150 702950 18170 703020
rect 18240 702950 18260 703020
rect 18330 702950 18350 703020
rect 18420 702950 18440 703020
rect 18510 702950 18530 703020
rect 18600 702950 18620 703020
rect 18690 702950 18710 703020
rect 18780 702950 18800 703020
rect 18870 702950 18890 703020
rect 18960 702950 18980 703020
rect 19050 702950 19070 703020
rect 19140 702950 19160 703020
rect 19230 702950 21194 703020
rect 16194 702930 21194 702950
rect 16194 702860 17270 702930
rect 17340 702860 17360 702930
rect 17430 702860 17450 702930
rect 17520 702860 17540 702930
rect 17610 702860 17630 702930
rect 17700 702860 17720 702930
rect 17790 702860 17810 702930
rect 17880 702860 17900 702930
rect 17970 702860 17990 702930
rect 18060 702860 18080 702930
rect 18150 702860 18170 702930
rect 18240 702860 18260 702930
rect 18330 702860 18350 702930
rect 18420 702860 18440 702930
rect 18510 702860 18530 702930
rect 18600 702860 18620 702930
rect 18690 702860 18710 702930
rect 18780 702860 18800 702930
rect 18870 702860 18890 702930
rect 18960 702860 18980 702930
rect 19050 702860 19070 702930
rect 19140 702860 19160 702930
rect 19230 702860 21194 702930
rect 16194 702840 21194 702860
rect 16194 702770 17270 702840
rect 17340 702770 17360 702840
rect 17430 702770 17450 702840
rect 17520 702770 17540 702840
rect 17610 702770 17630 702840
rect 17700 702770 17720 702840
rect 17790 702770 17810 702840
rect 17880 702770 17900 702840
rect 17970 702770 17990 702840
rect 18060 702770 18080 702840
rect 18150 702770 18170 702840
rect 18240 702770 18260 702840
rect 18330 702770 18350 702840
rect 18420 702770 18440 702840
rect 18510 702770 18530 702840
rect 18600 702770 18620 702840
rect 18690 702770 18710 702840
rect 18780 702770 18800 702840
rect 18870 702770 18890 702840
rect 18960 702770 18980 702840
rect 19050 702770 19070 702840
rect 19140 702770 19160 702840
rect 19230 702770 21194 702840
rect 16194 702750 21194 702770
rect 16194 702680 17270 702750
rect 17340 702680 17360 702750
rect 17430 702680 17450 702750
rect 17520 702680 17540 702750
rect 17610 702680 17630 702750
rect 17700 702680 17720 702750
rect 17790 702680 17810 702750
rect 17880 702680 17900 702750
rect 17970 702680 17990 702750
rect 18060 702680 18080 702750
rect 18150 702680 18170 702750
rect 18240 702680 18260 702750
rect 18330 702680 18350 702750
rect 18420 702680 18440 702750
rect 18510 702680 18530 702750
rect 18600 702680 18620 702750
rect 18690 702680 18710 702750
rect 18780 702680 18800 702750
rect 18870 702680 18890 702750
rect 18960 702680 18980 702750
rect 19050 702680 19070 702750
rect 19140 702680 19160 702750
rect 19230 702680 21194 702750
rect 16194 702660 21194 702680
rect 16194 702590 17270 702660
rect 17340 702590 17360 702660
rect 17430 702590 17450 702660
rect 17520 702590 17540 702660
rect 17610 702590 17630 702660
rect 17700 702590 17720 702660
rect 17790 702590 17810 702660
rect 17880 702590 17900 702660
rect 17970 702590 17990 702660
rect 18060 702590 18080 702660
rect 18150 702590 18170 702660
rect 18240 702590 18260 702660
rect 18330 702590 18350 702660
rect 18420 702590 18440 702660
rect 18510 702590 18530 702660
rect 18600 702590 18620 702660
rect 18690 702590 18710 702660
rect 18780 702590 18800 702660
rect 18870 702590 18890 702660
rect 18960 702590 18980 702660
rect 19050 702590 19070 702660
rect 19140 702590 19160 702660
rect 19230 702590 21194 702660
rect 16194 702570 21194 702590
rect 16194 702500 17270 702570
rect 17340 702500 17360 702570
rect 17430 702500 17450 702570
rect 17520 702500 17540 702570
rect 17610 702500 17630 702570
rect 17700 702500 17720 702570
rect 17790 702500 17810 702570
rect 17880 702500 17900 702570
rect 17970 702500 17990 702570
rect 18060 702500 18080 702570
rect 18150 702500 18170 702570
rect 18240 702500 18260 702570
rect 18330 702500 18350 702570
rect 18420 702500 18440 702570
rect 18510 702500 18530 702570
rect 18600 702500 18620 702570
rect 18690 702500 18710 702570
rect 18780 702500 18800 702570
rect 18870 702500 18890 702570
rect 18960 702500 18980 702570
rect 19050 702500 19070 702570
rect 19140 702500 19160 702570
rect 19230 702500 21194 702570
rect 16194 702480 21194 702500
rect 16194 702410 17270 702480
rect 17340 702410 17360 702480
rect 17430 702410 17450 702480
rect 17520 702410 17540 702480
rect 17610 702410 17630 702480
rect 17700 702410 17720 702480
rect 17790 702410 17810 702480
rect 17880 702410 17900 702480
rect 17970 702410 17990 702480
rect 18060 702410 18080 702480
rect 18150 702410 18170 702480
rect 18240 702410 18260 702480
rect 18330 702410 18350 702480
rect 18420 702410 18440 702480
rect 18510 702410 18530 702480
rect 18600 702410 18620 702480
rect 18690 702410 18710 702480
rect 18780 702410 18800 702480
rect 18870 702410 18890 702480
rect 18960 702410 18980 702480
rect 19050 702410 19070 702480
rect 19140 702410 19160 702480
rect 19230 702410 21194 702480
rect 16194 702390 21194 702410
rect 16194 702320 17270 702390
rect 17340 702320 17360 702390
rect 17430 702320 17450 702390
rect 17520 702320 17540 702390
rect 17610 702320 17630 702390
rect 17700 702320 17720 702390
rect 17790 702320 17810 702390
rect 17880 702320 17900 702390
rect 17970 702320 17990 702390
rect 18060 702320 18080 702390
rect 18150 702320 18170 702390
rect 18240 702320 18260 702390
rect 18330 702320 18350 702390
rect 18420 702320 18440 702390
rect 18510 702320 18530 702390
rect 18600 702320 18620 702390
rect 18690 702320 18710 702390
rect 18780 702320 18800 702390
rect 18870 702320 18890 702390
rect 18960 702320 18980 702390
rect 19050 702320 19070 702390
rect 19140 702320 19160 702390
rect 19230 702320 21194 702390
rect 16194 702300 21194 702320
rect 68194 703800 73194 704800
rect 68194 703500 68352 703800
rect 68652 703500 68852 703800
rect 69152 703500 69352 703800
rect 69652 703500 69852 703800
rect 70152 703500 70352 703800
rect 70652 703500 70852 703800
rect 71152 703500 71352 703800
rect 71652 703500 71852 703800
rect 72152 703500 72352 703800
rect 72652 703500 72852 703800
rect 73152 703500 73194 703800
rect 68194 703300 73194 703500
rect 68194 703000 68352 703300
rect 68652 703000 68852 703300
rect 69152 703000 69352 703300
rect 69652 703000 69852 703300
rect 70152 703000 70352 703300
rect 70652 703000 70852 703300
rect 71152 703000 71352 703300
rect 71652 703000 71852 703300
rect 72152 703000 72352 703300
rect 72652 703000 72852 703300
rect 73152 703000 73194 703300
rect 68194 702800 73194 703000
rect 68194 702500 68352 702800
rect 68652 702500 68852 702800
rect 69152 702500 69352 702800
rect 69652 702500 69852 702800
rect 70152 702500 70352 702800
rect 70652 702500 70852 702800
rect 71152 702500 71352 702800
rect 71652 702500 71852 702800
rect 72152 702500 72352 702800
rect 72652 702500 72852 702800
rect 73152 702500 73194 702800
rect 68194 702300 73194 702500
rect 120194 703800 125194 704800
rect 120194 703500 120352 703800
rect 120652 703500 120852 703800
rect 121152 703500 121352 703800
rect 121652 703500 121852 703800
rect 122152 703500 122352 703800
rect 122652 703500 122852 703800
rect 123152 703500 123352 703800
rect 123652 703500 123852 703800
rect 124152 703500 124352 703800
rect 124652 703500 124852 703800
rect 125152 703500 125194 703800
rect 120194 703300 125194 703500
rect 120194 703000 120352 703300
rect 120652 703000 120852 703300
rect 121152 703000 121352 703300
rect 121652 703000 121852 703300
rect 122152 703000 122352 703300
rect 122652 703000 122852 703300
rect 123152 703000 123352 703300
rect 123652 703000 123852 703300
rect 124152 703000 124352 703300
rect 124652 703000 124852 703300
rect 125152 703000 125194 703300
rect 120194 702800 125194 703000
rect 120194 702500 120352 702800
rect 120652 702500 120852 702800
rect 121152 702500 121352 702800
rect 121652 702500 121852 702800
rect 122152 702500 122352 702800
rect 122652 702500 122852 702800
rect 123152 702500 123352 702800
rect 123652 702500 123852 702800
rect 124152 702500 124352 702800
rect 124652 702500 124852 702800
rect 125152 702500 125194 702800
rect 120194 702300 125194 702500
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703110 418394 704800
rect 413394 703040 415760 703110
rect 415830 703040 415850 703110
rect 415920 703040 415940 703110
rect 416010 703040 416030 703110
rect 416100 703040 416120 703110
rect 416190 703040 418394 703110
rect 413394 703020 418394 703040
rect 413394 702950 415760 703020
rect 415830 702950 415850 703020
rect 415920 702950 415940 703020
rect 416010 702950 416030 703020
rect 416100 702950 416120 703020
rect 416190 702950 418394 703020
rect 413394 702930 418394 702950
rect 413394 702860 415760 702930
rect 415830 702860 415850 702930
rect 415920 702860 415940 702930
rect 416010 702860 416030 702930
rect 416100 702860 416120 702930
rect 416190 702860 418394 702930
rect 413394 702840 418394 702860
rect 413394 702770 415760 702840
rect 415830 702770 415850 702840
rect 415920 702770 415940 702840
rect 416010 702770 416030 702840
rect 416100 702770 416120 702840
rect 416190 702770 418394 702840
rect 413394 702750 418394 702770
rect 413394 702680 415760 702750
rect 415830 702680 415850 702750
rect 415920 702680 415940 702750
rect 416010 702680 416030 702750
rect 416100 702680 416120 702750
rect 416190 702680 418394 702750
rect 413394 702300 418394 702680
rect 465394 703110 470394 704800
rect 465394 703040 467010 703110
rect 467080 703040 467100 703110
rect 467170 703040 467190 703110
rect 467260 703040 467280 703110
rect 467350 703040 467370 703110
rect 467440 703040 470394 703110
rect 465394 703020 470394 703040
rect 465394 702950 467010 703020
rect 467080 702950 467100 703020
rect 467170 702950 467190 703020
rect 467260 702950 467280 703020
rect 467350 702950 467370 703020
rect 467440 702950 470394 703020
rect 465394 702930 470394 702950
rect 465394 702860 467010 702930
rect 467080 702860 467100 702930
rect 467170 702860 467190 702930
rect 467260 702860 467280 702930
rect 467350 702860 467370 702930
rect 467440 702860 470394 702930
rect 465394 702840 470394 702860
rect 465394 702770 467010 702840
rect 467080 702770 467100 702840
rect 467170 702770 467190 702840
rect 467260 702770 467280 702840
rect 467350 702770 467370 702840
rect 467440 702770 470394 702840
rect 465394 702750 470394 702770
rect 465394 702680 467010 702750
rect 467080 702680 467100 702750
rect 467170 702680 467190 702750
rect 467260 702680 467280 702750
rect 467350 702680 467370 702750
rect 467440 702680 470394 702750
rect 465394 702300 470394 702680
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 703110 571594 704800
rect 566594 703040 569140 703110
rect 569210 703040 569230 703110
rect 569300 703040 569320 703110
rect 569390 703040 569410 703110
rect 569480 703040 569500 703110
rect 569570 703040 571594 703110
rect 566594 703020 571594 703040
rect 566594 702950 569140 703020
rect 569210 702950 569230 703020
rect 569300 702950 569320 703020
rect 569390 702950 569410 703020
rect 569480 702950 569500 703020
rect 569570 702950 571594 703020
rect 566594 702930 571594 702950
rect 566594 702860 569140 702930
rect 569210 702860 569230 702930
rect 569300 702860 569320 702930
rect 569390 702860 569410 702930
rect 569480 702860 569500 702930
rect 569570 702860 571594 702930
rect 566594 702840 571594 702860
rect 566594 702770 569140 702840
rect 569210 702770 569230 702840
rect 569300 702770 569320 702840
rect 569390 702770 569410 702840
rect 569480 702770 569500 702840
rect 569570 702770 571594 702840
rect 566594 702750 571594 702770
rect 566594 702680 569140 702750
rect 569210 702680 569230 702750
rect 569300 702680 569320 702750
rect 569390 702680 569410 702750
rect 569480 702680 569500 702750
rect 569570 702680 571594 702750
rect 566594 702300 571594 702680
rect 224718 697420 235086 697448
rect 224718 697350 224744 697420
rect 224814 697350 224834 697420
rect 224904 697350 224924 697420
rect 224994 697350 225014 697420
rect 225084 697350 225104 697420
rect 225174 697350 234630 697420
rect 234700 697350 234720 697420
rect 234790 697350 234810 697420
rect 234880 697350 234900 697420
rect 234970 697350 234990 697420
rect 235060 697350 235086 697420
rect 224718 697330 235086 697350
rect 224718 697260 224744 697330
rect 224814 697260 224834 697330
rect 224904 697260 224924 697330
rect 224994 697260 225014 697330
rect 225084 697260 225104 697330
rect 225174 697260 234630 697330
rect 234700 697260 234720 697330
rect 234790 697260 234810 697330
rect 234880 697260 234900 697330
rect 234970 697260 234990 697330
rect 235060 697260 235086 697330
rect 224718 697240 235086 697260
rect 224718 697170 224744 697240
rect 224814 697170 224834 697240
rect 224904 697170 224924 697240
rect 224994 697170 225014 697240
rect 225084 697170 225104 697240
rect 225174 697170 234630 697240
rect 234700 697170 234720 697240
rect 234790 697170 234810 697240
rect 234880 697170 234900 697240
rect 234970 697170 234990 697240
rect 235060 697170 235086 697240
rect 224718 697150 235086 697170
rect 224718 697080 224744 697150
rect 224814 697080 224834 697150
rect 224904 697080 224924 697150
rect 224994 697080 225014 697150
rect 225084 697080 225104 697150
rect 225174 697080 234630 697150
rect 234700 697080 234720 697150
rect 234790 697080 234810 697150
rect 234880 697080 234900 697150
rect 234970 697080 234990 697150
rect 235060 697080 235086 697150
rect 224718 697060 235086 697080
rect 224718 696990 224744 697060
rect 224814 696990 224834 697060
rect 224904 696990 224924 697060
rect 224994 696990 225014 697060
rect 225084 696990 225104 697060
rect 225174 696990 234630 697060
rect 234700 696990 234720 697060
rect 234790 696990 234810 697060
rect 234880 696990 234900 697060
rect 234970 696990 234990 697060
rect 235060 696990 235086 697060
rect 224718 696968 235086 696990
rect 224718 696203 235086 696231
rect 224718 696133 224744 696203
rect 224814 696133 224834 696203
rect 224904 696133 224924 696203
rect 224994 696133 225014 696203
rect 225084 696133 225104 696203
rect 225174 696133 234630 696203
rect 234700 696133 234720 696203
rect 234790 696133 234810 696203
rect 234880 696133 234900 696203
rect 234970 696133 234990 696203
rect 235060 696133 235086 696203
rect 224718 696113 235086 696133
rect 224718 696043 224744 696113
rect 224814 696043 224834 696113
rect 224904 696043 224924 696113
rect 224994 696043 225014 696113
rect 225084 696043 225104 696113
rect 225174 696043 234630 696113
rect 234700 696043 234720 696113
rect 234790 696043 234810 696113
rect 234880 696043 234900 696113
rect 234970 696043 234990 696113
rect 235060 696043 235086 696113
rect 224718 696023 235086 696043
rect 224718 695953 224744 696023
rect 224814 695953 224834 696023
rect 224904 695953 224924 696023
rect 224994 695953 225014 696023
rect 225084 695953 225104 696023
rect 225174 695953 234630 696023
rect 234700 695953 234720 696023
rect 234790 695953 234810 696023
rect 234880 695953 234900 696023
rect 234970 695953 234990 696023
rect 235060 695953 235086 696023
rect 224718 695933 235086 695953
rect 224718 695863 224744 695933
rect 224814 695863 224834 695933
rect 224904 695863 224924 695933
rect 224994 695863 225014 695933
rect 225084 695863 225104 695933
rect 225174 695863 234630 695933
rect 234700 695863 234720 695933
rect 234790 695863 234810 695933
rect 234880 695863 234900 695933
rect 234970 695863 234990 695933
rect 235060 695863 235086 695933
rect 224718 695843 235086 695863
rect 224718 695773 224744 695843
rect 224814 695773 224834 695843
rect 224904 695773 224924 695843
rect 224994 695773 225014 695843
rect 225084 695773 225104 695843
rect 225174 695773 234630 695843
rect 234700 695773 234720 695843
rect 234790 695773 234810 695843
rect 234880 695773 234900 695843
rect 234970 695773 234990 695843
rect 235060 695773 235086 695843
rect 224718 695751 235086 695773
rect 224718 695138 235086 695166
rect 224718 695068 224744 695138
rect 224814 695068 224834 695138
rect 224904 695068 224924 695138
rect 224994 695068 225014 695138
rect 225084 695068 225104 695138
rect 225174 695068 234630 695138
rect 234700 695068 234720 695138
rect 234790 695068 234810 695138
rect 234880 695068 234900 695138
rect 234970 695068 234990 695138
rect 235060 695068 235086 695138
rect 224718 695048 235086 695068
rect 224718 694978 224744 695048
rect 224814 694978 224834 695048
rect 224904 694978 224924 695048
rect 224994 694978 225014 695048
rect 225084 694978 225104 695048
rect 225174 694978 234630 695048
rect 234700 694978 234720 695048
rect 234790 694978 234810 695048
rect 234880 694978 234900 695048
rect 234970 694978 234990 695048
rect 235060 694978 235086 695048
rect 224718 694958 235086 694978
rect 224718 694888 224744 694958
rect 224814 694888 224834 694958
rect 224904 694888 224924 694958
rect 224994 694888 225014 694958
rect 225084 694888 225104 694958
rect 225174 694888 234630 694958
rect 234700 694888 234720 694958
rect 234790 694888 234810 694958
rect 234880 694888 234900 694958
rect 234970 694888 234990 694958
rect 235060 694888 235086 694958
rect 224718 694868 235086 694888
rect 224718 694798 224744 694868
rect 224814 694798 224834 694868
rect 224904 694798 224924 694868
rect 224994 694798 225014 694868
rect 225084 694798 225104 694868
rect 225174 694798 234630 694868
rect 234700 694798 234720 694868
rect 234790 694798 234810 694868
rect 234880 694798 234900 694868
rect 234970 694798 234990 694868
rect 235060 694798 235086 694868
rect 224718 694778 235086 694798
rect 224718 694708 224744 694778
rect 224814 694708 224834 694778
rect 224904 694708 224924 694778
rect 224994 694708 225014 694778
rect 225084 694708 225104 694778
rect 225174 694708 234630 694778
rect 234700 694708 234720 694778
rect 234790 694708 234810 694778
rect 234880 694708 234900 694778
rect 234970 694708 234990 694778
rect 235060 694708 235086 694778
rect 224718 694686 235086 694708
rect 224718 693432 235086 693460
rect 224718 693362 224744 693432
rect 224814 693362 224834 693432
rect 224904 693362 224924 693432
rect 224994 693362 225014 693432
rect 225084 693362 225104 693432
rect 225174 693362 234630 693432
rect 234700 693362 234720 693432
rect 234790 693362 234810 693432
rect 234880 693362 234900 693432
rect 234970 693362 234990 693432
rect 235060 693362 235086 693432
rect 224718 693342 235086 693362
rect 224718 693272 224744 693342
rect 224814 693272 224834 693342
rect 224904 693272 224924 693342
rect 224994 693272 225014 693342
rect 225084 693272 225104 693342
rect 225174 693272 234630 693342
rect 234700 693272 234720 693342
rect 234790 693272 234810 693342
rect 234880 693272 234900 693342
rect 234970 693272 234990 693342
rect 235060 693272 235086 693342
rect 224718 693252 235086 693272
rect 224718 693182 224744 693252
rect 224814 693182 224834 693252
rect 224904 693182 224924 693252
rect 224994 693182 225014 693252
rect 225084 693182 225104 693252
rect 225174 693182 234630 693252
rect 234700 693182 234720 693252
rect 234790 693182 234810 693252
rect 234880 693182 234900 693252
rect 234970 693182 234990 693252
rect 235060 693182 235086 693252
rect 224718 693162 235086 693182
rect 224718 693092 224744 693162
rect 224814 693092 224834 693162
rect 224904 693092 224924 693162
rect 224994 693092 225014 693162
rect 225084 693092 225104 693162
rect 225174 693092 234630 693162
rect 234700 693092 234720 693162
rect 234790 693092 234810 693162
rect 234880 693092 234900 693162
rect 234970 693092 234990 693162
rect 235060 693092 235086 693162
rect 224718 693072 235086 693092
rect 224718 693002 224744 693072
rect 224814 693002 224834 693072
rect 224904 693002 224924 693072
rect 224994 693002 225014 693072
rect 225084 693002 225104 693072
rect 225174 693002 234630 693072
rect 234700 693002 234720 693072
rect 234790 693002 234810 693072
rect 234880 693002 234900 693072
rect 234970 693002 234990 693072
rect 235060 693002 235086 693072
rect 224718 692980 235086 693002
rect 224718 691718 235086 691746
rect 224718 691648 224744 691718
rect 224814 691648 224834 691718
rect 224904 691648 224924 691718
rect 224994 691648 225014 691718
rect 225084 691648 225104 691718
rect 225174 691648 234630 691718
rect 234700 691648 234720 691718
rect 234790 691648 234810 691718
rect 234880 691648 234900 691718
rect 234970 691648 234990 691718
rect 235060 691648 235086 691718
rect 165334 691580 170828 691635
rect 165334 691510 165360 691580
rect 165430 691510 165460 691580
rect 165530 691510 165560 691580
rect 165630 691510 165660 691580
rect 165730 691510 165760 691580
rect 165830 691510 165860 691580
rect 165930 691510 165960 691580
rect 166030 691510 166060 691580
rect 166130 691510 166160 691580
rect 166230 691510 166260 691580
rect 166330 691510 166360 691580
rect 166430 691510 166460 691580
rect 166530 691510 166560 691580
rect 166630 691510 166660 691580
rect 166730 691510 166760 691580
rect 166830 691510 166860 691580
rect 166930 691510 166960 691580
rect 167030 691510 167060 691580
rect 167130 691510 167160 691580
rect 167230 691510 167260 691580
rect 167330 691510 167360 691580
rect 167430 691510 167460 691580
rect 167530 691510 167560 691580
rect 167630 691510 167660 691580
rect 167730 691510 167760 691580
rect 167830 691510 167860 691580
rect 167930 691510 167960 691580
rect 168030 691510 168060 691580
rect 168130 691510 168160 691580
rect 168230 691510 168260 691580
rect 168330 691510 168360 691580
rect 168430 691510 168460 691580
rect 168530 691510 168560 691580
rect 168630 691510 168660 691580
rect 168730 691510 168760 691580
rect 168830 691510 168860 691580
rect 168930 691510 168960 691580
rect 169030 691510 169060 691580
rect 169130 691510 169160 691580
rect 169230 691510 169260 691580
rect 169330 691510 169360 691580
rect 169430 691510 169460 691580
rect 169530 691510 169560 691580
rect 169630 691510 169660 691580
rect 169730 691510 169760 691580
rect 169830 691510 169860 691580
rect 169930 691510 169960 691580
rect 170030 691510 170060 691580
rect 170130 691510 170160 691580
rect 170230 691510 170260 691580
rect 170330 691510 170360 691580
rect 170430 691510 170460 691580
rect 170530 691510 170828 691580
rect 165334 691470 170828 691510
rect 165334 691400 165360 691470
rect 165430 691400 165460 691470
rect 165530 691400 165560 691470
rect 165630 691400 165660 691470
rect 165730 691400 165760 691470
rect 165830 691400 165860 691470
rect 165930 691400 165960 691470
rect 166030 691400 166060 691470
rect 166130 691400 166160 691470
rect 166230 691400 166260 691470
rect 166330 691400 166360 691470
rect 166430 691400 166460 691470
rect 166530 691400 166560 691470
rect 166630 691400 166660 691470
rect 166730 691400 166760 691470
rect 166830 691400 166860 691470
rect 166930 691400 166960 691470
rect 167030 691400 167060 691470
rect 167130 691400 167160 691470
rect 167230 691400 167260 691470
rect 167330 691400 167360 691470
rect 167430 691400 167460 691470
rect 167530 691400 167560 691470
rect 167630 691400 167660 691470
rect 167730 691400 167760 691470
rect 167830 691400 167860 691470
rect 167930 691400 167960 691470
rect 168030 691400 168060 691470
rect 168130 691400 168160 691470
rect 168230 691400 168260 691470
rect 168330 691400 168360 691470
rect 168430 691400 168460 691470
rect 168530 691400 168560 691470
rect 168630 691400 168660 691470
rect 168730 691400 168760 691470
rect 168830 691400 168860 691470
rect 168930 691400 168960 691470
rect 169030 691400 169060 691470
rect 169130 691400 169160 691470
rect 169230 691400 169260 691470
rect 169330 691400 169360 691470
rect 169430 691400 169460 691470
rect 169530 691400 169560 691470
rect 169630 691400 169660 691470
rect 169730 691400 169760 691470
rect 169830 691400 169860 691470
rect 169930 691400 169960 691470
rect 170030 691400 170060 691470
rect 170130 691400 170160 691470
rect 170230 691400 170260 691470
rect 170330 691400 170360 691470
rect 170430 691400 170460 691470
rect 170530 691400 170828 691470
rect 165334 691360 170828 691400
rect 224718 691628 235086 691648
rect 224718 691558 224744 691628
rect 224814 691558 224834 691628
rect 224904 691558 224924 691628
rect 224994 691558 225014 691628
rect 225084 691558 225104 691628
rect 225174 691600 234630 691628
rect 225174 691558 227370 691600
rect 224718 691540 227370 691558
rect 227430 691540 227460 691600
rect 227520 691540 227550 691600
rect 227610 691540 227640 691600
rect 227700 691540 227730 691600
rect 227790 691540 227820 691600
rect 227880 691540 227910 691600
rect 227970 691540 228000 691600
rect 228060 691540 228090 691600
rect 228150 691540 228180 691600
rect 228240 691540 228270 691600
rect 228330 691540 228360 691600
rect 228420 691540 228450 691600
rect 228510 691540 228540 691600
rect 228600 691540 228630 691600
rect 228690 691540 228720 691600
rect 228780 691540 228810 691600
rect 228870 691540 228900 691600
rect 228960 691540 228990 691600
rect 229050 691540 229080 691600
rect 229140 691540 229170 691600
rect 229230 691540 229260 691600
rect 229320 691540 229350 691600
rect 229410 691540 229440 691600
rect 229500 691540 229530 691600
rect 229590 691540 229620 691600
rect 229680 691540 229710 691600
rect 229770 691540 229800 691600
rect 229860 691540 229890 691600
rect 229950 691540 229980 691600
rect 230040 691540 230070 691600
rect 230130 691540 230160 691600
rect 230220 691540 230250 691600
rect 230310 691540 230340 691600
rect 230400 691540 230430 691600
rect 230490 691540 230520 691600
rect 230580 691540 230610 691600
rect 230670 691540 230700 691600
rect 230760 691540 230790 691600
rect 230850 691540 230880 691600
rect 230940 691540 230970 691600
rect 231030 691540 231060 691600
rect 231120 691540 231150 691600
rect 231210 691540 231240 691600
rect 231300 691540 231330 691600
rect 231390 691540 231420 691600
rect 231480 691540 231510 691600
rect 231570 691540 231600 691600
rect 231660 691540 231690 691600
rect 231750 691540 231780 691600
rect 231840 691540 231870 691600
rect 231930 691540 231960 691600
rect 232020 691540 232050 691600
rect 232110 691540 232140 691600
rect 232200 691540 232230 691600
rect 232290 691540 232320 691600
rect 232380 691540 232410 691600
rect 232470 691540 232500 691600
rect 232560 691540 232590 691600
rect 232650 691540 232680 691600
rect 232740 691540 232770 691600
rect 232830 691558 234630 691600
rect 234700 691558 234720 691628
rect 234790 691558 234810 691628
rect 234880 691558 234900 691628
rect 234970 691558 234990 691628
rect 235060 691558 235086 691628
rect 232830 691540 235086 691558
rect 224718 691538 235086 691540
rect 224718 691468 224744 691538
rect 224814 691468 224834 691538
rect 224904 691468 224924 691538
rect 224994 691468 225014 691538
rect 225084 691468 225104 691538
rect 225174 691510 234630 691538
rect 225174 691468 227370 691510
rect 224718 691450 227370 691468
rect 227430 691450 227460 691510
rect 227520 691450 227550 691510
rect 227610 691450 227640 691510
rect 227700 691450 227730 691510
rect 227790 691450 227820 691510
rect 227880 691450 227910 691510
rect 227970 691450 228000 691510
rect 228060 691450 228090 691510
rect 228150 691450 228180 691510
rect 228240 691450 228270 691510
rect 228330 691450 228360 691510
rect 228420 691450 228450 691510
rect 228510 691450 228540 691510
rect 228600 691450 228630 691510
rect 228690 691450 228720 691510
rect 228780 691450 228810 691510
rect 228870 691450 228900 691510
rect 228960 691450 228990 691510
rect 229050 691450 229080 691510
rect 229140 691450 229170 691510
rect 229230 691450 229260 691510
rect 229320 691450 229350 691510
rect 229410 691450 229440 691510
rect 229500 691450 229530 691510
rect 229590 691450 229620 691510
rect 229680 691450 229710 691510
rect 229770 691450 229800 691510
rect 229860 691450 229890 691510
rect 229950 691450 229980 691510
rect 230040 691450 230070 691510
rect 230130 691450 230160 691510
rect 230220 691450 230250 691510
rect 230310 691450 230340 691510
rect 230400 691450 230430 691510
rect 230490 691450 230520 691510
rect 230580 691450 230610 691510
rect 230670 691450 230700 691510
rect 230760 691450 230790 691510
rect 230850 691450 230880 691510
rect 230940 691450 230970 691510
rect 231030 691450 231060 691510
rect 231120 691450 231150 691510
rect 231210 691450 231240 691510
rect 231300 691450 231330 691510
rect 231390 691450 231420 691510
rect 231480 691450 231510 691510
rect 231570 691450 231600 691510
rect 231660 691450 231690 691510
rect 231750 691450 231780 691510
rect 231840 691450 231870 691510
rect 231930 691450 231960 691510
rect 232020 691450 232050 691510
rect 232110 691450 232140 691510
rect 232200 691450 232230 691510
rect 232290 691450 232320 691510
rect 232380 691450 232410 691510
rect 232470 691450 232500 691510
rect 232560 691450 232590 691510
rect 232650 691450 232680 691510
rect 232740 691450 232770 691510
rect 232830 691468 234630 691510
rect 234700 691468 234720 691538
rect 234790 691468 234810 691538
rect 234880 691468 234900 691538
rect 234970 691468 234990 691538
rect 235060 691468 235086 691538
rect 232830 691450 235086 691468
rect 224718 691448 235086 691450
rect 224718 691378 224744 691448
rect 224814 691378 224834 691448
rect 224904 691378 224924 691448
rect 224994 691378 225014 691448
rect 225084 691378 225104 691448
rect 225174 691420 234630 691448
rect 225174 691378 227370 691420
rect 224718 691360 227370 691378
rect 227430 691360 227460 691420
rect 227520 691360 227550 691420
rect 227610 691360 227640 691420
rect 227700 691360 227730 691420
rect 227790 691360 227820 691420
rect 227880 691360 227910 691420
rect 227970 691360 228000 691420
rect 228060 691360 228090 691420
rect 228150 691360 228180 691420
rect 228240 691360 228270 691420
rect 228330 691360 228360 691420
rect 228420 691360 228450 691420
rect 228510 691360 228540 691420
rect 228600 691360 228630 691420
rect 228690 691360 228720 691420
rect 228780 691360 228810 691420
rect 228870 691360 228900 691420
rect 228960 691360 228990 691420
rect 229050 691360 229080 691420
rect 229140 691360 229170 691420
rect 229230 691360 229260 691420
rect 229320 691360 229350 691420
rect 229410 691360 229440 691420
rect 229500 691360 229530 691420
rect 229590 691360 229620 691420
rect 229680 691360 229710 691420
rect 229770 691360 229800 691420
rect 229860 691360 229890 691420
rect 229950 691360 229980 691420
rect 230040 691360 230070 691420
rect 230130 691360 230160 691420
rect 230220 691360 230250 691420
rect 230310 691360 230340 691420
rect 230400 691360 230430 691420
rect 230490 691360 230520 691420
rect 230580 691360 230610 691420
rect 230670 691360 230700 691420
rect 230760 691360 230790 691420
rect 230850 691360 230880 691420
rect 230940 691360 230970 691420
rect 231030 691360 231060 691420
rect 231120 691360 231150 691420
rect 231210 691360 231240 691420
rect 231300 691360 231330 691420
rect 231390 691360 231420 691420
rect 231480 691360 231510 691420
rect 231570 691360 231600 691420
rect 231660 691360 231690 691420
rect 231750 691360 231780 691420
rect 231840 691360 231870 691420
rect 231930 691360 231960 691420
rect 232020 691360 232050 691420
rect 232110 691360 232140 691420
rect 232200 691360 232230 691420
rect 232290 691360 232320 691420
rect 232380 691360 232410 691420
rect 232470 691360 232500 691420
rect 232560 691360 232590 691420
rect 232650 691360 232680 691420
rect 232740 691360 232770 691420
rect 232830 691378 234630 691420
rect 234700 691378 234720 691448
rect 234790 691378 234810 691448
rect 234880 691378 234900 691448
rect 234970 691378 234990 691448
rect 235060 691378 235086 691448
rect 232830 691360 235086 691378
rect 224718 691358 235086 691360
rect 224718 691288 224744 691358
rect 224814 691288 224834 691358
rect 224904 691288 224924 691358
rect 224994 691288 225014 691358
rect 225084 691288 225104 691358
rect 225174 691288 234630 691358
rect 234700 691288 234720 691358
rect 234790 691288 234810 691358
rect 234880 691288 234900 691358
rect 234970 691288 234990 691358
rect 235060 691288 235086 691358
rect 224718 691266 235086 691288
rect 165364 690070 170798 690104
rect 165364 690000 165620 690070
rect 165690 690000 165720 690070
rect 165790 690000 165820 690070
rect 165890 690000 165920 690070
rect 165990 690000 166020 690070
rect 166090 690000 166120 690070
rect 166190 690000 166220 690070
rect 166290 690000 166320 690070
rect 166390 690000 166420 690070
rect 166490 690000 166520 690070
rect 166590 690000 166620 690070
rect 166690 690000 166720 690070
rect 166790 690000 166820 690070
rect 166890 690000 166920 690070
rect 166990 690000 167020 690070
rect 167090 690000 167120 690070
rect 167190 690000 167220 690070
rect 167290 690000 167320 690070
rect 167390 690000 167420 690070
rect 167490 690000 167520 690070
rect 167590 690000 167620 690070
rect 167690 690000 167720 690070
rect 167790 690000 167820 690070
rect 167890 690000 167920 690070
rect 167990 690000 168020 690070
rect 168090 690000 168120 690070
rect 168190 690000 168220 690070
rect 168290 690000 168320 690070
rect 168390 690000 168420 690070
rect 168490 690000 168520 690070
rect 168590 690000 168620 690070
rect 168690 690000 168720 690070
rect 168790 690000 168820 690070
rect 168890 690000 168920 690070
rect 168990 690000 169020 690070
rect 169090 690000 169120 690070
rect 169190 690000 169220 690070
rect 169290 690000 169320 690070
rect 169390 690000 169420 690070
rect 169490 690000 169520 690070
rect 169590 690000 169620 690070
rect 169690 690000 169720 690070
rect 169790 690000 169820 690070
rect 169890 690000 169920 690070
rect 169990 690000 170020 690070
rect 170090 690000 170120 690070
rect 170190 690000 170220 690070
rect 170290 690000 170320 690070
rect 170390 690000 170420 690070
rect 170490 690000 170798 690070
rect 165364 689970 170798 690000
rect 165364 689900 165620 689970
rect 165690 689900 165720 689970
rect 165790 689900 165820 689970
rect 165890 689900 165920 689970
rect 165990 689900 166020 689970
rect 166090 689900 166120 689970
rect 166190 689900 166220 689970
rect 166290 689900 166320 689970
rect 166390 689900 166420 689970
rect 166490 689900 166520 689970
rect 166590 689900 166620 689970
rect 166690 689900 166720 689970
rect 166790 689900 166820 689970
rect 166890 689900 166920 689970
rect 166990 689900 167020 689970
rect 167090 689900 167120 689970
rect 167190 689900 167220 689970
rect 167290 689900 167320 689970
rect 167390 689900 167420 689970
rect 167490 689900 167520 689970
rect 167590 689900 167620 689970
rect 167690 689900 167720 689970
rect 167790 689900 167820 689970
rect 167890 689900 167920 689970
rect 167990 689900 168020 689970
rect 168090 689900 168120 689970
rect 168190 689900 168220 689970
rect 168290 689900 168320 689970
rect 168390 689900 168420 689970
rect 168490 689900 168520 689970
rect 168590 689900 168620 689970
rect 168690 689900 168720 689970
rect 168790 689900 168820 689970
rect 168890 689900 168920 689970
rect 168990 689900 169020 689970
rect 169090 689900 169120 689970
rect 169190 689900 169220 689970
rect 169290 689900 169320 689970
rect 169390 689900 169420 689970
rect 169490 689900 169520 689970
rect 169590 689900 169620 689970
rect 169690 689900 169720 689970
rect 169790 689900 169820 689970
rect 169890 689900 169920 689970
rect 169990 689900 170020 689970
rect 170090 689900 170120 689970
rect 170190 689900 170220 689970
rect 170290 689900 170320 689970
rect 170390 689900 170420 689970
rect 170490 689900 170798 689970
rect 165364 689877 170798 689900
rect 227386 690060 232820 690114
rect 227386 689990 227640 690060
rect 227710 689990 227740 690060
rect 227810 689990 227840 690060
rect 227910 689990 227940 690060
rect 228010 689990 228040 690060
rect 228110 689990 228140 690060
rect 228210 689990 228240 690060
rect 228310 689990 228340 690060
rect 228410 689990 228440 690060
rect 228510 689990 228540 690060
rect 228610 689990 228640 690060
rect 228710 689990 228740 690060
rect 228810 689990 228840 690060
rect 228910 689990 228940 690060
rect 229010 689990 229040 690060
rect 229110 689990 229140 690060
rect 229210 689990 229240 690060
rect 229310 689990 229340 690060
rect 229410 689990 229440 690060
rect 229510 689990 229540 690060
rect 229610 689990 229640 690060
rect 229710 689990 229740 690060
rect 229810 689990 229840 690060
rect 229910 689990 229940 690060
rect 230010 689990 230040 690060
rect 230110 689990 230140 690060
rect 230210 689990 230240 690060
rect 230310 689990 230340 690060
rect 230410 689990 230440 690060
rect 230510 689990 230540 690060
rect 230610 689990 230640 690060
rect 230710 689990 230740 690060
rect 230810 689990 230840 690060
rect 230910 689990 230940 690060
rect 231010 689990 231040 690060
rect 231110 689990 231140 690060
rect 231210 689990 231240 690060
rect 231310 689990 231340 690060
rect 231410 689990 231440 690060
rect 231510 689990 231540 690060
rect 231610 689990 231640 690060
rect 231710 689990 231740 690060
rect 231810 689990 231840 690060
rect 231910 689990 231940 690060
rect 232010 689990 232040 690060
rect 232110 689990 232140 690060
rect 232210 689990 232240 690060
rect 232310 689990 232340 690060
rect 232410 689990 232440 690060
rect 232510 689990 232820 690060
rect 227386 689960 232820 689990
rect 227386 689890 227640 689960
rect 227710 689890 227740 689960
rect 227810 689890 227840 689960
rect 227910 689890 227940 689960
rect 228010 689890 228040 689960
rect 228110 689890 228140 689960
rect 228210 689890 228240 689960
rect 228310 689890 228340 689960
rect 228410 689890 228440 689960
rect 228510 689890 228540 689960
rect 228610 689890 228640 689960
rect 228710 689890 228740 689960
rect 228810 689890 228840 689960
rect 228910 689890 228940 689960
rect 229010 689890 229040 689960
rect 229110 689890 229140 689960
rect 229210 689890 229240 689960
rect 229310 689890 229340 689960
rect 229410 689890 229440 689960
rect 229510 689890 229540 689960
rect 229610 689890 229640 689960
rect 229710 689890 229740 689960
rect 229810 689890 229840 689960
rect 229910 689890 229940 689960
rect 230010 689890 230040 689960
rect 230110 689890 230140 689960
rect 230210 689890 230240 689960
rect 230310 689890 230340 689960
rect 230410 689890 230440 689960
rect 230510 689890 230540 689960
rect 230610 689890 230640 689960
rect 230710 689890 230740 689960
rect 230810 689890 230840 689960
rect 230910 689890 230940 689960
rect 231010 689890 231040 689960
rect 231110 689890 231140 689960
rect 231210 689890 231240 689960
rect 231310 689890 231340 689960
rect 231410 689890 231440 689960
rect 231510 689890 231540 689960
rect 231610 689890 231640 689960
rect 231710 689890 231740 689960
rect 231810 689890 231840 689960
rect 231910 689890 231940 689960
rect 232010 689890 232040 689960
rect 232110 689890 232140 689960
rect 232210 689890 232240 689960
rect 232310 689890 232340 689960
rect 232410 689890 232440 689960
rect 232510 689890 232820 689960
rect 227386 689853 232820 689890
rect -800 683630 1700 685242
rect -800 683560 350 683630
rect 420 683560 440 683630
rect 510 683560 530 683630
rect 600 683560 620 683630
rect 690 683560 710 683630
rect 780 683560 800 683630
rect 870 683560 890 683630
rect 960 683560 980 683630
rect 1050 683560 1070 683630
rect 1140 683560 1160 683630
rect 1230 683560 1250 683630
rect 1320 683560 1340 683630
rect 1410 683560 1430 683630
rect 1500 683560 1520 683630
rect 1590 683560 1610 683630
rect 1680 683560 1700 683630
rect -800 683540 1700 683560
rect -800 683470 350 683540
rect 420 683470 440 683540
rect 510 683470 530 683540
rect 600 683470 620 683540
rect 690 683470 710 683540
rect 780 683470 800 683540
rect 870 683470 890 683540
rect 960 683470 980 683540
rect 1050 683470 1070 683540
rect 1140 683470 1160 683540
rect 1230 683470 1250 683540
rect 1320 683470 1340 683540
rect 1410 683470 1430 683540
rect 1500 683470 1520 683540
rect 1590 683470 1610 683540
rect 1680 683470 1700 683540
rect -800 683450 1700 683470
rect -800 683380 350 683450
rect 420 683380 440 683450
rect 510 683380 530 683450
rect 600 683380 620 683450
rect 690 683380 710 683450
rect 780 683380 800 683450
rect 870 683380 890 683450
rect 960 683380 980 683450
rect 1050 683380 1070 683450
rect 1140 683380 1160 683450
rect 1230 683380 1250 683450
rect 1320 683380 1340 683450
rect 1410 683380 1430 683450
rect 1500 683380 1520 683450
rect 1590 683380 1610 683450
rect 1680 683380 1700 683450
rect -800 683360 1700 683380
rect -800 683290 350 683360
rect 420 683290 440 683360
rect 510 683290 530 683360
rect 600 683290 620 683360
rect 690 683290 710 683360
rect 780 683290 800 683360
rect 870 683290 890 683360
rect 960 683290 980 683360
rect 1050 683290 1070 683360
rect 1140 683290 1160 683360
rect 1230 683290 1250 683360
rect 1320 683290 1340 683360
rect 1410 683290 1430 683360
rect 1500 683290 1520 683360
rect 1590 683290 1610 683360
rect 1680 683290 1700 683360
rect -800 683270 1700 683290
rect -800 683200 350 683270
rect 420 683200 440 683270
rect 510 683200 530 683270
rect 600 683200 620 683270
rect 690 683200 710 683270
rect 780 683200 800 683270
rect 870 683200 890 683270
rect 960 683200 980 683270
rect 1050 683200 1070 683270
rect 1140 683200 1160 683270
rect 1230 683200 1250 683270
rect 1320 683200 1340 683270
rect 1410 683200 1430 683270
rect 1500 683200 1520 683270
rect 1590 683200 1610 683270
rect 1680 683200 1700 683270
rect -800 683180 1700 683200
rect -800 683110 350 683180
rect 420 683110 440 683180
rect 510 683110 530 683180
rect 600 683110 620 683180
rect 690 683110 710 683180
rect 780 683110 800 683180
rect 870 683110 890 683180
rect 960 683110 980 683180
rect 1050 683110 1070 683180
rect 1140 683110 1160 683180
rect 1230 683110 1250 683180
rect 1320 683110 1340 683180
rect 1410 683110 1430 683180
rect 1500 683110 1520 683180
rect 1590 683110 1610 683180
rect 1680 683110 1700 683180
rect -800 683090 1700 683110
rect -800 683020 350 683090
rect 420 683020 440 683090
rect 510 683020 530 683090
rect 600 683020 620 683090
rect 690 683020 710 683090
rect 780 683020 800 683090
rect 870 683020 890 683090
rect 960 683020 980 683090
rect 1050 683020 1070 683090
rect 1140 683020 1160 683090
rect 1230 683020 1250 683090
rect 1320 683020 1340 683090
rect 1410 683020 1430 683090
rect 1500 683020 1520 683090
rect 1590 683020 1610 683090
rect 1680 683020 1700 683090
rect -800 683000 1700 683020
rect -800 682930 350 683000
rect 420 682930 440 683000
rect 510 682930 530 683000
rect 600 682930 620 683000
rect 690 682930 710 683000
rect 780 682930 800 683000
rect 870 682930 890 683000
rect 960 682930 980 683000
rect 1050 682930 1070 683000
rect 1140 682930 1160 683000
rect 1230 682930 1250 683000
rect 1320 682930 1340 683000
rect 1410 682930 1430 683000
rect 1500 682930 1520 683000
rect 1590 682930 1610 683000
rect 1680 682930 1700 683000
rect -800 682910 1700 682930
rect -800 682840 350 682910
rect 420 682840 440 682910
rect 510 682840 530 682910
rect 600 682840 620 682910
rect 690 682840 710 682910
rect 780 682840 800 682910
rect 870 682840 890 682910
rect 960 682840 980 682910
rect 1050 682840 1070 682910
rect 1140 682840 1160 682910
rect 1230 682840 1250 682910
rect 1320 682840 1340 682910
rect 1410 682840 1430 682910
rect 1500 682840 1520 682910
rect 1590 682840 1610 682910
rect 1680 682840 1700 682910
rect -800 682820 1700 682840
rect -800 682750 350 682820
rect 420 682750 440 682820
rect 510 682750 530 682820
rect 600 682750 620 682820
rect 690 682750 710 682820
rect 780 682750 800 682820
rect 870 682750 890 682820
rect 960 682750 980 682820
rect 1050 682750 1070 682820
rect 1140 682750 1160 682820
rect 1230 682750 1250 682820
rect 1320 682750 1340 682820
rect 1410 682750 1430 682820
rect 1500 682750 1520 682820
rect 1590 682750 1610 682820
rect 1680 682750 1700 682820
rect -800 682730 1700 682750
rect -800 682660 350 682730
rect 420 682660 440 682730
rect 510 682660 530 682730
rect 600 682660 620 682730
rect 690 682660 710 682730
rect 780 682660 800 682730
rect 870 682660 890 682730
rect 960 682660 980 682730
rect 1050 682660 1070 682730
rect 1140 682660 1160 682730
rect 1230 682660 1250 682730
rect 1320 682660 1340 682730
rect 1410 682660 1430 682730
rect 1500 682660 1520 682730
rect 1590 682660 1610 682730
rect 1680 682660 1700 682730
rect -800 682640 1700 682660
rect -800 682570 350 682640
rect 420 682570 440 682640
rect 510 682570 530 682640
rect 600 682570 620 682640
rect 690 682570 710 682640
rect 780 682570 800 682640
rect 870 682570 890 682640
rect 960 682570 980 682640
rect 1050 682570 1070 682640
rect 1140 682570 1160 682640
rect 1230 682570 1250 682640
rect 1320 682570 1340 682640
rect 1410 682570 1430 682640
rect 1500 682570 1520 682640
rect 1590 682570 1610 682640
rect 1680 682570 1700 682640
rect -800 682550 1700 682570
rect -800 682480 350 682550
rect 420 682480 440 682550
rect 510 682480 530 682550
rect 600 682480 620 682550
rect 690 682480 710 682550
rect 780 682480 800 682550
rect 870 682480 890 682550
rect 960 682480 980 682550
rect 1050 682480 1070 682550
rect 1140 682480 1160 682550
rect 1230 682480 1250 682550
rect 1320 682480 1340 682550
rect 1410 682480 1430 682550
rect 1500 682480 1520 682550
rect 1590 682480 1610 682550
rect 1680 682480 1700 682550
rect -800 682460 1700 682480
rect -800 682390 350 682460
rect 420 682390 440 682460
rect 510 682390 530 682460
rect 600 682390 620 682460
rect 690 682390 710 682460
rect 780 682390 800 682460
rect 870 682390 890 682460
rect 960 682390 980 682460
rect 1050 682390 1070 682460
rect 1140 682390 1160 682460
rect 1230 682390 1250 682460
rect 1320 682390 1340 682460
rect 1410 682390 1430 682460
rect 1500 682390 1520 682460
rect 1590 682390 1610 682460
rect 1680 682390 1700 682460
rect -800 682370 1700 682390
rect -800 682300 350 682370
rect 420 682300 440 682370
rect 510 682300 530 682370
rect 600 682300 620 682370
rect 690 682300 710 682370
rect 780 682300 800 682370
rect 870 682300 890 682370
rect 960 682300 980 682370
rect 1050 682300 1070 682370
rect 1140 682300 1160 682370
rect 1230 682300 1250 682370
rect 1320 682300 1340 682370
rect 1410 682300 1430 682370
rect 1500 682300 1520 682370
rect 1590 682300 1610 682370
rect 1680 682300 1700 682370
rect -800 682280 1700 682300
rect -800 682210 350 682280
rect 420 682210 440 682280
rect 510 682210 530 682280
rect 600 682210 620 682280
rect 690 682210 710 682280
rect 780 682210 800 682280
rect 870 682210 890 682280
rect 960 682210 980 682280
rect 1050 682210 1070 682280
rect 1140 682210 1160 682280
rect 1230 682210 1250 682280
rect 1320 682210 1340 682280
rect 1410 682210 1430 682280
rect 1500 682210 1520 682280
rect 1590 682210 1610 682280
rect 1680 682210 1700 682280
rect -800 682190 1700 682210
rect -800 682120 350 682190
rect 420 682120 440 682190
rect 510 682120 530 682190
rect 600 682120 620 682190
rect 690 682120 710 682190
rect 780 682120 800 682190
rect 870 682120 890 682190
rect 960 682120 980 682190
rect 1050 682120 1070 682190
rect 1140 682120 1160 682190
rect 1230 682120 1250 682190
rect 1320 682120 1340 682190
rect 1410 682120 1430 682190
rect 1500 682120 1520 682190
rect 1590 682120 1610 682190
rect 1680 682120 1700 682190
rect -800 682100 1700 682120
rect -800 682030 350 682100
rect 420 682030 440 682100
rect 510 682030 530 682100
rect 600 682030 620 682100
rect 690 682030 710 682100
rect 780 682030 800 682100
rect 870 682030 890 682100
rect 960 682030 980 682100
rect 1050 682030 1070 682100
rect 1140 682030 1160 682100
rect 1230 682030 1250 682100
rect 1320 682030 1340 682100
rect 1410 682030 1430 682100
rect 1500 682030 1520 682100
rect 1590 682030 1610 682100
rect 1680 682030 1700 682100
rect -800 682010 1700 682030
rect -800 681940 350 682010
rect 420 681940 440 682010
rect 510 681940 530 682010
rect 600 681940 620 682010
rect 690 681940 710 682010
rect 780 681940 800 682010
rect 870 681940 890 682010
rect 960 681940 980 682010
rect 1050 681940 1070 682010
rect 1140 681940 1160 682010
rect 1230 681940 1250 682010
rect 1320 681940 1340 682010
rect 1410 681940 1430 682010
rect 1500 681940 1520 682010
rect 1590 681940 1610 682010
rect 1680 681940 1700 682010
rect -800 681920 1700 681940
rect -800 681850 350 681920
rect 420 681850 440 681920
rect 510 681850 530 681920
rect 600 681850 620 681920
rect 690 681850 710 681920
rect 780 681850 800 681920
rect 870 681850 890 681920
rect 960 681850 980 681920
rect 1050 681850 1070 681920
rect 1140 681850 1160 681920
rect 1230 681850 1250 681920
rect 1320 681850 1340 681920
rect 1410 681850 1430 681920
rect 1500 681850 1520 681920
rect 1590 681850 1610 681920
rect 1680 681850 1700 681920
rect -800 681830 1700 681850
rect -800 681760 350 681830
rect 420 681760 440 681830
rect 510 681760 530 681830
rect 600 681760 620 681830
rect 690 681760 710 681830
rect 780 681760 800 681830
rect 870 681760 890 681830
rect 960 681760 980 681830
rect 1050 681760 1070 681830
rect 1140 681760 1160 681830
rect 1230 681760 1250 681830
rect 1320 681760 1340 681830
rect 1410 681760 1430 681830
rect 1500 681760 1520 681830
rect 1590 681760 1610 681830
rect 1680 681760 1700 681830
rect -800 681740 1700 681760
rect -800 681670 350 681740
rect 420 681670 440 681740
rect 510 681670 530 681740
rect 600 681670 620 681740
rect 690 681670 710 681740
rect 780 681670 800 681740
rect 870 681670 890 681740
rect 960 681670 980 681740
rect 1050 681670 1070 681740
rect 1140 681670 1160 681740
rect 1230 681670 1250 681740
rect 1320 681670 1340 681740
rect 1410 681670 1430 681740
rect 1500 681670 1520 681740
rect 1590 681670 1610 681740
rect 1680 681670 1700 681740
rect -800 680242 1700 681670
rect 582300 681110 584800 682984
rect 582300 681040 582680 681110
rect 582750 681040 582770 681110
rect 582840 681040 582860 681110
rect 582930 681040 582950 681110
rect 583020 681040 583040 681110
rect 583110 681040 584800 681110
rect 582300 681020 584800 681040
rect 582300 680950 582680 681020
rect 582750 680950 582770 681020
rect 582840 680950 582860 681020
rect 582930 680950 582950 681020
rect 583020 680950 583040 681020
rect 583110 680950 584800 681020
rect 582300 680930 584800 680950
rect 582300 680860 582680 680930
rect 582750 680860 582770 680930
rect 582840 680860 582860 680930
rect 582930 680860 582950 680930
rect 583020 680860 583040 680930
rect 583110 680860 584800 680930
rect 582300 680840 584800 680860
rect 582300 680770 582680 680840
rect 582750 680770 582770 680840
rect 582840 680770 582860 680840
rect 582930 680770 582950 680840
rect 583020 680770 583040 680840
rect 583110 680770 584800 680840
rect 582300 680750 584800 680770
rect 582300 680680 582680 680750
rect 582750 680680 582770 680750
rect 582840 680680 582860 680750
rect 582930 680680 582950 680750
rect 583020 680680 583040 680750
rect 583110 680680 584800 680750
rect 582300 677984 584800 680680
rect 94254 650470 94574 650690
rect 94254 650400 94280 650470
rect 94350 650400 94380 650470
rect 94450 650400 94480 650470
rect 94550 650400 94574 650470
rect 94254 650380 94574 650400
rect 94254 650310 94280 650380
rect 94350 650310 94380 650380
rect 94450 650310 94480 650380
rect 94550 650310 94574 650380
rect 94254 650280 94574 650310
rect 98814 650470 99134 650690
rect 98814 650400 98838 650470
rect 98908 650400 98938 650470
rect 99008 650400 99038 650470
rect 99108 650400 99134 650470
rect 98814 650380 99134 650400
rect 98814 650310 98838 650380
rect 98908 650310 98938 650380
rect 99008 650310 99038 650380
rect 99108 650310 99134 650380
rect 98814 650280 99134 650310
rect -800 643842 1660 648642
rect 582340 640642 584800 644584
rect 583832 639784 584800 640642
rect -800 636584 312 638642
rect -800 633842 1660 636584
rect 582340 635784 583832 636642
rect 312 632584 1660 633842
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 17270 703580 17340 703650
rect 17360 703580 17430 703650
rect 17450 703580 17520 703650
rect 17540 703580 17610 703650
rect 17630 703580 17700 703650
rect 17720 703580 17790 703650
rect 17810 703580 17880 703650
rect 17900 703580 17970 703650
rect 17990 703580 18060 703650
rect 18080 703580 18150 703650
rect 18170 703580 18240 703650
rect 18260 703580 18330 703650
rect 18350 703580 18420 703650
rect 18440 703580 18510 703650
rect 18530 703580 18600 703650
rect 18620 703580 18690 703650
rect 18710 703580 18780 703650
rect 18800 703580 18870 703650
rect 18890 703580 18960 703650
rect 18980 703580 19050 703650
rect 19070 703580 19140 703650
rect 19160 703580 19230 703650
rect 17270 703490 17340 703560
rect 17360 703490 17430 703560
rect 17450 703490 17520 703560
rect 17540 703490 17610 703560
rect 17630 703490 17700 703560
rect 17720 703490 17790 703560
rect 17810 703490 17880 703560
rect 17900 703490 17970 703560
rect 17990 703490 18060 703560
rect 18080 703490 18150 703560
rect 18170 703490 18240 703560
rect 18260 703490 18330 703560
rect 18350 703490 18420 703560
rect 18440 703490 18510 703560
rect 18530 703490 18600 703560
rect 18620 703490 18690 703560
rect 18710 703490 18780 703560
rect 18800 703490 18870 703560
rect 18890 703490 18960 703560
rect 18980 703490 19050 703560
rect 19070 703490 19140 703560
rect 19160 703490 19230 703560
rect 17270 703400 17340 703470
rect 17360 703400 17430 703470
rect 17450 703400 17520 703470
rect 17540 703400 17610 703470
rect 17630 703400 17700 703470
rect 17720 703400 17790 703470
rect 17810 703400 17880 703470
rect 17900 703400 17970 703470
rect 17990 703400 18060 703470
rect 18080 703400 18150 703470
rect 18170 703400 18240 703470
rect 18260 703400 18330 703470
rect 18350 703400 18420 703470
rect 18440 703400 18510 703470
rect 18530 703400 18600 703470
rect 18620 703400 18690 703470
rect 18710 703400 18780 703470
rect 18800 703400 18870 703470
rect 18890 703400 18960 703470
rect 18980 703400 19050 703470
rect 19070 703400 19140 703470
rect 19160 703400 19230 703470
rect 17270 703310 17340 703380
rect 17360 703310 17430 703380
rect 17450 703310 17520 703380
rect 17540 703310 17610 703380
rect 17630 703310 17700 703380
rect 17720 703310 17790 703380
rect 17810 703310 17880 703380
rect 17900 703310 17970 703380
rect 17990 703310 18060 703380
rect 18080 703310 18150 703380
rect 18170 703310 18240 703380
rect 18260 703310 18330 703380
rect 18350 703310 18420 703380
rect 18440 703310 18510 703380
rect 18530 703310 18600 703380
rect 18620 703310 18690 703380
rect 18710 703310 18780 703380
rect 18800 703310 18870 703380
rect 18890 703310 18960 703380
rect 18980 703310 19050 703380
rect 19070 703310 19140 703380
rect 19160 703310 19230 703380
rect 17270 703220 17340 703290
rect 17360 703220 17430 703290
rect 17450 703220 17520 703290
rect 17540 703220 17610 703290
rect 17630 703220 17700 703290
rect 17720 703220 17790 703290
rect 17810 703220 17880 703290
rect 17900 703220 17970 703290
rect 17990 703220 18060 703290
rect 18080 703220 18150 703290
rect 18170 703220 18240 703290
rect 18260 703220 18330 703290
rect 18350 703220 18420 703290
rect 18440 703220 18510 703290
rect 18530 703220 18600 703290
rect 18620 703220 18690 703290
rect 18710 703220 18780 703290
rect 18800 703220 18870 703290
rect 18890 703220 18960 703290
rect 18980 703220 19050 703290
rect 19070 703220 19140 703290
rect 19160 703220 19230 703290
rect 17270 703130 17340 703200
rect 17360 703130 17430 703200
rect 17450 703130 17520 703200
rect 17540 703130 17610 703200
rect 17630 703130 17700 703200
rect 17720 703130 17790 703200
rect 17810 703130 17880 703200
rect 17900 703130 17970 703200
rect 17990 703130 18060 703200
rect 18080 703130 18150 703200
rect 18170 703130 18240 703200
rect 18260 703130 18330 703200
rect 18350 703130 18420 703200
rect 18440 703130 18510 703200
rect 18530 703130 18600 703200
rect 18620 703130 18690 703200
rect 18710 703130 18780 703200
rect 18800 703130 18870 703200
rect 18890 703130 18960 703200
rect 18980 703130 19050 703200
rect 19070 703130 19140 703200
rect 19160 703130 19230 703200
rect 17270 703040 17340 703110
rect 17360 703040 17430 703110
rect 17450 703040 17520 703110
rect 17540 703040 17610 703110
rect 17630 703040 17700 703110
rect 17720 703040 17790 703110
rect 17810 703040 17880 703110
rect 17900 703040 17970 703110
rect 17990 703040 18060 703110
rect 18080 703040 18150 703110
rect 18170 703040 18240 703110
rect 18260 703040 18330 703110
rect 18350 703040 18420 703110
rect 18440 703040 18510 703110
rect 18530 703040 18600 703110
rect 18620 703040 18690 703110
rect 18710 703040 18780 703110
rect 18800 703040 18870 703110
rect 18890 703040 18960 703110
rect 18980 703040 19050 703110
rect 19070 703040 19140 703110
rect 19160 703040 19230 703110
rect 17270 702950 17340 703020
rect 17360 702950 17430 703020
rect 17450 702950 17520 703020
rect 17540 702950 17610 703020
rect 17630 702950 17700 703020
rect 17720 702950 17790 703020
rect 17810 702950 17880 703020
rect 17900 702950 17970 703020
rect 17990 702950 18060 703020
rect 18080 702950 18150 703020
rect 18170 702950 18240 703020
rect 18260 702950 18330 703020
rect 18350 702950 18420 703020
rect 18440 702950 18510 703020
rect 18530 702950 18600 703020
rect 18620 702950 18690 703020
rect 18710 702950 18780 703020
rect 18800 702950 18870 703020
rect 18890 702950 18960 703020
rect 18980 702950 19050 703020
rect 19070 702950 19140 703020
rect 19160 702950 19230 703020
rect 17270 702860 17340 702930
rect 17360 702860 17430 702930
rect 17450 702860 17520 702930
rect 17540 702860 17610 702930
rect 17630 702860 17700 702930
rect 17720 702860 17790 702930
rect 17810 702860 17880 702930
rect 17900 702860 17970 702930
rect 17990 702860 18060 702930
rect 18080 702860 18150 702930
rect 18170 702860 18240 702930
rect 18260 702860 18330 702930
rect 18350 702860 18420 702930
rect 18440 702860 18510 702930
rect 18530 702860 18600 702930
rect 18620 702860 18690 702930
rect 18710 702860 18780 702930
rect 18800 702860 18870 702930
rect 18890 702860 18960 702930
rect 18980 702860 19050 702930
rect 19070 702860 19140 702930
rect 19160 702860 19230 702930
rect 17270 702770 17340 702840
rect 17360 702770 17430 702840
rect 17450 702770 17520 702840
rect 17540 702770 17610 702840
rect 17630 702770 17700 702840
rect 17720 702770 17790 702840
rect 17810 702770 17880 702840
rect 17900 702770 17970 702840
rect 17990 702770 18060 702840
rect 18080 702770 18150 702840
rect 18170 702770 18240 702840
rect 18260 702770 18330 702840
rect 18350 702770 18420 702840
rect 18440 702770 18510 702840
rect 18530 702770 18600 702840
rect 18620 702770 18690 702840
rect 18710 702770 18780 702840
rect 18800 702770 18870 702840
rect 18890 702770 18960 702840
rect 18980 702770 19050 702840
rect 19070 702770 19140 702840
rect 19160 702770 19230 702840
rect 17270 702680 17340 702750
rect 17360 702680 17430 702750
rect 17450 702680 17520 702750
rect 17540 702680 17610 702750
rect 17630 702680 17700 702750
rect 17720 702680 17790 702750
rect 17810 702680 17880 702750
rect 17900 702680 17970 702750
rect 17990 702680 18060 702750
rect 18080 702680 18150 702750
rect 18170 702680 18240 702750
rect 18260 702680 18330 702750
rect 18350 702680 18420 702750
rect 18440 702680 18510 702750
rect 18530 702680 18600 702750
rect 18620 702680 18690 702750
rect 18710 702680 18780 702750
rect 18800 702680 18870 702750
rect 18890 702680 18960 702750
rect 18980 702680 19050 702750
rect 19070 702680 19140 702750
rect 19160 702680 19230 702750
rect 17270 702590 17340 702660
rect 17360 702590 17430 702660
rect 17450 702590 17520 702660
rect 17540 702590 17610 702660
rect 17630 702590 17700 702660
rect 17720 702590 17790 702660
rect 17810 702590 17880 702660
rect 17900 702590 17970 702660
rect 17990 702590 18060 702660
rect 18080 702590 18150 702660
rect 18170 702590 18240 702660
rect 18260 702590 18330 702660
rect 18350 702590 18420 702660
rect 18440 702590 18510 702660
rect 18530 702590 18600 702660
rect 18620 702590 18690 702660
rect 18710 702590 18780 702660
rect 18800 702590 18870 702660
rect 18890 702590 18960 702660
rect 18980 702590 19050 702660
rect 19070 702590 19140 702660
rect 19160 702590 19230 702660
rect 17270 702500 17340 702570
rect 17360 702500 17430 702570
rect 17450 702500 17520 702570
rect 17540 702500 17610 702570
rect 17630 702500 17700 702570
rect 17720 702500 17790 702570
rect 17810 702500 17880 702570
rect 17900 702500 17970 702570
rect 17990 702500 18060 702570
rect 18080 702500 18150 702570
rect 18170 702500 18240 702570
rect 18260 702500 18330 702570
rect 18350 702500 18420 702570
rect 18440 702500 18510 702570
rect 18530 702500 18600 702570
rect 18620 702500 18690 702570
rect 18710 702500 18780 702570
rect 18800 702500 18870 702570
rect 18890 702500 18960 702570
rect 18980 702500 19050 702570
rect 19070 702500 19140 702570
rect 19160 702500 19230 702570
rect 17270 702410 17340 702480
rect 17360 702410 17430 702480
rect 17450 702410 17520 702480
rect 17540 702410 17610 702480
rect 17630 702410 17700 702480
rect 17720 702410 17790 702480
rect 17810 702410 17880 702480
rect 17900 702410 17970 702480
rect 17990 702410 18060 702480
rect 18080 702410 18150 702480
rect 18170 702410 18240 702480
rect 18260 702410 18330 702480
rect 18350 702410 18420 702480
rect 18440 702410 18510 702480
rect 18530 702410 18600 702480
rect 18620 702410 18690 702480
rect 18710 702410 18780 702480
rect 18800 702410 18870 702480
rect 18890 702410 18960 702480
rect 18980 702410 19050 702480
rect 19070 702410 19140 702480
rect 19160 702410 19230 702480
rect 17270 702320 17340 702390
rect 17360 702320 17430 702390
rect 17450 702320 17520 702390
rect 17540 702320 17610 702390
rect 17630 702320 17700 702390
rect 17720 702320 17790 702390
rect 17810 702320 17880 702390
rect 17900 702320 17970 702390
rect 17990 702320 18060 702390
rect 18080 702320 18150 702390
rect 18170 702320 18240 702390
rect 18260 702320 18330 702390
rect 18350 702320 18420 702390
rect 18440 702320 18510 702390
rect 18530 702320 18600 702390
rect 18620 702320 18690 702390
rect 18710 702320 18780 702390
rect 18800 702320 18870 702390
rect 18890 702320 18960 702390
rect 18980 702320 19050 702390
rect 19070 702320 19140 702390
rect 19160 702320 19230 702390
rect 68352 703500 68652 703800
rect 68852 703500 69152 703800
rect 69352 703500 69652 703800
rect 69852 703500 70152 703800
rect 70352 703500 70652 703800
rect 70852 703500 71152 703800
rect 71352 703500 71652 703800
rect 71852 703500 72152 703800
rect 72352 703500 72652 703800
rect 72852 703500 73152 703800
rect 68352 703000 68652 703300
rect 68852 703000 69152 703300
rect 69352 703000 69652 703300
rect 69852 703000 70152 703300
rect 70352 703000 70652 703300
rect 70852 703000 71152 703300
rect 71352 703000 71652 703300
rect 71852 703000 72152 703300
rect 72352 703000 72652 703300
rect 72852 703000 73152 703300
rect 68352 702500 68652 702800
rect 68852 702500 69152 702800
rect 69352 702500 69652 702800
rect 69852 702500 70152 702800
rect 70352 702500 70652 702800
rect 70852 702500 71152 702800
rect 71352 702500 71652 702800
rect 71852 702500 72152 702800
rect 72352 702500 72652 702800
rect 72852 702500 73152 702800
rect 120352 703500 120652 703800
rect 120852 703500 121152 703800
rect 121352 703500 121652 703800
rect 121852 703500 122152 703800
rect 122352 703500 122652 703800
rect 122852 703500 123152 703800
rect 123352 703500 123652 703800
rect 123852 703500 124152 703800
rect 124352 703500 124652 703800
rect 124852 703500 125152 703800
rect 120352 703000 120652 703300
rect 120852 703000 121152 703300
rect 121352 703000 121652 703300
rect 121852 703000 122152 703300
rect 122352 703000 122652 703300
rect 122852 703000 123152 703300
rect 123352 703000 123652 703300
rect 123852 703000 124152 703300
rect 124352 703000 124652 703300
rect 124852 703000 125152 703300
rect 120352 702500 120652 702800
rect 120852 702500 121152 702800
rect 121352 702500 121652 702800
rect 121852 702500 122152 702800
rect 122352 702500 122652 702800
rect 122852 702500 123152 702800
rect 123352 702500 123652 702800
rect 123852 702500 124152 702800
rect 124352 702500 124652 702800
rect 124852 702500 125152 702800
rect 415760 703040 415830 703110
rect 415850 703040 415920 703110
rect 415940 703040 416010 703110
rect 416030 703040 416100 703110
rect 416120 703040 416190 703110
rect 415760 702950 415830 703020
rect 415850 702950 415920 703020
rect 415940 702950 416010 703020
rect 416030 702950 416100 703020
rect 416120 702950 416190 703020
rect 415760 702860 415830 702930
rect 415850 702860 415920 702930
rect 415940 702860 416010 702930
rect 416030 702860 416100 702930
rect 416120 702860 416190 702930
rect 415760 702770 415830 702840
rect 415850 702770 415920 702840
rect 415940 702770 416010 702840
rect 416030 702770 416100 702840
rect 416120 702770 416190 702840
rect 415760 702680 415830 702750
rect 415850 702680 415920 702750
rect 415940 702680 416010 702750
rect 416030 702680 416100 702750
rect 416120 702680 416190 702750
rect 467010 703040 467080 703110
rect 467100 703040 467170 703110
rect 467190 703040 467260 703110
rect 467280 703040 467350 703110
rect 467370 703040 467440 703110
rect 467010 702950 467080 703020
rect 467100 702950 467170 703020
rect 467190 702950 467260 703020
rect 467280 702950 467350 703020
rect 467370 702950 467440 703020
rect 467010 702860 467080 702930
rect 467100 702860 467170 702930
rect 467190 702860 467260 702930
rect 467280 702860 467350 702930
rect 467370 702860 467440 702930
rect 467010 702770 467080 702840
rect 467100 702770 467170 702840
rect 467190 702770 467260 702840
rect 467280 702770 467350 702840
rect 467370 702770 467440 702840
rect 467010 702680 467080 702750
rect 467100 702680 467170 702750
rect 467190 702680 467260 702750
rect 467280 702680 467350 702750
rect 467370 702680 467440 702750
rect 569140 703040 569210 703110
rect 569230 703040 569300 703110
rect 569320 703040 569390 703110
rect 569410 703040 569480 703110
rect 569500 703040 569570 703110
rect 569140 702950 569210 703020
rect 569230 702950 569300 703020
rect 569320 702950 569390 703020
rect 569410 702950 569480 703020
rect 569500 702950 569570 703020
rect 569140 702860 569210 702930
rect 569230 702860 569300 702930
rect 569320 702860 569390 702930
rect 569410 702860 569480 702930
rect 569500 702860 569570 702930
rect 569140 702770 569210 702840
rect 569230 702770 569300 702840
rect 569320 702770 569390 702840
rect 569410 702770 569480 702840
rect 569500 702770 569570 702840
rect 569140 702680 569210 702750
rect 569230 702680 569300 702750
rect 569320 702680 569390 702750
rect 569410 702680 569480 702750
rect 569500 702680 569570 702750
rect 224744 697350 224814 697420
rect 224834 697350 224904 697420
rect 224924 697350 224994 697420
rect 225014 697350 225084 697420
rect 225104 697350 225174 697420
rect 234630 697350 234700 697420
rect 234720 697350 234790 697420
rect 234810 697350 234880 697420
rect 234900 697350 234970 697420
rect 234990 697350 235060 697420
rect 224744 697260 224814 697330
rect 224834 697260 224904 697330
rect 224924 697260 224994 697330
rect 225014 697260 225084 697330
rect 225104 697260 225174 697330
rect 234630 697260 234700 697330
rect 234720 697260 234790 697330
rect 234810 697260 234880 697330
rect 234900 697260 234970 697330
rect 234990 697260 235060 697330
rect 224744 697170 224814 697240
rect 224834 697170 224904 697240
rect 224924 697170 224994 697240
rect 225014 697170 225084 697240
rect 225104 697170 225174 697240
rect 234630 697170 234700 697240
rect 234720 697170 234790 697240
rect 234810 697170 234880 697240
rect 234900 697170 234970 697240
rect 234990 697170 235060 697240
rect 224744 697080 224814 697150
rect 224834 697080 224904 697150
rect 224924 697080 224994 697150
rect 225014 697080 225084 697150
rect 225104 697080 225174 697150
rect 234630 697080 234700 697150
rect 234720 697080 234790 697150
rect 234810 697080 234880 697150
rect 234900 697080 234970 697150
rect 234990 697080 235060 697150
rect 224744 696990 224814 697060
rect 224834 696990 224904 697060
rect 224924 696990 224994 697060
rect 225014 696990 225084 697060
rect 225104 696990 225174 697060
rect 234630 696990 234700 697060
rect 234720 696990 234790 697060
rect 234810 696990 234880 697060
rect 234900 696990 234970 697060
rect 234990 696990 235060 697060
rect 224744 696133 224814 696203
rect 224834 696133 224904 696203
rect 224924 696133 224994 696203
rect 225014 696133 225084 696203
rect 225104 696133 225174 696203
rect 234630 696133 234700 696203
rect 234720 696133 234790 696203
rect 234810 696133 234880 696203
rect 234900 696133 234970 696203
rect 234990 696133 235060 696203
rect 224744 696043 224814 696113
rect 224834 696043 224904 696113
rect 224924 696043 224994 696113
rect 225014 696043 225084 696113
rect 225104 696043 225174 696113
rect 234630 696043 234700 696113
rect 234720 696043 234790 696113
rect 234810 696043 234880 696113
rect 234900 696043 234970 696113
rect 234990 696043 235060 696113
rect 224744 695953 224814 696023
rect 224834 695953 224904 696023
rect 224924 695953 224994 696023
rect 225014 695953 225084 696023
rect 225104 695953 225174 696023
rect 234630 695953 234700 696023
rect 234720 695953 234790 696023
rect 234810 695953 234880 696023
rect 234900 695953 234970 696023
rect 234990 695953 235060 696023
rect 224744 695863 224814 695933
rect 224834 695863 224904 695933
rect 224924 695863 224994 695933
rect 225014 695863 225084 695933
rect 225104 695863 225174 695933
rect 234630 695863 234700 695933
rect 234720 695863 234790 695933
rect 234810 695863 234880 695933
rect 234900 695863 234970 695933
rect 234990 695863 235060 695933
rect 224744 695773 224814 695843
rect 224834 695773 224904 695843
rect 224924 695773 224994 695843
rect 225014 695773 225084 695843
rect 225104 695773 225174 695843
rect 234630 695773 234700 695843
rect 234720 695773 234790 695843
rect 234810 695773 234880 695843
rect 234900 695773 234970 695843
rect 234990 695773 235060 695843
rect 224744 695068 224814 695138
rect 224834 695068 224904 695138
rect 224924 695068 224994 695138
rect 225014 695068 225084 695138
rect 225104 695068 225174 695138
rect 234630 695068 234700 695138
rect 234720 695068 234790 695138
rect 234810 695068 234880 695138
rect 234900 695068 234970 695138
rect 234990 695068 235060 695138
rect 224744 694978 224814 695048
rect 224834 694978 224904 695048
rect 224924 694978 224994 695048
rect 225014 694978 225084 695048
rect 225104 694978 225174 695048
rect 234630 694978 234700 695048
rect 234720 694978 234790 695048
rect 234810 694978 234880 695048
rect 234900 694978 234970 695048
rect 234990 694978 235060 695048
rect 224744 694888 224814 694958
rect 224834 694888 224904 694958
rect 224924 694888 224994 694958
rect 225014 694888 225084 694958
rect 225104 694888 225174 694958
rect 234630 694888 234700 694958
rect 234720 694888 234790 694958
rect 234810 694888 234880 694958
rect 234900 694888 234970 694958
rect 234990 694888 235060 694958
rect 224744 694798 224814 694868
rect 224834 694798 224904 694868
rect 224924 694798 224994 694868
rect 225014 694798 225084 694868
rect 225104 694798 225174 694868
rect 234630 694798 234700 694868
rect 234720 694798 234790 694868
rect 234810 694798 234880 694868
rect 234900 694798 234970 694868
rect 234990 694798 235060 694868
rect 224744 694708 224814 694778
rect 224834 694708 224904 694778
rect 224924 694708 224994 694778
rect 225014 694708 225084 694778
rect 225104 694708 225174 694778
rect 234630 694708 234700 694778
rect 234720 694708 234790 694778
rect 234810 694708 234880 694778
rect 234900 694708 234970 694778
rect 234990 694708 235060 694778
rect 224744 693362 224814 693432
rect 224834 693362 224904 693432
rect 224924 693362 224994 693432
rect 225014 693362 225084 693432
rect 225104 693362 225174 693432
rect 234630 693362 234700 693432
rect 234720 693362 234790 693432
rect 234810 693362 234880 693432
rect 234900 693362 234970 693432
rect 234990 693362 235060 693432
rect 224744 693272 224814 693342
rect 224834 693272 224904 693342
rect 224924 693272 224994 693342
rect 225014 693272 225084 693342
rect 225104 693272 225174 693342
rect 234630 693272 234700 693342
rect 234720 693272 234790 693342
rect 234810 693272 234880 693342
rect 234900 693272 234970 693342
rect 234990 693272 235060 693342
rect 224744 693182 224814 693252
rect 224834 693182 224904 693252
rect 224924 693182 224994 693252
rect 225014 693182 225084 693252
rect 225104 693182 225174 693252
rect 234630 693182 234700 693252
rect 234720 693182 234790 693252
rect 234810 693182 234880 693252
rect 234900 693182 234970 693252
rect 234990 693182 235060 693252
rect 224744 693092 224814 693162
rect 224834 693092 224904 693162
rect 224924 693092 224994 693162
rect 225014 693092 225084 693162
rect 225104 693092 225174 693162
rect 234630 693092 234700 693162
rect 234720 693092 234790 693162
rect 234810 693092 234880 693162
rect 234900 693092 234970 693162
rect 234990 693092 235060 693162
rect 224744 693002 224814 693072
rect 224834 693002 224904 693072
rect 224924 693002 224994 693072
rect 225014 693002 225084 693072
rect 225104 693002 225174 693072
rect 234630 693002 234700 693072
rect 234720 693002 234790 693072
rect 234810 693002 234880 693072
rect 234900 693002 234970 693072
rect 234990 693002 235060 693072
rect 224744 691648 224814 691718
rect 224834 691648 224904 691718
rect 224924 691648 224994 691718
rect 225014 691648 225084 691718
rect 225104 691648 225174 691718
rect 234630 691648 234700 691718
rect 234720 691648 234790 691718
rect 234810 691648 234880 691718
rect 234900 691648 234970 691718
rect 234990 691648 235060 691718
rect 165360 691510 165430 691580
rect 165460 691510 165530 691580
rect 165560 691510 165630 691580
rect 165660 691510 165730 691580
rect 165760 691510 165830 691580
rect 165860 691510 165930 691580
rect 165960 691510 166030 691580
rect 166060 691510 166130 691580
rect 166160 691510 166230 691580
rect 166260 691510 166330 691580
rect 166360 691510 166430 691580
rect 166460 691510 166530 691580
rect 166560 691510 166630 691580
rect 166660 691510 166730 691580
rect 166760 691510 166830 691580
rect 166860 691510 166930 691580
rect 166960 691510 167030 691580
rect 167060 691510 167130 691580
rect 167160 691510 167230 691580
rect 167260 691510 167330 691580
rect 167360 691510 167430 691580
rect 167460 691510 167530 691580
rect 167560 691510 167630 691580
rect 167660 691510 167730 691580
rect 167760 691510 167830 691580
rect 167860 691510 167930 691580
rect 167960 691510 168030 691580
rect 168060 691510 168130 691580
rect 168160 691510 168230 691580
rect 168260 691510 168330 691580
rect 168360 691510 168430 691580
rect 168460 691510 168530 691580
rect 168560 691510 168630 691580
rect 168660 691510 168730 691580
rect 168760 691510 168830 691580
rect 168860 691510 168930 691580
rect 168960 691510 169030 691580
rect 169060 691510 169130 691580
rect 169160 691510 169230 691580
rect 169260 691510 169330 691580
rect 169360 691510 169430 691580
rect 169460 691510 169530 691580
rect 169560 691510 169630 691580
rect 169660 691510 169730 691580
rect 169760 691510 169830 691580
rect 169860 691510 169930 691580
rect 169960 691510 170030 691580
rect 170060 691510 170130 691580
rect 170160 691510 170230 691580
rect 170260 691510 170330 691580
rect 170360 691510 170430 691580
rect 170460 691510 170530 691580
rect 165360 691400 165430 691470
rect 165460 691400 165530 691470
rect 165560 691400 165630 691470
rect 165660 691400 165730 691470
rect 165760 691400 165830 691470
rect 165860 691400 165930 691470
rect 165960 691400 166030 691470
rect 166060 691400 166130 691470
rect 166160 691400 166230 691470
rect 166260 691400 166330 691470
rect 166360 691400 166430 691470
rect 166460 691400 166530 691470
rect 166560 691400 166630 691470
rect 166660 691400 166730 691470
rect 166760 691400 166830 691470
rect 166860 691400 166930 691470
rect 166960 691400 167030 691470
rect 167060 691400 167130 691470
rect 167160 691400 167230 691470
rect 167260 691400 167330 691470
rect 167360 691400 167430 691470
rect 167460 691400 167530 691470
rect 167560 691400 167630 691470
rect 167660 691400 167730 691470
rect 167760 691400 167830 691470
rect 167860 691400 167930 691470
rect 167960 691400 168030 691470
rect 168060 691400 168130 691470
rect 168160 691400 168230 691470
rect 168260 691400 168330 691470
rect 168360 691400 168430 691470
rect 168460 691400 168530 691470
rect 168560 691400 168630 691470
rect 168660 691400 168730 691470
rect 168760 691400 168830 691470
rect 168860 691400 168930 691470
rect 168960 691400 169030 691470
rect 169060 691400 169130 691470
rect 169160 691400 169230 691470
rect 169260 691400 169330 691470
rect 169360 691400 169430 691470
rect 169460 691400 169530 691470
rect 169560 691400 169630 691470
rect 169660 691400 169730 691470
rect 169760 691400 169830 691470
rect 169860 691400 169930 691470
rect 169960 691400 170030 691470
rect 170060 691400 170130 691470
rect 170160 691400 170230 691470
rect 170260 691400 170330 691470
rect 170360 691400 170430 691470
rect 170460 691400 170530 691470
rect 224744 691558 224814 691628
rect 224834 691558 224904 691628
rect 224924 691558 224994 691628
rect 225014 691558 225084 691628
rect 225104 691558 225174 691628
rect 234630 691558 234700 691628
rect 234720 691558 234790 691628
rect 234810 691558 234880 691628
rect 234900 691558 234970 691628
rect 234990 691558 235060 691628
rect 224744 691468 224814 691538
rect 224834 691468 224904 691538
rect 224924 691468 224994 691538
rect 225014 691468 225084 691538
rect 225104 691468 225174 691538
rect 234630 691468 234700 691538
rect 234720 691468 234790 691538
rect 234810 691468 234880 691538
rect 234900 691468 234970 691538
rect 234990 691468 235060 691538
rect 224744 691378 224814 691448
rect 224834 691378 224904 691448
rect 224924 691378 224994 691448
rect 225014 691378 225084 691448
rect 225104 691378 225174 691448
rect 234630 691378 234700 691448
rect 234720 691378 234790 691448
rect 234810 691378 234880 691448
rect 234900 691378 234970 691448
rect 234990 691378 235060 691448
rect 224744 691288 224814 691358
rect 224834 691288 224904 691358
rect 224924 691288 224994 691358
rect 225014 691288 225084 691358
rect 225104 691288 225174 691358
rect 234630 691288 234700 691358
rect 234720 691288 234790 691358
rect 234810 691288 234880 691358
rect 234900 691288 234970 691358
rect 234990 691288 235060 691358
rect 165620 690000 165690 690070
rect 165720 690000 165790 690070
rect 165820 690000 165890 690070
rect 165920 690000 165990 690070
rect 166020 690000 166090 690070
rect 166120 690000 166190 690070
rect 166220 690000 166290 690070
rect 166320 690000 166390 690070
rect 166420 690000 166490 690070
rect 166520 690000 166590 690070
rect 166620 690000 166690 690070
rect 166720 690000 166790 690070
rect 166820 690000 166890 690070
rect 166920 690000 166990 690070
rect 167020 690000 167090 690070
rect 167120 690000 167190 690070
rect 167220 690000 167290 690070
rect 167320 690000 167390 690070
rect 167420 690000 167490 690070
rect 167520 690000 167590 690070
rect 167620 690000 167690 690070
rect 167720 690000 167790 690070
rect 167820 690000 167890 690070
rect 167920 690000 167990 690070
rect 168020 690000 168090 690070
rect 168120 690000 168190 690070
rect 168220 690000 168290 690070
rect 168320 690000 168390 690070
rect 168420 690000 168490 690070
rect 168520 690000 168590 690070
rect 168620 690000 168690 690070
rect 168720 690000 168790 690070
rect 168820 690000 168890 690070
rect 168920 690000 168990 690070
rect 169020 690000 169090 690070
rect 169120 690000 169190 690070
rect 169220 690000 169290 690070
rect 169320 690000 169390 690070
rect 169420 690000 169490 690070
rect 169520 690000 169590 690070
rect 169620 690000 169690 690070
rect 169720 690000 169790 690070
rect 169820 690000 169890 690070
rect 169920 690000 169990 690070
rect 170020 690000 170090 690070
rect 170120 690000 170190 690070
rect 170220 690000 170290 690070
rect 170320 690000 170390 690070
rect 170420 690000 170490 690070
rect 165620 689900 165690 689970
rect 165720 689900 165790 689970
rect 165820 689900 165890 689970
rect 165920 689900 165990 689970
rect 166020 689900 166090 689970
rect 166120 689900 166190 689970
rect 166220 689900 166290 689970
rect 166320 689900 166390 689970
rect 166420 689900 166490 689970
rect 166520 689900 166590 689970
rect 166620 689900 166690 689970
rect 166720 689900 166790 689970
rect 166820 689900 166890 689970
rect 166920 689900 166990 689970
rect 167020 689900 167090 689970
rect 167120 689900 167190 689970
rect 167220 689900 167290 689970
rect 167320 689900 167390 689970
rect 167420 689900 167490 689970
rect 167520 689900 167590 689970
rect 167620 689900 167690 689970
rect 167720 689900 167790 689970
rect 167820 689900 167890 689970
rect 167920 689900 167990 689970
rect 168020 689900 168090 689970
rect 168120 689900 168190 689970
rect 168220 689900 168290 689970
rect 168320 689900 168390 689970
rect 168420 689900 168490 689970
rect 168520 689900 168590 689970
rect 168620 689900 168690 689970
rect 168720 689900 168790 689970
rect 168820 689900 168890 689970
rect 168920 689900 168990 689970
rect 169020 689900 169090 689970
rect 169120 689900 169190 689970
rect 169220 689900 169290 689970
rect 169320 689900 169390 689970
rect 169420 689900 169490 689970
rect 169520 689900 169590 689970
rect 169620 689900 169690 689970
rect 169720 689900 169790 689970
rect 169820 689900 169890 689970
rect 169920 689900 169990 689970
rect 170020 689900 170090 689970
rect 170120 689900 170190 689970
rect 170220 689900 170290 689970
rect 170320 689900 170390 689970
rect 170420 689900 170490 689970
rect 227640 689990 227710 690060
rect 227740 689990 227810 690060
rect 227840 689990 227910 690060
rect 227940 689990 228010 690060
rect 228040 689990 228110 690060
rect 228140 689990 228210 690060
rect 228240 689990 228310 690060
rect 228340 689990 228410 690060
rect 228440 689990 228510 690060
rect 228540 689990 228610 690060
rect 228640 689990 228710 690060
rect 228740 689990 228810 690060
rect 228840 689990 228910 690060
rect 228940 689990 229010 690060
rect 229040 689990 229110 690060
rect 229140 689990 229210 690060
rect 229240 689990 229310 690060
rect 229340 689990 229410 690060
rect 229440 689990 229510 690060
rect 229540 689990 229610 690060
rect 229640 689990 229710 690060
rect 229740 689990 229810 690060
rect 229840 689990 229910 690060
rect 229940 689990 230010 690060
rect 230040 689990 230110 690060
rect 230140 689990 230210 690060
rect 230240 689990 230310 690060
rect 230340 689990 230410 690060
rect 230440 689990 230510 690060
rect 230540 689990 230610 690060
rect 230640 689990 230710 690060
rect 230740 689990 230810 690060
rect 230840 689990 230910 690060
rect 230940 689990 231010 690060
rect 231040 689990 231110 690060
rect 231140 689990 231210 690060
rect 231240 689990 231310 690060
rect 231340 689990 231410 690060
rect 231440 689990 231510 690060
rect 231540 689990 231610 690060
rect 231640 689990 231710 690060
rect 231740 689990 231810 690060
rect 231840 689990 231910 690060
rect 231940 689990 232010 690060
rect 232040 689990 232110 690060
rect 232140 689990 232210 690060
rect 232240 689990 232310 690060
rect 232340 689990 232410 690060
rect 232440 689990 232510 690060
rect 227640 689890 227710 689960
rect 227740 689890 227810 689960
rect 227840 689890 227910 689960
rect 227940 689890 228010 689960
rect 228040 689890 228110 689960
rect 228140 689890 228210 689960
rect 228240 689890 228310 689960
rect 228340 689890 228410 689960
rect 228440 689890 228510 689960
rect 228540 689890 228610 689960
rect 228640 689890 228710 689960
rect 228740 689890 228810 689960
rect 228840 689890 228910 689960
rect 228940 689890 229010 689960
rect 229040 689890 229110 689960
rect 229140 689890 229210 689960
rect 229240 689890 229310 689960
rect 229340 689890 229410 689960
rect 229440 689890 229510 689960
rect 229540 689890 229610 689960
rect 229640 689890 229710 689960
rect 229740 689890 229810 689960
rect 229840 689890 229910 689960
rect 229940 689890 230010 689960
rect 230040 689890 230110 689960
rect 230140 689890 230210 689960
rect 230240 689890 230310 689960
rect 230340 689890 230410 689960
rect 230440 689890 230510 689960
rect 230540 689890 230610 689960
rect 230640 689890 230710 689960
rect 230740 689890 230810 689960
rect 230840 689890 230910 689960
rect 230940 689890 231010 689960
rect 231040 689890 231110 689960
rect 231140 689890 231210 689960
rect 231240 689890 231310 689960
rect 231340 689890 231410 689960
rect 231440 689890 231510 689960
rect 231540 689890 231610 689960
rect 231640 689890 231710 689960
rect 231740 689890 231810 689960
rect 231840 689890 231910 689960
rect 231940 689890 232010 689960
rect 232040 689890 232110 689960
rect 232140 689890 232210 689960
rect 232240 689890 232310 689960
rect 232340 689890 232410 689960
rect 232440 689890 232510 689960
rect 350 683560 420 683630
rect 440 683560 510 683630
rect 530 683560 600 683630
rect 620 683560 690 683630
rect 710 683560 780 683630
rect 800 683560 870 683630
rect 890 683560 960 683630
rect 980 683560 1050 683630
rect 1070 683560 1140 683630
rect 1160 683560 1230 683630
rect 1250 683560 1320 683630
rect 1340 683560 1410 683630
rect 1430 683560 1500 683630
rect 1520 683560 1590 683630
rect 1610 683560 1680 683630
rect 350 683470 420 683540
rect 440 683470 510 683540
rect 530 683470 600 683540
rect 620 683470 690 683540
rect 710 683470 780 683540
rect 800 683470 870 683540
rect 890 683470 960 683540
rect 980 683470 1050 683540
rect 1070 683470 1140 683540
rect 1160 683470 1230 683540
rect 1250 683470 1320 683540
rect 1340 683470 1410 683540
rect 1430 683470 1500 683540
rect 1520 683470 1590 683540
rect 1610 683470 1680 683540
rect 350 683380 420 683450
rect 440 683380 510 683450
rect 530 683380 600 683450
rect 620 683380 690 683450
rect 710 683380 780 683450
rect 800 683380 870 683450
rect 890 683380 960 683450
rect 980 683380 1050 683450
rect 1070 683380 1140 683450
rect 1160 683380 1230 683450
rect 1250 683380 1320 683450
rect 1340 683380 1410 683450
rect 1430 683380 1500 683450
rect 1520 683380 1590 683450
rect 1610 683380 1680 683450
rect 350 683290 420 683360
rect 440 683290 510 683360
rect 530 683290 600 683360
rect 620 683290 690 683360
rect 710 683290 780 683360
rect 800 683290 870 683360
rect 890 683290 960 683360
rect 980 683290 1050 683360
rect 1070 683290 1140 683360
rect 1160 683290 1230 683360
rect 1250 683290 1320 683360
rect 1340 683290 1410 683360
rect 1430 683290 1500 683360
rect 1520 683290 1590 683360
rect 1610 683290 1680 683360
rect 350 683200 420 683270
rect 440 683200 510 683270
rect 530 683200 600 683270
rect 620 683200 690 683270
rect 710 683200 780 683270
rect 800 683200 870 683270
rect 890 683200 960 683270
rect 980 683200 1050 683270
rect 1070 683200 1140 683270
rect 1160 683200 1230 683270
rect 1250 683200 1320 683270
rect 1340 683200 1410 683270
rect 1430 683200 1500 683270
rect 1520 683200 1590 683270
rect 1610 683200 1680 683270
rect 350 683110 420 683180
rect 440 683110 510 683180
rect 530 683110 600 683180
rect 620 683110 690 683180
rect 710 683110 780 683180
rect 800 683110 870 683180
rect 890 683110 960 683180
rect 980 683110 1050 683180
rect 1070 683110 1140 683180
rect 1160 683110 1230 683180
rect 1250 683110 1320 683180
rect 1340 683110 1410 683180
rect 1430 683110 1500 683180
rect 1520 683110 1590 683180
rect 1610 683110 1680 683180
rect 350 683020 420 683090
rect 440 683020 510 683090
rect 530 683020 600 683090
rect 620 683020 690 683090
rect 710 683020 780 683090
rect 800 683020 870 683090
rect 890 683020 960 683090
rect 980 683020 1050 683090
rect 1070 683020 1140 683090
rect 1160 683020 1230 683090
rect 1250 683020 1320 683090
rect 1340 683020 1410 683090
rect 1430 683020 1500 683090
rect 1520 683020 1590 683090
rect 1610 683020 1680 683090
rect 350 682930 420 683000
rect 440 682930 510 683000
rect 530 682930 600 683000
rect 620 682930 690 683000
rect 710 682930 780 683000
rect 800 682930 870 683000
rect 890 682930 960 683000
rect 980 682930 1050 683000
rect 1070 682930 1140 683000
rect 1160 682930 1230 683000
rect 1250 682930 1320 683000
rect 1340 682930 1410 683000
rect 1430 682930 1500 683000
rect 1520 682930 1590 683000
rect 1610 682930 1680 683000
rect 350 682840 420 682910
rect 440 682840 510 682910
rect 530 682840 600 682910
rect 620 682840 690 682910
rect 710 682840 780 682910
rect 800 682840 870 682910
rect 890 682840 960 682910
rect 980 682840 1050 682910
rect 1070 682840 1140 682910
rect 1160 682840 1230 682910
rect 1250 682840 1320 682910
rect 1340 682840 1410 682910
rect 1430 682840 1500 682910
rect 1520 682840 1590 682910
rect 1610 682840 1680 682910
rect 350 682750 420 682820
rect 440 682750 510 682820
rect 530 682750 600 682820
rect 620 682750 690 682820
rect 710 682750 780 682820
rect 800 682750 870 682820
rect 890 682750 960 682820
rect 980 682750 1050 682820
rect 1070 682750 1140 682820
rect 1160 682750 1230 682820
rect 1250 682750 1320 682820
rect 1340 682750 1410 682820
rect 1430 682750 1500 682820
rect 1520 682750 1590 682820
rect 1610 682750 1680 682820
rect 350 682660 420 682730
rect 440 682660 510 682730
rect 530 682660 600 682730
rect 620 682660 690 682730
rect 710 682660 780 682730
rect 800 682660 870 682730
rect 890 682660 960 682730
rect 980 682660 1050 682730
rect 1070 682660 1140 682730
rect 1160 682660 1230 682730
rect 1250 682660 1320 682730
rect 1340 682660 1410 682730
rect 1430 682660 1500 682730
rect 1520 682660 1590 682730
rect 1610 682660 1680 682730
rect 350 682570 420 682640
rect 440 682570 510 682640
rect 530 682570 600 682640
rect 620 682570 690 682640
rect 710 682570 780 682640
rect 800 682570 870 682640
rect 890 682570 960 682640
rect 980 682570 1050 682640
rect 1070 682570 1140 682640
rect 1160 682570 1230 682640
rect 1250 682570 1320 682640
rect 1340 682570 1410 682640
rect 1430 682570 1500 682640
rect 1520 682570 1590 682640
rect 1610 682570 1680 682640
rect 350 682480 420 682550
rect 440 682480 510 682550
rect 530 682480 600 682550
rect 620 682480 690 682550
rect 710 682480 780 682550
rect 800 682480 870 682550
rect 890 682480 960 682550
rect 980 682480 1050 682550
rect 1070 682480 1140 682550
rect 1160 682480 1230 682550
rect 1250 682480 1320 682550
rect 1340 682480 1410 682550
rect 1430 682480 1500 682550
rect 1520 682480 1590 682550
rect 1610 682480 1680 682550
rect 350 682390 420 682460
rect 440 682390 510 682460
rect 530 682390 600 682460
rect 620 682390 690 682460
rect 710 682390 780 682460
rect 800 682390 870 682460
rect 890 682390 960 682460
rect 980 682390 1050 682460
rect 1070 682390 1140 682460
rect 1160 682390 1230 682460
rect 1250 682390 1320 682460
rect 1340 682390 1410 682460
rect 1430 682390 1500 682460
rect 1520 682390 1590 682460
rect 1610 682390 1680 682460
rect 350 682300 420 682370
rect 440 682300 510 682370
rect 530 682300 600 682370
rect 620 682300 690 682370
rect 710 682300 780 682370
rect 800 682300 870 682370
rect 890 682300 960 682370
rect 980 682300 1050 682370
rect 1070 682300 1140 682370
rect 1160 682300 1230 682370
rect 1250 682300 1320 682370
rect 1340 682300 1410 682370
rect 1430 682300 1500 682370
rect 1520 682300 1590 682370
rect 1610 682300 1680 682370
rect 350 682210 420 682280
rect 440 682210 510 682280
rect 530 682210 600 682280
rect 620 682210 690 682280
rect 710 682210 780 682280
rect 800 682210 870 682280
rect 890 682210 960 682280
rect 980 682210 1050 682280
rect 1070 682210 1140 682280
rect 1160 682210 1230 682280
rect 1250 682210 1320 682280
rect 1340 682210 1410 682280
rect 1430 682210 1500 682280
rect 1520 682210 1590 682280
rect 1610 682210 1680 682280
rect 350 682120 420 682190
rect 440 682120 510 682190
rect 530 682120 600 682190
rect 620 682120 690 682190
rect 710 682120 780 682190
rect 800 682120 870 682190
rect 890 682120 960 682190
rect 980 682120 1050 682190
rect 1070 682120 1140 682190
rect 1160 682120 1230 682190
rect 1250 682120 1320 682190
rect 1340 682120 1410 682190
rect 1430 682120 1500 682190
rect 1520 682120 1590 682190
rect 1610 682120 1680 682190
rect 350 682030 420 682100
rect 440 682030 510 682100
rect 530 682030 600 682100
rect 620 682030 690 682100
rect 710 682030 780 682100
rect 800 682030 870 682100
rect 890 682030 960 682100
rect 980 682030 1050 682100
rect 1070 682030 1140 682100
rect 1160 682030 1230 682100
rect 1250 682030 1320 682100
rect 1340 682030 1410 682100
rect 1430 682030 1500 682100
rect 1520 682030 1590 682100
rect 1610 682030 1680 682100
rect 350 681940 420 682010
rect 440 681940 510 682010
rect 530 681940 600 682010
rect 620 681940 690 682010
rect 710 681940 780 682010
rect 800 681940 870 682010
rect 890 681940 960 682010
rect 980 681940 1050 682010
rect 1070 681940 1140 682010
rect 1160 681940 1230 682010
rect 1250 681940 1320 682010
rect 1340 681940 1410 682010
rect 1430 681940 1500 682010
rect 1520 681940 1590 682010
rect 1610 681940 1680 682010
rect 350 681850 420 681920
rect 440 681850 510 681920
rect 530 681850 600 681920
rect 620 681850 690 681920
rect 710 681850 780 681920
rect 800 681850 870 681920
rect 890 681850 960 681920
rect 980 681850 1050 681920
rect 1070 681850 1140 681920
rect 1160 681850 1230 681920
rect 1250 681850 1320 681920
rect 1340 681850 1410 681920
rect 1430 681850 1500 681920
rect 1520 681850 1590 681920
rect 1610 681850 1680 681920
rect 350 681760 420 681830
rect 440 681760 510 681830
rect 530 681760 600 681830
rect 620 681760 690 681830
rect 710 681760 780 681830
rect 800 681760 870 681830
rect 890 681760 960 681830
rect 980 681760 1050 681830
rect 1070 681760 1140 681830
rect 1160 681760 1230 681830
rect 1250 681760 1320 681830
rect 1340 681760 1410 681830
rect 1430 681760 1500 681830
rect 1520 681760 1590 681830
rect 1610 681760 1680 681830
rect 350 681670 420 681740
rect 440 681670 510 681740
rect 530 681670 600 681740
rect 620 681670 690 681740
rect 710 681670 780 681740
rect 800 681670 870 681740
rect 890 681670 960 681740
rect 980 681670 1050 681740
rect 1070 681670 1140 681740
rect 1160 681670 1230 681740
rect 1250 681670 1320 681740
rect 1340 681670 1410 681740
rect 1430 681670 1500 681740
rect 1520 681670 1590 681740
rect 1610 681670 1680 681740
rect 582680 681040 582750 681110
rect 582770 681040 582840 681110
rect 582860 681040 582930 681110
rect 582950 681040 583020 681110
rect 583040 681040 583110 681110
rect 582680 680950 582750 681020
rect 582770 680950 582840 681020
rect 582860 680950 582930 681020
rect 582950 680950 583020 681020
rect 583040 680950 583110 681020
rect 582680 680860 582750 680930
rect 582770 680860 582840 680930
rect 582860 680860 582930 680930
rect 582950 680860 583020 680930
rect 583040 680860 583110 680930
rect 582680 680770 582750 680840
rect 582770 680770 582840 680840
rect 582860 680770 582930 680840
rect 582950 680770 583020 680840
rect 583040 680770 583110 680840
rect 582680 680680 582750 680750
rect 582770 680680 582840 680750
rect 582860 680680 582930 680750
rect 582950 680680 583020 680750
rect 583040 680680 583110 680750
rect 94280 650400 94350 650470
rect 94380 650400 94450 650470
rect 94480 650400 94550 650470
rect 94280 650310 94350 650380
rect 94380 650310 94450 650380
rect 94480 650310 94550 650380
rect 98838 650400 98908 650470
rect 98938 650400 99008 650470
rect 99038 650400 99108 650470
rect 98838 650310 98908 650380
rect 98938 650310 99008 650380
rect 99038 650310 99108 650380
<< metal4 >>
rect 68194 703800 73194 704000
rect 17246 703650 19246 703652
rect 17246 703580 17270 703650
rect 17340 703580 17360 703650
rect 17430 703580 17450 703650
rect 17520 703580 17540 703650
rect 17610 703580 17630 703650
rect 17700 703580 17720 703650
rect 17790 703580 17810 703650
rect 17880 703580 17900 703650
rect 17970 703580 17990 703650
rect 18060 703580 18080 703650
rect 18150 703580 18170 703650
rect 18240 703580 18260 703650
rect 18330 703580 18350 703650
rect 18420 703580 18440 703650
rect 18510 703580 18530 703650
rect 18600 703580 18620 703650
rect 18690 703580 18710 703650
rect 18780 703580 18800 703650
rect 18870 703580 18890 703650
rect 18960 703580 18980 703650
rect 19050 703580 19070 703650
rect 19140 703580 19160 703650
rect 19230 703580 19246 703650
rect 17246 703560 19246 703580
rect 17246 703490 17270 703560
rect 17340 703490 17360 703560
rect 17430 703490 17450 703560
rect 17520 703490 17540 703560
rect 17610 703490 17630 703560
rect 17700 703490 17720 703560
rect 17790 703490 17810 703560
rect 17880 703490 17900 703560
rect 17970 703490 17990 703560
rect 18060 703490 18080 703560
rect 18150 703490 18170 703560
rect 18240 703490 18260 703560
rect 18330 703490 18350 703560
rect 18420 703490 18440 703560
rect 18510 703490 18530 703560
rect 18600 703490 18620 703560
rect 18690 703490 18710 703560
rect 18780 703490 18800 703560
rect 18870 703490 18890 703560
rect 18960 703490 18980 703560
rect 19050 703490 19070 703560
rect 19140 703490 19160 703560
rect 19230 703490 19246 703560
rect 17246 703470 19246 703490
rect 17246 703400 17270 703470
rect 17340 703400 17360 703470
rect 17430 703400 17450 703470
rect 17520 703400 17540 703470
rect 17610 703400 17630 703470
rect 17700 703400 17720 703470
rect 17790 703400 17810 703470
rect 17880 703400 17900 703470
rect 17970 703400 17990 703470
rect 18060 703400 18080 703470
rect 18150 703400 18170 703470
rect 18240 703400 18260 703470
rect 18330 703400 18350 703470
rect 18420 703400 18440 703470
rect 18510 703400 18530 703470
rect 18600 703400 18620 703470
rect 18690 703400 18710 703470
rect 18780 703400 18800 703470
rect 18870 703400 18890 703470
rect 18960 703400 18980 703470
rect 19050 703400 19070 703470
rect 19140 703400 19160 703470
rect 19230 703400 19246 703470
rect 17246 703380 19246 703400
rect 17246 703310 17270 703380
rect 17340 703310 17360 703380
rect 17430 703310 17450 703380
rect 17520 703310 17540 703380
rect 17610 703310 17630 703380
rect 17700 703310 17720 703380
rect 17790 703310 17810 703380
rect 17880 703310 17900 703380
rect 17970 703310 17990 703380
rect 18060 703310 18080 703380
rect 18150 703310 18170 703380
rect 18240 703310 18260 703380
rect 18330 703310 18350 703380
rect 18420 703310 18440 703380
rect 18510 703310 18530 703380
rect 18600 703310 18620 703380
rect 18690 703310 18710 703380
rect 18780 703310 18800 703380
rect 18870 703310 18890 703380
rect 18960 703310 18980 703380
rect 19050 703310 19070 703380
rect 19140 703310 19160 703380
rect 19230 703310 19246 703380
rect 17246 703290 19246 703310
rect 17246 703220 17270 703290
rect 17340 703220 17360 703290
rect 17430 703220 17450 703290
rect 17520 703220 17540 703290
rect 17610 703220 17630 703290
rect 17700 703220 17720 703290
rect 17790 703220 17810 703290
rect 17880 703220 17900 703290
rect 17970 703220 17990 703290
rect 18060 703220 18080 703290
rect 18150 703220 18170 703290
rect 18240 703220 18260 703290
rect 18330 703220 18350 703290
rect 18420 703220 18440 703290
rect 18510 703220 18530 703290
rect 18600 703220 18620 703290
rect 18690 703220 18710 703290
rect 18780 703220 18800 703290
rect 18870 703220 18890 703290
rect 18960 703220 18980 703290
rect 19050 703220 19070 703290
rect 19140 703220 19160 703290
rect 19230 703220 19246 703290
rect 17246 703200 19246 703220
rect 17246 703130 17270 703200
rect 17340 703130 17360 703200
rect 17430 703130 17450 703200
rect 17520 703130 17540 703200
rect 17610 703130 17630 703200
rect 17700 703130 17720 703200
rect 17790 703130 17810 703200
rect 17880 703130 17900 703200
rect 17970 703130 17990 703200
rect 18060 703130 18080 703200
rect 18150 703130 18170 703200
rect 18240 703130 18260 703200
rect 18330 703130 18350 703200
rect 18420 703130 18440 703200
rect 18510 703130 18530 703200
rect 18600 703130 18620 703200
rect 18690 703130 18710 703200
rect 18780 703130 18800 703200
rect 18870 703130 18890 703200
rect 18960 703130 18980 703200
rect 19050 703130 19070 703200
rect 19140 703130 19160 703200
rect 19230 703130 19246 703200
rect 17246 703110 19246 703130
rect 17246 703040 17270 703110
rect 17340 703040 17360 703110
rect 17430 703040 17450 703110
rect 17520 703040 17540 703110
rect 17610 703040 17630 703110
rect 17700 703040 17720 703110
rect 17790 703040 17810 703110
rect 17880 703040 17900 703110
rect 17970 703040 17990 703110
rect 18060 703040 18080 703110
rect 18150 703040 18170 703110
rect 18240 703040 18260 703110
rect 18330 703040 18350 703110
rect 18420 703040 18440 703110
rect 18510 703040 18530 703110
rect 18600 703040 18620 703110
rect 18690 703040 18710 703110
rect 18780 703040 18800 703110
rect 18870 703040 18890 703110
rect 18960 703040 18980 703110
rect 19050 703040 19070 703110
rect 19140 703040 19160 703110
rect 19230 703040 19246 703110
rect 17246 703020 19246 703040
rect 17246 702950 17270 703020
rect 17340 702950 17360 703020
rect 17430 702950 17450 703020
rect 17520 702950 17540 703020
rect 17610 702950 17630 703020
rect 17700 702950 17720 703020
rect 17790 702950 17810 703020
rect 17880 702950 17900 703020
rect 17970 702950 17990 703020
rect 18060 702950 18080 703020
rect 18150 702950 18170 703020
rect 18240 702950 18260 703020
rect 18330 702950 18350 703020
rect 18420 702950 18440 703020
rect 18510 702950 18530 703020
rect 18600 702950 18620 703020
rect 18690 702950 18710 703020
rect 18780 702950 18800 703020
rect 18870 702950 18890 703020
rect 18960 702950 18980 703020
rect 19050 702950 19070 703020
rect 19140 702950 19160 703020
rect 19230 702950 19246 703020
rect 17246 702930 19246 702950
rect 17246 702860 17270 702930
rect 17340 702860 17360 702930
rect 17430 702860 17450 702930
rect 17520 702860 17540 702930
rect 17610 702860 17630 702930
rect 17700 702860 17720 702930
rect 17790 702860 17810 702930
rect 17880 702860 17900 702930
rect 17970 702860 17990 702930
rect 18060 702860 18080 702930
rect 18150 702860 18170 702930
rect 18240 702860 18260 702930
rect 18330 702860 18350 702930
rect 18420 702860 18440 702930
rect 18510 702860 18530 702930
rect 18600 702860 18620 702930
rect 18690 702860 18710 702930
rect 18780 702860 18800 702930
rect 18870 702860 18890 702930
rect 18960 702860 18980 702930
rect 19050 702860 19070 702930
rect 19140 702860 19160 702930
rect 19230 702860 19246 702930
rect 17246 702840 19246 702860
rect 17246 702770 17270 702840
rect 17340 702770 17360 702840
rect 17430 702770 17450 702840
rect 17520 702770 17540 702840
rect 17610 702770 17630 702840
rect 17700 702770 17720 702840
rect 17790 702770 17810 702840
rect 17880 702770 17900 702840
rect 17970 702770 17990 702840
rect 18060 702770 18080 702840
rect 18150 702770 18170 702840
rect 18240 702770 18260 702840
rect 18330 702770 18350 702840
rect 18420 702770 18440 702840
rect 18510 702770 18530 702840
rect 18600 702770 18620 702840
rect 18690 702770 18710 702840
rect 18780 702770 18800 702840
rect 18870 702770 18890 702840
rect 18960 702770 18980 702840
rect 19050 702770 19070 702840
rect 19140 702770 19160 702840
rect 19230 702770 19246 702840
rect 17246 702750 19246 702770
rect 17246 702680 17270 702750
rect 17340 702680 17360 702750
rect 17430 702680 17450 702750
rect 17520 702680 17540 702750
rect 17610 702680 17630 702750
rect 17700 702680 17720 702750
rect 17790 702680 17810 702750
rect 17880 702680 17900 702750
rect 17970 702680 17990 702750
rect 18060 702680 18080 702750
rect 18150 702680 18170 702750
rect 18240 702680 18260 702750
rect 18330 702680 18350 702750
rect 18420 702680 18440 702750
rect 18510 702680 18530 702750
rect 18600 702680 18620 702750
rect 18690 702680 18710 702750
rect 18780 702680 18800 702750
rect 18870 702680 18890 702750
rect 18960 702680 18980 702750
rect 19050 702680 19070 702750
rect 19140 702680 19160 702750
rect 19230 702680 19246 702750
rect 17246 702660 19246 702680
rect 17246 702590 17270 702660
rect 17340 702590 17360 702660
rect 17430 702590 17450 702660
rect 17520 702590 17540 702660
rect 17610 702590 17630 702660
rect 17700 702590 17720 702660
rect 17790 702590 17810 702660
rect 17880 702590 17900 702660
rect 17970 702590 17990 702660
rect 18060 702590 18080 702660
rect 18150 702590 18170 702660
rect 18240 702590 18260 702660
rect 18330 702590 18350 702660
rect 18420 702590 18440 702660
rect 18510 702590 18530 702660
rect 18600 702590 18620 702660
rect 18690 702590 18710 702660
rect 18780 702590 18800 702660
rect 18870 702590 18890 702660
rect 18960 702590 18980 702660
rect 19050 702590 19070 702660
rect 19140 702590 19160 702660
rect 19230 702590 19246 702660
rect 17246 702570 19246 702590
rect 17246 702500 17270 702570
rect 17340 702500 17360 702570
rect 17430 702500 17450 702570
rect 17520 702500 17540 702570
rect 17610 702500 17630 702570
rect 17700 702500 17720 702570
rect 17790 702500 17810 702570
rect 17880 702500 17900 702570
rect 17970 702500 17990 702570
rect 18060 702500 18080 702570
rect 18150 702500 18170 702570
rect 18240 702500 18260 702570
rect 18330 702500 18350 702570
rect 18420 702500 18440 702570
rect 18510 702500 18530 702570
rect 18600 702500 18620 702570
rect 18690 702500 18710 702570
rect 18780 702500 18800 702570
rect 18870 702500 18890 702570
rect 18960 702500 18980 702570
rect 19050 702500 19070 702570
rect 19140 702500 19160 702570
rect 19230 702500 19246 702570
rect 17246 702480 19246 702500
rect 17246 702410 17270 702480
rect 17340 702410 17360 702480
rect 17430 702410 17450 702480
rect 17520 702410 17540 702480
rect 17610 702410 17630 702480
rect 17700 702410 17720 702480
rect 17790 702410 17810 702480
rect 17880 702410 17900 702480
rect 17970 702410 17990 702480
rect 18060 702410 18080 702480
rect 18150 702410 18170 702480
rect 18240 702410 18260 702480
rect 18330 702410 18350 702480
rect 18420 702410 18440 702480
rect 18510 702410 18530 702480
rect 18600 702410 18620 702480
rect 18690 702410 18710 702480
rect 18780 702410 18800 702480
rect 18870 702410 18890 702480
rect 18960 702410 18980 702480
rect 19050 702410 19070 702480
rect 19140 702410 19160 702480
rect 19230 702410 19246 702480
rect 17246 702390 19246 702410
rect 17246 702320 17270 702390
rect 17340 702320 17360 702390
rect 17430 702320 17450 702390
rect 17520 702320 17540 702390
rect 17610 702320 17630 702390
rect 17700 702320 17720 702390
rect 17790 702320 17810 702390
rect 17880 702320 17900 702390
rect 17970 702320 17990 702390
rect 18060 702320 18080 702390
rect 18150 702320 18170 702390
rect 18240 702320 18260 702390
rect 18330 702320 18350 702390
rect 18420 702320 18440 702390
rect 18510 702320 18530 702390
rect 18600 702320 18620 702390
rect 18690 702320 18710 702390
rect 18780 702320 18800 702390
rect 18870 702320 18890 702390
rect 18960 702320 18980 702390
rect 19050 702320 19070 702390
rect 19140 702320 19160 702390
rect 19230 702320 19246 702390
rect 272 683630 14791 683653
rect 272 683560 350 683630
rect 420 683560 440 683630
rect 510 683560 530 683630
rect 600 683560 620 683630
rect 690 683560 710 683630
rect 780 683560 800 683630
rect 870 683560 890 683630
rect 960 683560 980 683630
rect 1050 683560 1070 683630
rect 1140 683560 1160 683630
rect 1230 683560 1250 683630
rect 1320 683560 1340 683630
rect 1410 683560 1430 683630
rect 1500 683560 1520 683630
rect 1590 683560 1610 683630
rect 1680 683560 14791 683630
rect 272 683540 14791 683560
rect 272 683470 350 683540
rect 420 683470 440 683540
rect 510 683470 530 683540
rect 600 683470 620 683540
rect 690 683470 710 683540
rect 780 683470 800 683540
rect 870 683470 890 683540
rect 960 683470 980 683540
rect 1050 683470 1070 683540
rect 1140 683470 1160 683540
rect 1230 683470 1250 683540
rect 1320 683470 1340 683540
rect 1410 683470 1430 683540
rect 1500 683470 1520 683540
rect 1590 683470 1610 683540
rect 1680 683470 14791 683540
rect 272 683450 14791 683470
rect 272 683380 350 683450
rect 420 683380 440 683450
rect 510 683380 530 683450
rect 600 683380 620 683450
rect 690 683380 710 683450
rect 780 683380 800 683450
rect 870 683380 890 683450
rect 960 683380 980 683450
rect 1050 683380 1070 683450
rect 1140 683380 1160 683450
rect 1230 683380 1250 683450
rect 1320 683380 1340 683450
rect 1410 683380 1430 683450
rect 1500 683380 1520 683450
rect 1590 683380 1610 683450
rect 1680 683380 14791 683450
rect 272 683360 14791 683380
rect 272 683290 350 683360
rect 420 683290 440 683360
rect 510 683290 530 683360
rect 600 683290 620 683360
rect 690 683290 710 683360
rect 780 683290 800 683360
rect 870 683290 890 683360
rect 960 683290 980 683360
rect 1050 683290 1070 683360
rect 1140 683290 1160 683360
rect 1230 683290 1250 683360
rect 1320 683290 1340 683360
rect 1410 683290 1430 683360
rect 1500 683290 1520 683360
rect 1590 683290 1610 683360
rect 1680 683290 14791 683360
rect 272 683270 14791 683290
rect 272 683200 350 683270
rect 420 683200 440 683270
rect 510 683200 530 683270
rect 600 683200 620 683270
rect 690 683200 710 683270
rect 780 683200 800 683270
rect 870 683200 890 683270
rect 960 683200 980 683270
rect 1050 683200 1070 683270
rect 1140 683200 1160 683270
rect 1230 683200 1250 683270
rect 1320 683200 1340 683270
rect 1410 683200 1430 683270
rect 1500 683200 1520 683270
rect 1590 683200 1610 683270
rect 1680 683200 14791 683270
rect 272 683180 14791 683200
rect 272 683110 350 683180
rect 420 683110 440 683180
rect 510 683110 530 683180
rect 600 683110 620 683180
rect 690 683110 710 683180
rect 780 683110 800 683180
rect 870 683110 890 683180
rect 960 683110 980 683180
rect 1050 683110 1070 683180
rect 1140 683110 1160 683180
rect 1230 683110 1250 683180
rect 1320 683110 1340 683180
rect 1410 683110 1430 683180
rect 1500 683110 1520 683180
rect 1590 683110 1610 683180
rect 1680 683110 14791 683180
rect 272 683090 14791 683110
rect 272 683020 350 683090
rect 420 683020 440 683090
rect 510 683020 530 683090
rect 600 683020 620 683090
rect 690 683020 710 683090
rect 780 683020 800 683090
rect 870 683020 890 683090
rect 960 683020 980 683090
rect 1050 683020 1070 683090
rect 1140 683020 1160 683090
rect 1230 683020 1250 683090
rect 1320 683020 1340 683090
rect 1410 683020 1430 683090
rect 1500 683020 1520 683090
rect 1590 683020 1610 683090
rect 1680 683020 14791 683090
rect 272 683000 14791 683020
rect 272 682930 350 683000
rect 420 682930 440 683000
rect 510 682930 530 683000
rect 600 682930 620 683000
rect 690 682930 710 683000
rect 780 682930 800 683000
rect 870 682930 890 683000
rect 960 682930 980 683000
rect 1050 682930 1070 683000
rect 1140 682930 1160 683000
rect 1230 682930 1250 683000
rect 1320 682930 1340 683000
rect 1410 682930 1430 683000
rect 1500 682930 1520 683000
rect 1590 682930 1610 683000
rect 1680 682930 14791 683000
rect 272 682910 14791 682930
rect 272 682840 350 682910
rect 420 682840 440 682910
rect 510 682840 530 682910
rect 600 682840 620 682910
rect 690 682840 710 682910
rect 780 682840 800 682910
rect 870 682840 890 682910
rect 960 682840 980 682910
rect 1050 682840 1070 682910
rect 1140 682840 1160 682910
rect 1230 682840 1250 682910
rect 1320 682840 1340 682910
rect 1410 682840 1430 682910
rect 1500 682840 1520 682910
rect 1590 682840 1610 682910
rect 1680 682840 14791 682910
rect 272 682820 14791 682840
rect 272 682750 350 682820
rect 420 682750 440 682820
rect 510 682750 530 682820
rect 600 682750 620 682820
rect 690 682750 710 682820
rect 780 682750 800 682820
rect 870 682750 890 682820
rect 960 682750 980 682820
rect 1050 682750 1070 682820
rect 1140 682750 1160 682820
rect 1230 682750 1250 682820
rect 1320 682750 1340 682820
rect 1410 682750 1430 682820
rect 1500 682750 1520 682820
rect 1590 682750 1610 682820
rect 1680 682750 14791 682820
rect 272 682730 14791 682750
rect 272 682660 350 682730
rect 420 682660 440 682730
rect 510 682660 530 682730
rect 600 682660 620 682730
rect 690 682660 710 682730
rect 780 682660 800 682730
rect 870 682660 890 682730
rect 960 682660 980 682730
rect 1050 682660 1070 682730
rect 1140 682660 1160 682730
rect 1230 682660 1250 682730
rect 1320 682660 1340 682730
rect 1410 682660 1430 682730
rect 1500 682660 1520 682730
rect 1590 682660 1610 682730
rect 1680 682660 14791 682730
rect 272 682640 14791 682660
rect 272 682570 350 682640
rect 420 682570 440 682640
rect 510 682570 530 682640
rect 600 682570 620 682640
rect 690 682570 710 682640
rect 780 682570 800 682640
rect 870 682570 890 682640
rect 960 682570 980 682640
rect 1050 682570 1070 682640
rect 1140 682570 1160 682640
rect 1230 682570 1250 682640
rect 1320 682570 1340 682640
rect 1410 682570 1430 682640
rect 1500 682570 1520 682640
rect 1590 682570 1610 682640
rect 1680 682570 14791 682640
rect 272 682550 14791 682570
rect 272 682480 350 682550
rect 420 682480 440 682550
rect 510 682480 530 682550
rect 600 682480 620 682550
rect 690 682480 710 682550
rect 780 682480 800 682550
rect 870 682480 890 682550
rect 960 682480 980 682550
rect 1050 682480 1070 682550
rect 1140 682480 1160 682550
rect 1230 682480 1250 682550
rect 1320 682480 1340 682550
rect 1410 682480 1430 682550
rect 1500 682480 1520 682550
rect 1590 682480 1610 682550
rect 1680 682480 14791 682550
rect 272 682460 14791 682480
rect 272 682390 350 682460
rect 420 682390 440 682460
rect 510 682390 530 682460
rect 600 682390 620 682460
rect 690 682390 710 682460
rect 780 682390 800 682460
rect 870 682390 890 682460
rect 960 682390 980 682460
rect 1050 682390 1070 682460
rect 1140 682390 1160 682460
rect 1230 682390 1250 682460
rect 1320 682390 1340 682460
rect 1410 682390 1430 682460
rect 1500 682390 1520 682460
rect 1590 682390 1610 682460
rect 1680 682390 14791 682460
rect 272 682370 14791 682390
rect 272 682300 350 682370
rect 420 682300 440 682370
rect 510 682300 530 682370
rect 600 682300 620 682370
rect 690 682300 710 682370
rect 780 682300 800 682370
rect 870 682300 890 682370
rect 960 682300 980 682370
rect 1050 682300 1070 682370
rect 1140 682300 1160 682370
rect 1230 682300 1250 682370
rect 1320 682300 1340 682370
rect 1410 682300 1430 682370
rect 1500 682300 1520 682370
rect 1590 682300 1610 682370
rect 1680 682300 14791 682370
rect 272 682280 14791 682300
rect 272 682210 350 682280
rect 420 682210 440 682280
rect 510 682210 530 682280
rect 600 682210 620 682280
rect 690 682210 710 682280
rect 780 682210 800 682280
rect 870 682210 890 682280
rect 960 682210 980 682280
rect 1050 682210 1070 682280
rect 1140 682210 1160 682280
rect 1230 682210 1250 682280
rect 1320 682210 1340 682280
rect 1410 682210 1430 682280
rect 1500 682210 1520 682280
rect 1590 682210 1610 682280
rect 1680 682210 14791 682280
rect 272 682190 14791 682210
rect 272 682120 350 682190
rect 420 682120 440 682190
rect 510 682120 530 682190
rect 600 682120 620 682190
rect 690 682120 710 682190
rect 780 682120 800 682190
rect 870 682120 890 682190
rect 960 682120 980 682190
rect 1050 682120 1070 682190
rect 1140 682120 1160 682190
rect 1230 682120 1250 682190
rect 1320 682120 1340 682190
rect 1410 682120 1430 682190
rect 1500 682120 1520 682190
rect 1590 682120 1610 682190
rect 1680 682120 14791 682190
rect 272 682100 14791 682120
rect 272 682030 350 682100
rect 420 682030 440 682100
rect 510 682030 530 682100
rect 600 682030 620 682100
rect 690 682030 710 682100
rect 780 682030 800 682100
rect 870 682030 890 682100
rect 960 682030 980 682100
rect 1050 682030 1070 682100
rect 1140 682030 1160 682100
rect 1230 682030 1250 682100
rect 1320 682030 1340 682100
rect 1410 682030 1430 682100
rect 1500 682030 1520 682100
rect 1590 682030 1610 682100
rect 1680 682030 14791 682100
rect 272 682010 14791 682030
rect 272 681940 350 682010
rect 420 681940 440 682010
rect 510 681940 530 682010
rect 600 681940 620 682010
rect 690 681940 710 682010
rect 780 681940 800 682010
rect 870 681940 890 682010
rect 960 681940 980 682010
rect 1050 681940 1070 682010
rect 1140 681940 1160 682010
rect 1230 681940 1250 682010
rect 1320 681940 1340 682010
rect 1410 681940 1430 682010
rect 1500 681940 1520 682010
rect 1590 681940 1610 682010
rect 1680 681940 14791 682010
rect 272 681920 14791 681940
rect 272 681850 350 681920
rect 420 681850 440 681920
rect 510 681850 530 681920
rect 600 681850 620 681920
rect 690 681850 710 681920
rect 780 681850 800 681920
rect 870 681850 890 681920
rect 960 681850 980 681920
rect 1050 681850 1070 681920
rect 1140 681850 1160 681920
rect 1230 681850 1250 681920
rect 1320 681850 1340 681920
rect 1410 681850 1430 681920
rect 1500 681850 1520 681920
rect 1590 681850 1610 681920
rect 1680 681850 14791 681920
rect 272 681830 14791 681850
rect 272 681760 350 681830
rect 420 681760 440 681830
rect 510 681760 530 681830
rect 600 681760 620 681830
rect 690 681760 710 681830
rect 780 681760 800 681830
rect 870 681760 890 681830
rect 960 681760 980 681830
rect 1050 681760 1070 681830
rect 1140 681760 1160 681830
rect 1230 681760 1250 681830
rect 1320 681760 1340 681830
rect 1410 681760 1430 681830
rect 1500 681760 1520 681830
rect 1590 681760 1610 681830
rect 1680 681760 14791 681830
rect 272 681740 14791 681760
rect 272 681670 350 681740
rect 420 681670 440 681740
rect 510 681670 530 681740
rect 600 681670 620 681740
rect 690 681670 710 681740
rect 780 681670 800 681740
rect 870 681670 890 681740
rect 960 681670 980 681740
rect 1050 681670 1070 681740
rect 1140 681670 1160 681740
rect 1230 681670 1250 681740
rect 1320 681670 1340 681740
rect 1410 681670 1430 681740
rect 1500 681670 1520 681740
rect 1590 681670 1610 681740
rect 1680 681670 14791 681740
rect 272 681653 14791 681670
rect 12791 643412 14791 681653
rect 17246 646861 19246 702320
rect 68194 703500 68352 703800
rect 68652 703500 68852 703800
rect 69152 703500 69352 703800
rect 69652 703500 69852 703800
rect 70152 703500 70352 703800
rect 70652 703500 70852 703800
rect 71152 703500 71352 703800
rect 71652 703500 71852 703800
rect 72152 703500 72352 703800
rect 72652 703500 72852 703800
rect 73152 703500 73194 703800
rect 68194 703300 73194 703500
rect 68194 703000 68352 703300
rect 68652 703000 68852 703300
rect 69152 703000 69352 703300
rect 69652 703000 69852 703300
rect 70152 703000 70352 703300
rect 70652 703000 70852 703300
rect 71152 703000 71352 703300
rect 71652 703000 71852 703300
rect 72152 703000 72352 703300
rect 72652 703000 72852 703300
rect 73152 703000 73194 703300
rect 68194 702800 73194 703000
rect 68194 702500 68352 702800
rect 68652 702500 68852 702800
rect 69152 702500 69352 702800
rect 69652 702500 69852 702800
rect 70152 702500 70352 702800
rect 70652 702500 70852 702800
rect 71152 702500 71352 702800
rect 71652 702500 71852 702800
rect 72152 702500 72352 702800
rect 72652 702500 72852 702800
rect 73152 702500 73194 702800
rect 68194 701060 73194 702500
rect 120194 703800 125194 704000
rect 120194 703500 120352 703800
rect 120652 703500 120852 703800
rect 121152 703500 121352 703800
rect 121652 703500 121852 703800
rect 122152 703500 122352 703800
rect 122652 703500 122852 703800
rect 123152 703500 123352 703800
rect 123652 703500 123852 703800
rect 124152 703500 124352 703800
rect 124652 703500 124852 703800
rect 125152 703500 125194 703800
rect 120194 703300 125194 703500
rect 120194 703000 120352 703300
rect 120652 703000 120852 703300
rect 121152 703000 121352 703300
rect 121652 703000 121852 703300
rect 122152 703000 122352 703300
rect 122652 703000 122852 703300
rect 123152 703000 123352 703300
rect 123652 703000 123852 703300
rect 124152 703000 124352 703300
rect 124652 703000 124852 703300
rect 125152 703000 125194 703300
rect 120194 702800 125194 703000
rect 120194 702500 120352 702800
rect 120652 702500 120852 702800
rect 121152 702500 121352 702800
rect 121652 702500 121852 702800
rect 122152 702500 122352 702800
rect 122652 702500 122852 702800
rect 123152 702500 123352 702800
rect 123652 702500 123852 702800
rect 124152 702500 124352 702800
rect 124652 702500 124852 702800
rect 125152 702500 125194 702800
rect 120194 701060 125194 702500
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 699884 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 415740 703110 416220 703170
rect 415740 703040 415760 703110
rect 415830 703040 415850 703110
rect 415920 703040 415940 703110
rect 416010 703040 416030 703110
rect 416100 703040 416120 703110
rect 416190 703040 416220 703110
rect 415740 703020 416220 703040
rect 415740 702950 415760 703020
rect 415830 702950 415850 703020
rect 415920 702950 415940 703020
rect 416010 702950 416030 703020
rect 416100 702950 416120 703020
rect 416190 702950 416220 703020
rect 415740 702930 416220 702950
rect 415740 702860 415760 702930
rect 415830 702860 415850 702930
rect 415920 702860 415940 702930
rect 416010 702860 416030 702930
rect 416100 702860 416120 702930
rect 416190 702860 416220 702930
rect 415740 702840 416220 702860
rect 415740 702770 415760 702840
rect 415830 702770 415850 702840
rect 415920 702770 415940 702840
rect 416010 702770 416030 702840
rect 416100 702770 416120 702840
rect 416190 702770 416220 702840
rect 415740 702750 416220 702770
rect 415740 702680 415760 702750
rect 415830 702680 415850 702750
rect 415920 702680 415940 702750
rect 416010 702680 416030 702750
rect 416100 702680 416120 702750
rect 416190 702680 416220 702750
rect 227594 699624 227767 699884
rect 228007 699624 228107 699884
rect 228347 699624 228447 699884
rect 228687 699624 228787 699884
rect 229027 699624 229127 699884
rect 229367 699624 229467 699884
rect 229707 699624 229807 699884
rect 230047 699624 230147 699884
rect 230387 699624 230487 699884
rect 230727 699624 230827 699884
rect 231067 699624 231167 699884
rect 231407 699624 231507 699884
rect 231747 699624 231847 699884
rect 232087 699624 232187 699884
rect 232427 699624 232594 699884
rect 227594 699524 232594 699624
rect 227594 699264 227767 699524
rect 228007 699264 228107 699524
rect 228347 699264 228447 699524
rect 228687 699264 228787 699524
rect 229027 699264 229127 699524
rect 229367 699264 229467 699524
rect 229707 699264 229807 699524
rect 230047 699264 230147 699524
rect 230387 699264 230487 699524
rect 230727 699264 230827 699524
rect 231067 699264 231167 699524
rect 231407 699264 231507 699524
rect 231747 699264 231847 699524
rect 232087 699264 232187 699524
rect 232427 699264 232594 699524
rect 227594 699164 232594 699264
rect 227594 698904 227767 699164
rect 228007 698904 228107 699164
rect 228347 698904 228447 699164
rect 228687 698904 228787 699164
rect 229027 698904 229127 699164
rect 229367 698904 229467 699164
rect 229707 698904 229807 699164
rect 230047 698904 230147 699164
rect 230387 698904 230487 699164
rect 230727 698904 230827 699164
rect 231067 698904 231167 699164
rect 231407 698904 231507 699164
rect 231747 698904 231847 699164
rect 232087 698904 232187 699164
rect 232427 698904 232594 699164
rect 227594 698804 232594 698904
rect 227594 698544 227767 698804
rect 228007 698544 228107 698804
rect 228347 698544 228447 698804
rect 228687 698544 228787 698804
rect 229027 698544 229127 698804
rect 229367 698544 229467 698804
rect 229707 698544 229807 698804
rect 230047 698544 230147 698804
rect 230387 698544 230487 698804
rect 230727 698544 230827 698804
rect 231067 698544 231167 698804
rect 231407 698544 231507 698804
rect 231747 698544 231847 698804
rect 232087 698544 232187 698804
rect 232427 698544 232594 698804
rect 131494 697420 225198 697448
rect 131494 697350 224744 697420
rect 224814 697350 224834 697420
rect 224904 697350 224924 697420
rect 224994 697350 225014 697420
rect 225084 697350 225104 697420
rect 225174 697350 225198 697420
rect 131494 697330 225198 697350
rect 131494 697260 224744 697330
rect 224814 697260 224834 697330
rect 224904 697260 224924 697330
rect 224994 697260 225014 697330
rect 225084 697260 225104 697330
rect 225174 697260 225198 697330
rect 131494 697240 225198 697260
rect 131494 697170 224744 697240
rect 224814 697170 224834 697240
rect 224904 697170 224924 697240
rect 224994 697170 225014 697240
rect 225084 697170 225104 697240
rect 225174 697170 225198 697240
rect 131494 697150 225198 697170
rect 131494 697080 224744 697150
rect 224814 697080 224834 697150
rect 224904 697080 224924 697150
rect 224994 697080 225014 697150
rect 225084 697080 225104 697150
rect 225174 697080 225198 697150
rect 131494 697060 225198 697080
rect 131494 696990 224744 697060
rect 224814 696990 224834 697060
rect 224904 696990 224924 697060
rect 224994 696990 225014 697060
rect 225084 696990 225104 697060
rect 225174 696990 225198 697060
rect 131494 696968 225198 696990
rect 131494 684650 131974 696968
rect 110364 684170 131974 684650
rect 132937 696203 225198 696231
rect 132937 696133 224744 696203
rect 224814 696133 224834 696203
rect 224904 696133 224924 696203
rect 224994 696133 225014 696203
rect 225084 696133 225104 696203
rect 225174 696133 225198 696203
rect 132937 696113 225198 696133
rect 132937 696043 224744 696113
rect 224814 696043 224834 696113
rect 224904 696043 224924 696113
rect 224994 696043 225014 696113
rect 225084 696043 225104 696113
rect 225174 696043 225198 696113
rect 132937 696023 225198 696043
rect 132937 695953 224744 696023
rect 224814 695953 224834 696023
rect 224904 695953 224924 696023
rect 224994 695953 225014 696023
rect 225084 695953 225104 696023
rect 225174 695953 225198 696023
rect 132937 695933 225198 695953
rect 132937 695863 224744 695933
rect 224814 695863 224834 695933
rect 224904 695863 224924 695933
rect 224994 695863 225014 695933
rect 225084 695863 225104 695933
rect 225174 695863 225198 695933
rect 132937 695843 225198 695863
rect 132937 695773 224744 695843
rect 224814 695773 224834 695843
rect 224904 695773 224924 695843
rect 224994 695773 225014 695843
rect 225084 695773 225104 695843
rect 225174 695773 225198 695843
rect 132937 695754 225198 695773
rect 110364 683130 110524 684170
rect 132937 682940 133414 695754
rect 224234 695751 225198 695754
rect 128410 682460 133414 682940
rect 134191 695138 225198 695166
rect 134191 695068 224744 695138
rect 224814 695068 224834 695138
rect 224904 695068 224924 695138
rect 224994 695068 225014 695138
rect 225084 695068 225104 695138
rect 225174 695068 225198 695138
rect 134191 695048 225198 695068
rect 134191 694978 224744 695048
rect 224814 694978 224834 695048
rect 224904 694978 224924 695048
rect 224994 694978 225014 695048
rect 225084 694978 225104 695048
rect 225174 694978 225198 695048
rect 134191 694958 225198 694978
rect 134191 694888 224744 694958
rect 224814 694888 224834 694958
rect 224904 694888 224924 694958
rect 224994 694888 225014 694958
rect 225084 694888 225104 694958
rect 225174 694888 225198 694958
rect 134191 694868 225198 694888
rect 134191 694798 224744 694868
rect 224814 694798 224834 694868
rect 224904 694798 224924 694868
rect 224994 694798 225014 694868
rect 225084 694798 225104 694868
rect 225174 694798 225198 694868
rect 134191 694778 225198 694798
rect 134191 694708 224744 694778
rect 224814 694708 224834 694778
rect 224904 694708 224924 694778
rect 224994 694708 225014 694778
rect 225084 694708 225104 694778
rect 225174 694708 225198 694778
rect 134191 694686 225198 694708
rect 134191 663940 134671 694686
rect 120014 663620 134671 663940
rect 135741 693432 225198 693460
rect 135741 693362 224744 693432
rect 224814 693362 224834 693432
rect 224904 693362 224924 693432
rect 224994 693362 225014 693432
rect 225084 693362 225104 693432
rect 225174 693362 225198 693432
rect 135741 693342 225198 693362
rect 135741 693272 224744 693342
rect 224814 693272 224834 693342
rect 224904 693272 224924 693342
rect 224994 693272 225014 693342
rect 225084 693272 225104 693342
rect 225174 693272 225198 693342
rect 135741 693252 225198 693272
rect 135741 693182 224744 693252
rect 224814 693182 224834 693252
rect 224904 693182 224924 693252
rect 224994 693182 225014 693252
rect 225084 693182 225104 693252
rect 225174 693182 225198 693252
rect 135741 693162 225198 693182
rect 135741 693092 224744 693162
rect 224814 693092 224834 693162
rect 224904 693092 224924 693162
rect 224994 693092 225014 693162
rect 225084 693092 225104 693162
rect 225174 693092 225198 693162
rect 135741 693072 225198 693092
rect 135741 693002 224744 693072
rect 224814 693002 224834 693072
rect 224904 693002 224924 693072
rect 224994 693002 225014 693072
rect 225084 693002 225104 693072
rect 225174 693002 225198 693072
rect 135741 692980 225198 693002
rect 135741 692969 224718 692980
rect 135741 658080 136232 692969
rect 227594 692568 232594 698544
rect 321017 697448 321497 702300
rect 234606 697420 321497 697448
rect 234606 697350 234630 697420
rect 234700 697350 234720 697420
rect 234790 697350 234810 697420
rect 234880 697350 234900 697420
rect 234970 697350 234990 697420
rect 235060 697350 321497 697420
rect 234606 697330 321497 697350
rect 234606 697260 234630 697330
rect 234700 697260 234720 697330
rect 234790 697260 234810 697330
rect 234880 697260 234900 697330
rect 234970 697260 234990 697330
rect 235060 697260 321497 697330
rect 234606 697240 321497 697260
rect 234606 697170 234630 697240
rect 234700 697170 234720 697240
rect 234790 697170 234810 697240
rect 234880 697170 234900 697240
rect 234970 697170 234990 697240
rect 235060 697170 321497 697240
rect 234606 697150 321497 697170
rect 234606 697080 234630 697150
rect 234700 697080 234720 697150
rect 234790 697080 234810 697150
rect 234880 697080 234900 697150
rect 234970 697080 234990 697150
rect 235060 697080 321497 697150
rect 234606 697060 321497 697080
rect 234606 696990 234630 697060
rect 234700 696990 234720 697060
rect 234790 696990 234810 697060
rect 234880 696990 234900 697060
rect 234970 696990 234990 697060
rect 235060 696990 321497 697060
rect 234606 696968 321497 696990
rect 415740 696231 416220 702680
rect 234606 696203 416220 696231
rect 234606 696133 234630 696203
rect 234700 696133 234720 696203
rect 234790 696133 234810 696203
rect 234880 696133 234900 696203
rect 234970 696133 234990 696203
rect 235060 696133 416220 696203
rect 234606 696113 416220 696133
rect 234606 696043 234630 696113
rect 234700 696043 234720 696113
rect 234790 696043 234810 696113
rect 234880 696043 234900 696113
rect 234970 696043 234990 696113
rect 235060 696043 416220 696113
rect 234606 696023 416220 696043
rect 234606 695953 234630 696023
rect 234700 695953 234720 696023
rect 234790 695953 234810 696023
rect 234880 695953 234900 696023
rect 234970 695953 234990 696023
rect 235060 695953 416220 696023
rect 234606 695933 416220 695953
rect 234606 695863 234630 695933
rect 234700 695863 234720 695933
rect 234790 695863 234810 695933
rect 234880 695863 234900 695933
rect 234970 695863 234990 695933
rect 235060 695863 416220 695933
rect 234606 695843 416220 695863
rect 234606 695773 234630 695843
rect 234700 695773 234720 695843
rect 234790 695773 234810 695843
rect 234880 695773 234900 695843
rect 234970 695773 234990 695843
rect 235060 695773 416220 695843
rect 234606 695754 416220 695773
rect 234606 695751 235570 695754
rect 415740 695752 416220 695754
rect 466990 703110 467470 703170
rect 466990 703040 467010 703110
rect 467080 703040 467100 703110
rect 467170 703040 467190 703110
rect 467260 703040 467280 703110
rect 467350 703040 467370 703110
rect 467440 703040 467470 703110
rect 466990 703020 467470 703040
rect 466990 702950 467010 703020
rect 467080 702950 467100 703020
rect 467170 702950 467190 703020
rect 467260 702950 467280 703020
rect 467350 702950 467370 703020
rect 467440 702950 467470 703020
rect 466990 702930 467470 702950
rect 466990 702860 467010 702930
rect 467080 702860 467100 702930
rect 467170 702860 467190 702930
rect 467260 702860 467280 702930
rect 467350 702860 467370 702930
rect 467440 702860 467470 702930
rect 466990 702840 467470 702860
rect 466990 702770 467010 702840
rect 467080 702770 467100 702840
rect 467170 702770 467190 702840
rect 467260 702770 467280 702840
rect 467350 702770 467370 702840
rect 467440 702770 467470 702840
rect 466990 702750 467470 702770
rect 466990 702680 467010 702750
rect 467080 702680 467100 702750
rect 467170 702680 467190 702750
rect 467260 702680 467280 702750
rect 467350 702680 467370 702750
rect 467440 702680 467470 702750
rect 466990 695166 467470 702680
rect 569120 703110 569600 703170
rect 569120 703040 569140 703110
rect 569210 703040 569230 703110
rect 569300 703040 569320 703110
rect 569390 703040 569410 703110
rect 569480 703040 569500 703110
rect 569570 703040 569600 703110
rect 569120 703020 569600 703040
rect 569120 702950 569140 703020
rect 569210 702950 569230 703020
rect 569300 702950 569320 703020
rect 569390 702950 569410 703020
rect 569480 702950 569500 703020
rect 569570 702950 569600 703020
rect 569120 702930 569600 702950
rect 569120 702860 569140 702930
rect 569210 702860 569230 702930
rect 569300 702860 569320 702930
rect 569390 702860 569410 702930
rect 569480 702860 569500 702930
rect 569570 702860 569600 702930
rect 569120 702840 569600 702860
rect 569120 702770 569140 702840
rect 569210 702770 569230 702840
rect 569300 702770 569320 702840
rect 569390 702770 569410 702840
rect 569480 702770 569500 702840
rect 569570 702770 569600 702840
rect 569120 702750 569600 702770
rect 569120 702680 569140 702750
rect 569210 702680 569230 702750
rect 569300 702680 569320 702750
rect 569390 702680 569410 702750
rect 569480 702680 569500 702750
rect 569570 702680 569600 702750
rect 569120 697324 569600 702680
rect 234606 695138 467470 695166
rect 234606 695068 234630 695138
rect 234700 695068 234720 695138
rect 234790 695068 234810 695138
rect 234880 695068 234900 695138
rect 234970 695068 234990 695138
rect 235060 695068 467470 695138
rect 234606 695048 467470 695068
rect 234606 694978 234630 695048
rect 234700 694978 234720 695048
rect 234790 694978 234810 695048
rect 234880 694978 234900 695048
rect 234970 694978 234990 695048
rect 235060 694978 467470 695048
rect 234606 694958 467470 694978
rect 234606 694888 234630 694958
rect 234700 694888 234720 694958
rect 234790 694888 234810 694958
rect 234880 694888 234900 694958
rect 234970 694888 234990 694958
rect 235060 694888 467470 694958
rect 234606 694868 467470 694888
rect 234606 694798 234630 694868
rect 234700 694798 234720 694868
rect 234790 694798 234810 694868
rect 234880 694798 234900 694868
rect 234970 694798 234990 694868
rect 235060 694798 467470 694868
rect 234606 694778 467470 694798
rect 234606 694708 234630 694778
rect 234700 694708 234720 694778
rect 234790 694708 234810 694778
rect 234880 694708 234900 694778
rect 234970 694708 234990 694778
rect 235060 694708 467470 694778
rect 234606 694686 467470 694708
rect 569115 693460 569606 697324
rect 234606 693432 569606 693460
rect 234606 693362 234630 693432
rect 234700 693362 234720 693432
rect 234790 693362 234810 693432
rect 234880 693362 234900 693432
rect 234970 693362 234990 693432
rect 235060 693362 569606 693432
rect 234606 693342 569606 693362
rect 234606 693272 234630 693342
rect 234700 693272 234720 693342
rect 234790 693272 234810 693342
rect 234880 693272 234900 693342
rect 234970 693272 234990 693342
rect 235060 693272 569606 693342
rect 234606 693252 569606 693272
rect 234606 693182 234630 693252
rect 234700 693182 234720 693252
rect 234790 693182 234810 693252
rect 234880 693182 234900 693252
rect 234970 693182 234990 693252
rect 235060 693182 569606 693252
rect 234606 693162 569606 693182
rect 234606 693092 234630 693162
rect 234700 693092 234720 693162
rect 234790 693092 234810 693162
rect 234880 693092 234900 693162
rect 234970 693092 234990 693162
rect 235060 693092 569606 693162
rect 234606 693072 569606 693092
rect 234606 693002 234630 693072
rect 234700 693002 234720 693072
rect 234790 693002 234810 693072
rect 234880 693002 234900 693072
rect 234970 693002 234990 693072
rect 235060 693002 569606 693072
rect 234606 692980 569606 693002
rect 235086 692969 569606 692980
rect 119854 657760 136232 658080
rect 137524 691718 225198 691746
rect 137524 691648 224744 691718
rect 224814 691648 224834 691718
rect 224904 691648 224924 691718
rect 224994 691648 225014 691718
rect 225084 691648 225104 691718
rect 225174 691648 225198 691718
rect 137524 691628 225198 691648
rect 137524 691580 224744 691628
rect 137524 691510 165360 691580
rect 165430 691510 165460 691580
rect 165530 691510 165560 691580
rect 165630 691510 165660 691580
rect 165730 691510 165760 691580
rect 165830 691510 165860 691580
rect 165930 691510 165960 691580
rect 166030 691510 166060 691580
rect 166130 691510 166160 691580
rect 166230 691510 166260 691580
rect 166330 691510 166360 691580
rect 166430 691510 166460 691580
rect 166530 691510 166560 691580
rect 166630 691510 166660 691580
rect 166730 691510 166760 691580
rect 166830 691510 166860 691580
rect 166930 691510 166960 691580
rect 167030 691510 167060 691580
rect 167130 691510 167160 691580
rect 167230 691510 167260 691580
rect 167330 691510 167360 691580
rect 167430 691510 167460 691580
rect 167530 691510 167560 691580
rect 167630 691510 167660 691580
rect 167730 691510 167760 691580
rect 167830 691510 167860 691580
rect 167930 691510 167960 691580
rect 168030 691510 168060 691580
rect 168130 691510 168160 691580
rect 168230 691510 168260 691580
rect 168330 691510 168360 691580
rect 168430 691510 168460 691580
rect 168530 691510 168560 691580
rect 168630 691510 168660 691580
rect 168730 691510 168760 691580
rect 168830 691510 168860 691580
rect 168930 691510 168960 691580
rect 169030 691510 169060 691580
rect 169130 691510 169160 691580
rect 169230 691510 169260 691580
rect 169330 691510 169360 691580
rect 169430 691510 169460 691580
rect 169530 691510 169560 691580
rect 169630 691510 169660 691580
rect 169730 691510 169760 691580
rect 169830 691510 169860 691580
rect 169930 691510 169960 691580
rect 170030 691510 170060 691580
rect 170130 691510 170160 691580
rect 170230 691510 170260 691580
rect 170330 691510 170360 691580
rect 170430 691510 170460 691580
rect 170530 691558 224744 691580
rect 224814 691558 224834 691628
rect 224904 691558 224924 691628
rect 224994 691558 225014 691628
rect 225084 691558 225104 691628
rect 225174 691558 225198 691628
rect 170530 691538 225198 691558
rect 170530 691510 224744 691538
rect 137524 691470 224744 691510
rect 137524 691400 165360 691470
rect 165430 691400 165460 691470
rect 165530 691400 165560 691470
rect 165630 691400 165660 691470
rect 165730 691400 165760 691470
rect 165830 691400 165860 691470
rect 165930 691400 165960 691470
rect 166030 691400 166060 691470
rect 166130 691400 166160 691470
rect 166230 691400 166260 691470
rect 166330 691400 166360 691470
rect 166430 691400 166460 691470
rect 166530 691400 166560 691470
rect 166630 691400 166660 691470
rect 166730 691400 166760 691470
rect 166830 691400 166860 691470
rect 166930 691400 166960 691470
rect 167030 691400 167060 691470
rect 167130 691400 167160 691470
rect 167230 691400 167260 691470
rect 167330 691400 167360 691470
rect 167430 691400 167460 691470
rect 167530 691400 167560 691470
rect 167630 691400 167660 691470
rect 167730 691400 167760 691470
rect 167830 691400 167860 691470
rect 167930 691400 167960 691470
rect 168030 691400 168060 691470
rect 168130 691400 168160 691470
rect 168230 691400 168260 691470
rect 168330 691400 168360 691470
rect 168430 691400 168460 691470
rect 168530 691400 168560 691470
rect 168630 691400 168660 691470
rect 168730 691400 168760 691470
rect 168830 691400 168860 691470
rect 168930 691400 168960 691470
rect 169030 691400 169060 691470
rect 169130 691400 169160 691470
rect 169230 691400 169260 691470
rect 169330 691400 169360 691470
rect 169430 691400 169460 691470
rect 169530 691400 169560 691470
rect 169630 691400 169660 691470
rect 169730 691400 169760 691470
rect 169830 691400 169860 691470
rect 169930 691400 169960 691470
rect 170030 691400 170060 691470
rect 170130 691400 170160 691470
rect 170230 691400 170260 691470
rect 170330 691400 170360 691470
rect 170430 691400 170460 691470
rect 170530 691468 224744 691470
rect 224814 691468 224834 691538
rect 224904 691468 224924 691538
rect 224994 691468 225014 691538
rect 225084 691468 225104 691538
rect 225174 691468 225198 691538
rect 170530 691448 225198 691468
rect 170530 691400 224744 691448
rect 137524 691378 224744 691400
rect 224814 691378 224834 691448
rect 224904 691378 224924 691448
rect 224994 691378 225014 691448
rect 225084 691378 225104 691448
rect 225174 691378 225198 691448
rect 137524 691358 225198 691378
rect 137524 691288 224744 691358
rect 224814 691288 224834 691358
rect 224904 691288 224924 691358
rect 224994 691288 225014 691358
rect 225084 691288 225104 691358
rect 225174 691288 225198 691358
rect 137524 691266 225198 691288
rect 137524 652221 138004 691266
rect 165364 690140 170800 690160
rect 165364 689900 165620 690140
rect 165860 690070 165950 690140
rect 166190 690070 166280 690140
rect 166520 690070 166610 690140
rect 166850 690070 166940 690140
rect 167180 690070 167270 690140
rect 167510 690070 167600 690140
rect 167840 690070 167930 690140
rect 168170 690070 168260 690140
rect 168500 690070 168590 690140
rect 168830 690070 168920 690140
rect 169160 690070 169250 690140
rect 169490 690070 169580 690140
rect 169820 690070 169910 690140
rect 170150 690070 170240 690140
rect 170480 690070 170800 690140
rect 165890 690000 165920 690070
rect 166190 690000 166220 690070
rect 166590 690000 166610 690070
rect 166890 690000 166920 690070
rect 167190 690000 167220 690070
rect 167510 690000 167520 690070
rect 167590 690000 167600 690070
rect 167890 690000 167920 690070
rect 168190 690000 168220 690070
rect 168500 690000 168520 690070
rect 168890 690000 168920 690070
rect 169190 690000 169220 690070
rect 169490 690000 169520 690070
rect 169890 690000 169910 690070
rect 170190 690000 170220 690070
rect 170490 690000 170800 690070
rect 165860 689970 165950 690000
rect 166190 689970 166280 690000
rect 166520 689970 166610 690000
rect 166850 689970 166940 690000
rect 167180 689970 167270 690000
rect 167510 689970 167600 690000
rect 167840 689970 167930 690000
rect 168170 689970 168260 690000
rect 168500 689970 168590 690000
rect 168830 689970 168920 690000
rect 169160 689970 169250 690000
rect 169490 689970 169580 690000
rect 169820 689970 169910 690000
rect 170150 689970 170240 690000
rect 170480 689970 170800 690000
rect 165890 689900 165920 689970
rect 166190 689900 166220 689970
rect 166590 689900 166610 689970
rect 166890 689900 166920 689970
rect 167190 689900 167220 689970
rect 167510 689900 167520 689970
rect 167590 689900 167600 689970
rect 167890 689900 167920 689970
rect 168190 689900 168220 689970
rect 168500 689900 168520 689970
rect 168890 689900 168920 689970
rect 169190 689900 169220 689970
rect 169490 689900 169520 689970
rect 169890 689900 169910 689970
rect 170190 689900 170220 689970
rect 170490 689900 170800 689970
rect 165364 689877 170800 689900
rect 227606 690060 232583 692568
rect 234606 691718 581422 691746
rect 234606 691648 234630 691718
rect 234700 691648 234720 691718
rect 234790 691648 234810 691718
rect 234880 691648 234900 691718
rect 234970 691648 234990 691718
rect 235060 691648 581422 691718
rect 234606 691628 581422 691648
rect 234606 691558 234630 691628
rect 234700 691558 234720 691628
rect 234790 691558 234810 691628
rect 234880 691558 234900 691628
rect 234970 691558 234990 691628
rect 235060 691558 581422 691628
rect 234606 691538 581422 691558
rect 234606 691468 234630 691538
rect 234700 691468 234720 691538
rect 234790 691468 234810 691538
rect 234880 691468 234900 691538
rect 234970 691468 234990 691538
rect 235060 691468 581422 691538
rect 234606 691448 581422 691468
rect 234606 691378 234630 691448
rect 234700 691378 234720 691448
rect 234790 691378 234810 691448
rect 234880 691378 234900 691448
rect 234970 691378 234990 691448
rect 235060 691378 581422 691448
rect 234606 691358 581422 691378
rect 234606 691288 234630 691358
rect 234700 691288 234720 691358
rect 234790 691288 234810 691358
rect 234880 691288 234900 691358
rect 234970 691288 234990 691358
rect 235060 691288 581422 691358
rect 234606 691266 581422 691288
rect 227606 689990 227640 690060
rect 227710 689990 227740 690060
rect 227810 689990 227840 690060
rect 227910 689990 227940 690060
rect 228010 689990 228040 690060
rect 228110 689990 228140 690060
rect 228210 689990 228240 690060
rect 228310 689990 228340 690060
rect 228410 689990 228440 690060
rect 228510 689990 228540 690060
rect 228610 689990 228640 690060
rect 228710 689990 228740 690060
rect 228810 689990 228840 690060
rect 228910 689990 228940 690060
rect 229010 689990 229040 690060
rect 229110 689990 229140 690060
rect 229210 689990 229240 690060
rect 229310 689990 229340 690060
rect 229410 689990 229440 690060
rect 229510 689990 229540 690060
rect 229610 689990 229640 690060
rect 229710 689990 229740 690060
rect 229810 689990 229840 690060
rect 229910 689990 229940 690060
rect 230010 689990 230040 690060
rect 230110 689990 230140 690060
rect 230210 689990 230240 690060
rect 230310 689990 230340 690060
rect 230410 689990 230440 690060
rect 230510 689990 230540 690060
rect 230610 689990 230640 690060
rect 230710 689990 230740 690060
rect 230810 689990 230840 690060
rect 230910 689990 230940 690060
rect 231010 689990 231040 690060
rect 231110 689990 231140 690060
rect 231210 689990 231240 690060
rect 231310 689990 231340 690060
rect 231410 689990 231440 690060
rect 231510 689990 231540 690060
rect 231610 689990 231640 690060
rect 231710 689990 231740 690060
rect 231810 689990 231840 690060
rect 231910 689990 231940 690060
rect 232010 689990 232040 690060
rect 232110 689990 232140 690060
rect 232210 689990 232240 690060
rect 232310 689990 232340 690060
rect 232410 689990 232440 690060
rect 232510 689990 232583 690060
rect 227606 689960 232583 689990
rect 227606 689890 227640 689960
rect 227710 689890 227740 689960
rect 227810 689890 227840 689960
rect 227910 689890 227940 689960
rect 228010 689890 228040 689960
rect 228110 689890 228140 689960
rect 228210 689890 228240 689960
rect 228310 689890 228340 689960
rect 228410 689890 228440 689960
rect 228510 689890 228540 689960
rect 228610 689890 228640 689960
rect 228710 689890 228740 689960
rect 228810 689890 228840 689960
rect 228910 689890 228940 689960
rect 229010 689890 229040 689960
rect 229110 689890 229140 689960
rect 229210 689890 229240 689960
rect 229310 689890 229340 689960
rect 229410 689890 229440 689960
rect 229510 689890 229540 689960
rect 229610 689890 229640 689960
rect 229710 689890 229740 689960
rect 229810 689890 229840 689960
rect 229910 689890 229940 689960
rect 230010 689890 230040 689960
rect 230110 689890 230140 689960
rect 230210 689890 230240 689960
rect 230310 689890 230340 689960
rect 230410 689890 230440 689960
rect 230510 689890 230540 689960
rect 230610 689890 230640 689960
rect 230710 689890 230740 689960
rect 230810 689890 230840 689960
rect 230910 689890 230940 689960
rect 231010 689890 231040 689960
rect 231110 689890 231140 689960
rect 231210 689890 231240 689960
rect 231310 689890 231340 689960
rect 231410 689890 231440 689960
rect 231510 689890 231540 689960
rect 231610 689890 231640 689960
rect 231710 689890 231740 689960
rect 231810 689890 231840 689960
rect 231910 689890 231940 689960
rect 232010 689890 232040 689960
rect 232110 689890 232140 689960
rect 232210 689890 232240 689960
rect 232310 689890 232340 689960
rect 232410 689890 232440 689960
rect 232510 689890 232583 689960
rect 227606 680746 232583 689890
rect 119500 651900 138004 652221
rect 173787 675750 232583 680746
rect 580942 681130 581422 691266
rect 580942 681110 583170 681130
rect 580942 681040 582680 681110
rect 582750 681040 582770 681110
rect 582840 681040 582860 681110
rect 582930 681040 582950 681110
rect 583020 681040 583040 681110
rect 583110 681040 583170 681110
rect 580942 681020 583170 681040
rect 580942 680950 582680 681020
rect 582750 680950 582770 681020
rect 582840 680950 582860 681020
rect 582930 680950 582950 681020
rect 583020 680950 583040 681020
rect 583110 680950 583170 681020
rect 580942 680930 583170 680950
rect 580942 680860 582680 680930
rect 582750 680860 582770 680930
rect 582840 680860 582860 680930
rect 582930 680860 582950 680930
rect 583020 680860 583040 680930
rect 583110 680860 583170 680930
rect 580942 680840 583170 680860
rect 580942 680770 582680 680840
rect 582750 680770 582770 680840
rect 582840 680770 582860 680840
rect 582930 680770 582950 680840
rect 583020 680770 583040 680840
rect 583110 680770 583170 680840
rect 580942 680750 583170 680770
rect 580942 680680 582680 680750
rect 582750 680680 582770 680750
rect 582840 680680 582860 680750
rect 582930 680680 582950 680750
rect 583020 680680 583040 680750
rect 583110 680680 583170 680750
rect 580942 680650 583170 680680
rect 173787 668865 178784 675750
rect 180904 668865 227118 668866
rect 227584 668865 232583 675750
rect 173787 667118 232583 668865
rect 173787 663870 232580 667118
rect 173787 660277 178784 663870
rect 227584 660277 232580 663870
rect 173787 655280 232580 660277
rect 93369 650470 95369 650507
rect 93369 650400 94280 650470
rect 94350 650400 94380 650470
rect 94450 650400 94480 650470
rect 94550 650400 95369 650470
rect 93369 650380 95369 650400
rect 93369 650310 94280 650380
rect 94350 650310 94380 650380
rect 94450 650310 94480 650380
rect 94550 650310 95369 650380
rect 93369 646861 95369 650310
rect 17246 644861 95369 646861
rect 97956 650470 99956 650493
rect 97956 650400 98838 650470
rect 98908 650400 98938 650470
rect 99008 650400 99038 650470
rect 99108 650400 99956 650470
rect 97956 650380 99956 650400
rect 97956 650310 98838 650380
rect 98908 650310 98938 650380
rect 99008 650310 99038 650380
rect 99108 650310 99956 650380
rect 97956 643412 99956 650310
rect 12791 641412 99956 643412
rect 173787 642452 178784 655280
rect 227584 642452 232580 655280
rect 156762 642285 232580 642452
rect 156762 642045 157818 642285
rect 158078 642045 158178 642285
rect 158438 642045 158538 642285
rect 158798 642045 158898 642285
rect 159158 642045 232580 642285
rect 156762 641945 232580 642045
rect 156762 641705 157818 641945
rect 158078 641705 158178 641945
rect 158438 641705 158538 641945
rect 158798 641705 158898 641945
rect 159158 641705 232580 641945
rect 156762 641605 232580 641705
rect 156762 641365 157818 641605
rect 158078 641365 158178 641605
rect 158438 641365 158538 641605
rect 158798 641365 158898 641605
rect 159158 641365 232580 641605
rect 156762 641265 232580 641365
rect 156762 641025 157818 641265
rect 158078 641025 158178 641265
rect 158438 641025 158538 641265
rect 158798 641025 158898 641265
rect 159158 641025 232580 641265
rect 156762 640925 232580 641025
rect 156762 640685 157818 640925
rect 158078 640685 158178 640925
rect 158438 640685 158538 640925
rect 158798 640685 158898 640925
rect 159158 640685 232580 640925
rect 156762 640585 232580 640685
rect 156762 640345 157818 640585
rect 158078 640345 158178 640585
rect 158438 640345 158538 640585
rect 158798 640345 158898 640585
rect 159158 640345 232580 640585
rect 156762 640245 232580 640345
rect 156762 640005 157818 640245
rect 158078 640005 158178 640245
rect 158438 640005 158538 640245
rect 158798 640005 158898 640245
rect 159158 640005 232580 640245
rect 156762 639905 232580 640005
rect 156762 639665 157818 639905
rect 158078 639665 158178 639905
rect 158438 639665 158538 639905
rect 158798 639665 158898 639905
rect 159158 639665 232580 639905
rect 156762 639565 232580 639665
rect 156762 639325 157818 639565
rect 158078 639325 158178 639565
rect 158438 639325 158538 639565
rect 158798 639325 158898 639565
rect 159158 639325 232580 639565
rect 156762 639225 232580 639325
rect 156762 638985 157818 639225
rect 158078 638985 158178 639225
rect 158438 638985 158538 639225
rect 158798 638985 158898 639225
rect 159158 638985 232580 639225
rect 156762 638885 232580 638985
rect 156762 638645 157818 638885
rect 158078 638645 158178 638885
rect 158438 638645 158538 638885
rect 158798 638645 158898 638885
rect 159158 638645 232580 638885
rect 156762 638545 232580 638645
rect 156762 638305 157818 638545
rect 158078 638305 158178 638545
rect 158438 638305 158538 638545
rect 158798 638305 158898 638545
rect 159158 638305 232580 638545
rect 156762 638205 232580 638305
rect 156762 637965 157818 638205
rect 158078 637965 158178 638205
rect 158438 637965 158538 638205
rect 158798 637965 158898 638205
rect 159158 637965 232580 638205
rect 156762 637865 232580 637965
rect 156762 637625 157818 637865
rect 158078 637625 158178 637865
rect 158438 637625 158538 637865
rect 158798 637625 158898 637865
rect 159158 637625 232580 637865
rect 156762 637452 232580 637625
<< via4 >>
rect 68352 703500 68652 703800
rect 68852 703500 69152 703800
rect 69352 703500 69652 703800
rect 69852 703500 70152 703800
rect 70352 703500 70652 703800
rect 70852 703500 71152 703800
rect 71352 703500 71652 703800
rect 71852 703500 72152 703800
rect 72352 703500 72652 703800
rect 72852 703500 73152 703800
rect 68352 703000 68652 703300
rect 68852 703000 69152 703300
rect 69352 703000 69652 703300
rect 69852 703000 70152 703300
rect 70352 703000 70652 703300
rect 70852 703000 71152 703300
rect 71352 703000 71652 703300
rect 71852 703000 72152 703300
rect 72352 703000 72652 703300
rect 72852 703000 73152 703300
rect 68352 702500 68652 702800
rect 68852 702500 69152 702800
rect 69352 702500 69652 702800
rect 69852 702500 70152 702800
rect 70352 702500 70652 702800
rect 70852 702500 71152 702800
rect 71352 702500 71652 702800
rect 71852 702500 72152 702800
rect 72352 702500 72652 702800
rect 72852 702500 73152 702800
rect 120352 703500 120652 703800
rect 120852 703500 121152 703800
rect 121352 703500 121652 703800
rect 121852 703500 122152 703800
rect 122352 703500 122652 703800
rect 122852 703500 123152 703800
rect 123352 703500 123652 703800
rect 123852 703500 124152 703800
rect 124352 703500 124652 703800
rect 124852 703500 125152 703800
rect 120352 703000 120652 703300
rect 120852 703000 121152 703300
rect 121352 703000 121652 703300
rect 121852 703000 122152 703300
rect 122352 703000 122652 703300
rect 122852 703000 123152 703300
rect 123352 703000 123652 703300
rect 123852 703000 124152 703300
rect 124352 703000 124652 703300
rect 124852 703000 125152 703300
rect 120352 702500 120652 702800
rect 120852 702500 121152 702800
rect 121352 702500 121652 702800
rect 121852 702500 122152 702800
rect 122352 702500 122652 702800
rect 122852 702500 123152 702800
rect 123352 702500 123652 702800
rect 123852 702500 124152 702800
rect 124352 702500 124652 702800
rect 124852 702500 125152 702800
rect 227767 699624 228007 699884
rect 228107 699624 228347 699884
rect 228447 699624 228687 699884
rect 228787 699624 229027 699884
rect 229127 699624 229367 699884
rect 229467 699624 229707 699884
rect 229807 699624 230047 699884
rect 230147 699624 230387 699884
rect 230487 699624 230727 699884
rect 230827 699624 231067 699884
rect 231167 699624 231407 699884
rect 231507 699624 231747 699884
rect 231847 699624 232087 699884
rect 232187 699624 232427 699884
rect 227767 699264 228007 699524
rect 228107 699264 228347 699524
rect 228447 699264 228687 699524
rect 228787 699264 229027 699524
rect 229127 699264 229367 699524
rect 229467 699264 229707 699524
rect 229807 699264 230047 699524
rect 230147 699264 230387 699524
rect 230487 699264 230727 699524
rect 230827 699264 231067 699524
rect 231167 699264 231407 699524
rect 231507 699264 231747 699524
rect 231847 699264 232087 699524
rect 232187 699264 232427 699524
rect 227767 698904 228007 699164
rect 228107 698904 228347 699164
rect 228447 698904 228687 699164
rect 228787 698904 229027 699164
rect 229127 698904 229367 699164
rect 229467 698904 229707 699164
rect 229807 698904 230047 699164
rect 230147 698904 230387 699164
rect 230487 698904 230727 699164
rect 230827 698904 231067 699164
rect 231167 698904 231407 699164
rect 231507 698904 231747 699164
rect 231847 698904 232087 699164
rect 232187 698904 232427 699164
rect 227767 698544 228007 698804
rect 228107 698544 228347 698804
rect 228447 698544 228687 698804
rect 228787 698544 229027 698804
rect 229127 698544 229367 698804
rect 229467 698544 229707 698804
rect 229807 698544 230047 698804
rect 230147 698544 230387 698804
rect 230487 698544 230727 698804
rect 230827 698544 231067 698804
rect 231167 698544 231407 698804
rect 231507 698544 231747 698804
rect 231847 698544 232087 698804
rect 232187 698544 232427 698804
rect 165620 690070 165860 690140
rect 165950 690070 166190 690140
rect 166280 690070 166520 690140
rect 166610 690070 166850 690140
rect 166940 690070 167180 690140
rect 167270 690070 167510 690140
rect 167600 690070 167840 690140
rect 167930 690070 168170 690140
rect 168260 690070 168500 690140
rect 168590 690070 168830 690140
rect 168920 690070 169160 690140
rect 169250 690070 169490 690140
rect 169580 690070 169820 690140
rect 169910 690070 170150 690140
rect 170240 690070 170480 690140
rect 165620 690000 165690 690070
rect 165690 690000 165720 690070
rect 165720 690000 165790 690070
rect 165790 690000 165820 690070
rect 165820 690000 165860 690070
rect 165950 690000 165990 690070
rect 165990 690000 166020 690070
rect 166020 690000 166090 690070
rect 166090 690000 166120 690070
rect 166120 690000 166190 690070
rect 166280 690000 166290 690070
rect 166290 690000 166320 690070
rect 166320 690000 166390 690070
rect 166390 690000 166420 690070
rect 166420 690000 166490 690070
rect 166490 690000 166520 690070
rect 166610 690000 166620 690070
rect 166620 690000 166690 690070
rect 166690 690000 166720 690070
rect 166720 690000 166790 690070
rect 166790 690000 166820 690070
rect 166820 690000 166850 690070
rect 166940 690000 166990 690070
rect 166990 690000 167020 690070
rect 167020 690000 167090 690070
rect 167090 690000 167120 690070
rect 167120 690000 167180 690070
rect 167270 690000 167290 690070
rect 167290 690000 167320 690070
rect 167320 690000 167390 690070
rect 167390 690000 167420 690070
rect 167420 690000 167490 690070
rect 167490 690000 167510 690070
rect 167600 690000 167620 690070
rect 167620 690000 167690 690070
rect 167690 690000 167720 690070
rect 167720 690000 167790 690070
rect 167790 690000 167820 690070
rect 167820 690000 167840 690070
rect 167930 690000 167990 690070
rect 167990 690000 168020 690070
rect 168020 690000 168090 690070
rect 168090 690000 168120 690070
rect 168120 690000 168170 690070
rect 168260 690000 168290 690070
rect 168290 690000 168320 690070
rect 168320 690000 168390 690070
rect 168390 690000 168420 690070
rect 168420 690000 168490 690070
rect 168490 690000 168500 690070
rect 168590 690000 168620 690070
rect 168620 690000 168690 690070
rect 168690 690000 168720 690070
rect 168720 690000 168790 690070
rect 168790 690000 168820 690070
rect 168820 690000 168830 690070
rect 168920 690000 168990 690070
rect 168990 690000 169020 690070
rect 169020 690000 169090 690070
rect 169090 690000 169120 690070
rect 169120 690000 169160 690070
rect 169250 690000 169290 690070
rect 169290 690000 169320 690070
rect 169320 690000 169390 690070
rect 169390 690000 169420 690070
rect 169420 690000 169490 690070
rect 169580 690000 169590 690070
rect 169590 690000 169620 690070
rect 169620 690000 169690 690070
rect 169690 690000 169720 690070
rect 169720 690000 169790 690070
rect 169790 690000 169820 690070
rect 169910 690000 169920 690070
rect 169920 690000 169990 690070
rect 169990 690000 170020 690070
rect 170020 690000 170090 690070
rect 170090 690000 170120 690070
rect 170120 690000 170150 690070
rect 170240 690000 170290 690070
rect 170290 690000 170320 690070
rect 170320 690000 170390 690070
rect 170390 690000 170420 690070
rect 170420 690000 170480 690070
rect 165620 689970 165860 690000
rect 165950 689970 166190 690000
rect 166280 689970 166520 690000
rect 166610 689970 166850 690000
rect 166940 689970 167180 690000
rect 167270 689970 167510 690000
rect 167600 689970 167840 690000
rect 167930 689970 168170 690000
rect 168260 689970 168500 690000
rect 168590 689970 168830 690000
rect 168920 689970 169160 690000
rect 169250 689970 169490 690000
rect 169580 689970 169820 690000
rect 169910 689970 170150 690000
rect 170240 689970 170480 690000
rect 165620 689900 165690 689970
rect 165690 689900 165720 689970
rect 165720 689900 165790 689970
rect 165790 689900 165820 689970
rect 165820 689900 165860 689970
rect 165950 689900 165990 689970
rect 165990 689900 166020 689970
rect 166020 689900 166090 689970
rect 166090 689900 166120 689970
rect 166120 689900 166190 689970
rect 166280 689900 166290 689970
rect 166290 689900 166320 689970
rect 166320 689900 166390 689970
rect 166390 689900 166420 689970
rect 166420 689900 166490 689970
rect 166490 689900 166520 689970
rect 166610 689900 166620 689970
rect 166620 689900 166690 689970
rect 166690 689900 166720 689970
rect 166720 689900 166790 689970
rect 166790 689900 166820 689970
rect 166820 689900 166850 689970
rect 166940 689900 166990 689970
rect 166990 689900 167020 689970
rect 167020 689900 167090 689970
rect 167090 689900 167120 689970
rect 167120 689900 167180 689970
rect 167270 689900 167290 689970
rect 167290 689900 167320 689970
rect 167320 689900 167390 689970
rect 167390 689900 167420 689970
rect 167420 689900 167490 689970
rect 167490 689900 167510 689970
rect 167600 689900 167620 689970
rect 167620 689900 167690 689970
rect 167690 689900 167720 689970
rect 167720 689900 167790 689970
rect 167790 689900 167820 689970
rect 167820 689900 167840 689970
rect 167930 689900 167990 689970
rect 167990 689900 168020 689970
rect 168020 689900 168090 689970
rect 168090 689900 168120 689970
rect 168120 689900 168170 689970
rect 168260 689900 168290 689970
rect 168290 689900 168320 689970
rect 168320 689900 168390 689970
rect 168390 689900 168420 689970
rect 168420 689900 168490 689970
rect 168490 689900 168500 689970
rect 168590 689900 168620 689970
rect 168620 689900 168690 689970
rect 168690 689900 168720 689970
rect 168720 689900 168790 689970
rect 168790 689900 168820 689970
rect 168820 689900 168830 689970
rect 168920 689900 168990 689970
rect 168990 689900 169020 689970
rect 169020 689900 169090 689970
rect 169090 689900 169120 689970
rect 169120 689900 169160 689970
rect 169250 689900 169290 689970
rect 169290 689900 169320 689970
rect 169320 689900 169390 689970
rect 169390 689900 169420 689970
rect 169420 689900 169490 689970
rect 169580 689900 169590 689970
rect 169590 689900 169620 689970
rect 169620 689900 169690 689970
rect 169690 689900 169720 689970
rect 169720 689900 169790 689970
rect 169790 689900 169820 689970
rect 169910 689900 169920 689970
rect 169920 689900 169990 689970
rect 169990 689900 170020 689970
rect 170020 689900 170090 689970
rect 170090 689900 170120 689970
rect 170120 689900 170150 689970
rect 170240 689900 170290 689970
rect 170290 689900 170320 689970
rect 170320 689900 170390 689970
rect 170390 689900 170420 689970
rect 170420 689900 170480 689970
rect 157818 642045 158078 642285
rect 158178 642045 158438 642285
rect 158538 642045 158798 642285
rect 158898 642045 159158 642285
rect 157818 641705 158078 641945
rect 158178 641705 158438 641945
rect 158538 641705 158798 641945
rect 158898 641705 159158 641945
rect 157818 641365 158078 641605
rect 158178 641365 158438 641605
rect 158538 641365 158798 641605
rect 158898 641365 159158 641605
rect 157818 641025 158078 641265
rect 158178 641025 158438 641265
rect 158538 641025 158798 641265
rect 158898 641025 159158 641265
rect 157818 640685 158078 640925
rect 158178 640685 158438 640925
rect 158538 640685 158798 640925
rect 158898 640685 159158 640925
rect 157818 640345 158078 640585
rect 158178 640345 158438 640585
rect 158538 640345 158798 640585
rect 158898 640345 159158 640585
rect 157818 640005 158078 640245
rect 158178 640005 158438 640245
rect 158538 640005 158798 640245
rect 158898 640005 159158 640245
rect 157818 639665 158078 639905
rect 158178 639665 158438 639905
rect 158538 639665 158798 639905
rect 158898 639665 159158 639905
rect 157818 639325 158078 639565
rect 158178 639325 158438 639565
rect 158538 639325 158798 639565
rect 158898 639325 159158 639565
rect 157818 638985 158078 639225
rect 158178 638985 158438 639225
rect 158538 638985 158798 639225
rect 158898 638985 159158 639225
rect 157818 638645 158078 638885
rect 158178 638645 158438 638885
rect 158538 638645 158798 638885
rect 158898 638645 159158 638885
rect 157818 638305 158078 638545
rect 158178 638305 158438 638545
rect 158538 638305 158798 638545
rect 158898 638305 159158 638545
rect 157818 637965 158078 638205
rect 158178 637965 158438 638205
rect 158538 637965 158798 638205
rect 158898 637965 159158 638205
rect 157818 637625 158078 637865
rect 158178 637625 158438 637865
rect 158538 637625 158798 637865
rect 158898 637625 159158 637865
<< metal5 >>
rect 68194 703800 73194 704000
rect 68194 703500 68352 703800
rect 68652 703500 68852 703800
rect 69152 703500 69352 703800
rect 69652 703500 69852 703800
rect 70152 703500 70352 703800
rect 70652 703500 70852 703800
rect 71152 703500 71352 703800
rect 71652 703500 71852 703800
rect 72152 703500 72352 703800
rect 72652 703500 72852 703800
rect 73152 703500 73194 703800
rect 68194 703300 73194 703500
rect 68194 703000 68352 703300
rect 68652 703000 68852 703300
rect 69152 703000 69352 703300
rect 69652 703000 69852 703300
rect 70152 703000 70352 703300
rect 70652 703000 70852 703300
rect 71152 703000 71352 703300
rect 71652 703000 71852 703300
rect 72152 703000 72352 703300
rect 72652 703000 72852 703300
rect 73152 703000 73194 703300
rect 68194 702800 73194 703000
rect 68194 702500 68352 702800
rect 68652 702500 68852 702800
rect 69152 702500 69352 702800
rect 69652 702500 69852 702800
rect 70152 702500 70352 702800
rect 70652 702500 70852 702800
rect 71152 702500 71352 702800
rect 71652 702500 71852 702800
rect 72152 702500 72352 702800
rect 72652 702500 72852 702800
rect 73152 702500 73194 702800
rect 68194 696090 73194 702500
rect 120194 703800 125194 704000
rect 120194 703500 120352 703800
rect 120652 703500 120852 703800
rect 121152 703500 121352 703800
rect 121652 703500 121852 703800
rect 122152 703500 122352 703800
rect 122652 703500 122852 703800
rect 123152 703500 123352 703800
rect 123652 703500 123852 703800
rect 124152 703500 124352 703800
rect 124652 703500 124852 703800
rect 125152 703500 125194 703800
rect 120194 703300 125194 703500
rect 120194 703000 120352 703300
rect 120652 703000 120852 703300
rect 121152 703000 121352 703300
rect 121652 703000 121852 703300
rect 122152 703000 122352 703300
rect 122652 703000 122852 703300
rect 123152 703000 123352 703300
rect 123652 703000 123852 703300
rect 124152 703000 124352 703300
rect 124652 703000 124852 703300
rect 125152 703000 125194 703300
rect 120194 702800 125194 703000
rect 120194 702500 120352 702800
rect 120652 702500 120852 702800
rect 121152 702500 121352 702800
rect 121652 702500 121852 702800
rect 122152 702500 122352 702800
rect 122652 702500 122852 702800
rect 123152 702500 123352 702800
rect 123652 702500 123852 702800
rect 124152 702500 124352 702800
rect 124652 702500 124852 702800
rect 125152 702500 125194 702800
rect 120194 696090 125194 702500
rect 68194 693190 84294 696090
rect 109094 693190 125194 696090
rect 165594 690140 170594 704800
rect 175894 701234 180894 704800
rect 217294 701234 222294 704800
rect 227594 699884 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 227594 699624 227767 699884
rect 228007 699624 228107 699884
rect 228347 699624 228447 699884
rect 228687 699624 228787 699884
rect 229027 699624 229127 699884
rect 229367 699624 229467 699884
rect 229707 699624 229807 699884
rect 230047 699624 230147 699884
rect 230387 699624 230487 699884
rect 230727 699624 230827 699884
rect 231067 699624 231167 699884
rect 231407 699624 231507 699884
rect 231747 699624 231847 699884
rect 232087 699624 232187 699884
rect 232427 699624 232594 699884
rect 227594 699524 232594 699624
rect 227594 699264 227767 699524
rect 228007 699264 228107 699524
rect 228347 699264 228447 699524
rect 228687 699264 228787 699524
rect 229027 699264 229127 699524
rect 229367 699264 229467 699524
rect 229707 699264 229807 699524
rect 230047 699264 230147 699524
rect 230387 699264 230487 699524
rect 230727 699264 230827 699524
rect 231067 699264 231167 699524
rect 231407 699264 231507 699524
rect 231747 699264 231847 699524
rect 232087 699264 232187 699524
rect 232427 699264 232594 699524
rect 227594 699164 232594 699264
rect 227594 698904 227767 699164
rect 228007 698904 228107 699164
rect 228347 698904 228447 699164
rect 228687 698904 228787 699164
rect 229027 698904 229127 699164
rect 229367 698904 229467 699164
rect 229707 698904 229807 699164
rect 230047 698904 230147 699164
rect 230387 698904 230487 699164
rect 230727 698904 230827 699164
rect 231067 698904 231167 699164
rect 231407 698904 231507 699164
rect 231747 698904 231847 699164
rect 232087 698904 232187 699164
rect 232427 698904 232594 699164
rect 227594 698804 232594 698904
rect 227594 698544 227767 698804
rect 228007 698544 228107 698804
rect 228347 698544 228447 698804
rect 228687 698544 228787 698804
rect 229027 698544 229127 698804
rect 229367 698544 229467 698804
rect 229707 698544 229807 698804
rect 230047 698544 230147 698804
rect 230387 698544 230487 698804
rect 230727 698544 230827 698804
rect 231067 698544 231167 698804
rect 231407 698544 231507 698804
rect 231747 698544 231847 698804
rect 232087 698544 232187 698804
rect 232427 698544 232594 698804
rect 227594 698464 232594 698544
rect 165594 689900 165620 690140
rect 165860 689900 165950 690140
rect 166190 689900 166280 690140
rect 166520 689900 166610 690140
rect 166850 689900 166940 690140
rect 167180 689900 167270 690140
rect 167510 689900 167600 690140
rect 167840 689900 167930 690140
rect 168170 689900 168260 690140
rect 168500 689900 168590 690140
rect 168830 689900 168920 690140
rect 169160 689900 169250 690140
rect 169490 689900 169580 690140
rect 169820 689900 169910 690140
rect 170150 689900 170240 690140
rect 170480 689900 170594 690140
rect 72330 676672 84314 682580
rect 72330 642452 77330 676672
rect 165594 675680 170594 689900
rect 165594 670680 225632 675680
rect 165594 651038 170594 670680
rect 82008 646038 226088 651038
rect 72330 642285 159238 642452
rect 72330 642045 157818 642285
rect 158078 642045 158178 642285
rect 158438 642045 158538 642285
rect 158798 642045 158898 642285
rect 159158 642045 159238 642285
rect 72330 641945 159238 642045
rect 72330 641705 157818 641945
rect 158078 641705 158178 641945
rect 158438 641705 158538 641945
rect 158798 641705 158898 641945
rect 159158 641705 159238 641945
rect 72330 641605 159238 641705
rect 72330 641365 157818 641605
rect 158078 641365 158178 641605
rect 158438 641365 158538 641605
rect 158798 641365 158898 641605
rect 159158 641365 159238 641605
rect 72330 641265 159238 641365
rect 72330 641025 157818 641265
rect 158078 641025 158178 641265
rect 158438 641025 158538 641265
rect 158798 641025 158898 641265
rect 159158 641025 159238 641265
rect 72330 640925 159238 641025
rect 72330 640685 157818 640925
rect 158078 640685 158178 640925
rect 158438 640685 158538 640925
rect 158798 640685 158898 640925
rect 159158 640685 159238 640925
rect 72330 640585 159238 640685
rect 72330 640345 157818 640585
rect 158078 640345 158178 640585
rect 158438 640345 158538 640585
rect 158798 640345 158898 640585
rect 159158 640345 159238 640585
rect 72330 640245 159238 640345
rect 72330 640005 157818 640245
rect 158078 640005 158178 640245
rect 158438 640005 158538 640245
rect 158798 640005 158898 640245
rect 159158 640005 159238 640245
rect 72330 639905 159238 640005
rect 72330 639665 157818 639905
rect 158078 639665 158178 639905
rect 158438 639665 158538 639905
rect 158798 639665 158898 639905
rect 159158 639665 159238 639905
rect 72330 639565 159238 639665
rect 72330 639325 157818 639565
rect 158078 639325 158178 639565
rect 158438 639325 158538 639565
rect 158798 639325 158898 639565
rect 159158 639325 159238 639565
rect 72330 639225 159238 639325
rect 72330 638985 157818 639225
rect 158078 638985 158178 639225
rect 158438 638985 158538 639225
rect 158798 638985 158898 639225
rect 159158 638985 159238 639225
rect 72330 638885 159238 638985
rect 72330 638645 157818 638885
rect 158078 638645 158178 638885
rect 158438 638645 158538 638885
rect 158798 638645 158898 638885
rect 159158 638645 159238 638885
rect 72330 638545 159238 638645
rect 72330 638305 157818 638545
rect 158078 638305 158178 638545
rect 158438 638305 158538 638545
rect 158798 638305 158898 638545
rect 159158 638305 159238 638545
rect 72330 638205 159238 638305
rect 72330 637965 157818 638205
rect 158078 637965 158178 638205
rect 158438 637965 158538 638205
rect 158798 637965 158898 638205
rect 159158 637965 159238 638205
rect 72330 637865 159238 637965
rect 72330 637625 157818 637865
rect 158078 637625 158178 637865
rect 158438 637625 158538 637865
rect 158798 637625 158898 637865
rect 159158 637625 159238 637865
rect 72330 637452 159238 637625
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 312 632584 583832 636642
rect 584000 0 584100 704000
rect -100 -100 584100 0
use big_cap  big_cap_1
timestamp 1636526374
transform 1 0 119364 0 1 670158
box 60730 -31110 106740 14450
use top  top_0
timestamp 1636213485
transform 1 0 89244 0 1 674450
box -6530 -24030 39650 21850
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
