magic
tech sky130A
magscale 1 2
timestamp 1637086603
<< nwell >>
rect 11630 16000 17124 17368
rect 17806 16000 23300 17368
<< pwell >>
rect 11630 12313 17124 13671
rect 17806 12313 23300 13671
<< pmoslvt >>
rect 11826 16220 12026 17220
rect 12084 16220 12284 17220
rect 12342 16220 12542 17220
rect 12600 16220 12800 17220
rect 12858 16220 13058 17220
rect 13116 16220 13316 17220
rect 13374 16220 13574 17220
rect 13632 16220 13832 17220
rect 13890 16220 14090 17220
rect 14148 16220 14348 17220
rect 14406 16220 14606 17220
rect 14664 16220 14864 17220
rect 14922 16220 15122 17220
rect 15180 16220 15380 17220
rect 15438 16220 15638 17220
rect 15696 16220 15896 17220
rect 15954 16220 16154 17220
rect 16212 16220 16412 17220
rect 16470 16220 16670 17220
rect 16728 16220 16928 17220
rect 18002 16220 18202 17220
rect 18260 16220 18460 17220
rect 18518 16220 18718 17220
rect 18776 16220 18976 17220
rect 19034 16220 19234 17220
rect 19292 16220 19492 17220
rect 19550 16220 19750 17220
rect 19808 16220 20008 17220
rect 20066 16220 20266 17220
rect 20324 16220 20524 17220
rect 20582 16220 20782 17220
rect 20840 16220 21040 17220
rect 21098 16220 21298 17220
rect 21356 16220 21556 17220
rect 21614 16220 21814 17220
rect 21872 16220 22072 17220
rect 22130 16220 22330 17220
rect 22388 16220 22588 17220
rect 22646 16220 22846 17220
rect 22904 16220 23104 17220
<< nmoslvt >>
rect 11826 12461 12026 13461
rect 12084 12461 12284 13461
rect 12342 12461 12542 13461
rect 12600 12461 12800 13461
rect 12858 12461 13058 13461
rect 13116 12461 13316 13461
rect 13374 12461 13574 13461
rect 13632 12461 13832 13461
rect 13890 12461 14090 13461
rect 14148 12461 14348 13461
rect 14406 12461 14606 13461
rect 14664 12461 14864 13461
rect 14922 12461 15122 13461
rect 15180 12461 15380 13461
rect 15438 12461 15638 13461
rect 15696 12461 15896 13461
rect 15954 12461 16154 13461
rect 16212 12461 16412 13461
rect 16470 12461 16670 13461
rect 16728 12461 16928 13461
rect 18002 12461 18202 13461
rect 18260 12461 18460 13461
rect 18518 12461 18718 13461
rect 18776 12461 18976 13461
rect 19034 12461 19234 13461
rect 19292 12461 19492 13461
rect 19550 12461 19750 13461
rect 19808 12461 20008 13461
rect 20066 12461 20266 13461
rect 20324 12461 20524 13461
rect 20582 12461 20782 13461
rect 20840 12461 21040 13461
rect 21098 12461 21298 13461
rect 21356 12461 21556 13461
rect 21614 12461 21814 13461
rect 21872 12461 22072 13461
rect 22130 12461 22330 13461
rect 22388 12461 22588 13461
rect 22646 12461 22846 13461
rect 22904 12461 23104 13461
<< ndiff >>
rect 11768 13449 11826 13461
rect 11768 12473 11780 13449
rect 11814 12473 11826 13449
rect 11768 12461 11826 12473
rect 12026 13449 12084 13461
rect 12026 12473 12038 13449
rect 12072 12473 12084 13449
rect 12026 12461 12084 12473
rect 12284 13449 12342 13461
rect 12284 12473 12296 13449
rect 12330 12473 12342 13449
rect 12284 12461 12342 12473
rect 12542 13449 12600 13461
rect 12542 12473 12554 13449
rect 12588 12473 12600 13449
rect 12542 12461 12600 12473
rect 12800 13449 12858 13461
rect 12800 12473 12812 13449
rect 12846 12473 12858 13449
rect 12800 12461 12858 12473
rect 13058 13449 13116 13461
rect 13058 12473 13070 13449
rect 13104 12473 13116 13449
rect 13058 12461 13116 12473
rect 13316 13449 13374 13461
rect 13316 12473 13328 13449
rect 13362 12473 13374 13449
rect 13316 12461 13374 12473
rect 13574 13449 13632 13461
rect 13574 12473 13586 13449
rect 13620 12473 13632 13449
rect 13574 12461 13632 12473
rect 13832 13449 13890 13461
rect 13832 12473 13844 13449
rect 13878 12473 13890 13449
rect 13832 12461 13890 12473
rect 14090 13449 14148 13461
rect 14090 12473 14102 13449
rect 14136 12473 14148 13449
rect 14090 12461 14148 12473
rect 14348 13449 14406 13461
rect 14348 12473 14360 13449
rect 14394 12473 14406 13449
rect 14348 12461 14406 12473
rect 14606 13449 14664 13461
rect 14606 12473 14618 13449
rect 14652 12473 14664 13449
rect 14606 12461 14664 12473
rect 14864 13449 14922 13461
rect 14864 12473 14876 13449
rect 14910 12473 14922 13449
rect 14864 12461 14922 12473
rect 15122 13449 15180 13461
rect 15122 12473 15134 13449
rect 15168 12473 15180 13449
rect 15122 12461 15180 12473
rect 15380 13449 15438 13461
rect 15380 12473 15392 13449
rect 15426 12473 15438 13449
rect 15380 12461 15438 12473
rect 15638 13449 15696 13461
rect 15638 12473 15650 13449
rect 15684 12473 15696 13449
rect 15638 12461 15696 12473
rect 15896 13449 15954 13461
rect 15896 12473 15908 13449
rect 15942 12473 15954 13449
rect 15896 12461 15954 12473
rect 16154 13449 16212 13461
rect 16154 12473 16166 13449
rect 16200 12473 16212 13449
rect 16154 12461 16212 12473
rect 16412 13449 16470 13461
rect 16412 12473 16424 13449
rect 16458 12473 16470 13449
rect 16412 12461 16470 12473
rect 16670 13449 16728 13461
rect 16670 12473 16682 13449
rect 16716 12473 16728 13449
rect 16670 12461 16728 12473
rect 16928 13449 16986 13461
rect 16928 12473 16940 13449
rect 16974 12473 16986 13449
rect 16928 12461 16986 12473
rect 17944 13449 18002 13461
rect 17944 12473 17956 13449
rect 17990 12473 18002 13449
rect 17944 12461 18002 12473
rect 18202 13449 18260 13461
rect 18202 12473 18214 13449
rect 18248 12473 18260 13449
rect 18202 12461 18260 12473
rect 18460 13449 18518 13461
rect 18460 12473 18472 13449
rect 18506 12473 18518 13449
rect 18460 12461 18518 12473
rect 18718 13449 18776 13461
rect 18718 12473 18730 13449
rect 18764 12473 18776 13449
rect 18718 12461 18776 12473
rect 18976 13449 19034 13461
rect 18976 12473 18988 13449
rect 19022 12473 19034 13449
rect 18976 12461 19034 12473
rect 19234 13449 19292 13461
rect 19234 12473 19246 13449
rect 19280 12473 19292 13449
rect 19234 12461 19292 12473
rect 19492 13449 19550 13461
rect 19492 12473 19504 13449
rect 19538 12473 19550 13449
rect 19492 12461 19550 12473
rect 19750 13449 19808 13461
rect 19750 12473 19762 13449
rect 19796 12473 19808 13449
rect 19750 12461 19808 12473
rect 20008 13449 20066 13461
rect 20008 12473 20020 13449
rect 20054 12473 20066 13449
rect 20008 12461 20066 12473
rect 20266 13449 20324 13461
rect 20266 12473 20278 13449
rect 20312 12473 20324 13449
rect 20266 12461 20324 12473
rect 20524 13449 20582 13461
rect 20524 12473 20536 13449
rect 20570 12473 20582 13449
rect 20524 12461 20582 12473
rect 20782 13449 20840 13461
rect 20782 12473 20794 13449
rect 20828 12473 20840 13449
rect 20782 12461 20840 12473
rect 21040 13449 21098 13461
rect 21040 12473 21052 13449
rect 21086 12473 21098 13449
rect 21040 12461 21098 12473
rect 21298 13449 21356 13461
rect 21298 12473 21310 13449
rect 21344 12473 21356 13449
rect 21298 12461 21356 12473
rect 21556 13449 21614 13461
rect 21556 12473 21568 13449
rect 21602 12473 21614 13449
rect 21556 12461 21614 12473
rect 21814 13449 21872 13461
rect 21814 12473 21826 13449
rect 21860 12473 21872 13449
rect 21814 12461 21872 12473
rect 22072 13449 22130 13461
rect 22072 12473 22084 13449
rect 22118 12473 22130 13449
rect 22072 12461 22130 12473
rect 22330 13449 22388 13461
rect 22330 12473 22342 13449
rect 22376 12473 22388 13449
rect 22330 12461 22388 12473
rect 22588 13449 22646 13461
rect 22588 12473 22600 13449
rect 22634 12473 22646 13449
rect 22588 12461 22646 12473
rect 22846 13449 22904 13461
rect 22846 12473 22858 13449
rect 22892 12473 22904 13449
rect 22846 12461 22904 12473
rect 23104 13449 23162 13461
rect 23104 12473 23116 13449
rect 23150 12473 23162 13449
rect 23104 12461 23162 12473
<< pdiff >>
rect 11768 17208 11826 17220
rect 11768 16232 11780 17208
rect 11814 16232 11826 17208
rect 11768 16220 11826 16232
rect 12026 17208 12084 17220
rect 12026 16232 12038 17208
rect 12072 16232 12084 17208
rect 12026 16220 12084 16232
rect 12284 17208 12342 17220
rect 12284 16232 12296 17208
rect 12330 16232 12342 17208
rect 12284 16220 12342 16232
rect 12542 17208 12600 17220
rect 12542 16232 12554 17208
rect 12588 16232 12600 17208
rect 12542 16220 12600 16232
rect 12800 17208 12858 17220
rect 12800 16232 12812 17208
rect 12846 16232 12858 17208
rect 12800 16220 12858 16232
rect 13058 17208 13116 17220
rect 13058 16232 13070 17208
rect 13104 16232 13116 17208
rect 13058 16220 13116 16232
rect 13316 17208 13374 17220
rect 13316 16232 13328 17208
rect 13362 16232 13374 17208
rect 13316 16220 13374 16232
rect 13574 17208 13632 17220
rect 13574 16232 13586 17208
rect 13620 16232 13632 17208
rect 13574 16220 13632 16232
rect 13832 17208 13890 17220
rect 13832 16232 13844 17208
rect 13878 16232 13890 17208
rect 13832 16220 13890 16232
rect 14090 17208 14148 17220
rect 14090 16232 14102 17208
rect 14136 16232 14148 17208
rect 14090 16220 14148 16232
rect 14348 17208 14406 17220
rect 14348 16232 14360 17208
rect 14394 16232 14406 17208
rect 14348 16220 14406 16232
rect 14606 17208 14664 17220
rect 14606 16232 14618 17208
rect 14652 16232 14664 17208
rect 14606 16220 14664 16232
rect 14864 17208 14922 17220
rect 14864 16232 14876 17208
rect 14910 16232 14922 17208
rect 14864 16220 14922 16232
rect 15122 17208 15180 17220
rect 15122 16232 15134 17208
rect 15168 16232 15180 17208
rect 15122 16220 15180 16232
rect 15380 17208 15438 17220
rect 15380 16232 15392 17208
rect 15426 16232 15438 17208
rect 15380 16220 15438 16232
rect 15638 17208 15696 17220
rect 15638 16232 15650 17208
rect 15684 16232 15696 17208
rect 15638 16220 15696 16232
rect 15896 17208 15954 17220
rect 15896 16232 15908 17208
rect 15942 16232 15954 17208
rect 15896 16220 15954 16232
rect 16154 17208 16212 17220
rect 16154 16232 16166 17208
rect 16200 16232 16212 17208
rect 16154 16220 16212 16232
rect 16412 17208 16470 17220
rect 16412 16232 16424 17208
rect 16458 16232 16470 17208
rect 16412 16220 16470 16232
rect 16670 17208 16728 17220
rect 16670 16232 16682 17208
rect 16716 16232 16728 17208
rect 16670 16220 16728 16232
rect 16928 17208 16986 17220
rect 16928 16232 16940 17208
rect 16974 16232 16986 17208
rect 16928 16220 16986 16232
rect 17944 17208 18002 17220
rect 17944 16232 17956 17208
rect 17990 16232 18002 17208
rect 17944 16220 18002 16232
rect 18202 17208 18260 17220
rect 18202 16232 18214 17208
rect 18248 16232 18260 17208
rect 18202 16220 18260 16232
rect 18460 17208 18518 17220
rect 18460 16232 18472 17208
rect 18506 16232 18518 17208
rect 18460 16220 18518 16232
rect 18718 17208 18776 17220
rect 18718 16232 18730 17208
rect 18764 16232 18776 17208
rect 18718 16220 18776 16232
rect 18976 17208 19034 17220
rect 18976 16232 18988 17208
rect 19022 16232 19034 17208
rect 18976 16220 19034 16232
rect 19234 17208 19292 17220
rect 19234 16232 19246 17208
rect 19280 16232 19292 17208
rect 19234 16220 19292 16232
rect 19492 17208 19550 17220
rect 19492 16232 19504 17208
rect 19538 16232 19550 17208
rect 19492 16220 19550 16232
rect 19750 17208 19808 17220
rect 19750 16232 19762 17208
rect 19796 16232 19808 17208
rect 19750 16220 19808 16232
rect 20008 17208 20066 17220
rect 20008 16232 20020 17208
rect 20054 16232 20066 17208
rect 20008 16220 20066 16232
rect 20266 17208 20324 17220
rect 20266 16232 20278 17208
rect 20312 16232 20324 17208
rect 20266 16220 20324 16232
rect 20524 17208 20582 17220
rect 20524 16232 20536 17208
rect 20570 16232 20582 17208
rect 20524 16220 20582 16232
rect 20782 17208 20840 17220
rect 20782 16232 20794 17208
rect 20828 16232 20840 17208
rect 20782 16220 20840 16232
rect 21040 17208 21098 17220
rect 21040 16232 21052 17208
rect 21086 16232 21098 17208
rect 21040 16220 21098 16232
rect 21298 17208 21356 17220
rect 21298 16232 21310 17208
rect 21344 16232 21356 17208
rect 21298 16220 21356 16232
rect 21556 17208 21614 17220
rect 21556 16232 21568 17208
rect 21602 16232 21614 17208
rect 21556 16220 21614 16232
rect 21814 17208 21872 17220
rect 21814 16232 21826 17208
rect 21860 16232 21872 17208
rect 21814 16220 21872 16232
rect 22072 17208 22130 17220
rect 22072 16232 22084 17208
rect 22118 16232 22130 17208
rect 22072 16220 22130 16232
rect 22330 17208 22388 17220
rect 22330 16232 22342 17208
rect 22376 16232 22388 17208
rect 22330 16220 22388 16232
rect 22588 17208 22646 17220
rect 22588 16232 22600 17208
rect 22634 16232 22646 17208
rect 22588 16220 22646 16232
rect 22846 17208 22904 17220
rect 22846 16232 22858 17208
rect 22892 16232 22904 17208
rect 22846 16220 22904 16232
rect 23104 17208 23162 17220
rect 23104 16232 23116 17208
rect 23150 16232 23162 17208
rect 23104 16220 23162 16232
<< ndiffc >>
rect 11780 12473 11814 13449
rect 12038 12473 12072 13449
rect 12296 12473 12330 13449
rect 12554 12473 12588 13449
rect 12812 12473 12846 13449
rect 13070 12473 13104 13449
rect 13328 12473 13362 13449
rect 13586 12473 13620 13449
rect 13844 12473 13878 13449
rect 14102 12473 14136 13449
rect 14360 12473 14394 13449
rect 14618 12473 14652 13449
rect 14876 12473 14910 13449
rect 15134 12473 15168 13449
rect 15392 12473 15426 13449
rect 15650 12473 15684 13449
rect 15908 12473 15942 13449
rect 16166 12473 16200 13449
rect 16424 12473 16458 13449
rect 16682 12473 16716 13449
rect 16940 12473 16974 13449
rect 17956 12473 17990 13449
rect 18214 12473 18248 13449
rect 18472 12473 18506 13449
rect 18730 12473 18764 13449
rect 18988 12473 19022 13449
rect 19246 12473 19280 13449
rect 19504 12473 19538 13449
rect 19762 12473 19796 13449
rect 20020 12473 20054 13449
rect 20278 12473 20312 13449
rect 20536 12473 20570 13449
rect 20794 12473 20828 13449
rect 21052 12473 21086 13449
rect 21310 12473 21344 13449
rect 21568 12473 21602 13449
rect 21826 12473 21860 13449
rect 22084 12473 22118 13449
rect 22342 12473 22376 13449
rect 22600 12473 22634 13449
rect 22858 12473 22892 13449
rect 23116 12473 23150 13449
<< pdiffc >>
rect 11780 16232 11814 17208
rect 12038 16232 12072 17208
rect 12296 16232 12330 17208
rect 12554 16232 12588 17208
rect 12812 16232 12846 17208
rect 13070 16232 13104 17208
rect 13328 16232 13362 17208
rect 13586 16232 13620 17208
rect 13844 16232 13878 17208
rect 14102 16232 14136 17208
rect 14360 16232 14394 17208
rect 14618 16232 14652 17208
rect 14876 16232 14910 17208
rect 15134 16232 15168 17208
rect 15392 16232 15426 17208
rect 15650 16232 15684 17208
rect 15908 16232 15942 17208
rect 16166 16232 16200 17208
rect 16424 16232 16458 17208
rect 16682 16232 16716 17208
rect 16940 16232 16974 17208
rect 17956 16232 17990 17208
rect 18214 16232 18248 17208
rect 18472 16232 18506 17208
rect 18730 16232 18764 17208
rect 18988 16232 19022 17208
rect 19246 16232 19280 17208
rect 19504 16232 19538 17208
rect 19762 16232 19796 17208
rect 20020 16232 20054 17208
rect 20278 16232 20312 17208
rect 20536 16232 20570 17208
rect 20794 16232 20828 17208
rect 21052 16232 21086 17208
rect 21310 16232 21344 17208
rect 21568 16232 21602 17208
rect 21826 16232 21860 17208
rect 22084 16232 22118 17208
rect 22342 16232 22376 17208
rect 22600 16232 22634 17208
rect 22858 16232 22892 17208
rect 23116 16232 23150 17208
<< psubdiff >>
rect 11666 13601 11762 13635
rect 16992 13601 17088 13635
rect 11666 13539 11700 13601
rect 17054 13539 17088 13601
rect 17842 13601 17938 13635
rect 23168 13601 23264 13635
rect 11666 12383 11700 12445
rect 17054 12383 17088 12445
rect 11666 12349 11762 12383
rect 16992 12349 17088 12383
rect 17842 13539 17876 13601
rect 23230 13539 23264 13601
rect 17842 12383 17876 12445
rect 23230 12383 23264 12445
rect 17842 12349 17938 12383
rect 23168 12349 23264 12383
<< nsubdiff >>
rect 11666 17298 11762 17332
rect 16992 17298 17088 17332
rect 11666 17235 11700 17298
rect 17054 17235 17088 17298
rect 11666 16070 11700 16133
rect 17054 16070 17088 16133
rect 17842 17298 17938 17332
rect 23168 17298 23264 17332
rect 17842 17235 17876 17298
rect 23230 17235 23264 17298
rect 11666 16036 11762 16070
rect 16992 16036 17088 16070
rect 17842 16070 17876 16133
rect 23230 16070 23264 16133
rect 17842 16036 17938 16070
rect 23168 16036 23264 16070
<< psubdiffcont >>
rect 11762 13601 16992 13635
rect 11666 12445 11700 13539
rect 17938 13601 23168 13635
rect 17054 12445 17088 13539
rect 11762 12349 16992 12383
rect 17842 12445 17876 13539
rect 23230 12445 23264 13539
rect 17938 12349 23168 12383
<< nsubdiffcont >>
rect 11762 17298 16992 17332
rect 11666 16133 11700 17235
rect 17054 16133 17088 17235
rect 17938 17298 23168 17332
rect 17842 16133 17876 17235
rect 11762 16036 16992 16070
rect 23230 16133 23264 17235
rect 17938 16036 23168 16070
<< poly >>
rect 11826 17220 12026 17246
rect 12084 17220 12284 17246
rect 12342 17220 12542 17246
rect 12600 17220 12800 17246
rect 12858 17220 13058 17246
rect 13116 17220 13316 17246
rect 13374 17220 13574 17246
rect 13632 17220 13832 17246
rect 13890 17220 14090 17246
rect 14148 17220 14348 17246
rect 14406 17220 14606 17246
rect 14664 17220 14864 17246
rect 14922 17220 15122 17246
rect 15180 17220 15380 17246
rect 15438 17220 15638 17246
rect 15696 17220 15896 17246
rect 15954 17220 16154 17246
rect 16212 17220 16412 17246
rect 16470 17220 16670 17246
rect 16728 17220 16928 17246
rect 11826 16173 12026 16220
rect 11826 16139 11842 16173
rect 12010 16139 12026 16173
rect 11826 16123 12026 16139
rect 12084 16173 12284 16220
rect 12084 16139 12100 16173
rect 12268 16139 12284 16173
rect 12084 16123 12284 16139
rect 12342 16173 12542 16220
rect 12342 16139 12358 16173
rect 12526 16139 12542 16173
rect 12342 16123 12542 16139
rect 12600 16173 12800 16220
rect 12600 16139 12616 16173
rect 12784 16139 12800 16173
rect 12600 16123 12800 16139
rect 12858 16173 13058 16220
rect 12858 16139 12874 16173
rect 13042 16139 13058 16173
rect 12858 16123 13058 16139
rect 13116 16173 13316 16220
rect 13116 16139 13132 16173
rect 13300 16139 13316 16173
rect 13116 16123 13316 16139
rect 13374 16173 13574 16220
rect 13374 16139 13390 16173
rect 13558 16139 13574 16173
rect 13374 16123 13574 16139
rect 13632 16173 13832 16220
rect 13632 16139 13648 16173
rect 13816 16139 13832 16173
rect 13632 16123 13832 16139
rect 13890 16173 14090 16220
rect 13890 16139 13906 16173
rect 14074 16139 14090 16173
rect 13890 16123 14090 16139
rect 14148 16173 14348 16220
rect 14148 16139 14164 16173
rect 14332 16139 14348 16173
rect 14148 16123 14348 16139
rect 14406 16173 14606 16220
rect 14406 16139 14422 16173
rect 14590 16139 14606 16173
rect 14406 16123 14606 16139
rect 14664 16173 14864 16220
rect 14664 16139 14680 16173
rect 14848 16139 14864 16173
rect 14664 16123 14864 16139
rect 14922 16173 15122 16220
rect 14922 16139 14938 16173
rect 15106 16139 15122 16173
rect 14922 16123 15122 16139
rect 15180 16173 15380 16220
rect 15180 16139 15196 16173
rect 15364 16139 15380 16173
rect 15180 16123 15380 16139
rect 15438 16173 15638 16220
rect 15438 16139 15454 16173
rect 15622 16139 15638 16173
rect 15438 16123 15638 16139
rect 15696 16173 15896 16220
rect 15696 16139 15712 16173
rect 15880 16139 15896 16173
rect 15696 16123 15896 16139
rect 15954 16173 16154 16220
rect 15954 16139 15970 16173
rect 16138 16139 16154 16173
rect 15954 16123 16154 16139
rect 16212 16173 16412 16220
rect 16212 16139 16228 16173
rect 16396 16139 16412 16173
rect 16212 16123 16412 16139
rect 16470 16173 16670 16220
rect 16470 16139 16486 16173
rect 16654 16139 16670 16173
rect 16470 16123 16670 16139
rect 16728 16173 16928 16220
rect 16728 16139 16744 16173
rect 16912 16139 16928 16173
rect 16728 16123 16928 16139
rect 18002 17220 18202 17246
rect 18260 17220 18460 17246
rect 18518 17220 18718 17246
rect 18776 17220 18976 17246
rect 19034 17220 19234 17246
rect 19292 17220 19492 17246
rect 19550 17220 19750 17246
rect 19808 17220 20008 17246
rect 20066 17220 20266 17246
rect 20324 17220 20524 17246
rect 20582 17220 20782 17246
rect 20840 17220 21040 17246
rect 21098 17220 21298 17246
rect 21356 17220 21556 17246
rect 21614 17220 21814 17246
rect 21872 17220 22072 17246
rect 22130 17220 22330 17246
rect 22388 17220 22588 17246
rect 22646 17220 22846 17246
rect 22904 17220 23104 17246
rect 17180 16090 17750 16100
rect 17180 16050 17200 16090
rect 17240 16050 17280 16090
rect 17320 16050 17360 16090
rect 17400 16050 17440 16090
rect 17480 16050 17520 16090
rect 17560 16050 17600 16090
rect 17640 16050 17680 16090
rect 17720 16050 17750 16090
rect 17180 16010 17750 16050
rect 18002 16173 18202 16220
rect 18002 16139 18018 16173
rect 18186 16139 18202 16173
rect 18002 16123 18202 16139
rect 18260 16173 18460 16220
rect 18260 16139 18276 16173
rect 18444 16139 18460 16173
rect 18260 16123 18460 16139
rect 18518 16173 18718 16220
rect 18518 16139 18534 16173
rect 18702 16139 18718 16173
rect 18518 16123 18718 16139
rect 18776 16173 18976 16220
rect 18776 16139 18792 16173
rect 18960 16139 18976 16173
rect 18776 16123 18976 16139
rect 19034 16173 19234 16220
rect 19034 16139 19050 16173
rect 19218 16139 19234 16173
rect 19034 16123 19234 16139
rect 19292 16173 19492 16220
rect 19292 16139 19308 16173
rect 19476 16139 19492 16173
rect 19292 16123 19492 16139
rect 19550 16173 19750 16220
rect 19550 16139 19566 16173
rect 19734 16139 19750 16173
rect 19550 16123 19750 16139
rect 19808 16173 20008 16220
rect 19808 16139 19824 16173
rect 19992 16139 20008 16173
rect 19808 16123 20008 16139
rect 20066 16173 20266 16220
rect 20066 16139 20082 16173
rect 20250 16139 20266 16173
rect 20066 16123 20266 16139
rect 20324 16173 20524 16220
rect 20324 16139 20340 16173
rect 20508 16139 20524 16173
rect 20324 16123 20524 16139
rect 20582 16173 20782 16220
rect 20582 16139 20598 16173
rect 20766 16139 20782 16173
rect 20582 16123 20782 16139
rect 20840 16173 21040 16220
rect 20840 16139 20856 16173
rect 21024 16139 21040 16173
rect 20840 16123 21040 16139
rect 21098 16173 21298 16220
rect 21098 16139 21114 16173
rect 21282 16139 21298 16173
rect 21098 16123 21298 16139
rect 21356 16173 21556 16220
rect 21356 16139 21372 16173
rect 21540 16139 21556 16173
rect 21356 16123 21556 16139
rect 21614 16173 21814 16220
rect 21614 16139 21630 16173
rect 21798 16139 21814 16173
rect 21614 16123 21814 16139
rect 21872 16173 22072 16220
rect 21872 16139 21888 16173
rect 22056 16139 22072 16173
rect 21872 16123 22072 16139
rect 22130 16173 22330 16220
rect 22130 16139 22146 16173
rect 22314 16139 22330 16173
rect 22130 16123 22330 16139
rect 22388 16173 22588 16220
rect 22388 16139 22404 16173
rect 22572 16139 22588 16173
rect 22388 16123 22588 16139
rect 22646 16173 22846 16220
rect 22646 16139 22662 16173
rect 22830 16139 22846 16173
rect 22646 16123 22846 16139
rect 22904 16173 23104 16220
rect 22904 16139 22920 16173
rect 23088 16139 23104 16173
rect 22904 16123 23104 16139
rect 17180 15970 17200 16010
rect 17240 15970 17280 16010
rect 17320 15970 17360 16010
rect 17400 15970 17440 16010
rect 17480 15970 17520 16010
rect 17560 15970 17600 16010
rect 17640 15970 17680 16010
rect 17720 15970 17750 16010
rect 17180 15930 17750 15970
rect 17180 15890 17200 15930
rect 17240 15890 17280 15930
rect 17320 15890 17360 15930
rect 17400 15890 17440 15930
rect 17480 15890 17520 15930
rect 17560 15890 17600 15930
rect 17640 15890 17680 15930
rect 17720 15890 17750 15930
rect 17180 15850 17750 15890
rect 17180 15810 17200 15850
rect 17240 15810 17280 15850
rect 17320 15810 17360 15850
rect 17400 15810 17440 15850
rect 17480 15810 17520 15850
rect 17560 15810 17600 15850
rect 17640 15810 17680 15850
rect 17720 15810 17750 15850
rect 17180 15770 17750 15810
rect 17180 15730 17200 15770
rect 17240 15730 17280 15770
rect 17320 15730 17360 15770
rect 17400 15730 17440 15770
rect 17480 15730 17520 15770
rect 17560 15730 17600 15770
rect 17640 15730 17680 15770
rect 17720 15730 17750 15770
rect 17180 15710 17750 15730
rect 17180 13980 17750 14000
rect 17180 13940 17200 13980
rect 17240 13940 17280 13980
rect 17320 13940 17360 13980
rect 17400 13940 17440 13980
rect 17480 13940 17520 13980
rect 17560 13940 17600 13980
rect 17640 13940 17680 13980
rect 17720 13940 17750 13980
rect 17180 13900 17750 13940
rect 17180 13860 17200 13900
rect 17240 13860 17280 13900
rect 17320 13860 17360 13900
rect 17400 13860 17440 13900
rect 17480 13860 17520 13900
rect 17560 13860 17600 13900
rect 17640 13860 17680 13900
rect 17720 13860 17750 13900
rect 17180 13820 17750 13860
rect 17180 13780 17200 13820
rect 17240 13780 17280 13820
rect 17320 13780 17360 13820
rect 17400 13780 17440 13820
rect 17480 13780 17520 13820
rect 17560 13780 17600 13820
rect 17640 13780 17680 13820
rect 17720 13780 17750 13820
rect 17180 13740 17750 13780
rect 17180 13700 17200 13740
rect 17240 13700 17280 13740
rect 17320 13700 17360 13740
rect 17400 13700 17440 13740
rect 17480 13700 17520 13740
rect 17560 13700 17600 13740
rect 17640 13700 17680 13740
rect 17720 13700 17750 13740
rect 17180 13660 17750 13700
rect 11826 13533 12026 13549
rect 11826 13499 11842 13533
rect 12010 13499 12026 13533
rect 11826 13461 12026 13499
rect 12084 13533 12284 13549
rect 12084 13499 12100 13533
rect 12268 13499 12284 13533
rect 12084 13461 12284 13499
rect 12342 13533 12542 13549
rect 12342 13499 12358 13533
rect 12526 13499 12542 13533
rect 12342 13461 12542 13499
rect 12600 13533 12800 13549
rect 12600 13499 12616 13533
rect 12784 13499 12800 13533
rect 12600 13461 12800 13499
rect 12858 13533 13058 13549
rect 12858 13499 12874 13533
rect 13042 13499 13058 13533
rect 12858 13461 13058 13499
rect 13116 13533 13316 13549
rect 13116 13499 13132 13533
rect 13300 13499 13316 13533
rect 13116 13461 13316 13499
rect 13374 13533 13574 13549
rect 13374 13499 13390 13533
rect 13558 13499 13574 13533
rect 13374 13461 13574 13499
rect 13632 13533 13832 13549
rect 13632 13499 13648 13533
rect 13816 13499 13832 13533
rect 13632 13461 13832 13499
rect 13890 13533 14090 13549
rect 13890 13499 13906 13533
rect 14074 13499 14090 13533
rect 13890 13461 14090 13499
rect 14148 13533 14348 13549
rect 14148 13499 14164 13533
rect 14332 13499 14348 13533
rect 14148 13461 14348 13499
rect 14406 13533 14606 13549
rect 14406 13499 14422 13533
rect 14590 13499 14606 13533
rect 14406 13461 14606 13499
rect 14664 13533 14864 13549
rect 14664 13499 14680 13533
rect 14848 13499 14864 13533
rect 14664 13461 14864 13499
rect 14922 13533 15122 13549
rect 14922 13499 14938 13533
rect 15106 13499 15122 13533
rect 14922 13461 15122 13499
rect 15180 13533 15380 13549
rect 15180 13499 15196 13533
rect 15364 13499 15380 13533
rect 15180 13461 15380 13499
rect 15438 13533 15638 13549
rect 15438 13499 15454 13533
rect 15622 13499 15638 13533
rect 15438 13461 15638 13499
rect 15696 13533 15896 13549
rect 15696 13499 15712 13533
rect 15880 13499 15896 13533
rect 15696 13461 15896 13499
rect 15954 13533 16154 13549
rect 15954 13499 15970 13533
rect 16138 13499 16154 13533
rect 15954 13461 16154 13499
rect 16212 13533 16412 13549
rect 16212 13499 16228 13533
rect 16396 13499 16412 13533
rect 16212 13461 16412 13499
rect 16470 13533 16670 13549
rect 16470 13499 16486 13533
rect 16654 13499 16670 13533
rect 16470 13461 16670 13499
rect 16728 13533 16928 13549
rect 16728 13499 16744 13533
rect 16912 13499 16928 13533
rect 16728 13461 16928 13499
rect 17180 13620 17200 13660
rect 17240 13620 17280 13660
rect 17320 13620 17360 13660
rect 17400 13620 17440 13660
rect 17480 13620 17520 13660
rect 17560 13620 17600 13660
rect 17640 13620 17680 13660
rect 17720 13620 17750 13660
rect 17180 13600 17750 13620
rect 11826 12435 12026 12461
rect 12084 12435 12284 12461
rect 12342 12435 12542 12461
rect 12600 12435 12800 12461
rect 12858 12435 13058 12461
rect 13116 12435 13316 12461
rect 13374 12435 13574 12461
rect 13632 12435 13832 12461
rect 13890 12435 14090 12461
rect 14148 12435 14348 12461
rect 14406 12435 14606 12461
rect 14664 12435 14864 12461
rect 14922 12435 15122 12461
rect 15180 12435 15380 12461
rect 15438 12435 15638 12461
rect 15696 12435 15896 12461
rect 15954 12435 16154 12461
rect 16212 12435 16412 12461
rect 16470 12435 16670 12461
rect 16728 12435 16928 12461
rect 18002 13533 18202 13549
rect 18002 13499 18018 13533
rect 18186 13499 18202 13533
rect 18002 13461 18202 13499
rect 18260 13533 18460 13549
rect 18260 13499 18276 13533
rect 18444 13499 18460 13533
rect 18260 13461 18460 13499
rect 18518 13533 18718 13549
rect 18518 13499 18534 13533
rect 18702 13499 18718 13533
rect 18518 13461 18718 13499
rect 18776 13533 18976 13549
rect 18776 13499 18792 13533
rect 18960 13499 18976 13533
rect 18776 13461 18976 13499
rect 19034 13533 19234 13549
rect 19034 13499 19050 13533
rect 19218 13499 19234 13533
rect 19034 13461 19234 13499
rect 19292 13533 19492 13549
rect 19292 13499 19308 13533
rect 19476 13499 19492 13533
rect 19292 13461 19492 13499
rect 19550 13533 19750 13549
rect 19550 13499 19566 13533
rect 19734 13499 19750 13533
rect 19550 13461 19750 13499
rect 19808 13533 20008 13549
rect 19808 13499 19824 13533
rect 19992 13499 20008 13533
rect 19808 13461 20008 13499
rect 20066 13533 20266 13549
rect 20066 13499 20082 13533
rect 20250 13499 20266 13533
rect 20066 13461 20266 13499
rect 20324 13533 20524 13549
rect 20324 13499 20340 13533
rect 20508 13499 20524 13533
rect 20324 13461 20524 13499
rect 20582 13533 20782 13549
rect 20582 13499 20598 13533
rect 20766 13499 20782 13533
rect 20582 13461 20782 13499
rect 20840 13533 21040 13549
rect 20840 13499 20856 13533
rect 21024 13499 21040 13533
rect 20840 13461 21040 13499
rect 21098 13533 21298 13549
rect 21098 13499 21114 13533
rect 21282 13499 21298 13533
rect 21098 13461 21298 13499
rect 21356 13533 21556 13549
rect 21356 13499 21372 13533
rect 21540 13499 21556 13533
rect 21356 13461 21556 13499
rect 21614 13533 21814 13549
rect 21614 13499 21630 13533
rect 21798 13499 21814 13533
rect 21614 13461 21814 13499
rect 21872 13533 22072 13549
rect 21872 13499 21888 13533
rect 22056 13499 22072 13533
rect 21872 13461 22072 13499
rect 22130 13533 22330 13549
rect 22130 13499 22146 13533
rect 22314 13499 22330 13533
rect 22130 13461 22330 13499
rect 22388 13533 22588 13549
rect 22388 13499 22404 13533
rect 22572 13499 22588 13533
rect 22388 13461 22588 13499
rect 22646 13533 22846 13549
rect 22646 13499 22662 13533
rect 22830 13499 22846 13533
rect 22646 13461 22846 13499
rect 22904 13533 23104 13549
rect 22904 13499 22920 13533
rect 23088 13499 23104 13533
rect 22904 13461 23104 13499
rect 18002 12435 18202 12461
rect 18260 12435 18460 12461
rect 18518 12435 18718 12461
rect 18776 12435 18976 12461
rect 19034 12435 19234 12461
rect 19292 12435 19492 12461
rect 19550 12435 19750 12461
rect 19808 12435 20008 12461
rect 20066 12435 20266 12461
rect 20324 12435 20524 12461
rect 20582 12435 20782 12461
rect 20840 12435 21040 12461
rect 21098 12435 21298 12461
rect 21356 12435 21556 12461
rect 21614 12435 21814 12461
rect 21872 12435 22072 12461
rect 22130 12435 22330 12461
rect 22388 12435 22588 12461
rect 22646 12435 22846 12461
rect 22904 12435 23104 12461
<< polycont >>
rect 11842 16139 12010 16173
rect 12100 16139 12268 16173
rect 12358 16139 12526 16173
rect 12616 16139 12784 16173
rect 12874 16139 13042 16173
rect 13132 16139 13300 16173
rect 13390 16139 13558 16173
rect 13648 16139 13816 16173
rect 13906 16139 14074 16173
rect 14164 16139 14332 16173
rect 14422 16139 14590 16173
rect 14680 16139 14848 16173
rect 14938 16139 15106 16173
rect 15196 16139 15364 16173
rect 15454 16139 15622 16173
rect 15712 16139 15880 16173
rect 15970 16139 16138 16173
rect 16228 16139 16396 16173
rect 16486 16139 16654 16173
rect 16744 16139 16912 16173
rect 17200 16050 17240 16090
rect 17280 16050 17320 16090
rect 17360 16050 17400 16090
rect 17440 16050 17480 16090
rect 17520 16050 17560 16090
rect 17600 16050 17640 16090
rect 17680 16050 17720 16090
rect 18018 16139 18186 16173
rect 18276 16139 18444 16173
rect 18534 16139 18702 16173
rect 18792 16139 18960 16173
rect 19050 16139 19218 16173
rect 19308 16139 19476 16173
rect 19566 16139 19734 16173
rect 19824 16139 19992 16173
rect 20082 16139 20250 16173
rect 20340 16139 20508 16173
rect 20598 16139 20766 16173
rect 20856 16139 21024 16173
rect 21114 16139 21282 16173
rect 21372 16139 21540 16173
rect 21630 16139 21798 16173
rect 21888 16139 22056 16173
rect 22146 16139 22314 16173
rect 22404 16139 22572 16173
rect 22662 16139 22830 16173
rect 22920 16139 23088 16173
rect 17200 15970 17240 16010
rect 17280 15970 17320 16010
rect 17360 15970 17400 16010
rect 17440 15970 17480 16010
rect 17520 15970 17560 16010
rect 17600 15970 17640 16010
rect 17680 15970 17720 16010
rect 17200 15890 17240 15930
rect 17280 15890 17320 15930
rect 17360 15890 17400 15930
rect 17440 15890 17480 15930
rect 17520 15890 17560 15930
rect 17600 15890 17640 15930
rect 17680 15890 17720 15930
rect 17200 15810 17240 15850
rect 17280 15810 17320 15850
rect 17360 15810 17400 15850
rect 17440 15810 17480 15850
rect 17520 15810 17560 15850
rect 17600 15810 17640 15850
rect 17680 15810 17720 15850
rect 17200 15730 17240 15770
rect 17280 15730 17320 15770
rect 17360 15730 17400 15770
rect 17440 15730 17480 15770
rect 17520 15730 17560 15770
rect 17600 15730 17640 15770
rect 17680 15730 17720 15770
rect 17200 13940 17240 13980
rect 17280 13940 17320 13980
rect 17360 13940 17400 13980
rect 17440 13940 17480 13980
rect 17520 13940 17560 13980
rect 17600 13940 17640 13980
rect 17680 13940 17720 13980
rect 17200 13860 17240 13900
rect 17280 13860 17320 13900
rect 17360 13860 17400 13900
rect 17440 13860 17480 13900
rect 17520 13860 17560 13900
rect 17600 13860 17640 13900
rect 17680 13860 17720 13900
rect 17200 13780 17240 13820
rect 17280 13780 17320 13820
rect 17360 13780 17400 13820
rect 17440 13780 17480 13820
rect 17520 13780 17560 13820
rect 17600 13780 17640 13820
rect 17680 13780 17720 13820
rect 17200 13700 17240 13740
rect 17280 13700 17320 13740
rect 17360 13700 17400 13740
rect 17440 13700 17480 13740
rect 17520 13700 17560 13740
rect 17600 13700 17640 13740
rect 17680 13700 17720 13740
rect 11842 13499 12010 13533
rect 12100 13499 12268 13533
rect 12358 13499 12526 13533
rect 12616 13499 12784 13533
rect 12874 13499 13042 13533
rect 13132 13499 13300 13533
rect 13390 13499 13558 13533
rect 13648 13499 13816 13533
rect 13906 13499 14074 13533
rect 14164 13499 14332 13533
rect 14422 13499 14590 13533
rect 14680 13499 14848 13533
rect 14938 13499 15106 13533
rect 15196 13499 15364 13533
rect 15454 13499 15622 13533
rect 15712 13499 15880 13533
rect 15970 13499 16138 13533
rect 16228 13499 16396 13533
rect 16486 13499 16654 13533
rect 16744 13499 16912 13533
rect 17200 13620 17240 13660
rect 17280 13620 17320 13660
rect 17360 13620 17400 13660
rect 17440 13620 17480 13660
rect 17520 13620 17560 13660
rect 17600 13620 17640 13660
rect 17680 13620 17720 13660
rect 18018 13499 18186 13533
rect 18276 13499 18444 13533
rect 18534 13499 18702 13533
rect 18792 13499 18960 13533
rect 19050 13499 19218 13533
rect 19308 13499 19476 13533
rect 19566 13499 19734 13533
rect 19824 13499 19992 13533
rect 20082 13499 20250 13533
rect 20340 13499 20508 13533
rect 20598 13499 20766 13533
rect 20856 13499 21024 13533
rect 21114 13499 21282 13533
rect 21372 13499 21540 13533
rect 21630 13499 21798 13533
rect 21888 13499 22056 13533
rect 22146 13499 22314 13533
rect 22404 13499 22572 13533
rect 22662 13499 22830 13533
rect 22920 13499 23088 13533
<< npolyres >>
rect 17180 14000 17750 15710
<< locali >>
rect 11666 17235 11700 17332
rect 17054 17235 17088 17332
rect 11780 17208 11814 17224
rect 11780 16216 11814 16232
rect 12038 17208 12072 17224
rect 12038 16173 12072 16232
rect 12296 17208 12330 17224
rect 12296 16216 12330 16232
rect 12554 17208 12588 17224
rect 12554 16173 12588 16232
rect 12812 17208 12846 17224
rect 12812 16216 12846 16232
rect 13070 17208 13104 17224
rect 13070 16173 13104 16232
rect 13328 17208 13362 17224
rect 13328 16216 13362 16232
rect 13586 17208 13620 17224
rect 13586 16173 13620 16232
rect 13844 17208 13878 17224
rect 13844 16216 13878 16232
rect 14102 17208 14136 17224
rect 14102 16173 14136 16232
rect 14360 17208 14394 17224
rect 14360 16216 14394 16232
rect 14618 17208 14652 17224
rect 14618 16173 14652 16232
rect 14876 17208 14910 17224
rect 14876 16216 14910 16232
rect 15134 17208 15168 17224
rect 15134 16173 15168 16232
rect 15392 17208 15426 17224
rect 15392 16216 15426 16232
rect 15650 17208 15684 17224
rect 15650 16173 15684 16232
rect 15908 17208 15942 17224
rect 15908 16216 15942 16232
rect 16166 17208 16200 17224
rect 16166 16173 16200 16232
rect 16424 17208 16458 17224
rect 16424 16216 16458 16232
rect 16682 17208 16716 17224
rect 16682 16173 16716 16232
rect 16940 17208 16974 17224
rect 16940 16216 16974 16232
rect 11780 16139 11842 16173
rect 12010 16139 12100 16173
rect 12268 16139 12358 16173
rect 12526 16139 12616 16173
rect 12784 16139 12874 16173
rect 13042 16139 13132 16173
rect 13300 16139 13390 16173
rect 13558 16139 13648 16173
rect 13816 16139 13906 16173
rect 14074 16139 14164 16173
rect 14332 16139 14422 16173
rect 14590 16139 14680 16173
rect 14848 16139 14938 16173
rect 15106 16139 15196 16173
rect 15364 16139 15454 16173
rect 15622 16139 15712 16173
rect 15880 16139 15970 16173
rect 16138 16139 16228 16173
rect 16396 16139 16486 16173
rect 16654 16139 16744 16173
rect 16912 16139 16974 16173
rect 11666 16070 11700 16133
rect 17054 16070 17088 16133
rect 17842 17235 17876 17332
rect 23230 17235 23264 17332
rect 17956 17208 17990 17224
rect 17956 16216 17990 16232
rect 18214 17208 18248 17224
rect 18214 16173 18248 16232
rect 18472 17208 18506 17224
rect 18472 16216 18506 16232
rect 18730 17208 18764 17224
rect 18730 16173 18764 16232
rect 18988 17208 19022 17224
rect 18988 16216 19022 16232
rect 19246 17208 19280 17224
rect 19246 16173 19280 16232
rect 19504 17208 19538 17224
rect 19504 16216 19538 16232
rect 19762 17208 19796 17224
rect 19762 16173 19796 16232
rect 20020 17208 20054 17224
rect 20020 16216 20054 16232
rect 20278 17208 20312 17224
rect 20278 16173 20312 16232
rect 20536 17208 20570 17224
rect 20536 16216 20570 16232
rect 20794 17208 20828 17224
rect 20794 16173 20828 16232
rect 21052 17208 21086 17224
rect 21052 16216 21086 16232
rect 21310 17208 21344 17224
rect 21310 16173 21344 16232
rect 21568 17208 21602 17224
rect 21568 16216 21602 16232
rect 21826 17208 21860 17224
rect 21826 16173 21860 16232
rect 22084 17208 22118 17224
rect 22084 16216 22118 16232
rect 22342 17208 22376 17224
rect 22342 16173 22376 16232
rect 22600 17208 22634 17224
rect 22600 16216 22634 16232
rect 22858 17208 22892 17224
rect 22858 16173 22892 16232
rect 23116 17208 23150 17224
rect 23116 16216 23150 16232
rect 17956 16139 18018 16173
rect 18186 16139 18276 16173
rect 18444 16139 18534 16173
rect 18702 16139 18792 16173
rect 18960 16139 19050 16173
rect 19218 16139 19308 16173
rect 19476 16139 19566 16173
rect 19734 16139 19824 16173
rect 19992 16139 20082 16173
rect 20250 16139 20340 16173
rect 20508 16139 20598 16173
rect 20766 16139 20856 16173
rect 21024 16139 21114 16173
rect 21282 16139 21372 16173
rect 21540 16139 21630 16173
rect 21798 16139 21888 16173
rect 22056 16139 22146 16173
rect 22314 16139 22404 16173
rect 22572 16139 22662 16173
rect 22830 16139 22920 16173
rect 23088 16139 23150 16173
rect 11666 16036 11762 16070
rect 16992 16036 17088 16070
rect 17180 16090 17750 16100
rect 17180 16050 17200 16090
rect 17240 16050 17280 16090
rect 17320 16050 17360 16090
rect 17400 16050 17440 16090
rect 17480 16050 17520 16090
rect 17560 16050 17600 16090
rect 17640 16050 17680 16090
rect 17720 16050 17750 16090
rect 17180 16010 17750 16050
rect 17842 16070 17876 16133
rect 23230 16070 23264 16133
rect 17842 16036 17938 16070
rect 23168 16036 23264 16070
rect 17180 15970 17200 16010
rect 17240 15970 17280 16010
rect 17320 15970 17360 16010
rect 17400 15970 17440 16010
rect 17480 15970 17520 16010
rect 17560 15970 17600 16010
rect 17640 15970 17680 16010
rect 17720 15970 17750 16010
rect 17180 15930 17750 15970
rect 17180 15890 17200 15930
rect 17240 15890 17280 15930
rect 17320 15890 17360 15930
rect 17400 15890 17440 15930
rect 17480 15890 17520 15930
rect 17560 15890 17600 15930
rect 17640 15890 17680 15930
rect 17720 15890 17750 15930
rect 17180 15850 17750 15890
rect 17180 15810 17200 15850
rect 17240 15810 17280 15850
rect 17320 15810 17360 15850
rect 17400 15810 17440 15850
rect 17480 15810 17520 15850
rect 17560 15810 17600 15850
rect 17640 15810 17680 15850
rect 17720 15810 17750 15850
rect 17180 15770 17750 15810
rect 17180 15730 17200 15770
rect 17240 15730 17280 15770
rect 17320 15730 17360 15770
rect 17400 15730 17440 15770
rect 17480 15730 17520 15770
rect 17560 15730 17600 15770
rect 17640 15730 17680 15770
rect 17720 15730 17750 15770
rect 17180 15710 17750 15730
rect 17180 13980 17750 14000
rect 17180 13940 17200 13980
rect 17240 13940 17280 13980
rect 17320 13940 17360 13980
rect 17400 13940 17440 13980
rect 17480 13940 17520 13980
rect 17560 13940 17600 13980
rect 17640 13940 17680 13980
rect 17720 13940 17750 13980
rect 17180 13900 17750 13940
rect 17180 13860 17200 13900
rect 17240 13860 17280 13900
rect 17320 13860 17360 13900
rect 17400 13860 17440 13900
rect 17480 13860 17520 13900
rect 17560 13860 17600 13900
rect 17640 13860 17680 13900
rect 17720 13860 17750 13900
rect 17180 13820 17750 13860
rect 17180 13780 17200 13820
rect 17240 13780 17280 13820
rect 17320 13780 17360 13820
rect 17400 13780 17440 13820
rect 17480 13780 17520 13820
rect 17560 13780 17600 13820
rect 17640 13780 17680 13820
rect 17720 13780 17750 13820
rect 17180 13740 17750 13780
rect 17180 13700 17200 13740
rect 17240 13700 17280 13740
rect 17320 13700 17360 13740
rect 17400 13700 17440 13740
rect 17480 13700 17520 13740
rect 17560 13700 17600 13740
rect 17640 13700 17680 13740
rect 17720 13700 17750 13740
rect 17180 13660 17750 13700
rect 11666 13601 11762 13635
rect 16992 13601 17088 13635
rect 11666 13539 11700 13601
rect 17054 13539 17088 13601
rect 17180 13620 17200 13660
rect 17240 13620 17280 13660
rect 17320 13620 17360 13660
rect 17400 13620 17440 13660
rect 17480 13620 17520 13660
rect 17560 13620 17600 13660
rect 17640 13620 17680 13660
rect 17720 13620 17750 13660
rect 17180 13600 17750 13620
rect 17842 13601 17938 13635
rect 23168 13601 23264 13635
rect 11778 13499 11842 13533
rect 12010 13499 12100 13533
rect 12268 13499 12358 13533
rect 12526 13499 12616 13533
rect 12784 13499 12874 13533
rect 13042 13499 13132 13533
rect 13300 13499 13390 13533
rect 13558 13499 13648 13533
rect 13816 13499 13906 13533
rect 14074 13499 14164 13533
rect 14332 13499 14422 13533
rect 14590 13499 14680 13533
rect 14848 13499 14938 13533
rect 15106 13499 15196 13533
rect 15364 13499 15454 13533
rect 15622 13499 15712 13533
rect 15880 13499 15970 13533
rect 16138 13499 16228 13533
rect 16396 13499 16486 13533
rect 16654 13499 16744 13533
rect 16912 13499 16975 13533
rect 11780 13449 11814 13465
rect 11780 12457 11814 12473
rect 12038 13449 12072 13499
rect 12038 12457 12072 12473
rect 12296 13449 12330 13465
rect 12296 12457 12330 12473
rect 12554 13449 12588 13499
rect 12554 12457 12588 12473
rect 12812 13449 12846 13465
rect 12812 12457 12846 12473
rect 13070 13449 13104 13499
rect 13070 12457 13104 12473
rect 13328 13449 13362 13465
rect 13328 12457 13362 12473
rect 13586 13449 13620 13499
rect 13586 12457 13620 12473
rect 13844 13449 13878 13465
rect 13844 12457 13878 12473
rect 14102 13449 14136 13499
rect 14102 12457 14136 12473
rect 14360 13449 14394 13465
rect 14360 12457 14394 12473
rect 14618 13449 14652 13499
rect 14618 12457 14652 12473
rect 14876 13449 14910 13465
rect 14876 12457 14910 12473
rect 15134 13449 15168 13499
rect 15134 12457 15168 12473
rect 15392 13449 15426 13465
rect 15392 12457 15426 12473
rect 15650 13449 15684 13499
rect 15650 12457 15684 12473
rect 15908 13449 15942 13465
rect 15908 12457 15942 12473
rect 16166 13449 16200 13499
rect 16166 12457 16200 12473
rect 16424 13449 16458 13465
rect 16424 12457 16458 12473
rect 16682 13449 16716 13499
rect 16682 12457 16716 12473
rect 16940 13449 16974 13465
rect 16940 12457 16974 12473
rect 11666 12349 11700 12445
rect 17054 12349 17088 12445
rect 17842 13539 17876 13601
rect 23230 13539 23264 13601
rect 17955 13499 18018 13533
rect 18186 13499 18276 13533
rect 18444 13499 18534 13533
rect 18702 13499 18792 13533
rect 18960 13499 19050 13533
rect 19218 13499 19308 13533
rect 19476 13499 19566 13533
rect 19734 13499 19824 13533
rect 19992 13499 20082 13533
rect 20250 13499 20340 13533
rect 20508 13499 20598 13533
rect 20766 13499 20856 13533
rect 21024 13499 21114 13533
rect 21282 13499 21372 13533
rect 21540 13499 21630 13533
rect 21798 13499 21888 13533
rect 22056 13499 22146 13533
rect 22314 13499 22404 13533
rect 22572 13499 22662 13533
rect 22830 13499 22920 13533
rect 23088 13499 23152 13533
rect 17956 13449 17990 13465
rect 17956 12457 17990 12473
rect 18214 13449 18248 13499
rect 18214 12457 18248 12473
rect 18472 13449 18506 13465
rect 18472 12457 18506 12473
rect 18730 13449 18764 13499
rect 18730 12457 18764 12473
rect 18988 13449 19022 13465
rect 18988 12457 19022 12473
rect 19246 13449 19280 13499
rect 19246 12457 19280 12473
rect 19504 13449 19538 13465
rect 19504 12457 19538 12473
rect 19762 13449 19796 13499
rect 19762 12457 19796 12473
rect 20020 13449 20054 13465
rect 20020 12457 20054 12473
rect 20278 13449 20312 13499
rect 20278 12457 20312 12473
rect 20536 13449 20570 13465
rect 20536 12457 20570 12473
rect 20794 13449 20828 13499
rect 20794 12457 20828 12473
rect 21052 13449 21086 13465
rect 21052 12457 21086 12473
rect 21310 13449 21344 13499
rect 21310 12457 21344 12473
rect 21568 13449 21602 13465
rect 21568 12457 21602 12473
rect 21826 13449 21860 13499
rect 21826 12457 21860 12473
rect 22084 13449 22118 13465
rect 22084 12457 22118 12473
rect 22342 13449 22376 13499
rect 22342 12457 22376 12473
rect 22600 13449 22634 13465
rect 22600 12457 22634 12473
rect 22858 13449 22892 13499
rect 22858 12457 22892 12473
rect 23116 13449 23150 13465
rect 23116 12457 23150 12473
rect 17842 12349 17876 12445
rect 23230 12349 23264 12445
<< viali >>
rect 11700 17298 11762 17332
rect 11762 17298 16992 17332
rect 16992 17298 17054 17332
rect 11666 16193 11700 17175
rect 11780 16232 11814 17208
rect 12038 16232 12072 17208
rect 12296 16232 12330 17208
rect 12554 16232 12588 17208
rect 12812 16232 12846 17208
rect 13070 16232 13104 17208
rect 13328 16232 13362 17208
rect 13586 16232 13620 17208
rect 13844 16232 13878 17208
rect 14102 16232 14136 17208
rect 14360 16232 14394 17208
rect 14618 16232 14652 17208
rect 14876 16232 14910 17208
rect 15134 16232 15168 17208
rect 15392 16232 15426 17208
rect 15650 16232 15684 17208
rect 15908 16232 15942 17208
rect 16166 16232 16200 17208
rect 16424 16232 16458 17208
rect 16682 16232 16716 17208
rect 16940 16232 16974 17208
rect 17054 16193 17088 17175
rect 11884 16139 11968 16173
rect 12142 16139 12226 16173
rect 12400 16139 12484 16173
rect 12658 16139 12742 16173
rect 12916 16139 13000 16173
rect 13174 16139 13258 16173
rect 13432 16139 13516 16173
rect 13690 16139 13774 16173
rect 13948 16139 14032 16173
rect 14206 16139 14290 16173
rect 14464 16139 14548 16173
rect 14722 16139 14806 16173
rect 14980 16139 15064 16173
rect 15238 16139 15322 16173
rect 15496 16139 15580 16173
rect 15754 16139 15838 16173
rect 16012 16139 16096 16173
rect 16270 16139 16354 16173
rect 16528 16139 16612 16173
rect 16786 16139 16870 16173
rect 17876 17298 17938 17332
rect 17938 17298 23168 17332
rect 23168 17298 23230 17332
rect 17842 16193 17876 17175
rect 17956 16232 17990 17208
rect 18214 16232 18248 17208
rect 18472 16232 18506 17208
rect 18730 16232 18764 17208
rect 18988 16232 19022 17208
rect 19246 16232 19280 17208
rect 19504 16232 19538 17208
rect 19762 16232 19796 17208
rect 20020 16232 20054 17208
rect 20278 16232 20312 17208
rect 20536 16232 20570 17208
rect 20794 16232 20828 17208
rect 21052 16232 21086 17208
rect 21310 16232 21344 17208
rect 21568 16232 21602 17208
rect 21826 16232 21860 17208
rect 22084 16232 22118 17208
rect 22342 16232 22376 17208
rect 22600 16232 22634 17208
rect 22858 16232 22892 17208
rect 23116 16232 23150 17208
rect 23230 16193 23264 17175
rect 18060 16139 18144 16173
rect 18318 16139 18402 16173
rect 18576 16139 18660 16173
rect 18834 16139 18918 16173
rect 19092 16139 19176 16173
rect 19350 16139 19434 16173
rect 19608 16139 19692 16173
rect 19866 16139 19950 16173
rect 20124 16139 20208 16173
rect 20382 16139 20466 16173
rect 20640 16139 20724 16173
rect 20898 16139 20982 16173
rect 21156 16139 21240 16173
rect 21414 16139 21498 16173
rect 21672 16139 21756 16173
rect 21930 16139 22014 16173
rect 22188 16139 22272 16173
rect 22446 16139 22530 16173
rect 22704 16139 22788 16173
rect 22962 16139 23046 16173
rect 17200 16050 17240 16090
rect 17280 16050 17320 16090
rect 17360 16050 17400 16090
rect 17440 16050 17480 16090
rect 17520 16050 17560 16090
rect 17600 16050 17640 16090
rect 17680 16050 17720 16090
rect 17200 15970 17240 16010
rect 17280 15970 17320 16010
rect 17360 15970 17400 16010
rect 17440 15970 17480 16010
rect 17520 15970 17560 16010
rect 17600 15970 17640 16010
rect 17680 15970 17720 16010
rect 17200 15890 17240 15930
rect 17280 15890 17320 15930
rect 17360 15890 17400 15930
rect 17440 15890 17480 15930
rect 17520 15890 17560 15930
rect 17600 15890 17640 15930
rect 17680 15890 17720 15930
rect 17200 13780 17240 13820
rect 17280 13780 17320 13820
rect 17360 13780 17400 13820
rect 17440 13780 17480 13820
rect 17520 13780 17560 13820
rect 17600 13780 17640 13820
rect 17680 13780 17720 13820
rect 17200 13700 17240 13740
rect 17280 13700 17320 13740
rect 17360 13700 17400 13740
rect 17440 13700 17480 13740
rect 17520 13700 17560 13740
rect 17600 13700 17640 13740
rect 17680 13700 17720 13740
rect 17200 13620 17240 13660
rect 17280 13620 17320 13660
rect 17360 13620 17400 13660
rect 17440 13620 17480 13660
rect 17520 13620 17560 13660
rect 17600 13620 17640 13660
rect 17680 13620 17720 13660
rect 11884 13499 11968 13533
rect 12142 13499 12226 13533
rect 12400 13499 12484 13533
rect 12658 13499 12742 13533
rect 12916 13499 13000 13533
rect 13174 13499 13258 13533
rect 13432 13499 13516 13533
rect 13690 13499 13774 13533
rect 13948 13499 14032 13533
rect 14206 13499 14290 13533
rect 14464 13499 14548 13533
rect 14722 13499 14806 13533
rect 14980 13499 15064 13533
rect 15238 13499 15322 13533
rect 15496 13499 15580 13533
rect 15754 13499 15838 13533
rect 16012 13499 16096 13533
rect 16270 13499 16354 13533
rect 16528 13499 16612 13533
rect 16786 13499 16870 13533
rect 11666 12505 11700 13479
rect 11780 12473 11814 13449
rect 12038 12473 12072 13449
rect 12296 12473 12330 13449
rect 12554 12473 12588 13449
rect 12812 12473 12846 13449
rect 13070 12473 13104 13449
rect 13328 12473 13362 13449
rect 13586 12473 13620 13449
rect 13844 12473 13878 13449
rect 14102 12473 14136 13449
rect 14360 12473 14394 13449
rect 14618 12473 14652 13449
rect 14876 12473 14910 13449
rect 15134 12473 15168 13449
rect 15392 12473 15426 13449
rect 15650 12473 15684 13449
rect 15908 12473 15942 13449
rect 16166 12473 16200 13449
rect 16424 12473 16458 13449
rect 16682 12473 16716 13449
rect 16940 12473 16974 13449
rect 17054 12505 17088 13479
rect 11700 12349 11762 12383
rect 11762 12349 16992 12383
rect 16992 12349 17054 12383
rect 18060 13499 18144 13533
rect 18318 13499 18402 13533
rect 18576 13499 18660 13533
rect 18834 13499 18918 13533
rect 19092 13499 19176 13533
rect 19350 13499 19434 13533
rect 19608 13499 19692 13533
rect 19866 13499 19950 13533
rect 20124 13499 20208 13533
rect 20382 13499 20466 13533
rect 20640 13499 20724 13533
rect 20898 13499 20982 13533
rect 21156 13499 21240 13533
rect 21414 13499 21498 13533
rect 21672 13499 21756 13533
rect 21930 13499 22014 13533
rect 22188 13499 22272 13533
rect 22446 13499 22530 13533
rect 22704 13499 22788 13533
rect 22962 13499 23046 13533
rect 17842 12505 17876 13479
rect 17956 12473 17990 13449
rect 18214 12473 18248 13449
rect 18472 12473 18506 13449
rect 18730 12473 18764 13449
rect 18988 12473 19022 13449
rect 19246 12473 19280 13449
rect 19504 12473 19538 13449
rect 19762 12473 19796 13449
rect 20020 12473 20054 13449
rect 20278 12473 20312 13449
rect 20536 12473 20570 13449
rect 20794 12473 20828 13449
rect 21052 12473 21086 13449
rect 21310 12473 21344 13449
rect 21568 12473 21602 13449
rect 21826 12473 21860 13449
rect 22084 12473 22118 13449
rect 22342 12473 22376 13449
rect 22600 12473 22634 13449
rect 22858 12473 22892 13449
rect 23116 12473 23150 13449
rect 23230 12505 23264 13479
rect 17876 12349 17938 12383
rect 17938 12349 23168 12383
rect 23168 12349 23230 12383
<< metal1 >>
rect 11690 17590 11930 17610
rect 12020 17590 12260 17610
rect 12350 17590 12590 17610
rect 12680 17590 12920 17610
rect 13010 17590 13250 17610
rect 13340 17590 13580 17610
rect 13670 17590 13910 17610
rect 14000 17590 14240 17610
rect 14330 17590 14570 17610
rect 14660 17590 14900 17610
rect 14990 17590 15230 17610
rect 15320 17590 15560 17610
rect 15650 17590 15890 17610
rect 15980 17590 16220 17610
rect 16310 17590 16550 17610
rect 16640 17590 16880 17610
rect 18050 17590 18290 17610
rect 18380 17590 18620 17610
rect 18710 17590 18950 17610
rect 19040 17590 19280 17610
rect 19370 17590 19610 17610
rect 19700 17590 19940 17610
rect 20030 17590 20270 17610
rect 20360 17590 20600 17610
rect 20690 17590 20930 17610
rect 21020 17590 21260 17610
rect 21350 17590 21590 17610
rect 21680 17590 21920 17610
rect 22010 17590 22250 17610
rect 22340 17590 22580 17610
rect 22670 17590 22910 17610
rect 23000 17590 23240 17610
rect 11660 17570 17094 17590
rect 11660 17560 14660 17570
rect 11660 17490 11690 17560
rect 11760 17490 11810 17560
rect 11880 17490 12020 17560
rect 12090 17490 12140 17560
rect 12210 17490 12350 17560
rect 12420 17490 12470 17560
rect 12540 17490 12680 17560
rect 12750 17490 12800 17560
rect 12870 17490 13010 17560
rect 13080 17490 13130 17560
rect 13200 17490 13340 17560
rect 13410 17490 13460 17560
rect 13530 17490 13670 17560
rect 13740 17490 13790 17560
rect 13860 17490 14000 17560
rect 14070 17490 14120 17560
rect 14190 17490 14330 17560
rect 14400 17490 14450 17560
rect 14520 17500 14660 17560
rect 14730 17500 14780 17570
rect 14850 17500 14990 17570
rect 15060 17500 15110 17570
rect 15180 17500 15320 17570
rect 15390 17500 15440 17570
rect 15510 17560 17094 17570
rect 15510 17500 15650 17560
rect 14520 17490 15650 17500
rect 15720 17490 15770 17560
rect 15840 17490 15980 17560
rect 16050 17490 16100 17560
rect 16170 17490 16310 17560
rect 16380 17490 16430 17560
rect 16500 17490 16640 17560
rect 16710 17490 16760 17560
rect 16830 17490 17094 17560
rect 11660 17450 17094 17490
rect 11660 17440 14660 17450
rect 11660 17370 11690 17440
rect 11760 17370 11810 17440
rect 11880 17370 12020 17440
rect 12090 17370 12140 17440
rect 12210 17370 12350 17440
rect 12420 17370 12470 17440
rect 12540 17370 12680 17440
rect 12750 17370 12800 17440
rect 12870 17370 13010 17440
rect 13080 17370 13130 17440
rect 13200 17370 13340 17440
rect 13410 17370 13460 17440
rect 13530 17370 13670 17440
rect 13740 17370 13790 17440
rect 13860 17370 14000 17440
rect 14070 17370 14120 17440
rect 14190 17370 14330 17440
rect 14400 17370 14450 17440
rect 14520 17380 14660 17440
rect 14730 17380 14780 17450
rect 14850 17380 14990 17450
rect 15060 17380 15110 17450
rect 15180 17380 15320 17450
rect 15390 17380 15440 17450
rect 15510 17440 17094 17450
rect 15510 17380 15650 17440
rect 14520 17370 15650 17380
rect 15720 17370 15770 17440
rect 15840 17370 15980 17440
rect 16050 17370 16100 17440
rect 16170 17370 16310 17440
rect 16380 17370 16430 17440
rect 16500 17370 16640 17440
rect 16710 17370 16760 17440
rect 16830 17370 17094 17440
rect 11660 17332 17094 17370
rect 11660 17298 11700 17332
rect 17054 17298 17094 17332
rect 11660 17292 17094 17298
rect 11660 17175 11706 17292
rect 11660 16193 11666 17175
rect 11700 16193 11706 17175
rect 11660 16181 11706 16193
rect 11774 17208 11820 17220
rect 11774 16232 11780 17208
rect 11814 16232 11820 17208
rect 11774 16100 11820 16232
rect 12032 17208 12078 17292
rect 12032 16232 12038 17208
rect 12072 16232 12078 17208
rect 12032 16220 12078 16232
rect 12290 17208 12336 17220
rect 12290 16232 12296 17208
rect 12330 16232 12336 17208
rect 11872 16173 11980 16179
rect 11872 16139 11884 16173
rect 11968 16139 11980 16173
rect 11872 16133 11980 16139
rect 12130 16173 12238 16179
rect 12130 16139 12142 16173
rect 12226 16139 12238 16173
rect 12130 16133 12238 16139
rect 12290 16100 12336 16232
rect 12548 17208 12594 17292
rect 12548 16232 12554 17208
rect 12588 16232 12594 17208
rect 12548 16220 12594 16232
rect 12806 17208 12852 17220
rect 12806 16232 12812 17208
rect 12846 16232 12852 17208
rect 12388 16173 12496 16179
rect 12388 16139 12400 16173
rect 12484 16139 12496 16173
rect 12388 16133 12496 16139
rect 12646 16173 12754 16179
rect 12646 16139 12658 16173
rect 12742 16139 12754 16173
rect 12646 16133 12754 16139
rect 12806 16100 12852 16232
rect 13064 17208 13110 17292
rect 13064 16232 13070 17208
rect 13104 16232 13110 17208
rect 13064 16220 13110 16232
rect 13322 17208 13368 17220
rect 13322 16232 13328 17208
rect 13362 16232 13368 17208
rect 12904 16173 13012 16179
rect 12904 16139 12916 16173
rect 13000 16139 13012 16173
rect 12904 16133 13012 16139
rect 13162 16173 13270 16179
rect 13162 16139 13174 16173
rect 13258 16139 13270 16173
rect 13162 16133 13270 16139
rect 13322 16100 13368 16232
rect 13580 17208 13626 17292
rect 13580 16232 13586 17208
rect 13620 16232 13626 17208
rect 13580 16220 13626 16232
rect 13838 17208 13884 17220
rect 13838 16232 13844 17208
rect 13878 16232 13884 17208
rect 13420 16173 13528 16179
rect 13420 16139 13432 16173
rect 13516 16139 13528 16173
rect 13420 16133 13528 16139
rect 13678 16173 13786 16179
rect 13678 16139 13690 16173
rect 13774 16139 13786 16173
rect 13678 16133 13786 16139
rect 13838 16100 13884 16232
rect 14096 17208 14142 17292
rect 14096 16232 14102 17208
rect 14136 16232 14142 17208
rect 14096 16220 14142 16232
rect 14354 17208 14400 17220
rect 14354 16232 14360 17208
rect 14394 16232 14400 17208
rect 13936 16173 14044 16179
rect 13936 16139 13948 16173
rect 14032 16139 14044 16173
rect 13936 16133 14044 16139
rect 14194 16173 14302 16179
rect 14194 16139 14206 16173
rect 14290 16139 14302 16173
rect 14194 16133 14302 16139
rect 14354 16100 14400 16232
rect 14612 17208 14658 17292
rect 14612 16232 14618 17208
rect 14652 16232 14658 17208
rect 14612 16220 14658 16232
rect 14870 17208 14916 17220
rect 14870 16232 14876 17208
rect 14910 16232 14916 17208
rect 14452 16173 14560 16179
rect 14452 16139 14464 16173
rect 14548 16139 14560 16173
rect 14452 16133 14560 16139
rect 14710 16173 14818 16179
rect 14710 16139 14722 16173
rect 14806 16139 14818 16173
rect 14710 16133 14818 16139
rect 14870 16100 14916 16232
rect 15128 17208 15174 17292
rect 15128 16232 15134 17208
rect 15168 16232 15174 17208
rect 15128 16220 15174 16232
rect 15386 17208 15432 17220
rect 15386 16232 15392 17208
rect 15426 16232 15432 17208
rect 14968 16173 15076 16179
rect 14968 16139 14980 16173
rect 15064 16139 15076 16173
rect 14968 16133 15076 16139
rect 15226 16173 15334 16179
rect 15226 16139 15238 16173
rect 15322 16139 15334 16173
rect 15226 16133 15334 16139
rect 15386 16100 15432 16232
rect 15644 17208 15690 17292
rect 15644 16232 15650 17208
rect 15684 16232 15690 17208
rect 15644 16220 15690 16232
rect 15902 17208 15948 17220
rect 15902 16232 15908 17208
rect 15942 16232 15948 17208
rect 15484 16173 15592 16179
rect 15484 16139 15496 16173
rect 15580 16139 15592 16173
rect 15484 16133 15592 16139
rect 15742 16173 15850 16179
rect 15742 16139 15754 16173
rect 15838 16139 15850 16173
rect 15742 16133 15850 16139
rect 15902 16100 15948 16232
rect 16160 17208 16206 17292
rect 16160 16232 16166 17208
rect 16200 16232 16206 17208
rect 16160 16220 16206 16232
rect 16418 17208 16464 17220
rect 16418 16232 16424 17208
rect 16458 16232 16464 17208
rect 16000 16173 16108 16179
rect 16000 16139 16012 16173
rect 16096 16139 16108 16173
rect 16000 16133 16108 16139
rect 16258 16173 16366 16179
rect 16258 16139 16270 16173
rect 16354 16139 16366 16173
rect 16258 16133 16366 16139
rect 16418 16100 16464 16232
rect 16676 17208 16722 17292
rect 16676 16232 16682 17208
rect 16716 16232 16722 17208
rect 16676 16220 16722 16232
rect 16934 17208 16980 17220
rect 16934 16232 16940 17208
rect 16974 16232 16980 17208
rect 16516 16173 16624 16179
rect 16516 16139 16528 16173
rect 16612 16139 16624 16173
rect 16516 16133 16624 16139
rect 16774 16173 16882 16179
rect 16774 16139 16786 16173
rect 16870 16139 16882 16173
rect 16774 16133 16882 16139
rect 16934 16100 16980 16232
rect 17048 17175 17094 17292
rect 17048 16193 17054 17175
rect 17088 16193 17094 17175
rect 17048 16181 17094 16193
rect 17836 17570 23270 17590
rect 17836 17560 19420 17570
rect 17836 17490 18100 17560
rect 18170 17490 18220 17560
rect 18290 17490 18430 17560
rect 18500 17490 18550 17560
rect 18620 17490 18760 17560
rect 18830 17490 18880 17560
rect 18950 17490 19090 17560
rect 19160 17490 19210 17560
rect 19280 17500 19420 17560
rect 19490 17500 19540 17570
rect 19610 17500 19750 17570
rect 19820 17500 19870 17570
rect 19940 17500 20080 17570
rect 20150 17500 20200 17570
rect 20270 17560 23270 17570
rect 20270 17500 20410 17560
rect 19280 17490 20410 17500
rect 20480 17490 20530 17560
rect 20600 17490 20740 17560
rect 20810 17490 20860 17560
rect 20930 17490 21070 17560
rect 21140 17490 21190 17560
rect 21260 17490 21400 17560
rect 21470 17490 21520 17560
rect 21590 17490 21730 17560
rect 21800 17490 21850 17560
rect 21920 17490 22060 17560
rect 22130 17490 22180 17560
rect 22250 17490 22390 17560
rect 22460 17490 22510 17560
rect 22580 17490 22720 17560
rect 22790 17490 22840 17560
rect 22910 17490 23050 17560
rect 23120 17490 23170 17560
rect 23240 17490 23270 17560
rect 17836 17450 23270 17490
rect 17836 17440 19420 17450
rect 17836 17370 18100 17440
rect 18170 17370 18220 17440
rect 18290 17370 18430 17440
rect 18500 17370 18550 17440
rect 18620 17370 18760 17440
rect 18830 17370 18880 17440
rect 18950 17370 19090 17440
rect 19160 17370 19210 17440
rect 19280 17380 19420 17440
rect 19490 17380 19540 17450
rect 19610 17380 19750 17450
rect 19820 17380 19870 17450
rect 19940 17380 20080 17450
rect 20150 17380 20200 17450
rect 20270 17440 23270 17450
rect 20270 17380 20410 17440
rect 19280 17370 20410 17380
rect 20480 17370 20530 17440
rect 20600 17370 20740 17440
rect 20810 17370 20860 17440
rect 20930 17370 21070 17440
rect 21140 17370 21190 17440
rect 21260 17370 21400 17440
rect 21470 17370 21520 17440
rect 21590 17370 21730 17440
rect 21800 17370 21850 17440
rect 21920 17370 22060 17440
rect 22130 17370 22180 17440
rect 22250 17370 22390 17440
rect 22460 17370 22510 17440
rect 22580 17370 22720 17440
rect 22790 17370 22840 17440
rect 22910 17370 23050 17440
rect 23120 17370 23170 17440
rect 23240 17370 23270 17440
rect 17836 17332 23270 17370
rect 17836 17298 17876 17332
rect 23230 17298 23270 17332
rect 17836 17292 23270 17298
rect 17836 17175 17882 17292
rect 17836 16193 17842 17175
rect 17876 16193 17882 17175
rect 17836 16181 17882 16193
rect 17950 17208 17996 17220
rect 17950 16232 17956 17208
rect 17990 16232 17996 17208
rect 17950 16100 17996 16232
rect 18208 17208 18254 17292
rect 18208 16232 18214 17208
rect 18248 16232 18254 17208
rect 18208 16220 18254 16232
rect 18466 17208 18512 17220
rect 18466 16232 18472 17208
rect 18506 16232 18512 17208
rect 18048 16173 18156 16179
rect 18048 16139 18060 16173
rect 18144 16139 18156 16173
rect 18048 16133 18156 16139
rect 18306 16173 18414 16179
rect 18306 16139 18318 16173
rect 18402 16139 18414 16173
rect 18306 16133 18414 16139
rect 18466 16100 18512 16232
rect 18724 17208 18770 17292
rect 18724 16232 18730 17208
rect 18764 16232 18770 17208
rect 18724 16220 18770 16232
rect 18982 17208 19028 17220
rect 18982 16232 18988 17208
rect 19022 16232 19028 17208
rect 18564 16173 18672 16179
rect 18564 16139 18576 16173
rect 18660 16139 18672 16173
rect 18564 16133 18672 16139
rect 18822 16173 18930 16179
rect 18822 16139 18834 16173
rect 18918 16139 18930 16173
rect 18822 16133 18930 16139
rect 18982 16100 19028 16232
rect 19240 17208 19286 17292
rect 19240 16232 19246 17208
rect 19280 16232 19286 17208
rect 19240 16220 19286 16232
rect 19498 17208 19544 17220
rect 19498 16232 19504 17208
rect 19538 16232 19544 17208
rect 19080 16173 19188 16179
rect 19080 16139 19092 16173
rect 19176 16139 19188 16173
rect 19080 16133 19188 16139
rect 19338 16173 19446 16179
rect 19338 16139 19350 16173
rect 19434 16139 19446 16173
rect 19338 16133 19446 16139
rect 19498 16100 19544 16232
rect 19756 17208 19802 17292
rect 19756 16232 19762 17208
rect 19796 16232 19802 17208
rect 19756 16220 19802 16232
rect 20014 17208 20060 17220
rect 20014 16232 20020 17208
rect 20054 16232 20060 17208
rect 19596 16173 19704 16179
rect 19596 16139 19608 16173
rect 19692 16139 19704 16173
rect 19596 16133 19704 16139
rect 19854 16173 19962 16179
rect 19854 16139 19866 16173
rect 19950 16139 19962 16173
rect 19854 16133 19962 16139
rect 20014 16100 20060 16232
rect 20272 17208 20318 17292
rect 20272 16232 20278 17208
rect 20312 16232 20318 17208
rect 20272 16220 20318 16232
rect 20530 17208 20576 17220
rect 20530 16232 20536 17208
rect 20570 16232 20576 17208
rect 20112 16173 20220 16179
rect 20112 16139 20124 16173
rect 20208 16139 20220 16173
rect 20112 16133 20220 16139
rect 20370 16173 20478 16179
rect 20370 16139 20382 16173
rect 20466 16139 20478 16173
rect 20370 16133 20478 16139
rect 20530 16100 20576 16232
rect 20788 17208 20834 17292
rect 20788 16232 20794 17208
rect 20828 16232 20834 17208
rect 20788 16220 20834 16232
rect 21046 17208 21092 17220
rect 21046 16232 21052 17208
rect 21086 16232 21092 17208
rect 20628 16173 20736 16179
rect 20628 16139 20640 16173
rect 20724 16139 20736 16173
rect 20628 16133 20736 16139
rect 20886 16173 20994 16179
rect 20886 16139 20898 16173
rect 20982 16139 20994 16173
rect 20886 16133 20994 16139
rect 21046 16100 21092 16232
rect 21304 17208 21350 17292
rect 21304 16232 21310 17208
rect 21344 16232 21350 17208
rect 21304 16220 21350 16232
rect 21562 17208 21608 17220
rect 21562 16232 21568 17208
rect 21602 16232 21608 17208
rect 21144 16173 21252 16179
rect 21144 16139 21156 16173
rect 21240 16139 21252 16173
rect 21144 16133 21252 16139
rect 21402 16173 21510 16179
rect 21402 16139 21414 16173
rect 21498 16139 21510 16173
rect 21402 16133 21510 16139
rect 21562 16100 21608 16232
rect 21820 17208 21866 17292
rect 21820 16232 21826 17208
rect 21860 16232 21866 17208
rect 21820 16220 21866 16232
rect 22078 17208 22124 17220
rect 22078 16232 22084 17208
rect 22118 16232 22124 17208
rect 21660 16173 21768 16179
rect 21660 16139 21672 16173
rect 21756 16139 21768 16173
rect 21660 16133 21768 16139
rect 21918 16173 22026 16179
rect 21918 16139 21930 16173
rect 22014 16139 22026 16173
rect 21918 16133 22026 16139
rect 22078 16100 22124 16232
rect 22336 17208 22382 17292
rect 22336 16232 22342 17208
rect 22376 16232 22382 17208
rect 22336 16220 22382 16232
rect 22594 17208 22640 17220
rect 22594 16232 22600 17208
rect 22634 16232 22640 17208
rect 22176 16173 22284 16179
rect 22176 16139 22188 16173
rect 22272 16139 22284 16173
rect 22176 16133 22284 16139
rect 22434 16173 22542 16179
rect 22434 16139 22446 16173
rect 22530 16139 22542 16173
rect 22434 16133 22542 16139
rect 22594 16100 22640 16232
rect 22852 17208 22898 17292
rect 22852 16232 22858 17208
rect 22892 16232 22898 17208
rect 22852 16220 22898 16232
rect 23110 17208 23156 17220
rect 23110 16232 23116 17208
rect 23150 16232 23156 17208
rect 22692 16173 22800 16179
rect 22692 16139 22704 16173
rect 22788 16139 22800 16173
rect 22692 16133 22800 16139
rect 22950 16173 23058 16179
rect 22950 16139 22962 16173
rect 23046 16139 23058 16173
rect 22950 16133 23058 16139
rect 23110 16100 23156 16232
rect 23224 17175 23270 17292
rect 23224 16193 23230 17175
rect 23264 16193 23270 17175
rect 23224 16181 23270 16193
rect 11630 16090 17750 16100
rect 11630 16050 17200 16090
rect 17240 16070 17280 16090
rect 17320 16070 17360 16090
rect 17400 16070 17440 16090
rect 17480 16070 17520 16090
rect 17560 16070 17600 16090
rect 17640 16070 17680 16090
rect 17320 16050 17330 16070
rect 11630 16010 17230 16050
rect 17300 16010 17330 16050
rect 11630 15990 17200 16010
rect 11630 15930 11650 15990
rect 11710 15930 11740 15990
rect 11800 15930 11830 15990
rect 11890 15930 11920 15990
rect 11980 15930 12010 15990
rect 12070 15930 12100 15990
rect 12160 15930 12190 15990
rect 12250 15930 12280 15990
rect 12340 15930 12370 15990
rect 12430 15930 12460 15990
rect 12520 15930 12550 15990
rect 12610 15930 12640 15990
rect 12700 15930 12730 15990
rect 12790 15930 12820 15990
rect 12880 15930 12910 15990
rect 12970 15930 13000 15990
rect 13060 15930 13090 15990
rect 13150 15930 13180 15990
rect 13240 15930 13270 15990
rect 13330 15930 13360 15990
rect 13420 15930 13450 15990
rect 13510 15930 13540 15990
rect 13600 15930 13630 15990
rect 13690 15930 13720 15990
rect 13780 15930 13810 15990
rect 13870 15930 13900 15990
rect 13960 15930 13990 15990
rect 14050 15930 14080 15990
rect 14140 15930 14170 15990
rect 14230 15930 14260 15990
rect 14320 15930 14350 15990
rect 14410 15930 14440 15990
rect 14500 15930 14530 15990
rect 14590 15930 14620 15990
rect 14680 15930 14710 15990
rect 14770 15930 14800 15990
rect 14860 15930 14890 15990
rect 14950 15930 14980 15990
rect 15040 15930 15070 15990
rect 15130 15930 15160 15990
rect 15220 15930 15250 15990
rect 15310 15930 15340 15990
rect 15400 15930 15430 15990
rect 15490 15930 15520 15990
rect 15580 15930 15610 15990
rect 15670 15930 15700 15990
rect 15760 15930 15790 15990
rect 15850 15930 15880 15990
rect 15940 15930 15970 15990
rect 16030 15930 16060 15990
rect 16120 15930 16150 15990
rect 16210 15930 16240 15990
rect 16300 15930 16330 15990
rect 16390 15930 16420 15990
rect 16480 15930 16510 15990
rect 16570 15930 16600 15990
rect 16660 15930 16690 15990
rect 16750 15930 16780 15990
rect 16840 15930 16870 15990
rect 16930 15930 16960 15990
rect 17020 15930 17050 15990
rect 17110 15970 17200 15990
rect 17320 15980 17330 16010
rect 17400 15980 17430 16070
rect 17500 16050 17520 16070
rect 17720 16050 17750 16090
rect 17500 16010 17530 16050
rect 17600 16010 17630 16050
rect 17700 16010 17750 16050
rect 17500 15980 17520 16010
rect 17240 15970 17280 15980
rect 17320 15970 17360 15980
rect 17400 15970 17440 15980
rect 17480 15970 17520 15980
rect 17560 15970 17600 15980
rect 17640 15970 17680 15980
rect 17720 15970 17750 16010
rect 17110 15940 17750 15970
rect 17110 15930 17230 15940
rect 17300 15930 17330 15940
rect 11630 15900 17200 15930
rect 11630 15840 11650 15900
rect 11710 15840 11740 15900
rect 11800 15840 11830 15900
rect 11890 15840 11920 15900
rect 11980 15840 12010 15900
rect 12070 15840 12100 15900
rect 12160 15840 12190 15900
rect 12250 15840 12280 15900
rect 12340 15840 12370 15900
rect 12430 15840 12460 15900
rect 12520 15840 12550 15900
rect 12610 15840 12640 15900
rect 12700 15840 12730 15900
rect 12790 15840 12820 15900
rect 12880 15840 12910 15900
rect 12970 15840 13000 15900
rect 13060 15840 13090 15900
rect 13150 15840 13180 15900
rect 13240 15840 13270 15900
rect 13330 15840 13360 15900
rect 13420 15840 13450 15900
rect 13510 15840 13540 15900
rect 13600 15840 13630 15900
rect 13690 15840 13720 15900
rect 13780 15840 13810 15900
rect 13870 15840 13900 15900
rect 13960 15840 13990 15900
rect 14050 15840 14080 15900
rect 14140 15840 14170 15900
rect 14230 15840 14260 15900
rect 14320 15840 14350 15900
rect 14410 15840 14440 15900
rect 14500 15840 14530 15900
rect 14590 15840 14620 15900
rect 14680 15840 14710 15900
rect 14770 15840 14800 15900
rect 14860 15840 14890 15900
rect 14950 15840 14980 15900
rect 15040 15840 15070 15900
rect 15130 15840 15160 15900
rect 15220 15840 15250 15900
rect 15310 15840 15340 15900
rect 15400 15840 15430 15900
rect 15490 15840 15520 15900
rect 15580 15840 15610 15900
rect 15670 15840 15700 15900
rect 15760 15840 15790 15900
rect 15850 15840 15880 15900
rect 15940 15840 15970 15900
rect 16030 15840 16060 15900
rect 16120 15840 16150 15900
rect 16210 15840 16240 15900
rect 16300 15840 16330 15900
rect 16390 15840 16420 15900
rect 16480 15840 16510 15900
rect 16570 15840 16600 15900
rect 16660 15840 16690 15900
rect 16750 15840 16780 15900
rect 16840 15840 16870 15900
rect 16930 15840 16960 15900
rect 17020 15840 17050 15900
rect 17110 15890 17200 15900
rect 17320 15890 17330 15930
rect 17110 15850 17230 15890
rect 17300 15850 17330 15890
rect 17400 15850 17430 15940
rect 17500 15930 17530 15940
rect 17600 15930 17630 15940
rect 17700 15930 17750 15940
rect 17500 15890 17520 15930
rect 17720 15890 17750 15930
rect 17500 15850 17530 15890
rect 17600 15850 17630 15890
rect 17700 15850 17750 15890
rect 17110 15840 17750 15850
rect 11630 15820 17750 15840
rect 17950 15990 23300 16100
rect 17950 15930 18000 15990
rect 18060 15930 18090 15990
rect 18150 15930 18180 15990
rect 18240 15930 18270 15990
rect 18330 15930 18360 15990
rect 18420 15930 18450 15990
rect 18510 15930 18540 15990
rect 18600 15930 18630 15990
rect 18690 15930 18720 15990
rect 18780 15930 18810 15990
rect 18870 15930 18900 15990
rect 18960 15930 18990 15990
rect 19050 15930 19080 15990
rect 19140 15930 19170 15990
rect 19230 15930 19260 15990
rect 19320 15930 19350 15990
rect 19410 15930 19440 15990
rect 19500 15930 19530 15990
rect 19590 15930 19620 15990
rect 19680 15930 19710 15990
rect 19770 15930 19800 15990
rect 19860 15930 19890 15990
rect 19950 15930 19980 15990
rect 20040 15930 20070 15990
rect 20130 15930 20160 15990
rect 20220 15930 20250 15990
rect 20310 15930 20340 15990
rect 20400 15930 20430 15990
rect 20490 15930 20520 15990
rect 20580 15930 20610 15990
rect 20670 15930 20700 15990
rect 20760 15930 20790 15990
rect 20850 15930 20880 15990
rect 20940 15930 20970 15990
rect 21030 15930 21060 15990
rect 21120 15930 21150 15990
rect 21210 15930 21240 15990
rect 21300 15930 21330 15990
rect 21390 15930 21420 15990
rect 21480 15930 21510 15990
rect 21570 15930 21600 15990
rect 21660 15930 21690 15990
rect 21750 15930 21780 15990
rect 21840 15930 21870 15990
rect 21930 15930 21960 15990
rect 22020 15930 22050 15990
rect 22110 15930 22140 15990
rect 22200 15930 22230 15990
rect 22290 15930 22320 15990
rect 22380 15930 22410 15990
rect 22470 15930 22500 15990
rect 22560 15930 22590 15990
rect 22650 15930 22680 15990
rect 22740 15930 22770 15990
rect 22830 15930 22860 15990
rect 22920 15930 22950 15990
rect 23010 15930 23040 15990
rect 23100 15930 23130 15990
rect 23190 15930 23220 15990
rect 23280 15930 23300 15990
rect 17950 15900 23300 15930
rect 17950 15840 18000 15900
rect 18060 15840 18090 15900
rect 18150 15840 18180 15900
rect 18240 15840 18270 15900
rect 18330 15840 18360 15900
rect 18420 15840 18450 15900
rect 18510 15840 18540 15900
rect 18600 15840 18630 15900
rect 18690 15840 18720 15900
rect 18780 15840 18810 15900
rect 18870 15840 18900 15900
rect 18960 15840 18990 15900
rect 19050 15840 19080 15900
rect 19140 15840 19170 15900
rect 19230 15840 19260 15900
rect 19320 15840 19350 15900
rect 19410 15840 19440 15900
rect 19500 15840 19530 15900
rect 19590 15840 19620 15900
rect 19680 15840 19710 15900
rect 19770 15840 19800 15900
rect 19860 15840 19890 15900
rect 19950 15840 19980 15900
rect 20040 15840 20070 15900
rect 20130 15840 20160 15900
rect 20220 15840 20250 15900
rect 20310 15840 20340 15900
rect 20400 15840 20430 15900
rect 20490 15840 20520 15900
rect 20580 15840 20610 15900
rect 20670 15840 20700 15900
rect 20760 15840 20790 15900
rect 20850 15840 20880 15900
rect 20940 15840 20970 15900
rect 21030 15840 21060 15900
rect 21120 15840 21150 15900
rect 21210 15840 21240 15900
rect 21300 15840 21330 15900
rect 21390 15840 21420 15900
rect 21480 15840 21510 15900
rect 21570 15840 21600 15900
rect 21660 15840 21690 15900
rect 21750 15840 21780 15900
rect 21840 15840 21870 15900
rect 21930 15840 21960 15900
rect 22020 15840 22050 15900
rect 22110 15840 22140 15900
rect 22200 15840 22230 15900
rect 22290 15840 22320 15900
rect 22380 15840 22410 15900
rect 22470 15840 22500 15900
rect 22560 15840 22590 15900
rect 22650 15840 22680 15900
rect 22740 15840 22770 15900
rect 22830 15840 22860 15900
rect 22920 15840 22950 15900
rect 23010 15840 23040 15900
rect 23100 15840 23130 15900
rect 23190 15840 23220 15900
rect 23280 15840 23300 15900
rect 17950 15820 23300 15840
rect 11630 13860 16980 13880
rect 11630 13800 11650 13860
rect 11710 13800 11740 13860
rect 11800 13800 11830 13860
rect 11890 13800 11920 13860
rect 11980 13800 12010 13860
rect 12070 13800 12100 13860
rect 12160 13800 12190 13860
rect 12250 13800 12280 13860
rect 12340 13800 12370 13860
rect 12430 13800 12460 13860
rect 12520 13800 12550 13860
rect 12610 13800 12640 13860
rect 12700 13800 12730 13860
rect 12790 13800 12820 13860
rect 12880 13800 12910 13860
rect 12970 13800 13000 13860
rect 13060 13800 13090 13860
rect 13150 13800 13180 13860
rect 13240 13800 13270 13860
rect 13330 13800 13360 13860
rect 13420 13800 13450 13860
rect 13510 13800 13540 13860
rect 13600 13800 13630 13860
rect 13690 13800 13720 13860
rect 13780 13800 13810 13860
rect 13870 13800 13900 13860
rect 13960 13800 13990 13860
rect 14050 13800 14080 13860
rect 14140 13800 14170 13860
rect 14230 13800 14260 13860
rect 14320 13800 14350 13860
rect 14410 13800 14440 13860
rect 14500 13800 14530 13860
rect 14590 13800 14620 13860
rect 14680 13800 14710 13860
rect 14770 13800 14800 13860
rect 14860 13800 14890 13860
rect 14950 13800 14980 13860
rect 15040 13800 15070 13860
rect 15130 13800 15160 13860
rect 15220 13800 15250 13860
rect 15310 13800 15340 13860
rect 15400 13800 15430 13860
rect 15490 13800 15520 13860
rect 15580 13800 15610 13860
rect 15670 13800 15700 13860
rect 15760 13800 15790 13860
rect 15850 13800 15880 13860
rect 15940 13800 15970 13860
rect 16030 13800 16060 13860
rect 16120 13800 16150 13860
rect 16210 13800 16240 13860
rect 16300 13800 16330 13860
rect 16390 13800 16420 13860
rect 16480 13800 16510 13860
rect 16570 13800 16600 13860
rect 16660 13800 16690 13860
rect 16750 13800 16780 13860
rect 16840 13800 16870 13860
rect 16930 13800 16980 13860
rect 11630 13770 16980 13800
rect 11630 13710 11650 13770
rect 11710 13710 11740 13770
rect 11800 13710 11830 13770
rect 11890 13710 11920 13770
rect 11980 13710 12010 13770
rect 12070 13710 12100 13770
rect 12160 13710 12190 13770
rect 12250 13710 12280 13770
rect 12340 13710 12370 13770
rect 12430 13710 12460 13770
rect 12520 13710 12550 13770
rect 12610 13710 12640 13770
rect 12700 13710 12730 13770
rect 12790 13710 12820 13770
rect 12880 13710 12910 13770
rect 12970 13710 13000 13770
rect 13060 13710 13090 13770
rect 13150 13710 13180 13770
rect 13240 13710 13270 13770
rect 13330 13710 13360 13770
rect 13420 13710 13450 13770
rect 13510 13710 13540 13770
rect 13600 13710 13630 13770
rect 13690 13710 13720 13770
rect 13780 13710 13810 13770
rect 13870 13710 13900 13770
rect 13960 13710 13990 13770
rect 14050 13710 14080 13770
rect 14140 13710 14170 13770
rect 14230 13710 14260 13770
rect 14320 13710 14350 13770
rect 14410 13710 14440 13770
rect 14500 13710 14530 13770
rect 14590 13710 14620 13770
rect 14680 13710 14710 13770
rect 14770 13710 14800 13770
rect 14860 13710 14890 13770
rect 14950 13710 14980 13770
rect 15040 13710 15070 13770
rect 15130 13710 15160 13770
rect 15220 13710 15250 13770
rect 15310 13710 15340 13770
rect 15400 13710 15430 13770
rect 15490 13710 15520 13770
rect 15580 13710 15610 13770
rect 15670 13710 15700 13770
rect 15760 13710 15790 13770
rect 15850 13710 15880 13770
rect 15940 13710 15970 13770
rect 16030 13710 16060 13770
rect 16120 13710 16150 13770
rect 16210 13710 16240 13770
rect 16300 13710 16330 13770
rect 16390 13710 16420 13770
rect 16480 13710 16510 13770
rect 16570 13710 16600 13770
rect 16660 13710 16690 13770
rect 16750 13710 16780 13770
rect 16840 13710 16870 13770
rect 16930 13710 16980 13770
rect 11630 13600 16980 13710
rect 17180 13860 23300 13880
rect 17180 13850 17820 13860
rect 17180 13820 17230 13850
rect 17300 13820 17330 13850
rect 17180 13780 17200 13820
rect 17320 13780 17330 13820
rect 17180 13760 17230 13780
rect 17300 13760 17330 13780
rect 17400 13760 17430 13850
rect 17500 13820 17530 13850
rect 17600 13820 17630 13850
rect 17700 13820 17820 13850
rect 17500 13780 17520 13820
rect 17720 13800 17820 13820
rect 17880 13800 17910 13860
rect 17970 13800 18000 13860
rect 18060 13800 18090 13860
rect 18150 13800 18180 13860
rect 18240 13800 18270 13860
rect 18330 13800 18360 13860
rect 18420 13800 18450 13860
rect 18510 13800 18540 13860
rect 18600 13800 18630 13860
rect 18690 13800 18720 13860
rect 18780 13800 18810 13860
rect 18870 13800 18900 13860
rect 18960 13800 18990 13860
rect 19050 13800 19080 13860
rect 19140 13800 19170 13860
rect 19230 13800 19260 13860
rect 19320 13800 19350 13860
rect 19410 13800 19440 13860
rect 19500 13800 19530 13860
rect 19590 13800 19620 13860
rect 19680 13800 19710 13860
rect 19770 13800 19800 13860
rect 19860 13800 19890 13860
rect 19950 13800 19980 13860
rect 20040 13800 20070 13860
rect 20130 13800 20160 13860
rect 20220 13800 20250 13860
rect 20310 13800 20340 13860
rect 20400 13800 20430 13860
rect 20490 13800 20520 13860
rect 20580 13800 20610 13860
rect 20670 13800 20700 13860
rect 20760 13800 20790 13860
rect 20850 13800 20880 13860
rect 20940 13800 20970 13860
rect 21030 13800 21060 13860
rect 21120 13800 21150 13860
rect 21210 13800 21240 13860
rect 21300 13800 21330 13860
rect 21390 13800 21420 13860
rect 21480 13800 21510 13860
rect 21570 13800 21600 13860
rect 21660 13800 21690 13860
rect 21750 13800 21780 13860
rect 21840 13800 21870 13860
rect 21930 13800 21960 13860
rect 22020 13800 22050 13860
rect 22110 13800 22140 13860
rect 22200 13800 22230 13860
rect 22290 13800 22320 13860
rect 22380 13800 22410 13860
rect 22470 13800 22500 13860
rect 22560 13800 22590 13860
rect 22650 13800 22680 13860
rect 22740 13800 22770 13860
rect 22830 13800 22860 13860
rect 22920 13800 22950 13860
rect 23010 13800 23040 13860
rect 23100 13800 23130 13860
rect 23190 13800 23220 13860
rect 23280 13800 23300 13860
rect 17720 13780 23300 13800
rect 17500 13760 17530 13780
rect 17600 13760 17630 13780
rect 17700 13770 23300 13780
rect 17700 13760 17820 13770
rect 17180 13740 17820 13760
rect 17180 13700 17200 13740
rect 17240 13720 17280 13740
rect 17320 13720 17360 13740
rect 17400 13720 17440 13740
rect 17480 13720 17520 13740
rect 17560 13720 17600 13740
rect 17640 13720 17680 13740
rect 17320 13700 17330 13720
rect 17180 13660 17230 13700
rect 17300 13660 17330 13700
rect 17180 13620 17200 13660
rect 17320 13630 17330 13660
rect 17400 13630 17430 13720
rect 17500 13700 17520 13720
rect 17720 13710 17820 13740
rect 17880 13710 17910 13770
rect 17970 13710 18000 13770
rect 18060 13710 18090 13770
rect 18150 13710 18180 13770
rect 18240 13710 18270 13770
rect 18330 13710 18360 13770
rect 18420 13710 18450 13770
rect 18510 13710 18540 13770
rect 18600 13710 18630 13770
rect 18690 13710 18720 13770
rect 18780 13710 18810 13770
rect 18870 13710 18900 13770
rect 18960 13710 18990 13770
rect 19050 13710 19080 13770
rect 19140 13710 19170 13770
rect 19230 13710 19260 13770
rect 19320 13710 19350 13770
rect 19410 13710 19440 13770
rect 19500 13710 19530 13770
rect 19590 13710 19620 13770
rect 19680 13710 19710 13770
rect 19770 13710 19800 13770
rect 19860 13710 19890 13770
rect 19950 13710 19980 13770
rect 20040 13710 20070 13770
rect 20130 13710 20160 13770
rect 20220 13710 20250 13770
rect 20310 13710 20340 13770
rect 20400 13710 20430 13770
rect 20490 13710 20520 13770
rect 20580 13710 20610 13770
rect 20670 13710 20700 13770
rect 20760 13710 20790 13770
rect 20850 13710 20880 13770
rect 20940 13710 20970 13770
rect 21030 13710 21060 13770
rect 21120 13710 21150 13770
rect 21210 13710 21240 13770
rect 21300 13710 21330 13770
rect 21390 13710 21420 13770
rect 21480 13710 21510 13770
rect 21570 13710 21600 13770
rect 21660 13710 21690 13770
rect 21750 13710 21780 13770
rect 21840 13710 21870 13770
rect 21930 13710 21960 13770
rect 22020 13710 22050 13770
rect 22110 13710 22140 13770
rect 22200 13710 22230 13770
rect 22290 13710 22320 13770
rect 22380 13710 22410 13770
rect 22470 13710 22500 13770
rect 22560 13710 22590 13770
rect 22650 13710 22680 13770
rect 22740 13710 22770 13770
rect 22830 13710 22860 13770
rect 22920 13710 22950 13770
rect 23010 13710 23040 13770
rect 23100 13710 23130 13770
rect 23190 13710 23220 13770
rect 23280 13710 23300 13770
rect 17720 13700 23300 13710
rect 17500 13660 17530 13700
rect 17600 13660 17630 13700
rect 17700 13660 23300 13700
rect 17500 13630 17520 13660
rect 17240 13620 17280 13630
rect 17320 13620 17360 13630
rect 17400 13620 17440 13630
rect 17480 13620 17520 13630
rect 17560 13620 17600 13630
rect 17640 13620 17680 13630
rect 17720 13620 23300 13660
rect 17180 13600 23300 13620
rect 11660 13479 11706 13491
rect 11660 12505 11666 13479
rect 11700 12505 11706 13479
rect 11660 12423 11706 12505
rect 11774 13449 11820 13600
rect 11872 13533 11980 13539
rect 11872 13499 11884 13533
rect 11968 13499 11980 13533
rect 11872 13493 11980 13499
rect 12130 13533 12238 13539
rect 12130 13499 12142 13533
rect 12226 13499 12238 13533
rect 12130 13493 12238 13499
rect 11774 12473 11780 13449
rect 11814 12473 11820 13449
rect 11774 12461 11820 12473
rect 12032 13449 12078 13461
rect 12032 12473 12038 13449
rect 12072 12473 12078 13449
rect 12032 12461 12078 12473
rect 12290 13449 12336 13600
rect 12388 13533 12496 13539
rect 12388 13499 12400 13533
rect 12484 13499 12496 13533
rect 12388 13493 12496 13499
rect 12646 13533 12754 13539
rect 12646 13499 12658 13533
rect 12742 13499 12754 13533
rect 12646 13493 12754 13499
rect 12290 12473 12296 13449
rect 12330 12473 12336 13449
rect 12290 12461 12336 12473
rect 12548 13449 12594 13461
rect 12548 12473 12554 13449
rect 12588 12473 12594 13449
rect 12548 12461 12594 12473
rect 12806 13449 12852 13600
rect 12904 13533 13012 13539
rect 12904 13499 12916 13533
rect 13000 13499 13012 13533
rect 12904 13493 13012 13499
rect 13162 13533 13270 13539
rect 13162 13499 13174 13533
rect 13258 13499 13270 13533
rect 13162 13493 13270 13499
rect 12806 12473 12812 13449
rect 12846 12473 12852 13449
rect 12806 12461 12852 12473
rect 13064 13449 13110 13461
rect 13064 12473 13070 13449
rect 13104 12473 13110 13449
rect 13064 12461 13110 12473
rect 13322 13449 13368 13600
rect 13420 13533 13528 13539
rect 13420 13499 13432 13533
rect 13516 13499 13528 13533
rect 13420 13493 13528 13499
rect 13678 13533 13786 13539
rect 13678 13499 13690 13533
rect 13774 13499 13786 13533
rect 13678 13493 13786 13499
rect 13322 12473 13328 13449
rect 13362 12473 13368 13449
rect 13322 12461 13368 12473
rect 13580 13449 13626 13461
rect 13580 12473 13586 13449
rect 13620 12473 13626 13449
rect 13580 12461 13626 12473
rect 13838 13449 13884 13600
rect 13936 13533 14044 13539
rect 13936 13499 13948 13533
rect 14032 13499 14044 13533
rect 13936 13493 14044 13499
rect 14194 13533 14302 13539
rect 14194 13499 14206 13533
rect 14290 13499 14302 13533
rect 14194 13493 14302 13499
rect 13838 12473 13844 13449
rect 13878 12473 13884 13449
rect 13838 12461 13884 12473
rect 14096 13449 14142 13461
rect 14096 12473 14102 13449
rect 14136 12473 14142 13449
rect 14096 12461 14142 12473
rect 14354 13449 14400 13600
rect 14452 13533 14560 13539
rect 14452 13499 14464 13533
rect 14548 13499 14560 13533
rect 14452 13493 14560 13499
rect 14710 13533 14818 13539
rect 14710 13499 14722 13533
rect 14806 13499 14818 13533
rect 14710 13493 14818 13499
rect 14354 12473 14360 13449
rect 14394 12473 14400 13449
rect 14354 12461 14400 12473
rect 14612 13449 14658 13461
rect 14612 12473 14618 13449
rect 14652 12473 14658 13449
rect 14612 12461 14658 12473
rect 14870 13449 14916 13600
rect 14968 13533 15076 13539
rect 14968 13499 14980 13533
rect 15064 13499 15076 13533
rect 14968 13493 15076 13499
rect 15226 13533 15334 13539
rect 15226 13499 15238 13533
rect 15322 13499 15334 13533
rect 15226 13493 15334 13499
rect 14870 12473 14876 13449
rect 14910 12473 14916 13449
rect 14870 12461 14916 12473
rect 15128 13449 15174 13461
rect 15128 12473 15134 13449
rect 15168 12473 15174 13449
rect 15128 12461 15174 12473
rect 15386 13449 15432 13600
rect 15484 13533 15592 13539
rect 15484 13499 15496 13533
rect 15580 13499 15592 13533
rect 15484 13493 15592 13499
rect 15742 13533 15850 13539
rect 15742 13499 15754 13533
rect 15838 13499 15850 13533
rect 15742 13493 15850 13499
rect 15386 12473 15392 13449
rect 15426 12473 15432 13449
rect 15386 12461 15432 12473
rect 15644 13449 15690 13461
rect 15644 12473 15650 13449
rect 15684 12473 15690 13449
rect 15644 12461 15690 12473
rect 15902 13449 15948 13600
rect 16000 13533 16108 13539
rect 16000 13499 16012 13533
rect 16096 13499 16108 13533
rect 16000 13493 16108 13499
rect 16258 13533 16366 13539
rect 16258 13499 16270 13533
rect 16354 13499 16366 13533
rect 16258 13493 16366 13499
rect 15902 12473 15908 13449
rect 15942 12473 15948 13449
rect 15902 12461 15948 12473
rect 16160 13449 16206 13461
rect 16160 12473 16166 13449
rect 16200 12473 16206 13449
rect 16160 12461 16206 12473
rect 16418 13449 16464 13600
rect 16516 13533 16624 13539
rect 16516 13499 16528 13533
rect 16612 13499 16624 13533
rect 16516 13493 16624 13499
rect 16774 13533 16882 13539
rect 16774 13499 16786 13533
rect 16870 13499 16882 13533
rect 16774 13493 16882 13499
rect 16418 12473 16424 13449
rect 16458 12473 16464 13449
rect 16418 12461 16464 12473
rect 16676 13449 16722 13461
rect 16676 12473 16682 13449
rect 16716 12473 16722 13449
rect 16676 12461 16722 12473
rect 16934 13449 16980 13600
rect 16934 12473 16940 13449
rect 16974 12473 16980 13449
rect 16934 12461 16980 12473
rect 17048 13479 17094 13491
rect 17048 12505 17054 13479
rect 17088 12505 17094 13479
rect 12038 12423 12072 12461
rect 12554 12423 12588 12461
rect 13070 12423 13104 12461
rect 13586 12423 13620 12461
rect 14102 12423 14136 12461
rect 14618 12423 14652 12461
rect 15134 12423 15168 12461
rect 15650 12423 15684 12461
rect 16166 12423 16200 12461
rect 16682 12423 16716 12461
rect 17048 12423 17094 12505
rect 11660 12383 17094 12423
rect 11660 12349 11700 12383
rect 17054 12349 17094 12383
rect 11660 12310 17094 12349
rect 11660 12240 11690 12310
rect 11760 12240 11810 12310
rect 11880 12240 12020 12310
rect 12090 12240 12140 12310
rect 12210 12240 12350 12310
rect 12420 12240 12470 12310
rect 12540 12240 12680 12310
rect 12750 12240 12800 12310
rect 12870 12240 13010 12310
rect 13080 12240 13130 12310
rect 13200 12240 13340 12310
rect 13410 12240 13460 12310
rect 13530 12240 13670 12310
rect 13740 12240 13790 12310
rect 13860 12240 14000 12310
rect 14070 12240 14120 12310
rect 14190 12240 14330 12310
rect 14400 12240 14450 12310
rect 14520 12300 15650 12310
rect 14520 12240 14660 12300
rect 11660 12230 14660 12240
rect 14730 12230 14780 12300
rect 14850 12230 14990 12300
rect 15060 12230 15110 12300
rect 15180 12230 15320 12300
rect 15390 12230 15440 12300
rect 15510 12240 15650 12300
rect 15720 12240 15770 12310
rect 15840 12240 15980 12310
rect 16050 12240 16100 12310
rect 16170 12240 16310 12310
rect 16380 12240 16430 12310
rect 16500 12240 16640 12310
rect 16710 12240 16760 12310
rect 16830 12240 17094 12310
rect 15510 12230 17094 12240
rect 11660 12190 17094 12230
rect 11660 12120 11690 12190
rect 11760 12120 11810 12190
rect 11880 12120 12020 12190
rect 12090 12120 12140 12190
rect 12210 12120 12350 12190
rect 12420 12120 12470 12190
rect 12540 12120 12680 12190
rect 12750 12120 12800 12190
rect 12870 12120 13010 12190
rect 13080 12120 13130 12190
rect 13200 12120 13340 12190
rect 13410 12120 13460 12190
rect 13530 12120 13670 12190
rect 13740 12120 13790 12190
rect 13860 12120 14000 12190
rect 14070 12120 14120 12190
rect 14190 12120 14330 12190
rect 14400 12120 14450 12190
rect 14520 12180 15650 12190
rect 14520 12120 14660 12180
rect 11660 12110 14660 12120
rect 14730 12110 14780 12180
rect 14850 12110 14990 12180
rect 15060 12110 15110 12180
rect 15180 12110 15320 12180
rect 15390 12110 15440 12180
rect 15510 12120 15650 12180
rect 15720 12120 15770 12190
rect 15840 12120 15980 12190
rect 16050 12120 16100 12190
rect 16170 12120 16310 12190
rect 16380 12120 16430 12190
rect 16500 12120 16640 12190
rect 16710 12120 16760 12190
rect 16830 12130 17094 12190
rect 17836 13479 17882 13491
rect 17836 12505 17842 13479
rect 17876 12505 17882 13479
rect 17836 12423 17882 12505
rect 17950 13449 17996 13600
rect 18048 13533 18156 13539
rect 18048 13499 18060 13533
rect 18144 13499 18156 13533
rect 18048 13493 18156 13499
rect 18306 13533 18414 13539
rect 18306 13499 18318 13533
rect 18402 13499 18414 13533
rect 18306 13493 18414 13499
rect 17950 12473 17956 13449
rect 17990 12473 17996 13449
rect 17950 12461 17996 12473
rect 18208 13449 18254 13461
rect 18208 12473 18214 13449
rect 18248 12473 18254 13449
rect 18208 12461 18254 12473
rect 18466 13449 18512 13600
rect 18564 13533 18672 13539
rect 18564 13499 18576 13533
rect 18660 13499 18672 13533
rect 18564 13493 18672 13499
rect 18822 13533 18930 13539
rect 18822 13499 18834 13533
rect 18918 13499 18930 13533
rect 18822 13493 18930 13499
rect 18466 12473 18472 13449
rect 18506 12473 18512 13449
rect 18466 12461 18512 12473
rect 18724 13449 18770 13461
rect 18724 12473 18730 13449
rect 18764 12473 18770 13449
rect 18724 12461 18770 12473
rect 18982 13449 19028 13600
rect 19080 13533 19188 13539
rect 19080 13499 19092 13533
rect 19176 13499 19188 13533
rect 19080 13493 19188 13499
rect 19338 13533 19446 13539
rect 19338 13499 19350 13533
rect 19434 13499 19446 13533
rect 19338 13493 19446 13499
rect 18982 12473 18988 13449
rect 19022 12473 19028 13449
rect 18982 12461 19028 12473
rect 19240 13449 19286 13461
rect 19240 12473 19246 13449
rect 19280 12473 19286 13449
rect 19240 12461 19286 12473
rect 19498 13449 19544 13600
rect 19596 13533 19704 13539
rect 19596 13499 19608 13533
rect 19692 13499 19704 13533
rect 19596 13493 19704 13499
rect 19854 13533 19962 13539
rect 19854 13499 19866 13533
rect 19950 13499 19962 13533
rect 19854 13493 19962 13499
rect 19498 12473 19504 13449
rect 19538 12473 19544 13449
rect 19498 12461 19544 12473
rect 19756 13449 19802 13461
rect 19756 12473 19762 13449
rect 19796 12473 19802 13449
rect 19756 12461 19802 12473
rect 20014 13449 20060 13600
rect 20112 13533 20220 13539
rect 20112 13499 20124 13533
rect 20208 13499 20220 13533
rect 20112 13493 20220 13499
rect 20370 13533 20478 13539
rect 20370 13499 20382 13533
rect 20466 13499 20478 13533
rect 20370 13493 20478 13499
rect 20014 12473 20020 13449
rect 20054 12473 20060 13449
rect 20014 12461 20060 12473
rect 20272 13449 20318 13461
rect 20272 12473 20278 13449
rect 20312 12473 20318 13449
rect 20272 12461 20318 12473
rect 20530 13449 20576 13600
rect 20628 13533 20736 13539
rect 20628 13499 20640 13533
rect 20724 13499 20736 13533
rect 20628 13493 20736 13499
rect 20886 13533 20994 13539
rect 20886 13499 20898 13533
rect 20982 13499 20994 13533
rect 20886 13493 20994 13499
rect 20530 12473 20536 13449
rect 20570 12473 20576 13449
rect 20530 12461 20576 12473
rect 20788 13449 20834 13461
rect 20788 12473 20794 13449
rect 20828 12473 20834 13449
rect 20788 12461 20834 12473
rect 21046 13449 21092 13600
rect 21144 13533 21252 13539
rect 21144 13499 21156 13533
rect 21240 13499 21252 13533
rect 21144 13493 21252 13499
rect 21402 13533 21510 13539
rect 21402 13499 21414 13533
rect 21498 13499 21510 13533
rect 21402 13493 21510 13499
rect 21046 12473 21052 13449
rect 21086 12473 21092 13449
rect 21046 12461 21092 12473
rect 21304 13449 21350 13461
rect 21304 12473 21310 13449
rect 21344 12473 21350 13449
rect 21304 12461 21350 12473
rect 21562 13449 21608 13600
rect 21660 13533 21768 13539
rect 21660 13499 21672 13533
rect 21756 13499 21768 13533
rect 21660 13493 21768 13499
rect 21918 13533 22026 13539
rect 21918 13499 21930 13533
rect 22014 13499 22026 13533
rect 21918 13493 22026 13499
rect 21562 12473 21568 13449
rect 21602 12473 21608 13449
rect 21562 12461 21608 12473
rect 21820 13449 21866 13461
rect 21820 12473 21826 13449
rect 21860 12473 21866 13449
rect 21820 12461 21866 12473
rect 22078 13449 22124 13600
rect 22176 13533 22284 13539
rect 22176 13499 22188 13533
rect 22272 13499 22284 13533
rect 22176 13493 22284 13499
rect 22434 13533 22542 13539
rect 22434 13499 22446 13533
rect 22530 13499 22542 13533
rect 22434 13493 22542 13499
rect 22078 12473 22084 13449
rect 22118 12473 22124 13449
rect 22078 12461 22124 12473
rect 22336 13449 22382 13461
rect 22336 12473 22342 13449
rect 22376 12473 22382 13449
rect 22336 12461 22382 12473
rect 22594 13449 22640 13600
rect 22692 13533 22800 13539
rect 22692 13499 22704 13533
rect 22788 13499 22800 13533
rect 22692 13493 22800 13499
rect 22950 13533 23058 13539
rect 22950 13499 22962 13533
rect 23046 13499 23058 13533
rect 22950 13493 23058 13499
rect 22594 12473 22600 13449
rect 22634 12473 22640 13449
rect 22594 12461 22640 12473
rect 22852 13449 22898 13461
rect 22852 12473 22858 13449
rect 22892 12473 22898 13449
rect 22852 12461 22898 12473
rect 23110 13449 23156 13600
rect 23110 12473 23116 13449
rect 23150 12473 23156 13449
rect 23110 12461 23156 12473
rect 23224 13479 23270 13491
rect 23224 12505 23230 13479
rect 23264 12505 23270 13479
rect 18214 12423 18248 12461
rect 18730 12423 18764 12461
rect 19246 12423 19280 12461
rect 19762 12423 19796 12461
rect 20278 12423 20312 12461
rect 20794 12423 20828 12461
rect 21310 12423 21344 12461
rect 21826 12423 21860 12461
rect 22342 12423 22376 12461
rect 22858 12423 22892 12461
rect 23224 12423 23270 12505
rect 17836 12383 23270 12423
rect 17836 12349 17876 12383
rect 23230 12349 23270 12383
rect 17836 12310 23270 12349
rect 17836 12240 18100 12310
rect 18170 12240 18220 12310
rect 18290 12240 18430 12310
rect 18500 12240 18550 12310
rect 18620 12240 18760 12310
rect 18830 12240 18880 12310
rect 18950 12240 19090 12310
rect 19160 12240 19210 12310
rect 19280 12300 20410 12310
rect 19280 12240 19420 12300
rect 17836 12230 19420 12240
rect 19490 12230 19540 12300
rect 19610 12230 19750 12300
rect 19820 12230 19870 12300
rect 19940 12230 20080 12300
rect 20150 12230 20200 12300
rect 20270 12240 20410 12300
rect 20480 12240 20530 12310
rect 20600 12240 20740 12310
rect 20810 12240 20860 12310
rect 20930 12240 21070 12310
rect 21140 12240 21190 12310
rect 21260 12240 21400 12310
rect 21470 12240 21520 12310
rect 21590 12240 21730 12310
rect 21800 12240 21850 12310
rect 21920 12240 22060 12310
rect 22130 12240 22180 12310
rect 22250 12240 22390 12310
rect 22460 12240 22510 12310
rect 22580 12240 22720 12310
rect 22790 12240 22840 12310
rect 22910 12240 23050 12310
rect 23120 12240 23170 12310
rect 23240 12240 23270 12310
rect 20270 12230 23270 12240
rect 17836 12190 23270 12230
rect 17836 12130 18100 12190
rect 16830 12120 17090 12130
rect 15510 12110 17090 12120
rect 11660 12090 17090 12110
rect 17840 12120 18100 12130
rect 18170 12120 18220 12190
rect 18290 12120 18430 12190
rect 18500 12120 18550 12190
rect 18620 12120 18760 12190
rect 18830 12120 18880 12190
rect 18950 12120 19090 12190
rect 19160 12120 19210 12190
rect 19280 12180 20410 12190
rect 19280 12120 19420 12180
rect 17840 12110 19420 12120
rect 19490 12110 19540 12180
rect 19610 12110 19750 12180
rect 19820 12110 19870 12180
rect 19940 12110 20080 12180
rect 20150 12110 20200 12180
rect 20270 12120 20410 12180
rect 20480 12120 20530 12190
rect 20600 12120 20740 12190
rect 20810 12120 20860 12190
rect 20930 12120 21070 12190
rect 21140 12120 21190 12190
rect 21260 12120 21400 12190
rect 21470 12120 21520 12190
rect 21590 12120 21730 12190
rect 21800 12120 21850 12190
rect 21920 12120 22060 12190
rect 22130 12120 22180 12190
rect 22250 12120 22390 12190
rect 22460 12120 22510 12190
rect 22580 12120 22720 12190
rect 22790 12120 22840 12190
rect 22910 12120 23050 12190
rect 23120 12120 23170 12190
rect 23240 12120 23270 12190
rect 20270 12110 23270 12120
rect 17840 12090 23270 12110
rect 11690 12070 11930 12090
rect 12020 12070 12260 12090
rect 12350 12070 12590 12090
rect 12680 12070 12920 12090
rect 13010 12070 13250 12090
rect 13340 12070 13580 12090
rect 13670 12070 13910 12090
rect 14000 12070 14240 12090
rect 14330 12070 14570 12090
rect 14660 12070 14900 12090
rect 14990 12070 15230 12090
rect 15320 12070 15560 12090
rect 15650 12070 15890 12090
rect 15980 12070 16220 12090
rect 16310 12070 16550 12090
rect 16640 12070 16880 12090
rect 18050 12070 18290 12090
rect 18380 12070 18620 12090
rect 18710 12070 18950 12090
rect 19040 12070 19280 12090
rect 19370 12070 19610 12090
rect 19700 12070 19940 12090
rect 20030 12070 20270 12090
rect 20360 12070 20600 12090
rect 20690 12070 20930 12090
rect 21020 12070 21260 12090
rect 21350 12070 21590 12090
rect 21680 12070 21920 12090
rect 22010 12070 22250 12090
rect 22340 12070 22580 12090
rect 22670 12070 22910 12090
rect 23000 12070 23240 12090
<< via1 >>
rect 11690 17490 11760 17560
rect 11810 17490 11880 17560
rect 12020 17490 12090 17560
rect 12140 17490 12210 17560
rect 12350 17490 12420 17560
rect 12470 17490 12540 17560
rect 12680 17490 12750 17560
rect 12800 17490 12870 17560
rect 13010 17490 13080 17560
rect 13130 17490 13200 17560
rect 13340 17490 13410 17560
rect 13460 17490 13530 17560
rect 13670 17490 13740 17560
rect 13790 17490 13860 17560
rect 14000 17490 14070 17560
rect 14120 17490 14190 17560
rect 14330 17490 14400 17560
rect 14450 17490 14520 17560
rect 14660 17500 14730 17570
rect 14780 17500 14850 17570
rect 14990 17500 15060 17570
rect 15110 17500 15180 17570
rect 15320 17500 15390 17570
rect 15440 17500 15510 17570
rect 15650 17490 15720 17560
rect 15770 17490 15840 17560
rect 15980 17490 16050 17560
rect 16100 17490 16170 17560
rect 16310 17490 16380 17560
rect 16430 17490 16500 17560
rect 16640 17490 16710 17560
rect 16760 17490 16830 17560
rect 11690 17370 11760 17440
rect 11810 17370 11880 17440
rect 12020 17370 12090 17440
rect 12140 17370 12210 17440
rect 12350 17370 12420 17440
rect 12470 17370 12540 17440
rect 12680 17370 12750 17440
rect 12800 17370 12870 17440
rect 13010 17370 13080 17440
rect 13130 17370 13200 17440
rect 13340 17370 13410 17440
rect 13460 17370 13530 17440
rect 13670 17370 13740 17440
rect 13790 17370 13860 17440
rect 14000 17370 14070 17440
rect 14120 17370 14190 17440
rect 14330 17370 14400 17440
rect 14450 17370 14520 17440
rect 14660 17380 14730 17450
rect 14780 17380 14850 17450
rect 14990 17380 15060 17450
rect 15110 17380 15180 17450
rect 15320 17380 15390 17450
rect 15440 17380 15510 17450
rect 15650 17370 15720 17440
rect 15770 17370 15840 17440
rect 15980 17370 16050 17440
rect 16100 17370 16170 17440
rect 16310 17370 16380 17440
rect 16430 17370 16500 17440
rect 16640 17370 16710 17440
rect 16760 17370 16830 17440
rect 18100 17490 18170 17560
rect 18220 17490 18290 17560
rect 18430 17490 18500 17560
rect 18550 17490 18620 17560
rect 18760 17490 18830 17560
rect 18880 17490 18950 17560
rect 19090 17490 19160 17560
rect 19210 17490 19280 17560
rect 19420 17500 19490 17570
rect 19540 17500 19610 17570
rect 19750 17500 19820 17570
rect 19870 17500 19940 17570
rect 20080 17500 20150 17570
rect 20200 17500 20270 17570
rect 20410 17490 20480 17560
rect 20530 17490 20600 17560
rect 20740 17490 20810 17560
rect 20860 17490 20930 17560
rect 21070 17490 21140 17560
rect 21190 17490 21260 17560
rect 21400 17490 21470 17560
rect 21520 17490 21590 17560
rect 21730 17490 21800 17560
rect 21850 17490 21920 17560
rect 22060 17490 22130 17560
rect 22180 17490 22250 17560
rect 22390 17490 22460 17560
rect 22510 17490 22580 17560
rect 22720 17490 22790 17560
rect 22840 17490 22910 17560
rect 23050 17490 23120 17560
rect 23170 17490 23240 17560
rect 18100 17370 18170 17440
rect 18220 17370 18290 17440
rect 18430 17370 18500 17440
rect 18550 17370 18620 17440
rect 18760 17370 18830 17440
rect 18880 17370 18950 17440
rect 19090 17370 19160 17440
rect 19210 17370 19280 17440
rect 19420 17380 19490 17450
rect 19540 17380 19610 17450
rect 19750 17380 19820 17450
rect 19870 17380 19940 17450
rect 20080 17380 20150 17450
rect 20200 17380 20270 17450
rect 20410 17370 20480 17440
rect 20530 17370 20600 17440
rect 20740 17370 20810 17440
rect 20860 17370 20930 17440
rect 21070 17370 21140 17440
rect 21190 17370 21260 17440
rect 21400 17370 21470 17440
rect 21520 17370 21590 17440
rect 21730 17370 21800 17440
rect 21850 17370 21920 17440
rect 22060 17370 22130 17440
rect 22180 17370 22250 17440
rect 22390 17370 22460 17440
rect 22510 17370 22580 17440
rect 22720 17370 22790 17440
rect 22840 17370 22910 17440
rect 23050 17370 23120 17440
rect 23170 17370 23240 17440
rect 17230 16050 17240 16070
rect 17240 16050 17280 16070
rect 17280 16050 17300 16070
rect 17330 16050 17360 16070
rect 17360 16050 17400 16070
rect 17230 16010 17300 16050
rect 17330 16010 17400 16050
rect 11650 15930 11710 15990
rect 11740 15930 11800 15990
rect 11830 15930 11890 15990
rect 11920 15930 11980 15990
rect 12010 15930 12070 15990
rect 12100 15930 12160 15990
rect 12190 15930 12250 15990
rect 12280 15930 12340 15990
rect 12370 15930 12430 15990
rect 12460 15930 12520 15990
rect 12550 15930 12610 15990
rect 12640 15930 12700 15990
rect 12730 15930 12790 15990
rect 12820 15930 12880 15990
rect 12910 15930 12970 15990
rect 13000 15930 13060 15990
rect 13090 15930 13150 15990
rect 13180 15930 13240 15990
rect 13270 15930 13330 15990
rect 13360 15930 13420 15990
rect 13450 15930 13510 15990
rect 13540 15930 13600 15990
rect 13630 15930 13690 15990
rect 13720 15930 13780 15990
rect 13810 15930 13870 15990
rect 13900 15930 13960 15990
rect 13990 15930 14050 15990
rect 14080 15930 14140 15990
rect 14170 15930 14230 15990
rect 14260 15930 14320 15990
rect 14350 15930 14410 15990
rect 14440 15930 14500 15990
rect 14530 15930 14590 15990
rect 14620 15930 14680 15990
rect 14710 15930 14770 15990
rect 14800 15930 14860 15990
rect 14890 15930 14950 15990
rect 14980 15930 15040 15990
rect 15070 15930 15130 15990
rect 15160 15930 15220 15990
rect 15250 15930 15310 15990
rect 15340 15930 15400 15990
rect 15430 15930 15490 15990
rect 15520 15930 15580 15990
rect 15610 15930 15670 15990
rect 15700 15930 15760 15990
rect 15790 15930 15850 15990
rect 15880 15930 15940 15990
rect 15970 15930 16030 15990
rect 16060 15930 16120 15990
rect 16150 15930 16210 15990
rect 16240 15930 16300 15990
rect 16330 15930 16390 15990
rect 16420 15930 16480 15990
rect 16510 15930 16570 15990
rect 16600 15930 16660 15990
rect 16690 15930 16750 15990
rect 16780 15930 16840 15990
rect 16870 15930 16930 15990
rect 16960 15930 17020 15990
rect 17050 15930 17110 15990
rect 17230 15980 17240 16010
rect 17240 15980 17280 16010
rect 17280 15980 17300 16010
rect 17330 15980 17360 16010
rect 17360 15980 17400 16010
rect 17430 16050 17440 16070
rect 17440 16050 17480 16070
rect 17480 16050 17500 16070
rect 17530 16050 17560 16070
rect 17560 16050 17600 16070
rect 17630 16050 17640 16070
rect 17640 16050 17680 16070
rect 17680 16050 17700 16070
rect 17430 16010 17500 16050
rect 17530 16010 17600 16050
rect 17630 16010 17700 16050
rect 17430 15980 17440 16010
rect 17440 15980 17480 16010
rect 17480 15980 17500 16010
rect 17530 15980 17560 16010
rect 17560 15980 17600 16010
rect 17630 15980 17640 16010
rect 17640 15980 17680 16010
rect 17680 15980 17700 16010
rect 17230 15930 17300 15940
rect 17330 15930 17400 15940
rect 11650 15840 11710 15900
rect 11740 15840 11800 15900
rect 11830 15840 11890 15900
rect 11920 15840 11980 15900
rect 12010 15840 12070 15900
rect 12100 15840 12160 15900
rect 12190 15840 12250 15900
rect 12280 15840 12340 15900
rect 12370 15840 12430 15900
rect 12460 15840 12520 15900
rect 12550 15840 12610 15900
rect 12640 15840 12700 15900
rect 12730 15840 12790 15900
rect 12820 15840 12880 15900
rect 12910 15840 12970 15900
rect 13000 15840 13060 15900
rect 13090 15840 13150 15900
rect 13180 15840 13240 15900
rect 13270 15840 13330 15900
rect 13360 15840 13420 15900
rect 13450 15840 13510 15900
rect 13540 15840 13600 15900
rect 13630 15840 13690 15900
rect 13720 15840 13780 15900
rect 13810 15840 13870 15900
rect 13900 15840 13960 15900
rect 13990 15840 14050 15900
rect 14080 15840 14140 15900
rect 14170 15840 14230 15900
rect 14260 15840 14320 15900
rect 14350 15840 14410 15900
rect 14440 15840 14500 15900
rect 14530 15840 14590 15900
rect 14620 15840 14680 15900
rect 14710 15840 14770 15900
rect 14800 15840 14860 15900
rect 14890 15840 14950 15900
rect 14980 15840 15040 15900
rect 15070 15840 15130 15900
rect 15160 15840 15220 15900
rect 15250 15840 15310 15900
rect 15340 15840 15400 15900
rect 15430 15840 15490 15900
rect 15520 15840 15580 15900
rect 15610 15840 15670 15900
rect 15700 15840 15760 15900
rect 15790 15840 15850 15900
rect 15880 15840 15940 15900
rect 15970 15840 16030 15900
rect 16060 15840 16120 15900
rect 16150 15840 16210 15900
rect 16240 15840 16300 15900
rect 16330 15840 16390 15900
rect 16420 15840 16480 15900
rect 16510 15840 16570 15900
rect 16600 15840 16660 15900
rect 16690 15840 16750 15900
rect 16780 15840 16840 15900
rect 16870 15840 16930 15900
rect 16960 15840 17020 15900
rect 17050 15840 17110 15900
rect 17230 15890 17240 15930
rect 17240 15890 17280 15930
rect 17280 15890 17300 15930
rect 17330 15890 17360 15930
rect 17360 15890 17400 15930
rect 17230 15850 17300 15890
rect 17330 15850 17400 15890
rect 17430 15930 17500 15940
rect 17530 15930 17600 15940
rect 17630 15930 17700 15940
rect 17430 15890 17440 15930
rect 17440 15890 17480 15930
rect 17480 15890 17500 15930
rect 17530 15890 17560 15930
rect 17560 15890 17600 15930
rect 17630 15890 17640 15930
rect 17640 15890 17680 15930
rect 17680 15890 17700 15930
rect 17430 15850 17500 15890
rect 17530 15850 17600 15890
rect 17630 15850 17700 15890
rect 18000 15930 18060 15990
rect 18090 15930 18150 15990
rect 18180 15930 18240 15990
rect 18270 15930 18330 15990
rect 18360 15930 18420 15990
rect 18450 15930 18510 15990
rect 18540 15930 18600 15990
rect 18630 15930 18690 15990
rect 18720 15930 18780 15990
rect 18810 15930 18870 15990
rect 18900 15930 18960 15990
rect 18990 15930 19050 15990
rect 19080 15930 19140 15990
rect 19170 15930 19230 15990
rect 19260 15930 19320 15990
rect 19350 15930 19410 15990
rect 19440 15930 19500 15990
rect 19530 15930 19590 15990
rect 19620 15930 19680 15990
rect 19710 15930 19770 15990
rect 19800 15930 19860 15990
rect 19890 15930 19950 15990
rect 19980 15930 20040 15990
rect 20070 15930 20130 15990
rect 20160 15930 20220 15990
rect 20250 15930 20310 15990
rect 20340 15930 20400 15990
rect 20430 15930 20490 15990
rect 20520 15930 20580 15990
rect 20610 15930 20670 15990
rect 20700 15930 20760 15990
rect 20790 15930 20850 15990
rect 20880 15930 20940 15990
rect 20970 15930 21030 15990
rect 21060 15930 21120 15990
rect 21150 15930 21210 15990
rect 21240 15930 21300 15990
rect 21330 15930 21390 15990
rect 21420 15930 21480 15990
rect 21510 15930 21570 15990
rect 21600 15930 21660 15990
rect 21690 15930 21750 15990
rect 21780 15930 21840 15990
rect 21870 15930 21930 15990
rect 21960 15930 22020 15990
rect 22050 15930 22110 15990
rect 22140 15930 22200 15990
rect 22230 15930 22290 15990
rect 22320 15930 22380 15990
rect 22410 15930 22470 15990
rect 22500 15930 22560 15990
rect 22590 15930 22650 15990
rect 22680 15930 22740 15990
rect 22770 15930 22830 15990
rect 22860 15930 22920 15990
rect 22950 15930 23010 15990
rect 23040 15930 23100 15990
rect 23130 15930 23190 15990
rect 23220 15930 23280 15990
rect 18000 15840 18060 15900
rect 18090 15840 18150 15900
rect 18180 15840 18240 15900
rect 18270 15840 18330 15900
rect 18360 15840 18420 15900
rect 18450 15840 18510 15900
rect 18540 15840 18600 15900
rect 18630 15840 18690 15900
rect 18720 15840 18780 15900
rect 18810 15840 18870 15900
rect 18900 15840 18960 15900
rect 18990 15840 19050 15900
rect 19080 15840 19140 15900
rect 19170 15840 19230 15900
rect 19260 15840 19320 15900
rect 19350 15840 19410 15900
rect 19440 15840 19500 15900
rect 19530 15840 19590 15900
rect 19620 15840 19680 15900
rect 19710 15840 19770 15900
rect 19800 15840 19860 15900
rect 19890 15840 19950 15900
rect 19980 15840 20040 15900
rect 20070 15840 20130 15900
rect 20160 15840 20220 15900
rect 20250 15840 20310 15900
rect 20340 15840 20400 15900
rect 20430 15840 20490 15900
rect 20520 15840 20580 15900
rect 20610 15840 20670 15900
rect 20700 15840 20760 15900
rect 20790 15840 20850 15900
rect 20880 15840 20940 15900
rect 20970 15840 21030 15900
rect 21060 15840 21120 15900
rect 21150 15840 21210 15900
rect 21240 15840 21300 15900
rect 21330 15840 21390 15900
rect 21420 15840 21480 15900
rect 21510 15840 21570 15900
rect 21600 15840 21660 15900
rect 21690 15840 21750 15900
rect 21780 15840 21840 15900
rect 21870 15840 21930 15900
rect 21960 15840 22020 15900
rect 22050 15840 22110 15900
rect 22140 15840 22200 15900
rect 22230 15840 22290 15900
rect 22320 15840 22380 15900
rect 22410 15840 22470 15900
rect 22500 15840 22560 15900
rect 22590 15840 22650 15900
rect 22680 15840 22740 15900
rect 22770 15840 22830 15900
rect 22860 15840 22920 15900
rect 22950 15840 23010 15900
rect 23040 15840 23100 15900
rect 23130 15840 23190 15900
rect 23220 15840 23280 15900
rect 11650 13800 11710 13860
rect 11740 13800 11800 13860
rect 11830 13800 11890 13860
rect 11920 13800 11980 13860
rect 12010 13800 12070 13860
rect 12100 13800 12160 13860
rect 12190 13800 12250 13860
rect 12280 13800 12340 13860
rect 12370 13800 12430 13860
rect 12460 13800 12520 13860
rect 12550 13800 12610 13860
rect 12640 13800 12700 13860
rect 12730 13800 12790 13860
rect 12820 13800 12880 13860
rect 12910 13800 12970 13860
rect 13000 13800 13060 13860
rect 13090 13800 13150 13860
rect 13180 13800 13240 13860
rect 13270 13800 13330 13860
rect 13360 13800 13420 13860
rect 13450 13800 13510 13860
rect 13540 13800 13600 13860
rect 13630 13800 13690 13860
rect 13720 13800 13780 13860
rect 13810 13800 13870 13860
rect 13900 13800 13960 13860
rect 13990 13800 14050 13860
rect 14080 13800 14140 13860
rect 14170 13800 14230 13860
rect 14260 13800 14320 13860
rect 14350 13800 14410 13860
rect 14440 13800 14500 13860
rect 14530 13800 14590 13860
rect 14620 13800 14680 13860
rect 14710 13800 14770 13860
rect 14800 13800 14860 13860
rect 14890 13800 14950 13860
rect 14980 13800 15040 13860
rect 15070 13800 15130 13860
rect 15160 13800 15220 13860
rect 15250 13800 15310 13860
rect 15340 13800 15400 13860
rect 15430 13800 15490 13860
rect 15520 13800 15580 13860
rect 15610 13800 15670 13860
rect 15700 13800 15760 13860
rect 15790 13800 15850 13860
rect 15880 13800 15940 13860
rect 15970 13800 16030 13860
rect 16060 13800 16120 13860
rect 16150 13800 16210 13860
rect 16240 13800 16300 13860
rect 16330 13800 16390 13860
rect 16420 13800 16480 13860
rect 16510 13800 16570 13860
rect 16600 13800 16660 13860
rect 16690 13800 16750 13860
rect 16780 13800 16840 13860
rect 16870 13800 16930 13860
rect 11650 13710 11710 13770
rect 11740 13710 11800 13770
rect 11830 13710 11890 13770
rect 11920 13710 11980 13770
rect 12010 13710 12070 13770
rect 12100 13710 12160 13770
rect 12190 13710 12250 13770
rect 12280 13710 12340 13770
rect 12370 13710 12430 13770
rect 12460 13710 12520 13770
rect 12550 13710 12610 13770
rect 12640 13710 12700 13770
rect 12730 13710 12790 13770
rect 12820 13710 12880 13770
rect 12910 13710 12970 13770
rect 13000 13710 13060 13770
rect 13090 13710 13150 13770
rect 13180 13710 13240 13770
rect 13270 13710 13330 13770
rect 13360 13710 13420 13770
rect 13450 13710 13510 13770
rect 13540 13710 13600 13770
rect 13630 13710 13690 13770
rect 13720 13710 13780 13770
rect 13810 13710 13870 13770
rect 13900 13710 13960 13770
rect 13990 13710 14050 13770
rect 14080 13710 14140 13770
rect 14170 13710 14230 13770
rect 14260 13710 14320 13770
rect 14350 13710 14410 13770
rect 14440 13710 14500 13770
rect 14530 13710 14590 13770
rect 14620 13710 14680 13770
rect 14710 13710 14770 13770
rect 14800 13710 14860 13770
rect 14890 13710 14950 13770
rect 14980 13710 15040 13770
rect 15070 13710 15130 13770
rect 15160 13710 15220 13770
rect 15250 13710 15310 13770
rect 15340 13710 15400 13770
rect 15430 13710 15490 13770
rect 15520 13710 15580 13770
rect 15610 13710 15670 13770
rect 15700 13710 15760 13770
rect 15790 13710 15850 13770
rect 15880 13710 15940 13770
rect 15970 13710 16030 13770
rect 16060 13710 16120 13770
rect 16150 13710 16210 13770
rect 16240 13710 16300 13770
rect 16330 13710 16390 13770
rect 16420 13710 16480 13770
rect 16510 13710 16570 13770
rect 16600 13710 16660 13770
rect 16690 13710 16750 13770
rect 16780 13710 16840 13770
rect 16870 13710 16930 13770
rect 17230 13820 17300 13850
rect 17330 13820 17400 13850
rect 17230 13780 17240 13820
rect 17240 13780 17280 13820
rect 17280 13780 17300 13820
rect 17330 13780 17360 13820
rect 17360 13780 17400 13820
rect 17230 13760 17300 13780
rect 17330 13760 17400 13780
rect 17430 13820 17500 13850
rect 17530 13820 17600 13850
rect 17630 13820 17700 13850
rect 17430 13780 17440 13820
rect 17440 13780 17480 13820
rect 17480 13780 17500 13820
rect 17530 13780 17560 13820
rect 17560 13780 17600 13820
rect 17630 13780 17640 13820
rect 17640 13780 17680 13820
rect 17680 13780 17700 13820
rect 17820 13800 17880 13860
rect 17910 13800 17970 13860
rect 18000 13800 18060 13860
rect 18090 13800 18150 13860
rect 18180 13800 18240 13860
rect 18270 13800 18330 13860
rect 18360 13800 18420 13860
rect 18450 13800 18510 13860
rect 18540 13800 18600 13860
rect 18630 13800 18690 13860
rect 18720 13800 18780 13860
rect 18810 13800 18870 13860
rect 18900 13800 18960 13860
rect 18990 13800 19050 13860
rect 19080 13800 19140 13860
rect 19170 13800 19230 13860
rect 19260 13800 19320 13860
rect 19350 13800 19410 13860
rect 19440 13800 19500 13860
rect 19530 13800 19590 13860
rect 19620 13800 19680 13860
rect 19710 13800 19770 13860
rect 19800 13800 19860 13860
rect 19890 13800 19950 13860
rect 19980 13800 20040 13860
rect 20070 13800 20130 13860
rect 20160 13800 20220 13860
rect 20250 13800 20310 13860
rect 20340 13800 20400 13860
rect 20430 13800 20490 13860
rect 20520 13800 20580 13860
rect 20610 13800 20670 13860
rect 20700 13800 20760 13860
rect 20790 13800 20850 13860
rect 20880 13800 20940 13860
rect 20970 13800 21030 13860
rect 21060 13800 21120 13860
rect 21150 13800 21210 13860
rect 21240 13800 21300 13860
rect 21330 13800 21390 13860
rect 21420 13800 21480 13860
rect 21510 13800 21570 13860
rect 21600 13800 21660 13860
rect 21690 13800 21750 13860
rect 21780 13800 21840 13860
rect 21870 13800 21930 13860
rect 21960 13800 22020 13860
rect 22050 13800 22110 13860
rect 22140 13800 22200 13860
rect 22230 13800 22290 13860
rect 22320 13800 22380 13860
rect 22410 13800 22470 13860
rect 22500 13800 22560 13860
rect 22590 13800 22650 13860
rect 22680 13800 22740 13860
rect 22770 13800 22830 13860
rect 22860 13800 22920 13860
rect 22950 13800 23010 13860
rect 23040 13800 23100 13860
rect 23130 13800 23190 13860
rect 23220 13800 23280 13860
rect 17430 13760 17500 13780
rect 17530 13760 17600 13780
rect 17630 13760 17700 13780
rect 17230 13700 17240 13720
rect 17240 13700 17280 13720
rect 17280 13700 17300 13720
rect 17330 13700 17360 13720
rect 17360 13700 17400 13720
rect 17230 13660 17300 13700
rect 17330 13660 17400 13700
rect 17230 13630 17240 13660
rect 17240 13630 17280 13660
rect 17280 13630 17300 13660
rect 17330 13630 17360 13660
rect 17360 13630 17400 13660
rect 17430 13700 17440 13720
rect 17440 13700 17480 13720
rect 17480 13700 17500 13720
rect 17530 13700 17560 13720
rect 17560 13700 17600 13720
rect 17630 13700 17640 13720
rect 17640 13700 17680 13720
rect 17680 13700 17700 13720
rect 17820 13710 17880 13770
rect 17910 13710 17970 13770
rect 18000 13710 18060 13770
rect 18090 13710 18150 13770
rect 18180 13710 18240 13770
rect 18270 13710 18330 13770
rect 18360 13710 18420 13770
rect 18450 13710 18510 13770
rect 18540 13710 18600 13770
rect 18630 13710 18690 13770
rect 18720 13710 18780 13770
rect 18810 13710 18870 13770
rect 18900 13710 18960 13770
rect 18990 13710 19050 13770
rect 19080 13710 19140 13770
rect 19170 13710 19230 13770
rect 19260 13710 19320 13770
rect 19350 13710 19410 13770
rect 19440 13710 19500 13770
rect 19530 13710 19590 13770
rect 19620 13710 19680 13770
rect 19710 13710 19770 13770
rect 19800 13710 19860 13770
rect 19890 13710 19950 13770
rect 19980 13710 20040 13770
rect 20070 13710 20130 13770
rect 20160 13710 20220 13770
rect 20250 13710 20310 13770
rect 20340 13710 20400 13770
rect 20430 13710 20490 13770
rect 20520 13710 20580 13770
rect 20610 13710 20670 13770
rect 20700 13710 20760 13770
rect 20790 13710 20850 13770
rect 20880 13710 20940 13770
rect 20970 13710 21030 13770
rect 21060 13710 21120 13770
rect 21150 13710 21210 13770
rect 21240 13710 21300 13770
rect 21330 13710 21390 13770
rect 21420 13710 21480 13770
rect 21510 13710 21570 13770
rect 21600 13710 21660 13770
rect 21690 13710 21750 13770
rect 21780 13710 21840 13770
rect 21870 13710 21930 13770
rect 21960 13710 22020 13770
rect 22050 13710 22110 13770
rect 22140 13710 22200 13770
rect 22230 13710 22290 13770
rect 22320 13710 22380 13770
rect 22410 13710 22470 13770
rect 22500 13710 22560 13770
rect 22590 13710 22650 13770
rect 22680 13710 22740 13770
rect 22770 13710 22830 13770
rect 22860 13710 22920 13770
rect 22950 13710 23010 13770
rect 23040 13710 23100 13770
rect 23130 13710 23190 13770
rect 23220 13710 23280 13770
rect 17430 13660 17500 13700
rect 17530 13660 17600 13700
rect 17630 13660 17700 13700
rect 17430 13630 17440 13660
rect 17440 13630 17480 13660
rect 17480 13630 17500 13660
rect 17530 13630 17560 13660
rect 17560 13630 17600 13660
rect 17630 13630 17640 13660
rect 17640 13630 17680 13660
rect 17680 13630 17700 13660
rect 11690 12240 11760 12310
rect 11810 12240 11880 12310
rect 12020 12240 12090 12310
rect 12140 12240 12210 12310
rect 12350 12240 12420 12310
rect 12470 12240 12540 12310
rect 12680 12240 12750 12310
rect 12800 12240 12870 12310
rect 13010 12240 13080 12310
rect 13130 12240 13200 12310
rect 13340 12240 13410 12310
rect 13460 12240 13530 12310
rect 13670 12240 13740 12310
rect 13790 12240 13860 12310
rect 14000 12240 14070 12310
rect 14120 12240 14190 12310
rect 14330 12240 14400 12310
rect 14450 12240 14520 12310
rect 14660 12230 14730 12300
rect 14780 12230 14850 12300
rect 14990 12230 15060 12300
rect 15110 12230 15180 12300
rect 15320 12230 15390 12300
rect 15440 12230 15510 12300
rect 15650 12240 15720 12310
rect 15770 12240 15840 12310
rect 15980 12240 16050 12310
rect 16100 12240 16170 12310
rect 16310 12240 16380 12310
rect 16430 12240 16500 12310
rect 16640 12240 16710 12310
rect 16760 12240 16830 12310
rect 11690 12120 11760 12190
rect 11810 12120 11880 12190
rect 12020 12120 12090 12190
rect 12140 12120 12210 12190
rect 12350 12120 12420 12190
rect 12470 12120 12540 12190
rect 12680 12120 12750 12190
rect 12800 12120 12870 12190
rect 13010 12120 13080 12190
rect 13130 12120 13200 12190
rect 13340 12120 13410 12190
rect 13460 12120 13530 12190
rect 13670 12120 13740 12190
rect 13790 12120 13860 12190
rect 14000 12120 14070 12190
rect 14120 12120 14190 12190
rect 14330 12120 14400 12190
rect 14450 12120 14520 12190
rect 14660 12110 14730 12180
rect 14780 12110 14850 12180
rect 14990 12110 15060 12180
rect 15110 12110 15180 12180
rect 15320 12110 15390 12180
rect 15440 12110 15510 12180
rect 15650 12120 15720 12190
rect 15770 12120 15840 12190
rect 15980 12120 16050 12190
rect 16100 12120 16170 12190
rect 16310 12120 16380 12190
rect 16430 12120 16500 12190
rect 16640 12120 16710 12190
rect 16760 12120 16830 12190
rect 18100 12240 18170 12310
rect 18220 12240 18290 12310
rect 18430 12240 18500 12310
rect 18550 12240 18620 12310
rect 18760 12240 18830 12310
rect 18880 12240 18950 12310
rect 19090 12240 19160 12310
rect 19210 12240 19280 12310
rect 19420 12230 19490 12300
rect 19540 12230 19610 12300
rect 19750 12230 19820 12300
rect 19870 12230 19940 12300
rect 20080 12230 20150 12300
rect 20200 12230 20270 12300
rect 20410 12240 20480 12310
rect 20530 12240 20600 12310
rect 20740 12240 20810 12310
rect 20860 12240 20930 12310
rect 21070 12240 21140 12310
rect 21190 12240 21260 12310
rect 21400 12240 21470 12310
rect 21520 12240 21590 12310
rect 21730 12240 21800 12310
rect 21850 12240 21920 12310
rect 22060 12240 22130 12310
rect 22180 12240 22250 12310
rect 22390 12240 22460 12310
rect 22510 12240 22580 12310
rect 22720 12240 22790 12310
rect 22840 12240 22910 12310
rect 23050 12240 23120 12310
rect 23170 12240 23240 12310
rect 18100 12120 18170 12190
rect 18220 12120 18290 12190
rect 18430 12120 18500 12190
rect 18550 12120 18620 12190
rect 18760 12120 18830 12190
rect 18880 12120 18950 12190
rect 19090 12120 19160 12190
rect 19210 12120 19280 12190
rect 19420 12110 19490 12180
rect 19540 12110 19610 12180
rect 19750 12110 19820 12180
rect 19870 12110 19940 12180
rect 20080 12110 20150 12180
rect 20200 12110 20270 12180
rect 20410 12120 20480 12190
rect 20530 12120 20600 12190
rect 20740 12120 20810 12190
rect 20860 12120 20930 12190
rect 21070 12120 21140 12190
rect 21190 12120 21260 12190
rect 21400 12120 21470 12190
rect 21520 12120 21590 12190
rect 21730 12120 21800 12190
rect 21850 12120 21920 12190
rect 22060 12120 22130 12190
rect 22180 12120 22250 12190
rect 22390 12120 22460 12190
rect 22510 12120 22580 12190
rect 22720 12120 22790 12190
rect 22840 12120 22910 12190
rect 23050 12120 23120 12190
rect 23170 12120 23240 12190
<< metal2 >>
rect 11690 17590 11930 17610
rect 12020 17590 12260 17610
rect 12350 17590 12590 17610
rect 12680 17590 12920 17610
rect 13010 17590 13250 17610
rect 13340 17590 13580 17610
rect 13670 17590 13910 17610
rect 14000 17590 14240 17610
rect 14330 17590 14570 17610
rect 14660 17590 14900 17610
rect 14990 17590 15230 17610
rect 15320 17590 15560 17610
rect 15650 17590 15890 17610
rect 15980 17590 16220 17610
rect 16310 17590 16550 17610
rect 16640 17590 16880 17610
rect 18050 17590 18290 17610
rect 18380 17590 18620 17610
rect 18710 17590 18950 17610
rect 19040 17590 19280 17610
rect 19370 17590 19610 17610
rect 19700 17590 19940 17610
rect 20030 17590 20270 17610
rect 20360 17590 20600 17610
rect 20690 17590 20930 17610
rect 21020 17590 21260 17610
rect 21350 17590 21590 17610
rect 21680 17590 21920 17610
rect 22010 17590 22250 17610
rect 22340 17590 22580 17610
rect 22670 17590 22910 17610
rect 23000 17590 23240 17610
rect 11660 17570 17090 17590
rect 11660 17560 14660 17570
rect 11660 17490 11690 17560
rect 11760 17490 11810 17560
rect 11880 17490 12020 17560
rect 12090 17490 12140 17560
rect 12210 17490 12350 17560
rect 12420 17490 12470 17560
rect 12540 17490 12680 17560
rect 12750 17490 12800 17560
rect 12870 17490 13010 17560
rect 13080 17490 13130 17560
rect 13200 17490 13340 17560
rect 13410 17490 13460 17560
rect 13530 17490 13670 17560
rect 13740 17490 13790 17560
rect 13860 17490 14000 17560
rect 14070 17490 14120 17560
rect 14190 17490 14330 17560
rect 14400 17490 14450 17560
rect 14520 17500 14660 17560
rect 14730 17500 14780 17570
rect 14850 17500 14990 17570
rect 15060 17500 15110 17570
rect 15180 17500 15320 17570
rect 15390 17500 15440 17570
rect 15510 17560 17090 17570
rect 15510 17500 15650 17560
rect 14520 17490 15650 17500
rect 15720 17490 15770 17560
rect 15840 17490 15980 17560
rect 16050 17490 16100 17560
rect 16170 17490 16310 17560
rect 16380 17490 16430 17560
rect 16500 17490 16640 17560
rect 16710 17490 16760 17560
rect 16830 17490 17090 17560
rect 11660 17450 17090 17490
rect 11660 17440 14660 17450
rect 11660 17370 11690 17440
rect 11760 17370 11810 17440
rect 11880 17370 12020 17440
rect 12090 17370 12140 17440
rect 12210 17370 12350 17440
rect 12420 17370 12470 17440
rect 12540 17370 12680 17440
rect 12750 17370 12800 17440
rect 12870 17370 13010 17440
rect 13080 17370 13130 17440
rect 13200 17370 13340 17440
rect 13410 17370 13460 17440
rect 13530 17370 13670 17440
rect 13740 17370 13790 17440
rect 13860 17370 14000 17440
rect 14070 17370 14120 17440
rect 14190 17370 14330 17440
rect 14400 17370 14450 17440
rect 14520 17380 14660 17440
rect 14730 17380 14780 17450
rect 14850 17380 14990 17450
rect 15060 17380 15110 17450
rect 15180 17380 15320 17450
rect 15390 17380 15440 17450
rect 15510 17440 17090 17450
rect 15510 17380 15650 17440
rect 14520 17370 15650 17380
rect 15720 17370 15770 17440
rect 15840 17370 15980 17440
rect 16050 17370 16100 17440
rect 16170 17370 16310 17440
rect 16380 17370 16430 17440
rect 16500 17370 16640 17440
rect 16710 17370 16760 17440
rect 16830 17370 17090 17440
rect 11660 17340 17090 17370
rect 17840 17570 23270 17590
rect 17840 17560 19420 17570
rect 17840 17490 18100 17560
rect 18170 17490 18220 17560
rect 18290 17490 18430 17560
rect 18500 17490 18550 17560
rect 18620 17490 18760 17560
rect 18830 17490 18880 17560
rect 18950 17490 19090 17560
rect 19160 17490 19210 17560
rect 19280 17500 19420 17560
rect 19490 17500 19540 17570
rect 19610 17500 19750 17570
rect 19820 17500 19870 17570
rect 19940 17500 20080 17570
rect 20150 17500 20200 17570
rect 20270 17560 23270 17570
rect 20270 17500 20410 17560
rect 19280 17490 20410 17500
rect 20480 17490 20530 17560
rect 20600 17490 20740 17560
rect 20810 17490 20860 17560
rect 20930 17490 21070 17560
rect 21140 17490 21190 17560
rect 21260 17490 21400 17560
rect 21470 17490 21520 17560
rect 21590 17490 21730 17560
rect 21800 17490 21850 17560
rect 21920 17490 22060 17560
rect 22130 17490 22180 17560
rect 22250 17490 22390 17560
rect 22460 17490 22510 17560
rect 22580 17490 22720 17560
rect 22790 17490 22840 17560
rect 22910 17490 23050 17560
rect 23120 17490 23170 17560
rect 23240 17490 23270 17560
rect 17840 17450 23270 17490
rect 17840 17440 19420 17450
rect 17840 17370 18100 17440
rect 18170 17370 18220 17440
rect 18290 17370 18430 17440
rect 18500 17370 18550 17440
rect 18620 17370 18760 17440
rect 18830 17370 18880 17440
rect 18950 17370 19090 17440
rect 19160 17370 19210 17440
rect 19280 17380 19420 17440
rect 19490 17380 19540 17450
rect 19610 17380 19750 17450
rect 19820 17380 19870 17450
rect 19940 17380 20080 17450
rect 20150 17380 20200 17450
rect 20270 17440 23270 17450
rect 20270 17380 20410 17440
rect 19280 17370 20410 17380
rect 20480 17370 20530 17440
rect 20600 17370 20740 17440
rect 20810 17370 20860 17440
rect 20930 17370 21070 17440
rect 21140 17370 21190 17440
rect 21260 17370 21400 17440
rect 21470 17370 21520 17440
rect 21590 17370 21730 17440
rect 21800 17370 21850 17440
rect 21920 17370 22060 17440
rect 22130 17370 22180 17440
rect 22250 17370 22390 17440
rect 22460 17370 22510 17440
rect 22580 17370 22720 17440
rect 22790 17370 22840 17440
rect 22910 17370 23050 17440
rect 23120 17370 23170 17440
rect 23240 17370 23270 17440
rect 17840 17340 23270 17370
rect 17180 16070 17750 16100
rect 17180 16000 17230 16070
rect 11630 15990 17230 16000
rect 11630 15930 11650 15990
rect 11710 15930 11740 15990
rect 11800 15930 11830 15990
rect 11890 15930 11920 15990
rect 11980 15930 12010 15990
rect 12070 15930 12100 15990
rect 12160 15930 12190 15990
rect 12250 15930 12280 15990
rect 12340 15930 12370 15990
rect 12430 15930 12460 15990
rect 12520 15930 12550 15990
rect 12610 15930 12640 15990
rect 12700 15930 12730 15990
rect 12790 15930 12820 15990
rect 12880 15930 12910 15990
rect 12970 15930 13000 15990
rect 13060 15930 13090 15990
rect 13150 15930 13180 15990
rect 13240 15930 13270 15990
rect 13330 15930 13360 15990
rect 13420 15930 13450 15990
rect 13510 15930 13540 15990
rect 13600 15930 13630 15990
rect 13690 15930 13720 15990
rect 13780 15930 13810 15990
rect 13870 15930 13900 15990
rect 13960 15930 13990 15990
rect 14050 15930 14080 15990
rect 14140 15930 14170 15990
rect 14230 15930 14260 15990
rect 14320 15930 14350 15990
rect 14410 15930 14440 15990
rect 14500 15930 14530 15990
rect 14590 15930 14620 15990
rect 14680 15930 14710 15990
rect 14770 15930 14800 15990
rect 14860 15930 14890 15990
rect 14950 15930 14980 15990
rect 15040 15930 15070 15990
rect 15130 15930 15160 15990
rect 15220 15930 15250 15990
rect 15310 15930 15340 15990
rect 15400 15930 15430 15990
rect 15490 15930 15520 15990
rect 15580 15930 15610 15990
rect 15670 15930 15700 15990
rect 15760 15930 15790 15990
rect 15850 15930 15880 15990
rect 15940 15930 15970 15990
rect 16030 15930 16060 15990
rect 16120 15930 16150 15990
rect 16210 15930 16240 15990
rect 16300 15930 16330 15990
rect 16390 15930 16420 15990
rect 16480 15930 16510 15990
rect 16570 15930 16600 15990
rect 16660 15930 16690 15990
rect 16750 15930 16780 15990
rect 16840 15930 16870 15990
rect 16930 15930 16960 15990
rect 17020 15930 17050 15990
rect 17110 15980 17230 15990
rect 17300 15980 17330 16070
rect 17400 15980 17430 16070
rect 17500 15980 17530 16070
rect 17600 15980 17630 16070
rect 17700 15980 17750 16070
rect 17110 15940 17750 15980
rect 17110 15930 17230 15940
rect 11630 15900 17230 15930
rect 11630 15840 11650 15900
rect 11710 15840 11740 15900
rect 11800 15840 11830 15900
rect 11890 15840 11920 15900
rect 11980 15840 12010 15900
rect 12070 15840 12100 15900
rect 12160 15840 12190 15900
rect 12250 15840 12280 15900
rect 12340 15840 12370 15900
rect 12430 15840 12460 15900
rect 12520 15840 12550 15900
rect 12610 15840 12640 15900
rect 12700 15840 12730 15900
rect 12790 15840 12820 15900
rect 12880 15840 12910 15900
rect 12970 15840 13000 15900
rect 13060 15840 13090 15900
rect 13150 15840 13180 15900
rect 13240 15840 13270 15900
rect 13330 15840 13360 15900
rect 13420 15840 13450 15900
rect 13510 15840 13540 15900
rect 13600 15840 13630 15900
rect 13690 15840 13720 15900
rect 13780 15840 13810 15900
rect 13870 15840 13900 15900
rect 13960 15840 13990 15900
rect 14050 15840 14080 15900
rect 14140 15840 14170 15900
rect 14230 15840 14260 15900
rect 14320 15840 14350 15900
rect 14410 15840 14440 15900
rect 14500 15840 14530 15900
rect 14590 15840 14620 15900
rect 14680 15840 14710 15900
rect 14770 15840 14800 15900
rect 14860 15840 14890 15900
rect 14950 15840 14980 15900
rect 15040 15840 15070 15900
rect 15130 15840 15160 15900
rect 15220 15840 15250 15900
rect 15310 15840 15340 15900
rect 15400 15840 15430 15900
rect 15490 15840 15520 15900
rect 15580 15840 15610 15900
rect 15670 15840 15700 15900
rect 15760 15840 15790 15900
rect 15850 15840 15880 15900
rect 15940 15840 15970 15900
rect 16030 15840 16060 15900
rect 16120 15840 16150 15900
rect 16210 15840 16240 15900
rect 16300 15840 16330 15900
rect 16390 15840 16420 15900
rect 16480 15840 16510 15900
rect 16570 15840 16600 15900
rect 16660 15840 16690 15900
rect 16750 15840 16780 15900
rect 16840 15840 16870 15900
rect 16930 15840 16960 15900
rect 17020 15840 17050 15900
rect 17110 15850 17230 15900
rect 17300 15850 17330 15940
rect 17400 15850 17430 15940
rect 17500 15850 17530 15940
rect 17600 15850 17630 15940
rect 17700 15850 17750 15940
rect 17110 15840 17750 15850
rect 11630 15820 17750 15840
rect 17950 15990 23300 16000
rect 17950 15930 18000 15990
rect 18060 15930 18090 15990
rect 18150 15930 18180 15990
rect 18240 15930 18270 15990
rect 18330 15930 18360 15990
rect 18420 15930 18450 15990
rect 18510 15930 18540 15990
rect 18600 15930 18630 15990
rect 18690 15930 18720 15990
rect 18780 15930 18810 15990
rect 18870 15930 18900 15990
rect 18960 15930 18990 15990
rect 19050 15930 19080 15990
rect 19140 15930 19170 15990
rect 19230 15930 19260 15990
rect 19320 15930 19350 15990
rect 19410 15930 19440 15990
rect 19500 15930 19530 15990
rect 19590 15930 19620 15990
rect 19680 15930 19710 15990
rect 19770 15930 19800 15990
rect 19860 15930 19890 15990
rect 19950 15930 19980 15990
rect 20040 15930 20070 15990
rect 20130 15930 20160 15990
rect 20220 15930 20250 15990
rect 20310 15930 20340 15990
rect 20400 15930 20430 15990
rect 20490 15930 20520 15990
rect 20580 15930 20610 15990
rect 20670 15930 20700 15990
rect 20760 15930 20790 15990
rect 20850 15930 20880 15990
rect 20940 15930 20970 15990
rect 21030 15930 21060 15990
rect 21120 15930 21150 15990
rect 21210 15930 21240 15990
rect 21300 15930 21330 15990
rect 21390 15930 21420 15990
rect 21480 15930 21510 15990
rect 21570 15930 21600 15990
rect 21660 15930 21690 15990
rect 21750 15930 21780 15990
rect 21840 15930 21870 15990
rect 21930 15930 21960 15990
rect 22020 15930 22050 15990
rect 22110 15930 22140 15990
rect 22200 15930 22230 15990
rect 22290 15930 22320 15990
rect 22380 15930 22410 15990
rect 22470 15930 22500 15990
rect 22560 15930 22590 15990
rect 22650 15930 22680 15990
rect 22740 15930 22770 15990
rect 22830 15930 22860 15990
rect 22920 15930 22950 15990
rect 23010 15930 23040 15990
rect 23100 15930 23130 15990
rect 23190 15930 23220 15990
rect 23280 15930 23300 15990
rect 17950 15900 23300 15930
rect 17950 15840 18000 15900
rect 18060 15840 18090 15900
rect 18150 15840 18180 15900
rect 18240 15840 18270 15900
rect 18330 15840 18360 15900
rect 18420 15840 18450 15900
rect 18510 15840 18540 15900
rect 18600 15840 18630 15900
rect 18690 15840 18720 15900
rect 18780 15840 18810 15900
rect 18870 15840 18900 15900
rect 18960 15840 18990 15900
rect 19050 15840 19080 15900
rect 19140 15840 19170 15900
rect 19230 15840 19260 15900
rect 19320 15840 19350 15900
rect 19410 15840 19440 15900
rect 19500 15840 19530 15900
rect 19590 15840 19620 15900
rect 19680 15840 19710 15900
rect 19770 15840 19800 15900
rect 19860 15840 19890 15900
rect 19950 15840 19980 15900
rect 20040 15840 20070 15900
rect 20130 15840 20160 15900
rect 20220 15840 20250 15900
rect 20310 15840 20340 15900
rect 20400 15840 20430 15900
rect 20490 15840 20520 15900
rect 20580 15840 20610 15900
rect 20670 15840 20700 15900
rect 20760 15840 20790 15900
rect 20850 15840 20880 15900
rect 20940 15840 20970 15900
rect 21030 15840 21060 15900
rect 21120 15840 21150 15900
rect 21210 15840 21240 15900
rect 21300 15840 21330 15900
rect 21390 15840 21420 15900
rect 21480 15840 21510 15900
rect 21570 15840 21600 15900
rect 21660 15840 21690 15900
rect 21750 15840 21780 15900
rect 21840 15840 21870 15900
rect 21930 15840 21960 15900
rect 22020 15840 22050 15900
rect 22110 15840 22140 15900
rect 22200 15840 22230 15900
rect 22290 15840 22320 15900
rect 22380 15840 22410 15900
rect 22470 15840 22500 15900
rect 22560 15840 22590 15900
rect 22650 15840 22680 15900
rect 22740 15840 22770 15900
rect 22830 15840 22860 15900
rect 22920 15840 22950 15900
rect 23010 15840 23040 15900
rect 23100 15840 23130 15900
rect 23190 15840 23220 15900
rect 23280 15840 23300 15900
rect 17950 15820 23300 15840
rect 11630 13860 16980 13880
rect 11630 13800 11650 13860
rect 11710 13800 11740 13860
rect 11800 13800 11830 13860
rect 11890 13800 11920 13860
rect 11980 13800 12010 13860
rect 12070 13800 12100 13860
rect 12160 13800 12190 13860
rect 12250 13800 12280 13860
rect 12340 13800 12370 13860
rect 12430 13800 12460 13860
rect 12520 13800 12550 13860
rect 12610 13800 12640 13860
rect 12700 13800 12730 13860
rect 12790 13800 12820 13860
rect 12880 13800 12910 13860
rect 12970 13800 13000 13860
rect 13060 13800 13090 13860
rect 13150 13800 13180 13860
rect 13240 13800 13270 13860
rect 13330 13800 13360 13860
rect 13420 13800 13450 13860
rect 13510 13800 13540 13860
rect 13600 13800 13630 13860
rect 13690 13800 13720 13860
rect 13780 13800 13810 13860
rect 13870 13800 13900 13860
rect 13960 13800 13990 13860
rect 14050 13800 14080 13860
rect 14140 13800 14170 13860
rect 14230 13800 14260 13860
rect 14320 13800 14350 13860
rect 14410 13800 14440 13860
rect 14500 13800 14530 13860
rect 14590 13800 14620 13860
rect 14680 13800 14710 13860
rect 14770 13800 14800 13860
rect 14860 13800 14890 13860
rect 14950 13800 14980 13860
rect 15040 13800 15070 13860
rect 15130 13800 15160 13860
rect 15220 13800 15250 13860
rect 15310 13800 15340 13860
rect 15400 13800 15430 13860
rect 15490 13800 15520 13860
rect 15580 13800 15610 13860
rect 15670 13800 15700 13860
rect 15760 13800 15790 13860
rect 15850 13800 15880 13860
rect 15940 13800 15970 13860
rect 16030 13800 16060 13860
rect 16120 13800 16150 13860
rect 16210 13800 16240 13860
rect 16300 13800 16330 13860
rect 16390 13800 16420 13860
rect 16480 13800 16510 13860
rect 16570 13800 16600 13860
rect 16660 13800 16690 13860
rect 16750 13800 16780 13860
rect 16840 13800 16870 13860
rect 16930 13800 16980 13860
rect 11630 13770 16980 13800
rect 11630 13710 11650 13770
rect 11710 13710 11740 13770
rect 11800 13710 11830 13770
rect 11890 13710 11920 13770
rect 11980 13710 12010 13770
rect 12070 13710 12100 13770
rect 12160 13710 12190 13770
rect 12250 13710 12280 13770
rect 12340 13710 12370 13770
rect 12430 13710 12460 13770
rect 12520 13710 12550 13770
rect 12610 13710 12640 13770
rect 12700 13710 12730 13770
rect 12790 13710 12820 13770
rect 12880 13710 12910 13770
rect 12970 13710 13000 13770
rect 13060 13710 13090 13770
rect 13150 13710 13180 13770
rect 13240 13710 13270 13770
rect 13330 13710 13360 13770
rect 13420 13710 13450 13770
rect 13510 13710 13540 13770
rect 13600 13710 13630 13770
rect 13690 13710 13720 13770
rect 13780 13710 13810 13770
rect 13870 13710 13900 13770
rect 13960 13710 13990 13770
rect 14050 13710 14080 13770
rect 14140 13710 14170 13770
rect 14230 13710 14260 13770
rect 14320 13710 14350 13770
rect 14410 13710 14440 13770
rect 14500 13710 14530 13770
rect 14590 13710 14620 13770
rect 14680 13710 14710 13770
rect 14770 13710 14800 13770
rect 14860 13710 14890 13770
rect 14950 13710 14980 13770
rect 15040 13710 15070 13770
rect 15130 13710 15160 13770
rect 15220 13710 15250 13770
rect 15310 13710 15340 13770
rect 15400 13710 15430 13770
rect 15490 13710 15520 13770
rect 15580 13710 15610 13770
rect 15670 13710 15700 13770
rect 15760 13710 15790 13770
rect 15850 13710 15880 13770
rect 15940 13710 15970 13770
rect 16030 13710 16060 13770
rect 16120 13710 16150 13770
rect 16210 13710 16240 13770
rect 16300 13710 16330 13770
rect 16390 13710 16420 13770
rect 16480 13710 16510 13770
rect 16570 13710 16600 13770
rect 16660 13710 16690 13770
rect 16750 13710 16780 13770
rect 16840 13710 16870 13770
rect 16930 13710 16980 13770
rect 11630 13700 16980 13710
rect 17180 13860 23300 13880
rect 17180 13850 17820 13860
rect 17180 13760 17230 13850
rect 17300 13760 17330 13850
rect 17400 13760 17430 13850
rect 17500 13760 17530 13850
rect 17600 13760 17630 13850
rect 17700 13800 17820 13850
rect 17880 13800 17910 13860
rect 17970 13800 18000 13860
rect 18060 13800 18090 13860
rect 18150 13800 18180 13860
rect 18240 13800 18270 13860
rect 18330 13800 18360 13860
rect 18420 13800 18450 13860
rect 18510 13800 18540 13860
rect 18600 13800 18630 13860
rect 18690 13800 18720 13860
rect 18780 13800 18810 13860
rect 18870 13800 18900 13860
rect 18960 13800 18990 13860
rect 19050 13800 19080 13860
rect 19140 13800 19170 13860
rect 19230 13800 19260 13860
rect 19320 13800 19350 13860
rect 19410 13800 19440 13860
rect 19500 13800 19530 13860
rect 19590 13800 19620 13860
rect 19680 13800 19710 13860
rect 19770 13800 19800 13860
rect 19860 13800 19890 13860
rect 19950 13800 19980 13860
rect 20040 13800 20070 13860
rect 20130 13800 20160 13860
rect 20220 13800 20250 13860
rect 20310 13800 20340 13860
rect 20400 13800 20430 13860
rect 20490 13800 20520 13860
rect 20580 13800 20610 13860
rect 20670 13800 20700 13860
rect 20760 13800 20790 13860
rect 20850 13800 20880 13860
rect 20940 13800 20970 13860
rect 21030 13800 21060 13860
rect 21120 13800 21150 13860
rect 21210 13800 21240 13860
rect 21300 13800 21330 13860
rect 21390 13800 21420 13860
rect 21480 13800 21510 13860
rect 21570 13800 21600 13860
rect 21660 13800 21690 13860
rect 21750 13800 21780 13860
rect 21840 13800 21870 13860
rect 21930 13800 21960 13860
rect 22020 13800 22050 13860
rect 22110 13800 22140 13860
rect 22200 13800 22230 13860
rect 22290 13800 22320 13860
rect 22380 13800 22410 13860
rect 22470 13800 22500 13860
rect 22560 13800 22590 13860
rect 22650 13800 22680 13860
rect 22740 13800 22770 13860
rect 22830 13800 22860 13860
rect 22920 13800 22950 13860
rect 23010 13800 23040 13860
rect 23100 13800 23130 13860
rect 23190 13800 23220 13860
rect 23280 13800 23300 13860
rect 17700 13770 23300 13800
rect 17700 13760 17820 13770
rect 17180 13720 17820 13760
rect 17180 13630 17230 13720
rect 17300 13630 17330 13720
rect 17400 13630 17430 13720
rect 17500 13630 17530 13720
rect 17600 13630 17630 13720
rect 17700 13710 17820 13720
rect 17880 13710 17910 13770
rect 17970 13710 18000 13770
rect 18060 13710 18090 13770
rect 18150 13710 18180 13770
rect 18240 13710 18270 13770
rect 18330 13710 18360 13770
rect 18420 13710 18450 13770
rect 18510 13710 18540 13770
rect 18600 13710 18630 13770
rect 18690 13710 18720 13770
rect 18780 13710 18810 13770
rect 18870 13710 18900 13770
rect 18960 13710 18990 13770
rect 19050 13710 19080 13770
rect 19140 13710 19170 13770
rect 19230 13710 19260 13770
rect 19320 13710 19350 13770
rect 19410 13710 19440 13770
rect 19500 13710 19530 13770
rect 19590 13710 19620 13770
rect 19680 13710 19710 13770
rect 19770 13710 19800 13770
rect 19860 13710 19890 13770
rect 19950 13710 19980 13770
rect 20040 13710 20070 13770
rect 20130 13710 20160 13770
rect 20220 13710 20250 13770
rect 20310 13710 20340 13770
rect 20400 13710 20430 13770
rect 20490 13710 20520 13770
rect 20580 13710 20610 13770
rect 20670 13710 20700 13770
rect 20760 13710 20790 13770
rect 20850 13710 20880 13770
rect 20940 13710 20970 13770
rect 21030 13710 21060 13770
rect 21120 13710 21150 13770
rect 21210 13710 21240 13770
rect 21300 13710 21330 13770
rect 21390 13710 21420 13770
rect 21480 13710 21510 13770
rect 21570 13710 21600 13770
rect 21660 13710 21690 13770
rect 21750 13710 21780 13770
rect 21840 13710 21870 13770
rect 21930 13710 21960 13770
rect 22020 13710 22050 13770
rect 22110 13710 22140 13770
rect 22200 13710 22230 13770
rect 22290 13710 22320 13770
rect 22380 13710 22410 13770
rect 22470 13710 22500 13770
rect 22560 13710 22590 13770
rect 22650 13710 22680 13770
rect 22740 13710 22770 13770
rect 22830 13710 22860 13770
rect 22920 13710 22950 13770
rect 23010 13710 23040 13770
rect 23100 13710 23130 13770
rect 23190 13710 23220 13770
rect 23280 13710 23300 13770
rect 17700 13700 23300 13710
rect 17700 13630 17750 13700
rect 17180 13600 17750 13630
rect 11660 12310 17090 12340
rect 11660 12240 11690 12310
rect 11760 12240 11810 12310
rect 11880 12240 12020 12310
rect 12090 12240 12140 12310
rect 12210 12240 12350 12310
rect 12420 12240 12470 12310
rect 12540 12240 12680 12310
rect 12750 12240 12800 12310
rect 12870 12240 13010 12310
rect 13080 12240 13130 12310
rect 13200 12240 13340 12310
rect 13410 12240 13460 12310
rect 13530 12240 13670 12310
rect 13740 12240 13790 12310
rect 13860 12240 14000 12310
rect 14070 12240 14120 12310
rect 14190 12240 14330 12310
rect 14400 12240 14450 12310
rect 14520 12300 15650 12310
rect 14520 12240 14660 12300
rect 11660 12230 14660 12240
rect 14730 12230 14780 12300
rect 14850 12230 14990 12300
rect 15060 12230 15110 12300
rect 15180 12230 15320 12300
rect 15390 12230 15440 12300
rect 15510 12240 15650 12300
rect 15720 12240 15770 12310
rect 15840 12240 15980 12310
rect 16050 12240 16100 12310
rect 16170 12240 16310 12310
rect 16380 12240 16430 12310
rect 16500 12240 16640 12310
rect 16710 12240 16760 12310
rect 16830 12240 17090 12310
rect 15510 12230 17090 12240
rect 11660 12190 17090 12230
rect 11660 12120 11690 12190
rect 11760 12120 11810 12190
rect 11880 12120 12020 12190
rect 12090 12120 12140 12190
rect 12210 12120 12350 12190
rect 12420 12120 12470 12190
rect 12540 12120 12680 12190
rect 12750 12120 12800 12190
rect 12870 12120 13010 12190
rect 13080 12120 13130 12190
rect 13200 12120 13340 12190
rect 13410 12120 13460 12190
rect 13530 12120 13670 12190
rect 13740 12120 13790 12190
rect 13860 12120 14000 12190
rect 14070 12120 14120 12190
rect 14190 12120 14330 12190
rect 14400 12120 14450 12190
rect 14520 12180 15650 12190
rect 14520 12120 14660 12180
rect 11660 12110 14660 12120
rect 14730 12110 14780 12180
rect 14850 12110 14990 12180
rect 15060 12110 15110 12180
rect 15180 12110 15320 12180
rect 15390 12110 15440 12180
rect 15510 12120 15650 12180
rect 15720 12120 15770 12190
rect 15840 12120 15980 12190
rect 16050 12120 16100 12190
rect 16170 12120 16310 12190
rect 16380 12120 16430 12190
rect 16500 12120 16640 12190
rect 16710 12120 16760 12190
rect 16830 12120 17090 12190
rect 15510 12110 17090 12120
rect 11660 12090 17090 12110
rect 17840 12310 23270 12340
rect 17840 12240 18100 12310
rect 18170 12240 18220 12310
rect 18290 12240 18430 12310
rect 18500 12240 18550 12310
rect 18620 12240 18760 12310
rect 18830 12240 18880 12310
rect 18950 12240 19090 12310
rect 19160 12240 19210 12310
rect 19280 12300 20410 12310
rect 19280 12240 19420 12300
rect 17840 12230 19420 12240
rect 19490 12230 19540 12300
rect 19610 12230 19750 12300
rect 19820 12230 19870 12300
rect 19940 12230 20080 12300
rect 20150 12230 20200 12300
rect 20270 12240 20410 12300
rect 20480 12240 20530 12310
rect 20600 12240 20740 12310
rect 20810 12240 20860 12310
rect 20930 12240 21070 12310
rect 21140 12240 21190 12310
rect 21260 12240 21400 12310
rect 21470 12240 21520 12310
rect 21590 12240 21730 12310
rect 21800 12240 21850 12310
rect 21920 12240 22060 12310
rect 22130 12240 22180 12310
rect 22250 12240 22390 12310
rect 22460 12240 22510 12310
rect 22580 12240 22720 12310
rect 22790 12240 22840 12310
rect 22910 12240 23050 12310
rect 23120 12240 23170 12310
rect 23240 12240 23270 12310
rect 20270 12230 23270 12240
rect 17840 12190 23270 12230
rect 17840 12120 18100 12190
rect 18170 12120 18220 12190
rect 18290 12120 18430 12190
rect 18500 12120 18550 12190
rect 18620 12120 18760 12190
rect 18830 12120 18880 12190
rect 18950 12120 19090 12190
rect 19160 12120 19210 12190
rect 19280 12180 20410 12190
rect 19280 12120 19420 12180
rect 17840 12110 19420 12120
rect 19490 12110 19540 12180
rect 19610 12110 19750 12180
rect 19820 12110 19870 12180
rect 19940 12110 20080 12180
rect 20150 12110 20200 12180
rect 20270 12120 20410 12180
rect 20480 12120 20530 12190
rect 20600 12120 20740 12190
rect 20810 12120 20860 12190
rect 20930 12120 21070 12190
rect 21140 12120 21190 12190
rect 21260 12120 21400 12190
rect 21470 12120 21520 12190
rect 21590 12120 21730 12190
rect 21800 12120 21850 12190
rect 21920 12120 22060 12190
rect 22130 12120 22180 12190
rect 22250 12120 22390 12190
rect 22460 12120 22510 12190
rect 22580 12120 22720 12190
rect 22790 12120 22840 12190
rect 22910 12120 23050 12190
rect 23120 12120 23170 12190
rect 23240 12120 23270 12190
rect 20270 12110 23270 12120
rect 17840 12090 23270 12110
rect 11690 12070 11930 12090
rect 12020 12070 12260 12090
rect 12350 12070 12590 12090
rect 12680 12070 12920 12090
rect 13010 12070 13250 12090
rect 13340 12070 13580 12090
rect 13670 12070 13910 12090
rect 14000 12070 14240 12090
rect 14330 12070 14570 12090
rect 14660 12070 14900 12090
rect 14990 12070 15230 12090
rect 15320 12070 15560 12090
rect 15650 12070 15890 12090
rect 15980 12070 16220 12090
rect 16310 12070 16550 12090
rect 16640 12070 16880 12090
rect 18050 12070 18290 12090
rect 18380 12070 18620 12090
rect 18710 12070 18950 12090
rect 19040 12070 19280 12090
rect 19370 12070 19610 12090
rect 19700 12070 19940 12090
rect 20030 12070 20270 12090
rect 20360 12070 20600 12090
rect 20690 12070 20930 12090
rect 21020 12070 21260 12090
rect 21350 12070 21590 12090
rect 21680 12070 21920 12090
rect 22010 12070 22250 12090
rect 22340 12070 22580 12090
rect 22670 12070 22910 12090
rect 23000 12070 23240 12090
<< via2 >>
rect 11690 17490 11760 17560
rect 11810 17490 11880 17560
rect 12020 17490 12090 17560
rect 12140 17490 12210 17560
rect 12350 17490 12420 17560
rect 12470 17490 12540 17560
rect 12680 17490 12750 17560
rect 12800 17490 12870 17560
rect 13010 17490 13080 17560
rect 13130 17490 13200 17560
rect 13340 17490 13410 17560
rect 13460 17490 13530 17560
rect 13670 17490 13740 17560
rect 13790 17490 13860 17560
rect 14000 17490 14070 17560
rect 14120 17490 14190 17560
rect 14330 17490 14400 17560
rect 14450 17490 14520 17560
rect 14660 17500 14730 17570
rect 14780 17500 14850 17570
rect 14990 17500 15060 17570
rect 15110 17500 15180 17570
rect 15320 17500 15390 17570
rect 15440 17500 15510 17570
rect 15650 17490 15720 17560
rect 15770 17490 15840 17560
rect 15980 17490 16050 17560
rect 16100 17490 16170 17560
rect 16310 17490 16380 17560
rect 16430 17490 16500 17560
rect 16640 17490 16710 17560
rect 16760 17490 16830 17560
rect 11690 17370 11760 17440
rect 11810 17370 11880 17440
rect 12020 17370 12090 17440
rect 12140 17370 12210 17440
rect 12350 17370 12420 17440
rect 12470 17370 12540 17440
rect 12680 17370 12750 17440
rect 12800 17370 12870 17440
rect 13010 17370 13080 17440
rect 13130 17370 13200 17440
rect 13340 17370 13410 17440
rect 13460 17370 13530 17440
rect 13670 17370 13740 17440
rect 13790 17370 13860 17440
rect 14000 17370 14070 17440
rect 14120 17370 14190 17440
rect 14330 17370 14400 17440
rect 14450 17370 14520 17440
rect 14660 17380 14730 17450
rect 14780 17380 14850 17450
rect 14990 17380 15060 17450
rect 15110 17380 15180 17450
rect 15320 17380 15390 17450
rect 15440 17380 15510 17450
rect 15650 17370 15720 17440
rect 15770 17370 15840 17440
rect 15980 17370 16050 17440
rect 16100 17370 16170 17440
rect 16310 17370 16380 17440
rect 16430 17370 16500 17440
rect 16640 17370 16710 17440
rect 16760 17370 16830 17440
rect 18100 17490 18170 17560
rect 18220 17490 18290 17560
rect 18430 17490 18500 17560
rect 18550 17490 18620 17560
rect 18760 17490 18830 17560
rect 18880 17490 18950 17560
rect 19090 17490 19160 17560
rect 19210 17490 19280 17560
rect 19420 17500 19490 17570
rect 19540 17500 19610 17570
rect 19750 17500 19820 17570
rect 19870 17500 19940 17570
rect 20080 17500 20150 17570
rect 20200 17500 20270 17570
rect 20410 17490 20480 17560
rect 20530 17490 20600 17560
rect 20740 17490 20810 17560
rect 20860 17490 20930 17560
rect 21070 17490 21140 17560
rect 21190 17490 21260 17560
rect 21400 17490 21470 17560
rect 21520 17490 21590 17560
rect 21730 17490 21800 17560
rect 21850 17490 21920 17560
rect 22060 17490 22130 17560
rect 22180 17490 22250 17560
rect 22390 17490 22460 17560
rect 22510 17490 22580 17560
rect 22720 17490 22790 17560
rect 22840 17490 22910 17560
rect 23050 17490 23120 17560
rect 23170 17490 23240 17560
rect 18100 17370 18170 17440
rect 18220 17370 18290 17440
rect 18430 17370 18500 17440
rect 18550 17370 18620 17440
rect 18760 17370 18830 17440
rect 18880 17370 18950 17440
rect 19090 17370 19160 17440
rect 19210 17370 19280 17440
rect 19420 17380 19490 17450
rect 19540 17380 19610 17450
rect 19750 17380 19820 17450
rect 19870 17380 19940 17450
rect 20080 17380 20150 17450
rect 20200 17380 20270 17450
rect 20410 17370 20480 17440
rect 20530 17370 20600 17440
rect 20740 17370 20810 17440
rect 20860 17370 20930 17440
rect 21070 17370 21140 17440
rect 21190 17370 21260 17440
rect 21400 17370 21470 17440
rect 21520 17370 21590 17440
rect 21730 17370 21800 17440
rect 21850 17370 21920 17440
rect 22060 17370 22130 17440
rect 22180 17370 22250 17440
rect 22390 17370 22460 17440
rect 22510 17370 22580 17440
rect 22720 17370 22790 17440
rect 22840 17370 22910 17440
rect 23050 17370 23120 17440
rect 23170 17370 23240 17440
rect 11650 15930 11710 15990
rect 11740 15930 11800 15990
rect 11830 15930 11890 15990
rect 11920 15930 11980 15990
rect 12010 15930 12070 15990
rect 12100 15930 12160 15990
rect 12190 15930 12250 15990
rect 12280 15930 12340 15990
rect 12370 15930 12430 15990
rect 12460 15930 12520 15990
rect 12550 15930 12610 15990
rect 12640 15930 12700 15990
rect 12730 15930 12790 15990
rect 12820 15930 12880 15990
rect 12910 15930 12970 15990
rect 13000 15930 13060 15990
rect 13090 15930 13150 15990
rect 13180 15930 13240 15990
rect 13270 15930 13330 15990
rect 13360 15930 13420 15990
rect 13450 15930 13510 15990
rect 13540 15930 13600 15990
rect 13630 15930 13690 15990
rect 13720 15930 13780 15990
rect 13810 15930 13870 15990
rect 13900 15930 13960 15990
rect 13990 15930 14050 15990
rect 14080 15930 14140 15990
rect 14170 15930 14230 15990
rect 14260 15930 14320 15990
rect 14350 15930 14410 15990
rect 14440 15930 14500 15990
rect 14530 15930 14590 15990
rect 14620 15930 14680 15990
rect 14710 15930 14770 15990
rect 14800 15930 14860 15990
rect 14890 15930 14950 15990
rect 14980 15930 15040 15990
rect 15070 15930 15130 15990
rect 15160 15930 15220 15990
rect 15250 15930 15310 15990
rect 15340 15930 15400 15990
rect 15430 15930 15490 15990
rect 15520 15930 15580 15990
rect 15610 15930 15670 15990
rect 15700 15930 15760 15990
rect 15790 15930 15850 15990
rect 15880 15930 15940 15990
rect 15970 15930 16030 15990
rect 16060 15930 16120 15990
rect 16150 15930 16210 15990
rect 16240 15930 16300 15990
rect 16330 15930 16390 15990
rect 16420 15930 16480 15990
rect 16510 15930 16570 15990
rect 16600 15930 16660 15990
rect 16690 15930 16750 15990
rect 16780 15930 16840 15990
rect 16870 15930 16930 15990
rect 16960 15930 17020 15990
rect 17050 15930 17110 15990
rect 17230 15980 17300 16070
rect 17330 15980 17400 16070
rect 17430 15980 17500 16070
rect 17530 15980 17600 16070
rect 17630 15980 17700 16070
rect 11650 15840 11710 15900
rect 11740 15840 11800 15900
rect 11830 15840 11890 15900
rect 11920 15840 11980 15900
rect 12010 15840 12070 15900
rect 12100 15840 12160 15900
rect 12190 15840 12250 15900
rect 12280 15840 12340 15900
rect 12370 15840 12430 15900
rect 12460 15840 12520 15900
rect 12550 15840 12610 15900
rect 12640 15840 12700 15900
rect 12730 15840 12790 15900
rect 12820 15840 12880 15900
rect 12910 15840 12970 15900
rect 13000 15840 13060 15900
rect 13090 15840 13150 15900
rect 13180 15840 13240 15900
rect 13270 15840 13330 15900
rect 13360 15840 13420 15900
rect 13450 15840 13510 15900
rect 13540 15840 13600 15900
rect 13630 15840 13690 15900
rect 13720 15840 13780 15900
rect 13810 15840 13870 15900
rect 13900 15840 13960 15900
rect 13990 15840 14050 15900
rect 14080 15840 14140 15900
rect 14170 15840 14230 15900
rect 14260 15840 14320 15900
rect 14350 15840 14410 15900
rect 14440 15840 14500 15900
rect 14530 15840 14590 15900
rect 14620 15840 14680 15900
rect 14710 15840 14770 15900
rect 14800 15840 14860 15900
rect 14890 15840 14950 15900
rect 14980 15840 15040 15900
rect 15070 15840 15130 15900
rect 15160 15840 15220 15900
rect 15250 15840 15310 15900
rect 15340 15840 15400 15900
rect 15430 15840 15490 15900
rect 15520 15840 15580 15900
rect 15610 15840 15670 15900
rect 15700 15840 15760 15900
rect 15790 15840 15850 15900
rect 15880 15840 15940 15900
rect 15970 15840 16030 15900
rect 16060 15840 16120 15900
rect 16150 15840 16210 15900
rect 16240 15840 16300 15900
rect 16330 15840 16390 15900
rect 16420 15840 16480 15900
rect 16510 15840 16570 15900
rect 16600 15840 16660 15900
rect 16690 15840 16750 15900
rect 16780 15840 16840 15900
rect 16870 15840 16930 15900
rect 16960 15840 17020 15900
rect 17050 15840 17110 15900
rect 17230 15850 17300 15940
rect 17330 15850 17400 15940
rect 17430 15850 17500 15940
rect 17530 15850 17600 15940
rect 17630 15850 17700 15940
rect 18000 15930 18060 15990
rect 18090 15930 18150 15990
rect 18180 15930 18240 15990
rect 18270 15930 18330 15990
rect 18360 15930 18420 15990
rect 18450 15930 18510 15990
rect 18540 15930 18600 15990
rect 18630 15930 18690 15990
rect 18720 15930 18780 15990
rect 18810 15930 18870 15990
rect 18900 15930 18960 15990
rect 18990 15930 19050 15990
rect 19080 15930 19140 15990
rect 19170 15930 19230 15990
rect 19260 15930 19320 15990
rect 19350 15930 19410 15990
rect 19440 15930 19500 15990
rect 19530 15930 19590 15990
rect 19620 15930 19680 15990
rect 19710 15930 19770 15990
rect 19800 15930 19860 15990
rect 19890 15930 19950 15990
rect 19980 15930 20040 15990
rect 20070 15930 20130 15990
rect 20160 15930 20220 15990
rect 20250 15930 20310 15990
rect 20340 15930 20400 15990
rect 20430 15930 20490 15990
rect 20520 15930 20580 15990
rect 20610 15930 20670 15990
rect 20700 15930 20760 15990
rect 20790 15930 20850 15990
rect 20880 15930 20940 15990
rect 20970 15930 21030 15990
rect 21060 15930 21120 15990
rect 21150 15930 21210 15990
rect 21240 15930 21300 15990
rect 21330 15930 21390 15990
rect 21420 15930 21480 15990
rect 21510 15930 21570 15990
rect 21600 15930 21660 15990
rect 21690 15930 21750 15990
rect 21780 15930 21840 15990
rect 21870 15930 21930 15990
rect 21960 15930 22020 15990
rect 22050 15930 22110 15990
rect 22140 15930 22200 15990
rect 22230 15930 22290 15990
rect 22320 15930 22380 15990
rect 22410 15930 22470 15990
rect 22500 15930 22560 15990
rect 22590 15930 22650 15990
rect 22680 15930 22740 15990
rect 22770 15930 22830 15990
rect 22860 15930 22920 15990
rect 22950 15930 23010 15990
rect 23040 15930 23100 15990
rect 23130 15930 23190 15990
rect 23220 15930 23280 15990
rect 18000 15840 18060 15900
rect 18090 15840 18150 15900
rect 18180 15840 18240 15900
rect 18270 15840 18330 15900
rect 18360 15840 18420 15900
rect 18450 15840 18510 15900
rect 18540 15840 18600 15900
rect 18630 15840 18690 15900
rect 18720 15840 18780 15900
rect 18810 15840 18870 15900
rect 18900 15840 18960 15900
rect 18990 15840 19050 15900
rect 19080 15840 19140 15900
rect 19170 15840 19230 15900
rect 19260 15840 19320 15900
rect 19350 15840 19410 15900
rect 19440 15840 19500 15900
rect 19530 15840 19590 15900
rect 19620 15840 19680 15900
rect 19710 15840 19770 15900
rect 19800 15840 19860 15900
rect 19890 15840 19950 15900
rect 19980 15840 20040 15900
rect 20070 15840 20130 15900
rect 20160 15840 20220 15900
rect 20250 15840 20310 15900
rect 20340 15840 20400 15900
rect 20430 15840 20490 15900
rect 20520 15840 20580 15900
rect 20610 15840 20670 15900
rect 20700 15840 20760 15900
rect 20790 15840 20850 15900
rect 20880 15840 20940 15900
rect 20970 15840 21030 15900
rect 21060 15840 21120 15900
rect 21150 15840 21210 15900
rect 21240 15840 21300 15900
rect 21330 15840 21390 15900
rect 21420 15840 21480 15900
rect 21510 15840 21570 15900
rect 21600 15840 21660 15900
rect 21690 15840 21750 15900
rect 21780 15840 21840 15900
rect 21870 15840 21930 15900
rect 21960 15840 22020 15900
rect 22050 15840 22110 15900
rect 22140 15840 22200 15900
rect 22230 15840 22290 15900
rect 22320 15840 22380 15900
rect 22410 15840 22470 15900
rect 22500 15840 22560 15900
rect 22590 15840 22650 15900
rect 22680 15840 22740 15900
rect 22770 15840 22830 15900
rect 22860 15840 22920 15900
rect 22950 15840 23010 15900
rect 23040 15840 23100 15900
rect 23130 15840 23190 15900
rect 23220 15840 23280 15900
rect 11650 13800 11710 13860
rect 11740 13800 11800 13860
rect 11830 13800 11890 13860
rect 11920 13800 11980 13860
rect 12010 13800 12070 13860
rect 12100 13800 12160 13860
rect 12190 13800 12250 13860
rect 12280 13800 12340 13860
rect 12370 13800 12430 13860
rect 12460 13800 12520 13860
rect 12550 13800 12610 13860
rect 12640 13800 12700 13860
rect 12730 13800 12790 13860
rect 12820 13800 12880 13860
rect 12910 13800 12970 13860
rect 13000 13800 13060 13860
rect 13090 13800 13150 13860
rect 13180 13800 13240 13860
rect 13270 13800 13330 13860
rect 13360 13800 13420 13860
rect 13450 13800 13510 13860
rect 13540 13800 13600 13860
rect 13630 13800 13690 13860
rect 13720 13800 13780 13860
rect 13810 13800 13870 13860
rect 13900 13800 13960 13860
rect 13990 13800 14050 13860
rect 14080 13800 14140 13860
rect 14170 13800 14230 13860
rect 14260 13800 14320 13860
rect 14350 13800 14410 13860
rect 14440 13800 14500 13860
rect 14530 13800 14590 13860
rect 14620 13800 14680 13860
rect 14710 13800 14770 13860
rect 14800 13800 14860 13860
rect 14890 13800 14950 13860
rect 14980 13800 15040 13860
rect 15070 13800 15130 13860
rect 15160 13800 15220 13860
rect 15250 13800 15310 13860
rect 15340 13800 15400 13860
rect 15430 13800 15490 13860
rect 15520 13800 15580 13860
rect 15610 13800 15670 13860
rect 15700 13800 15760 13860
rect 15790 13800 15850 13860
rect 15880 13800 15940 13860
rect 15970 13800 16030 13860
rect 16060 13800 16120 13860
rect 16150 13800 16210 13860
rect 16240 13800 16300 13860
rect 16330 13800 16390 13860
rect 16420 13800 16480 13860
rect 16510 13800 16570 13860
rect 16600 13800 16660 13860
rect 16690 13800 16750 13860
rect 16780 13800 16840 13860
rect 16870 13800 16930 13860
rect 11650 13710 11710 13770
rect 11740 13710 11800 13770
rect 11830 13710 11890 13770
rect 11920 13710 11980 13770
rect 12010 13710 12070 13770
rect 12100 13710 12160 13770
rect 12190 13710 12250 13770
rect 12280 13710 12340 13770
rect 12370 13710 12430 13770
rect 12460 13710 12520 13770
rect 12550 13710 12610 13770
rect 12640 13710 12700 13770
rect 12730 13710 12790 13770
rect 12820 13710 12880 13770
rect 12910 13710 12970 13770
rect 13000 13710 13060 13770
rect 13090 13710 13150 13770
rect 13180 13710 13240 13770
rect 13270 13710 13330 13770
rect 13360 13710 13420 13770
rect 13450 13710 13510 13770
rect 13540 13710 13600 13770
rect 13630 13710 13690 13770
rect 13720 13710 13780 13770
rect 13810 13710 13870 13770
rect 13900 13710 13960 13770
rect 13990 13710 14050 13770
rect 14080 13710 14140 13770
rect 14170 13710 14230 13770
rect 14260 13710 14320 13770
rect 14350 13710 14410 13770
rect 14440 13710 14500 13770
rect 14530 13710 14590 13770
rect 14620 13710 14680 13770
rect 14710 13710 14770 13770
rect 14800 13710 14860 13770
rect 14890 13710 14950 13770
rect 14980 13710 15040 13770
rect 15070 13710 15130 13770
rect 15160 13710 15220 13770
rect 15250 13710 15310 13770
rect 15340 13710 15400 13770
rect 15430 13710 15490 13770
rect 15520 13710 15580 13770
rect 15610 13710 15670 13770
rect 15700 13710 15760 13770
rect 15790 13710 15850 13770
rect 15880 13710 15940 13770
rect 15970 13710 16030 13770
rect 16060 13710 16120 13770
rect 16150 13710 16210 13770
rect 16240 13710 16300 13770
rect 16330 13710 16390 13770
rect 16420 13710 16480 13770
rect 16510 13710 16570 13770
rect 16600 13710 16660 13770
rect 16690 13710 16750 13770
rect 16780 13710 16840 13770
rect 16870 13710 16930 13770
rect 17230 13760 17300 13850
rect 17330 13760 17400 13850
rect 17430 13760 17500 13850
rect 17530 13760 17600 13850
rect 17630 13760 17700 13850
rect 17820 13800 17880 13860
rect 17910 13800 17970 13860
rect 18000 13800 18060 13860
rect 18090 13800 18150 13860
rect 18180 13800 18240 13860
rect 18270 13800 18330 13860
rect 18360 13800 18420 13860
rect 18450 13800 18510 13860
rect 18540 13800 18600 13860
rect 18630 13800 18690 13860
rect 18720 13800 18780 13860
rect 18810 13800 18870 13860
rect 18900 13800 18960 13860
rect 18990 13800 19050 13860
rect 19080 13800 19140 13860
rect 19170 13800 19230 13860
rect 19260 13800 19320 13860
rect 19350 13800 19410 13860
rect 19440 13800 19500 13860
rect 19530 13800 19590 13860
rect 19620 13800 19680 13860
rect 19710 13800 19770 13860
rect 19800 13800 19860 13860
rect 19890 13800 19950 13860
rect 19980 13800 20040 13860
rect 20070 13800 20130 13860
rect 20160 13800 20220 13860
rect 20250 13800 20310 13860
rect 20340 13800 20400 13860
rect 20430 13800 20490 13860
rect 20520 13800 20580 13860
rect 20610 13800 20670 13860
rect 20700 13800 20760 13860
rect 20790 13800 20850 13860
rect 20880 13800 20940 13860
rect 20970 13800 21030 13860
rect 21060 13800 21120 13860
rect 21150 13800 21210 13860
rect 21240 13800 21300 13860
rect 21330 13800 21390 13860
rect 21420 13800 21480 13860
rect 21510 13800 21570 13860
rect 21600 13800 21660 13860
rect 21690 13800 21750 13860
rect 21780 13800 21840 13860
rect 21870 13800 21930 13860
rect 21960 13800 22020 13860
rect 22050 13800 22110 13860
rect 22140 13800 22200 13860
rect 22230 13800 22290 13860
rect 22320 13800 22380 13860
rect 22410 13800 22470 13860
rect 22500 13800 22560 13860
rect 22590 13800 22650 13860
rect 22680 13800 22740 13860
rect 22770 13800 22830 13860
rect 22860 13800 22920 13860
rect 22950 13800 23010 13860
rect 23040 13800 23100 13860
rect 23130 13800 23190 13860
rect 23220 13800 23280 13860
rect 17230 13630 17300 13720
rect 17330 13630 17400 13720
rect 17430 13630 17500 13720
rect 17530 13630 17600 13720
rect 17630 13630 17700 13720
rect 17820 13710 17880 13770
rect 17910 13710 17970 13770
rect 18000 13710 18060 13770
rect 18090 13710 18150 13770
rect 18180 13710 18240 13770
rect 18270 13710 18330 13770
rect 18360 13710 18420 13770
rect 18450 13710 18510 13770
rect 18540 13710 18600 13770
rect 18630 13710 18690 13770
rect 18720 13710 18780 13770
rect 18810 13710 18870 13770
rect 18900 13710 18960 13770
rect 18990 13710 19050 13770
rect 19080 13710 19140 13770
rect 19170 13710 19230 13770
rect 19260 13710 19320 13770
rect 19350 13710 19410 13770
rect 19440 13710 19500 13770
rect 19530 13710 19590 13770
rect 19620 13710 19680 13770
rect 19710 13710 19770 13770
rect 19800 13710 19860 13770
rect 19890 13710 19950 13770
rect 19980 13710 20040 13770
rect 20070 13710 20130 13770
rect 20160 13710 20220 13770
rect 20250 13710 20310 13770
rect 20340 13710 20400 13770
rect 20430 13710 20490 13770
rect 20520 13710 20580 13770
rect 20610 13710 20670 13770
rect 20700 13710 20760 13770
rect 20790 13710 20850 13770
rect 20880 13710 20940 13770
rect 20970 13710 21030 13770
rect 21060 13710 21120 13770
rect 21150 13710 21210 13770
rect 21240 13710 21300 13770
rect 21330 13710 21390 13770
rect 21420 13710 21480 13770
rect 21510 13710 21570 13770
rect 21600 13710 21660 13770
rect 21690 13710 21750 13770
rect 21780 13710 21840 13770
rect 21870 13710 21930 13770
rect 21960 13710 22020 13770
rect 22050 13710 22110 13770
rect 22140 13710 22200 13770
rect 22230 13710 22290 13770
rect 22320 13710 22380 13770
rect 22410 13710 22470 13770
rect 22500 13710 22560 13770
rect 22590 13710 22650 13770
rect 22680 13710 22740 13770
rect 22770 13710 22830 13770
rect 22860 13710 22920 13770
rect 22950 13710 23010 13770
rect 23040 13710 23100 13770
rect 23130 13710 23190 13770
rect 23220 13710 23280 13770
rect 11690 12240 11760 12310
rect 11810 12240 11880 12310
rect 12020 12240 12090 12310
rect 12140 12240 12210 12310
rect 12350 12240 12420 12310
rect 12470 12240 12540 12310
rect 12680 12240 12750 12310
rect 12800 12240 12870 12310
rect 13010 12240 13080 12310
rect 13130 12240 13200 12310
rect 13340 12240 13410 12310
rect 13460 12240 13530 12310
rect 13670 12240 13740 12310
rect 13790 12240 13860 12310
rect 14000 12240 14070 12310
rect 14120 12240 14190 12310
rect 14330 12240 14400 12310
rect 14450 12240 14520 12310
rect 14660 12230 14730 12300
rect 14780 12230 14850 12300
rect 14990 12230 15060 12300
rect 15110 12230 15180 12300
rect 15320 12230 15390 12300
rect 15440 12230 15510 12300
rect 15650 12240 15720 12310
rect 15770 12240 15840 12310
rect 15980 12240 16050 12310
rect 16100 12240 16170 12310
rect 16310 12240 16380 12310
rect 16430 12240 16500 12310
rect 16640 12240 16710 12310
rect 16760 12240 16830 12310
rect 11690 12120 11760 12190
rect 11810 12120 11880 12190
rect 12020 12120 12090 12190
rect 12140 12120 12210 12190
rect 12350 12120 12420 12190
rect 12470 12120 12540 12190
rect 12680 12120 12750 12190
rect 12800 12120 12870 12190
rect 13010 12120 13080 12190
rect 13130 12120 13200 12190
rect 13340 12120 13410 12190
rect 13460 12120 13530 12190
rect 13670 12120 13740 12190
rect 13790 12120 13860 12190
rect 14000 12120 14070 12190
rect 14120 12120 14190 12190
rect 14330 12120 14400 12190
rect 14450 12120 14520 12190
rect 14660 12110 14730 12180
rect 14780 12110 14850 12180
rect 14990 12110 15060 12180
rect 15110 12110 15180 12180
rect 15320 12110 15390 12180
rect 15440 12110 15510 12180
rect 15650 12120 15720 12190
rect 15770 12120 15840 12190
rect 15980 12120 16050 12190
rect 16100 12120 16170 12190
rect 16310 12120 16380 12190
rect 16430 12120 16500 12190
rect 16640 12120 16710 12190
rect 16760 12120 16830 12190
rect 18100 12240 18170 12310
rect 18220 12240 18290 12310
rect 18430 12240 18500 12310
rect 18550 12240 18620 12310
rect 18760 12240 18830 12310
rect 18880 12240 18950 12310
rect 19090 12240 19160 12310
rect 19210 12240 19280 12310
rect 19420 12230 19490 12300
rect 19540 12230 19610 12300
rect 19750 12230 19820 12300
rect 19870 12230 19940 12300
rect 20080 12230 20150 12300
rect 20200 12230 20270 12300
rect 20410 12240 20480 12310
rect 20530 12240 20600 12310
rect 20740 12240 20810 12310
rect 20860 12240 20930 12310
rect 21070 12240 21140 12310
rect 21190 12240 21260 12310
rect 21400 12240 21470 12310
rect 21520 12240 21590 12310
rect 21730 12240 21800 12310
rect 21850 12240 21920 12310
rect 22060 12240 22130 12310
rect 22180 12240 22250 12310
rect 22390 12240 22460 12310
rect 22510 12240 22580 12310
rect 22720 12240 22790 12310
rect 22840 12240 22910 12310
rect 23050 12240 23120 12310
rect 23170 12240 23240 12310
rect 18100 12120 18170 12190
rect 18220 12120 18290 12190
rect 18430 12120 18500 12190
rect 18550 12120 18620 12190
rect 18760 12120 18830 12190
rect 18880 12120 18950 12190
rect 19090 12120 19160 12190
rect 19210 12120 19280 12190
rect 19420 12110 19490 12180
rect 19540 12110 19610 12180
rect 19750 12110 19820 12180
rect 19870 12110 19940 12180
rect 20080 12110 20150 12180
rect 20200 12110 20270 12180
rect 20410 12120 20480 12190
rect 20530 12120 20600 12190
rect 20740 12120 20810 12190
rect 20860 12120 20930 12190
rect 21070 12120 21140 12190
rect 21190 12120 21260 12190
rect 21400 12120 21470 12190
rect 21520 12120 21590 12190
rect 21730 12120 21800 12190
rect 21850 12120 21920 12190
rect 22060 12120 22130 12190
rect 22180 12120 22250 12190
rect 22390 12120 22460 12190
rect 22510 12120 22580 12190
rect 22720 12120 22790 12190
rect 22840 12120 22910 12190
rect 23050 12120 23120 12190
rect 23170 12120 23240 12190
<< metal3 >>
rect 11690 17590 11930 17610
rect 12020 17590 12260 17610
rect 12350 17590 12590 17610
rect 12680 17590 12920 17610
rect 13010 17590 13250 17610
rect 13340 17590 13580 17610
rect 13670 17590 13910 17610
rect 14000 17590 14240 17610
rect 14330 17590 14570 17610
rect 14660 17590 14900 17610
rect 14990 17590 15230 17610
rect 15320 17590 15560 17610
rect 15650 17590 15890 17610
rect 15980 17590 16220 17610
rect 16310 17590 16550 17610
rect 16640 17590 16880 17610
rect 18050 17590 18290 17610
rect 18380 17590 18620 17610
rect 18710 17590 18950 17610
rect 19040 17590 19280 17610
rect 19370 17590 19610 17610
rect 19700 17590 19940 17610
rect 20030 17590 20270 17610
rect 20360 17590 20600 17610
rect 20690 17590 20930 17610
rect 21020 17590 21260 17610
rect 21350 17590 21590 17610
rect 21680 17590 21920 17610
rect 22010 17590 22250 17610
rect 22340 17590 22580 17610
rect 22670 17590 22910 17610
rect 23000 17590 23240 17610
rect 11660 17570 17090 17590
rect 11660 17560 14660 17570
rect 11660 17490 11690 17560
rect 11760 17490 11810 17560
rect 11880 17490 12020 17560
rect 12090 17490 12140 17560
rect 12210 17490 12350 17560
rect 12420 17490 12470 17560
rect 12540 17490 12680 17560
rect 12750 17490 12800 17560
rect 12870 17490 13010 17560
rect 13080 17490 13130 17560
rect 13200 17490 13340 17560
rect 13410 17490 13460 17560
rect 13530 17490 13670 17560
rect 13740 17490 13790 17560
rect 13860 17490 14000 17560
rect 14070 17490 14120 17560
rect 14190 17490 14330 17560
rect 14400 17490 14450 17560
rect 14520 17500 14660 17560
rect 14730 17500 14780 17570
rect 14850 17500 14990 17570
rect 15060 17500 15110 17570
rect 15180 17500 15320 17570
rect 15390 17500 15440 17570
rect 15510 17560 17090 17570
rect 15510 17500 15650 17560
rect 14520 17490 15650 17500
rect 15720 17490 15770 17560
rect 15840 17490 15980 17560
rect 16050 17490 16100 17560
rect 16170 17490 16310 17560
rect 16380 17490 16430 17560
rect 16500 17490 16640 17560
rect 16710 17490 16760 17560
rect 16830 17490 17090 17560
rect 11660 17450 17090 17490
rect 11660 17440 14660 17450
rect 11660 17370 11690 17440
rect 11760 17370 11810 17440
rect 11880 17370 12020 17440
rect 12090 17370 12140 17440
rect 12210 17370 12350 17440
rect 12420 17370 12470 17440
rect 12540 17370 12680 17440
rect 12750 17370 12800 17440
rect 12870 17370 13010 17440
rect 13080 17370 13130 17440
rect 13200 17370 13340 17440
rect 13410 17370 13460 17440
rect 13530 17370 13670 17440
rect 13740 17370 13790 17440
rect 13860 17370 14000 17440
rect 14070 17370 14120 17440
rect 14190 17370 14330 17440
rect 14400 17370 14450 17440
rect 14520 17380 14660 17440
rect 14730 17380 14780 17450
rect 14850 17380 14990 17450
rect 15060 17380 15110 17450
rect 15180 17380 15320 17450
rect 15390 17380 15440 17450
rect 15510 17440 17090 17450
rect 15510 17380 15650 17440
rect 14520 17370 15650 17380
rect 15720 17370 15770 17440
rect 15840 17370 15980 17440
rect 16050 17370 16100 17440
rect 16170 17370 16310 17440
rect 16380 17370 16430 17440
rect 16500 17370 16640 17440
rect 16710 17370 16760 17440
rect 16830 17370 17090 17440
rect 11660 17340 17090 17370
rect 17840 17570 23270 17590
rect 17840 17560 19420 17570
rect 17840 17490 18100 17560
rect 18170 17490 18220 17560
rect 18290 17490 18430 17560
rect 18500 17490 18550 17560
rect 18620 17490 18760 17560
rect 18830 17490 18880 17560
rect 18950 17490 19090 17560
rect 19160 17490 19210 17560
rect 19280 17500 19420 17560
rect 19490 17500 19540 17570
rect 19610 17500 19750 17570
rect 19820 17500 19870 17570
rect 19940 17500 20080 17570
rect 20150 17500 20200 17570
rect 20270 17560 23270 17570
rect 20270 17500 20410 17560
rect 19280 17490 20410 17500
rect 20480 17490 20530 17560
rect 20600 17490 20740 17560
rect 20810 17490 20860 17560
rect 20930 17490 21070 17560
rect 21140 17490 21190 17560
rect 21260 17490 21400 17560
rect 21470 17490 21520 17560
rect 21590 17490 21730 17560
rect 21800 17490 21850 17560
rect 21920 17490 22060 17560
rect 22130 17490 22180 17560
rect 22250 17490 22390 17560
rect 22460 17490 22510 17560
rect 22580 17490 22720 17560
rect 22790 17490 22840 17560
rect 22910 17490 23050 17560
rect 23120 17490 23170 17560
rect 23240 17490 23270 17560
rect 17840 17450 23270 17490
rect 17840 17440 19420 17450
rect 17840 17370 18100 17440
rect 18170 17370 18220 17440
rect 18290 17370 18430 17440
rect 18500 17370 18550 17440
rect 18620 17370 18760 17440
rect 18830 17370 18880 17440
rect 18950 17370 19090 17440
rect 19160 17370 19210 17440
rect 19280 17380 19420 17440
rect 19490 17380 19540 17450
rect 19610 17380 19750 17450
rect 19820 17380 19870 17450
rect 19940 17380 20080 17450
rect 20150 17380 20200 17450
rect 20270 17440 23270 17450
rect 20270 17380 20410 17440
rect 19280 17370 20410 17380
rect 20480 17370 20530 17440
rect 20600 17370 20740 17440
rect 20810 17370 20860 17440
rect 20930 17370 21070 17440
rect 21140 17370 21190 17440
rect 21260 17370 21400 17440
rect 21470 17370 21520 17440
rect 21590 17370 21730 17440
rect 21800 17370 21850 17440
rect 21920 17370 22060 17440
rect 22130 17370 22180 17440
rect 22250 17370 22390 17440
rect 22460 17370 22510 17440
rect 22580 17370 22720 17440
rect 22790 17370 22840 17440
rect 22910 17370 23050 17440
rect 23120 17370 23170 17440
rect 23240 17370 23270 17440
rect 17840 17340 23270 17370
rect 17180 16070 17750 16100
rect 17180 16000 17230 16070
rect 11630 15990 17230 16000
rect 11630 15930 11650 15990
rect 11710 15930 11740 15990
rect 11800 15930 11830 15990
rect 11890 15930 11920 15990
rect 11980 15930 12010 15990
rect 12070 15930 12100 15990
rect 12160 15930 12190 15990
rect 12250 15930 12280 15990
rect 12340 15930 12370 15990
rect 12430 15930 12460 15990
rect 12520 15930 12550 15990
rect 12610 15930 12640 15990
rect 12700 15930 12730 15990
rect 12790 15930 12820 15990
rect 12880 15930 12910 15990
rect 12970 15930 13000 15990
rect 13060 15930 13090 15990
rect 13150 15930 13180 15990
rect 13240 15930 13270 15990
rect 13330 15930 13360 15990
rect 13420 15930 13450 15990
rect 13510 15930 13540 15990
rect 13600 15930 13630 15990
rect 13690 15930 13720 15990
rect 13780 15930 13810 15990
rect 13870 15930 13900 15990
rect 13960 15930 13990 15990
rect 14050 15930 14080 15990
rect 14140 15930 14170 15990
rect 14230 15930 14260 15990
rect 14320 15930 14350 15990
rect 14410 15930 14440 15990
rect 14500 15930 14530 15990
rect 14590 15930 14620 15990
rect 14680 15930 14710 15990
rect 14770 15930 14800 15990
rect 14860 15930 14890 15990
rect 14950 15930 14980 15990
rect 15040 15930 15070 15990
rect 15130 15930 15160 15990
rect 15220 15930 15250 15990
rect 15310 15930 15340 15990
rect 15400 15930 15430 15990
rect 15490 15930 15520 15990
rect 15580 15930 15610 15990
rect 15670 15930 15700 15990
rect 15760 15930 15790 15990
rect 15850 15930 15880 15990
rect 15940 15930 15970 15990
rect 16030 15930 16060 15990
rect 16120 15930 16150 15990
rect 16210 15930 16240 15990
rect 16300 15930 16330 15990
rect 16390 15930 16420 15990
rect 16480 15930 16510 15990
rect 16570 15930 16600 15990
rect 16660 15930 16690 15990
rect 16750 15930 16780 15990
rect 16840 15930 16870 15990
rect 16930 15930 16960 15990
rect 17020 15930 17050 15990
rect 17110 15980 17230 15990
rect 17300 15980 17330 16070
rect 17400 15980 17430 16070
rect 17500 15980 17530 16070
rect 17600 15980 17630 16070
rect 17700 15980 17750 16070
rect 17110 15940 17750 15980
rect 17110 15930 17230 15940
rect 11630 15900 17230 15930
rect 11630 15840 11650 15900
rect 11710 15840 11740 15900
rect 11800 15840 11830 15900
rect 11890 15840 11920 15900
rect 11980 15840 12010 15900
rect 12070 15840 12100 15900
rect 12160 15840 12190 15900
rect 12250 15840 12280 15900
rect 12340 15840 12370 15900
rect 12430 15840 12460 15900
rect 12520 15840 12550 15900
rect 12610 15840 12640 15900
rect 12700 15840 12730 15900
rect 12790 15840 12820 15900
rect 12880 15840 12910 15900
rect 12970 15840 13000 15900
rect 13060 15840 13090 15900
rect 13150 15840 13180 15900
rect 13240 15840 13270 15900
rect 13330 15840 13360 15900
rect 13420 15840 13450 15900
rect 13510 15840 13540 15900
rect 13600 15840 13630 15900
rect 13690 15840 13720 15900
rect 13780 15840 13810 15900
rect 13870 15840 13900 15900
rect 13960 15840 13990 15900
rect 14050 15840 14080 15900
rect 14140 15840 14170 15900
rect 14230 15840 14260 15900
rect 14320 15840 14350 15900
rect 14410 15840 14440 15900
rect 14500 15840 14530 15900
rect 14590 15840 14620 15900
rect 14680 15840 14710 15900
rect 14770 15840 14800 15900
rect 14860 15840 14890 15900
rect 14950 15840 14980 15900
rect 15040 15840 15070 15900
rect 15130 15840 15160 15900
rect 15220 15840 15250 15900
rect 15310 15840 15340 15900
rect 15400 15840 15430 15900
rect 15490 15840 15520 15900
rect 15580 15840 15610 15900
rect 15670 15840 15700 15900
rect 15760 15840 15790 15900
rect 15850 15840 15880 15900
rect 15940 15840 15970 15900
rect 16030 15840 16060 15900
rect 16120 15840 16150 15900
rect 16210 15840 16240 15900
rect 16300 15840 16330 15900
rect 16390 15840 16420 15900
rect 16480 15840 16510 15900
rect 16570 15840 16600 15900
rect 16660 15840 16690 15900
rect 16750 15840 16780 15900
rect 16840 15840 16870 15900
rect 16930 15840 16960 15900
rect 17020 15840 17050 15900
rect 17110 15850 17230 15900
rect 17300 15850 17330 15940
rect 17400 15850 17430 15940
rect 17500 15850 17530 15940
rect 17600 15850 17630 15940
rect 17700 15850 17750 15940
rect 17110 15840 17750 15850
rect 11630 15820 17750 15840
rect 17950 15990 23300 16000
rect 17950 15930 18000 15990
rect 18060 15930 18090 15990
rect 18150 15930 18180 15990
rect 18240 15930 18270 15990
rect 18330 15930 18360 15990
rect 18420 15930 18450 15990
rect 18510 15930 18540 15990
rect 18600 15930 18630 15990
rect 18690 15930 18720 15990
rect 18780 15930 18810 15990
rect 18870 15930 18900 15990
rect 18960 15930 18990 15990
rect 19050 15930 19080 15990
rect 19140 15930 19170 15990
rect 19230 15930 19260 15990
rect 19320 15930 19350 15990
rect 19410 15930 19440 15990
rect 19500 15930 19530 15990
rect 19590 15930 19620 15990
rect 19680 15930 19710 15990
rect 19770 15930 19800 15990
rect 19860 15930 19890 15990
rect 19950 15930 19980 15990
rect 20040 15930 20070 15990
rect 20130 15930 20160 15990
rect 20220 15930 20250 15990
rect 20310 15930 20340 15990
rect 20400 15930 20430 15990
rect 20490 15930 20520 15990
rect 20580 15930 20610 15990
rect 20670 15930 20700 15990
rect 20760 15930 20790 15990
rect 20850 15930 20880 15990
rect 20940 15930 20970 15990
rect 21030 15930 21060 15990
rect 21120 15930 21150 15990
rect 21210 15930 21240 15990
rect 21300 15930 21330 15990
rect 21390 15930 21420 15990
rect 21480 15930 21510 15990
rect 21570 15930 21600 15990
rect 21660 15930 21690 15990
rect 21750 15930 21780 15990
rect 21840 15930 21870 15990
rect 21930 15930 21960 15990
rect 22020 15930 22050 15990
rect 22110 15930 22140 15990
rect 22200 15930 22230 15990
rect 22290 15930 22320 15990
rect 22380 15930 22410 15990
rect 22470 15930 22500 15990
rect 22560 15930 22590 15990
rect 22650 15930 22680 15990
rect 22740 15930 22770 15990
rect 22830 15930 22860 15990
rect 22920 15930 22950 15990
rect 23010 15930 23040 15990
rect 23100 15930 23130 15990
rect 23190 15930 23220 15990
rect 23280 15930 23300 15990
rect 17950 15900 23300 15930
rect 17950 15840 18000 15900
rect 18060 15840 18090 15900
rect 18150 15840 18180 15900
rect 18240 15840 18270 15900
rect 18330 15840 18360 15900
rect 18420 15840 18450 15900
rect 18510 15840 18540 15900
rect 18600 15840 18630 15900
rect 18690 15840 18720 15900
rect 18780 15840 18810 15900
rect 18870 15840 18900 15900
rect 18960 15840 18990 15900
rect 19050 15840 19080 15900
rect 19140 15840 19170 15900
rect 19230 15840 19260 15900
rect 19320 15840 19350 15900
rect 19410 15840 19440 15900
rect 19500 15840 19530 15900
rect 19590 15840 19620 15900
rect 19680 15840 19710 15900
rect 19770 15840 19800 15900
rect 19860 15840 19890 15900
rect 19950 15840 19980 15900
rect 20040 15840 20070 15900
rect 20130 15840 20160 15900
rect 20220 15840 20250 15900
rect 20310 15840 20340 15900
rect 20400 15840 20430 15900
rect 20490 15840 20520 15900
rect 20580 15840 20610 15900
rect 20670 15840 20700 15900
rect 20760 15840 20790 15900
rect 20850 15840 20880 15900
rect 20940 15840 20970 15900
rect 21030 15840 21060 15900
rect 21120 15840 21150 15900
rect 21210 15840 21240 15900
rect 21300 15840 21330 15900
rect 21390 15840 21420 15900
rect 21480 15840 21510 15900
rect 21570 15840 21600 15900
rect 21660 15840 21690 15900
rect 21750 15840 21780 15900
rect 21840 15840 21870 15900
rect 21930 15840 21960 15900
rect 22020 15840 22050 15900
rect 22110 15840 22140 15900
rect 22200 15840 22230 15900
rect 22290 15840 22320 15900
rect 22380 15840 22410 15900
rect 22470 15840 22500 15900
rect 22560 15840 22590 15900
rect 22650 15840 22680 15900
rect 22740 15840 22770 15900
rect 22830 15840 22860 15900
rect 22920 15840 22950 15900
rect 23010 15840 23040 15900
rect 23100 15840 23130 15900
rect 23190 15840 23220 15900
rect 23280 15840 23300 15900
rect 11630 13860 16980 15820
rect 17950 13880 23300 15840
rect 11630 13800 11650 13860
rect 11710 13800 11740 13860
rect 11800 13800 11830 13860
rect 11890 13800 11920 13860
rect 11980 13800 12010 13860
rect 12070 13800 12100 13860
rect 12160 13800 12190 13860
rect 12250 13800 12280 13860
rect 12340 13800 12370 13860
rect 12430 13800 12460 13860
rect 12520 13800 12550 13860
rect 12610 13800 12640 13860
rect 12700 13800 12730 13860
rect 12790 13800 12820 13860
rect 12880 13800 12910 13860
rect 12970 13800 13000 13860
rect 13060 13800 13090 13860
rect 13150 13800 13180 13860
rect 13240 13800 13270 13860
rect 13330 13800 13360 13860
rect 13420 13800 13450 13860
rect 13510 13800 13540 13860
rect 13600 13800 13630 13860
rect 13690 13800 13720 13860
rect 13780 13800 13810 13860
rect 13870 13800 13900 13860
rect 13960 13800 13990 13860
rect 14050 13800 14080 13860
rect 14140 13800 14170 13860
rect 14230 13800 14260 13860
rect 14320 13800 14350 13860
rect 14410 13800 14440 13860
rect 14500 13800 14530 13860
rect 14590 13800 14620 13860
rect 14680 13800 14710 13860
rect 14770 13800 14800 13860
rect 14860 13800 14890 13860
rect 14950 13800 14980 13860
rect 15040 13800 15070 13860
rect 15130 13800 15160 13860
rect 15220 13800 15250 13860
rect 15310 13800 15340 13860
rect 15400 13800 15430 13860
rect 15490 13800 15520 13860
rect 15580 13800 15610 13860
rect 15670 13800 15700 13860
rect 15760 13800 15790 13860
rect 15850 13800 15880 13860
rect 15940 13800 15970 13860
rect 16030 13800 16060 13860
rect 16120 13800 16150 13860
rect 16210 13800 16240 13860
rect 16300 13800 16330 13860
rect 16390 13800 16420 13860
rect 16480 13800 16510 13860
rect 16570 13800 16600 13860
rect 16660 13800 16690 13860
rect 16750 13800 16780 13860
rect 16840 13800 16870 13860
rect 16930 13800 16980 13860
rect 11630 13770 16980 13800
rect 11630 13710 11650 13770
rect 11710 13710 11740 13770
rect 11800 13710 11830 13770
rect 11890 13710 11920 13770
rect 11980 13710 12010 13770
rect 12070 13710 12100 13770
rect 12160 13710 12190 13770
rect 12250 13710 12280 13770
rect 12340 13710 12370 13770
rect 12430 13710 12460 13770
rect 12520 13710 12550 13770
rect 12610 13710 12640 13770
rect 12700 13710 12730 13770
rect 12790 13710 12820 13770
rect 12880 13710 12910 13770
rect 12970 13710 13000 13770
rect 13060 13710 13090 13770
rect 13150 13710 13180 13770
rect 13240 13710 13270 13770
rect 13330 13710 13360 13770
rect 13420 13710 13450 13770
rect 13510 13710 13540 13770
rect 13600 13710 13630 13770
rect 13690 13710 13720 13770
rect 13780 13710 13810 13770
rect 13870 13710 13900 13770
rect 13960 13710 13990 13770
rect 14050 13710 14080 13770
rect 14140 13710 14170 13770
rect 14230 13710 14260 13770
rect 14320 13710 14350 13770
rect 14410 13710 14440 13770
rect 14500 13710 14530 13770
rect 14590 13710 14620 13770
rect 14680 13710 14710 13770
rect 14770 13710 14800 13770
rect 14860 13710 14890 13770
rect 14950 13710 14980 13770
rect 15040 13710 15070 13770
rect 15130 13710 15160 13770
rect 15220 13710 15250 13770
rect 15310 13710 15340 13770
rect 15400 13710 15430 13770
rect 15490 13710 15520 13770
rect 15580 13710 15610 13770
rect 15670 13710 15700 13770
rect 15760 13710 15790 13770
rect 15850 13710 15880 13770
rect 15940 13710 15970 13770
rect 16030 13710 16060 13770
rect 16120 13710 16150 13770
rect 16210 13710 16240 13770
rect 16300 13710 16330 13770
rect 16390 13710 16420 13770
rect 16480 13710 16510 13770
rect 16570 13710 16600 13770
rect 16660 13710 16690 13770
rect 16750 13710 16780 13770
rect 16840 13710 16870 13770
rect 16930 13710 16980 13770
rect 11630 13700 16980 13710
rect 17180 13860 23300 13880
rect 17180 13850 17820 13860
rect 17180 13760 17230 13850
rect 17300 13760 17330 13850
rect 17400 13760 17430 13850
rect 17500 13760 17530 13850
rect 17600 13760 17630 13850
rect 17700 13800 17820 13850
rect 17880 13800 17910 13860
rect 17970 13800 18000 13860
rect 18060 13800 18090 13860
rect 18150 13800 18180 13860
rect 18240 13800 18270 13860
rect 18330 13800 18360 13860
rect 18420 13800 18450 13860
rect 18510 13800 18540 13860
rect 18600 13800 18630 13860
rect 18690 13800 18720 13860
rect 18780 13800 18810 13860
rect 18870 13800 18900 13860
rect 18960 13800 18990 13860
rect 19050 13800 19080 13860
rect 19140 13800 19170 13860
rect 19230 13800 19260 13860
rect 19320 13800 19350 13860
rect 19410 13800 19440 13860
rect 19500 13800 19530 13860
rect 19590 13800 19620 13860
rect 19680 13800 19710 13860
rect 19770 13800 19800 13860
rect 19860 13800 19890 13860
rect 19950 13800 19980 13860
rect 20040 13800 20070 13860
rect 20130 13800 20160 13860
rect 20220 13800 20250 13860
rect 20310 13800 20340 13860
rect 20400 13800 20430 13860
rect 20490 13800 20520 13860
rect 20580 13800 20610 13860
rect 20670 13800 20700 13860
rect 20760 13800 20790 13860
rect 20850 13800 20880 13860
rect 20940 13800 20970 13860
rect 21030 13800 21060 13860
rect 21120 13800 21150 13860
rect 21210 13800 21240 13860
rect 21300 13800 21330 13860
rect 21390 13800 21420 13860
rect 21480 13800 21510 13860
rect 21570 13800 21600 13860
rect 21660 13800 21690 13860
rect 21750 13800 21780 13860
rect 21840 13800 21870 13860
rect 21930 13800 21960 13860
rect 22020 13800 22050 13860
rect 22110 13800 22140 13860
rect 22200 13800 22230 13860
rect 22290 13800 22320 13860
rect 22380 13800 22410 13860
rect 22470 13800 22500 13860
rect 22560 13800 22590 13860
rect 22650 13800 22680 13860
rect 22740 13800 22770 13860
rect 22830 13800 22860 13860
rect 22920 13800 22950 13860
rect 23010 13800 23040 13860
rect 23100 13800 23130 13860
rect 23190 13800 23220 13860
rect 23280 13800 23300 13860
rect 17700 13770 23300 13800
rect 17700 13760 17820 13770
rect 17180 13720 17820 13760
rect 17180 13630 17230 13720
rect 17300 13630 17330 13720
rect 17400 13630 17430 13720
rect 17500 13630 17530 13720
rect 17600 13630 17630 13720
rect 17700 13710 17820 13720
rect 17880 13710 17910 13770
rect 17970 13710 18000 13770
rect 18060 13710 18090 13770
rect 18150 13710 18180 13770
rect 18240 13710 18270 13770
rect 18330 13710 18360 13770
rect 18420 13710 18450 13770
rect 18510 13710 18540 13770
rect 18600 13710 18630 13770
rect 18690 13710 18720 13770
rect 18780 13710 18810 13770
rect 18870 13710 18900 13770
rect 18960 13710 18990 13770
rect 19050 13710 19080 13770
rect 19140 13710 19170 13770
rect 19230 13710 19260 13770
rect 19320 13710 19350 13770
rect 19410 13710 19440 13770
rect 19500 13710 19530 13770
rect 19590 13710 19620 13770
rect 19680 13710 19710 13770
rect 19770 13710 19800 13770
rect 19860 13710 19890 13770
rect 19950 13710 19980 13770
rect 20040 13710 20070 13770
rect 20130 13710 20160 13770
rect 20220 13710 20250 13770
rect 20310 13710 20340 13770
rect 20400 13710 20430 13770
rect 20490 13710 20520 13770
rect 20580 13710 20610 13770
rect 20670 13710 20700 13770
rect 20760 13710 20790 13770
rect 20850 13710 20880 13770
rect 20940 13710 20970 13770
rect 21030 13710 21060 13770
rect 21120 13710 21150 13770
rect 21210 13710 21240 13770
rect 21300 13710 21330 13770
rect 21390 13710 21420 13770
rect 21480 13710 21510 13770
rect 21570 13710 21600 13770
rect 21660 13710 21690 13770
rect 21750 13710 21780 13770
rect 21840 13710 21870 13770
rect 21930 13710 21960 13770
rect 22020 13710 22050 13770
rect 22110 13710 22140 13770
rect 22200 13710 22230 13770
rect 22290 13710 22320 13770
rect 22380 13710 22410 13770
rect 22470 13710 22500 13770
rect 22560 13710 22590 13770
rect 22650 13710 22680 13770
rect 22740 13710 22770 13770
rect 22830 13710 22860 13770
rect 22920 13710 22950 13770
rect 23010 13710 23040 13770
rect 23100 13710 23130 13770
rect 23190 13710 23220 13770
rect 23280 13710 23300 13770
rect 17700 13700 23300 13710
rect 17700 13630 17750 13700
rect 17180 13600 17750 13630
rect 11660 12310 17090 12340
rect 11660 12240 11690 12310
rect 11760 12240 11810 12310
rect 11880 12240 12020 12310
rect 12090 12240 12140 12310
rect 12210 12240 12350 12310
rect 12420 12240 12470 12310
rect 12540 12240 12680 12310
rect 12750 12240 12800 12310
rect 12870 12240 13010 12310
rect 13080 12240 13130 12310
rect 13200 12240 13340 12310
rect 13410 12240 13460 12310
rect 13530 12240 13670 12310
rect 13740 12240 13790 12310
rect 13860 12240 14000 12310
rect 14070 12240 14120 12310
rect 14190 12240 14330 12310
rect 14400 12240 14450 12310
rect 14520 12300 15650 12310
rect 14520 12240 14660 12300
rect 11660 12230 14660 12240
rect 14730 12230 14780 12300
rect 14850 12230 14990 12300
rect 15060 12230 15110 12300
rect 15180 12230 15320 12300
rect 15390 12230 15440 12300
rect 15510 12240 15650 12300
rect 15720 12240 15770 12310
rect 15840 12240 15980 12310
rect 16050 12240 16100 12310
rect 16170 12240 16310 12310
rect 16380 12240 16430 12310
rect 16500 12240 16640 12310
rect 16710 12240 16760 12310
rect 16830 12240 17090 12310
rect 15510 12230 17090 12240
rect 11660 12190 17090 12230
rect 11660 12120 11690 12190
rect 11760 12120 11810 12190
rect 11880 12120 12020 12190
rect 12090 12120 12140 12190
rect 12210 12120 12350 12190
rect 12420 12120 12470 12190
rect 12540 12120 12680 12190
rect 12750 12120 12800 12190
rect 12870 12120 13010 12190
rect 13080 12120 13130 12190
rect 13200 12120 13340 12190
rect 13410 12120 13460 12190
rect 13530 12120 13670 12190
rect 13740 12120 13790 12190
rect 13860 12120 14000 12190
rect 14070 12120 14120 12190
rect 14190 12120 14330 12190
rect 14400 12120 14450 12190
rect 14520 12180 15650 12190
rect 14520 12120 14660 12180
rect 11660 12110 14660 12120
rect 14730 12110 14780 12180
rect 14850 12110 14990 12180
rect 15060 12110 15110 12180
rect 15180 12110 15320 12180
rect 15390 12110 15440 12180
rect 15510 12120 15650 12180
rect 15720 12120 15770 12190
rect 15840 12120 15980 12190
rect 16050 12120 16100 12190
rect 16170 12120 16310 12190
rect 16380 12120 16430 12190
rect 16500 12120 16640 12190
rect 16710 12120 16760 12190
rect 16830 12120 17090 12190
rect 15510 12110 17090 12120
rect 11660 12090 17090 12110
rect 17840 12310 23270 12340
rect 17840 12240 18100 12310
rect 18170 12240 18220 12310
rect 18290 12240 18430 12310
rect 18500 12240 18550 12310
rect 18620 12240 18760 12310
rect 18830 12240 18880 12310
rect 18950 12240 19090 12310
rect 19160 12240 19210 12310
rect 19280 12300 20410 12310
rect 19280 12240 19420 12300
rect 17840 12230 19420 12240
rect 19490 12230 19540 12300
rect 19610 12230 19750 12300
rect 19820 12230 19870 12300
rect 19940 12230 20080 12300
rect 20150 12230 20200 12300
rect 20270 12240 20410 12300
rect 20480 12240 20530 12310
rect 20600 12240 20740 12310
rect 20810 12240 20860 12310
rect 20930 12240 21070 12310
rect 21140 12240 21190 12310
rect 21260 12240 21400 12310
rect 21470 12240 21520 12310
rect 21590 12240 21730 12310
rect 21800 12240 21850 12310
rect 21920 12240 22060 12310
rect 22130 12240 22180 12310
rect 22250 12240 22390 12310
rect 22460 12240 22510 12310
rect 22580 12240 22720 12310
rect 22790 12240 22840 12310
rect 22910 12240 23050 12310
rect 23120 12240 23170 12310
rect 23240 12240 23270 12310
rect 20270 12230 23270 12240
rect 17840 12190 23270 12230
rect 17840 12120 18100 12190
rect 18170 12120 18220 12190
rect 18290 12120 18430 12190
rect 18500 12120 18550 12190
rect 18620 12120 18760 12190
rect 18830 12120 18880 12190
rect 18950 12120 19090 12190
rect 19160 12120 19210 12190
rect 19280 12180 20410 12190
rect 19280 12120 19420 12180
rect 17840 12110 19420 12120
rect 19490 12110 19540 12180
rect 19610 12110 19750 12180
rect 19820 12110 19870 12180
rect 19940 12110 20080 12180
rect 20150 12110 20200 12180
rect 20270 12120 20410 12180
rect 20480 12120 20530 12190
rect 20600 12120 20740 12190
rect 20810 12120 20860 12190
rect 20930 12120 21070 12190
rect 21140 12120 21190 12190
rect 21260 12120 21400 12190
rect 21470 12120 21520 12190
rect 21590 12120 21730 12190
rect 21800 12120 21850 12190
rect 21920 12120 22060 12190
rect 22130 12120 22180 12190
rect 22250 12120 22390 12190
rect 22460 12120 22510 12190
rect 22580 12120 22720 12190
rect 22790 12120 22840 12190
rect 22910 12120 23050 12190
rect 23120 12120 23170 12190
rect 23240 12120 23270 12190
rect 20270 12110 23270 12120
rect 17840 12090 23270 12110
rect 11690 12070 11930 12090
rect 12020 12070 12260 12090
rect 12350 12070 12590 12090
rect 12680 12070 12920 12090
rect 13010 12070 13250 12090
rect 13340 12070 13580 12090
rect 13670 12070 13910 12090
rect 14000 12070 14240 12090
rect 14330 12070 14570 12090
rect 14660 12070 14900 12090
rect 14990 12070 15230 12090
rect 15320 12070 15560 12090
rect 15650 12070 15890 12090
rect 15980 12070 16220 12090
rect 16310 12070 16550 12090
rect 16640 12070 16880 12090
rect 18050 12070 18290 12090
rect 18380 12070 18620 12090
rect 18710 12070 18950 12090
rect 19040 12070 19280 12090
rect 19370 12070 19610 12090
rect 19700 12070 19940 12090
rect 20030 12070 20270 12090
rect 20360 12070 20600 12090
rect 20690 12070 20930 12090
rect 21020 12070 21260 12090
rect 21350 12070 21590 12090
rect 21680 12070 21920 12090
rect 22010 12070 22250 12090
rect 22340 12070 22580 12090
rect 22670 12070 22910 12090
rect 23000 12070 23240 12090
<< via3 >>
rect 11690 17490 11760 17560
rect 11810 17490 11880 17560
rect 12020 17490 12090 17560
rect 12140 17490 12210 17560
rect 12350 17490 12420 17560
rect 12470 17490 12540 17560
rect 12680 17490 12750 17560
rect 12800 17490 12870 17560
rect 13010 17490 13080 17560
rect 13130 17490 13200 17560
rect 13340 17490 13410 17560
rect 13460 17490 13530 17560
rect 13670 17490 13740 17560
rect 13790 17490 13860 17560
rect 14000 17490 14070 17560
rect 14120 17490 14190 17560
rect 14330 17490 14400 17560
rect 14450 17490 14520 17560
rect 14660 17500 14730 17570
rect 14780 17500 14850 17570
rect 14990 17500 15060 17570
rect 15110 17500 15180 17570
rect 15320 17500 15390 17570
rect 15440 17500 15510 17570
rect 15650 17490 15720 17560
rect 15770 17490 15840 17560
rect 15980 17490 16050 17560
rect 16100 17490 16170 17560
rect 16310 17490 16380 17560
rect 16430 17490 16500 17560
rect 16640 17490 16710 17560
rect 16760 17490 16830 17560
rect 11690 17370 11760 17440
rect 11810 17370 11880 17440
rect 12020 17370 12090 17440
rect 12140 17370 12210 17440
rect 12350 17370 12420 17440
rect 12470 17370 12540 17440
rect 12680 17370 12750 17440
rect 12800 17370 12870 17440
rect 13010 17370 13080 17440
rect 13130 17370 13200 17440
rect 13340 17370 13410 17440
rect 13460 17370 13530 17440
rect 13670 17370 13740 17440
rect 13790 17370 13860 17440
rect 14000 17370 14070 17440
rect 14120 17370 14190 17440
rect 14330 17370 14400 17440
rect 14450 17370 14520 17440
rect 14660 17380 14730 17450
rect 14780 17380 14850 17450
rect 14990 17380 15060 17450
rect 15110 17380 15180 17450
rect 15320 17380 15390 17450
rect 15440 17380 15510 17450
rect 15650 17370 15720 17440
rect 15770 17370 15840 17440
rect 15980 17370 16050 17440
rect 16100 17370 16170 17440
rect 16310 17370 16380 17440
rect 16430 17370 16500 17440
rect 16640 17370 16710 17440
rect 16760 17370 16830 17440
rect 18100 17490 18170 17560
rect 18220 17490 18290 17560
rect 18430 17490 18500 17560
rect 18550 17490 18620 17560
rect 18760 17490 18830 17560
rect 18880 17490 18950 17560
rect 19090 17490 19160 17560
rect 19210 17490 19280 17560
rect 19420 17500 19490 17570
rect 19540 17500 19610 17570
rect 19750 17500 19820 17570
rect 19870 17500 19940 17570
rect 20080 17500 20150 17570
rect 20200 17500 20270 17570
rect 20410 17490 20480 17560
rect 20530 17490 20600 17560
rect 20740 17490 20810 17560
rect 20860 17490 20930 17560
rect 21070 17490 21140 17560
rect 21190 17490 21260 17560
rect 21400 17490 21470 17560
rect 21520 17490 21590 17560
rect 21730 17490 21800 17560
rect 21850 17490 21920 17560
rect 22060 17490 22130 17560
rect 22180 17490 22250 17560
rect 22390 17490 22460 17560
rect 22510 17490 22580 17560
rect 22720 17490 22790 17560
rect 22840 17490 22910 17560
rect 23050 17490 23120 17560
rect 23170 17490 23240 17560
rect 18100 17370 18170 17440
rect 18220 17370 18290 17440
rect 18430 17370 18500 17440
rect 18550 17370 18620 17440
rect 18760 17370 18830 17440
rect 18880 17370 18950 17440
rect 19090 17370 19160 17440
rect 19210 17370 19280 17440
rect 19420 17380 19490 17450
rect 19540 17380 19610 17450
rect 19750 17380 19820 17450
rect 19870 17380 19940 17450
rect 20080 17380 20150 17450
rect 20200 17380 20270 17450
rect 20410 17370 20480 17440
rect 20530 17370 20600 17440
rect 20740 17370 20810 17440
rect 20860 17370 20930 17440
rect 21070 17370 21140 17440
rect 21190 17370 21260 17440
rect 21400 17370 21470 17440
rect 21520 17370 21590 17440
rect 21730 17370 21800 17440
rect 21850 17370 21920 17440
rect 22060 17370 22130 17440
rect 22180 17370 22250 17440
rect 22390 17370 22460 17440
rect 22510 17370 22580 17440
rect 22720 17370 22790 17440
rect 22840 17370 22910 17440
rect 23050 17370 23120 17440
rect 23170 17370 23240 17440
rect 17230 15980 17300 16070
rect 17330 15980 17400 16070
rect 17430 15980 17500 16070
rect 17530 15980 17600 16070
rect 17630 15980 17700 16070
rect 17230 15850 17300 15940
rect 17330 15850 17400 15940
rect 17430 15850 17500 15940
rect 17530 15850 17600 15940
rect 17630 15850 17700 15940
rect 17230 13760 17300 13850
rect 17330 13760 17400 13850
rect 17430 13760 17500 13850
rect 17530 13760 17600 13850
rect 17630 13760 17700 13850
rect 17230 13630 17300 13720
rect 17330 13630 17400 13720
rect 17430 13630 17500 13720
rect 17530 13630 17600 13720
rect 17630 13630 17700 13720
rect 11690 12240 11760 12310
rect 11810 12240 11880 12310
rect 12020 12240 12090 12310
rect 12140 12240 12210 12310
rect 12350 12240 12420 12310
rect 12470 12240 12540 12310
rect 12680 12240 12750 12310
rect 12800 12240 12870 12310
rect 13010 12240 13080 12310
rect 13130 12240 13200 12310
rect 13340 12240 13410 12310
rect 13460 12240 13530 12310
rect 13670 12240 13740 12310
rect 13790 12240 13860 12310
rect 14000 12240 14070 12310
rect 14120 12240 14190 12310
rect 14330 12240 14400 12310
rect 14450 12240 14520 12310
rect 14660 12230 14730 12300
rect 14780 12230 14850 12300
rect 14990 12230 15060 12300
rect 15110 12230 15180 12300
rect 15320 12230 15390 12300
rect 15440 12230 15510 12300
rect 15650 12240 15720 12310
rect 15770 12240 15840 12310
rect 15980 12240 16050 12310
rect 16100 12240 16170 12310
rect 16310 12240 16380 12310
rect 16430 12240 16500 12310
rect 16640 12240 16710 12310
rect 16760 12240 16830 12310
rect 11690 12120 11760 12190
rect 11810 12120 11880 12190
rect 12020 12120 12090 12190
rect 12140 12120 12210 12190
rect 12350 12120 12420 12190
rect 12470 12120 12540 12190
rect 12680 12120 12750 12190
rect 12800 12120 12870 12190
rect 13010 12120 13080 12190
rect 13130 12120 13200 12190
rect 13340 12120 13410 12190
rect 13460 12120 13530 12190
rect 13670 12120 13740 12190
rect 13790 12120 13860 12190
rect 14000 12120 14070 12190
rect 14120 12120 14190 12190
rect 14330 12120 14400 12190
rect 14450 12120 14520 12190
rect 14660 12110 14730 12180
rect 14780 12110 14850 12180
rect 14990 12110 15060 12180
rect 15110 12110 15180 12180
rect 15320 12110 15390 12180
rect 15440 12110 15510 12180
rect 15650 12120 15720 12190
rect 15770 12120 15840 12190
rect 15980 12120 16050 12190
rect 16100 12120 16170 12190
rect 16310 12120 16380 12190
rect 16430 12120 16500 12190
rect 16640 12120 16710 12190
rect 16760 12120 16830 12190
rect 18100 12240 18170 12310
rect 18220 12240 18290 12310
rect 18430 12240 18500 12310
rect 18550 12240 18620 12310
rect 18760 12240 18830 12310
rect 18880 12240 18950 12310
rect 19090 12240 19160 12310
rect 19210 12240 19280 12310
rect 19420 12230 19490 12300
rect 19540 12230 19610 12300
rect 19750 12230 19820 12300
rect 19870 12230 19940 12300
rect 20080 12230 20150 12300
rect 20200 12230 20270 12300
rect 20410 12240 20480 12310
rect 20530 12240 20600 12310
rect 20740 12240 20810 12310
rect 20860 12240 20930 12310
rect 21070 12240 21140 12310
rect 21190 12240 21260 12310
rect 21400 12240 21470 12310
rect 21520 12240 21590 12310
rect 21730 12240 21800 12310
rect 21850 12240 21920 12310
rect 22060 12240 22130 12310
rect 22180 12240 22250 12310
rect 22390 12240 22460 12310
rect 22510 12240 22580 12310
rect 22720 12240 22790 12310
rect 22840 12240 22910 12310
rect 23050 12240 23120 12310
rect 23170 12240 23240 12310
rect 18100 12120 18170 12190
rect 18220 12120 18290 12190
rect 18430 12120 18500 12190
rect 18550 12120 18620 12190
rect 18760 12120 18830 12190
rect 18880 12120 18950 12190
rect 19090 12120 19160 12190
rect 19210 12120 19280 12190
rect 19420 12110 19490 12180
rect 19540 12110 19610 12180
rect 19750 12110 19820 12180
rect 19870 12110 19940 12180
rect 20080 12110 20150 12180
rect 20200 12110 20270 12180
rect 20410 12120 20480 12190
rect 20530 12120 20600 12190
rect 20740 12120 20810 12190
rect 20860 12120 20930 12190
rect 21070 12120 21140 12190
rect 21190 12120 21260 12190
rect 21400 12120 21470 12190
rect 21520 12120 21590 12190
rect 21730 12120 21800 12190
rect 21850 12120 21920 12190
rect 22060 12120 22130 12190
rect 22180 12120 22250 12190
rect 22390 12120 22460 12190
rect 22510 12120 22580 12190
rect 22720 12120 22790 12190
rect 22840 12120 22910 12190
rect 23050 12120 23120 12190
rect 23170 12120 23240 12190
<< metal4 >>
rect 11660 17610 17090 17660
rect 11660 17370 11690 17610
rect 11930 17370 12020 17610
rect 12260 17370 12350 17610
rect 12590 17370 12680 17610
rect 12920 17370 13010 17610
rect 13250 17370 13340 17610
rect 13580 17370 13670 17610
rect 13910 17370 14000 17610
rect 14240 17370 14330 17610
rect 14570 17370 14660 17610
rect 14900 17370 14990 17610
rect 15230 17370 15320 17610
rect 15560 17370 15650 17610
rect 15890 17370 15980 17610
rect 16220 17370 16310 17610
rect 16550 17370 16640 17610
rect 16880 17370 17090 17610
rect 11660 17340 17090 17370
rect 17180 16070 17750 18230
rect 17840 17610 23270 17660
rect 17840 17370 18050 17610
rect 18290 17370 18380 17610
rect 18620 17370 18710 17610
rect 18950 17370 19040 17610
rect 19280 17370 19370 17610
rect 19610 17370 19700 17610
rect 19940 17370 20030 17610
rect 20270 17370 20360 17610
rect 20600 17370 20690 17610
rect 20930 17370 21020 17610
rect 21260 17370 21350 17610
rect 21590 17370 21680 17610
rect 21920 17370 22010 17610
rect 22250 17370 22340 17610
rect 22580 17370 22670 17610
rect 22910 17370 23000 17610
rect 23240 17370 23270 17610
rect 17840 17340 23270 17370
rect 17180 15980 17230 16070
rect 17300 15980 17330 16070
rect 17400 15980 17430 16070
rect 17500 15980 17530 16070
rect 17600 15980 17630 16070
rect 17700 15980 17750 16070
rect 17180 15940 17750 15980
rect 17180 15850 17230 15940
rect 17300 15850 17330 15940
rect 17400 15850 17430 15940
rect 17500 15850 17530 15940
rect 17600 15850 17630 15940
rect 17700 15850 17750 15940
rect 17180 15820 17750 15850
rect 17180 13850 17750 13880
rect 17180 13760 17230 13850
rect 17300 13760 17330 13850
rect 17400 13760 17430 13850
rect 17500 13760 17530 13850
rect 17600 13760 17630 13850
rect 17700 13760 17750 13850
rect 17180 13720 17750 13760
rect 17180 13630 17230 13720
rect 17300 13630 17330 13720
rect 17400 13630 17430 13720
rect 17500 13630 17530 13720
rect 17600 13630 17630 13720
rect 17700 13630 17750 13720
rect 11660 12310 17090 12340
rect 11660 12070 11690 12310
rect 11930 12070 12020 12310
rect 12260 12070 12350 12310
rect 12590 12070 12680 12310
rect 12920 12070 13010 12310
rect 13250 12070 13340 12310
rect 13580 12070 13670 12310
rect 13910 12070 14000 12310
rect 14240 12070 14330 12310
rect 14570 12070 14660 12310
rect 14900 12070 14990 12310
rect 15230 12070 15320 12310
rect 15560 12070 15650 12310
rect 15890 12070 15980 12310
rect 16220 12070 16310 12310
rect 16550 12070 16640 12310
rect 16880 12070 17090 12310
rect 11660 12020 17090 12070
rect 17180 11470 17750 13630
rect 17840 12310 23270 12340
rect 17840 12070 18050 12310
rect 18290 12070 18380 12310
rect 18620 12070 18710 12310
rect 18950 12070 19040 12310
rect 19280 12070 19370 12310
rect 19610 12070 19700 12310
rect 19940 12070 20030 12310
rect 20270 12070 20360 12310
rect 20600 12070 20690 12310
rect 20930 12070 21020 12310
rect 21260 12070 21350 12310
rect 21590 12070 21680 12310
rect 21920 12070 22010 12310
rect 22250 12070 22340 12310
rect 22580 12070 22670 12310
rect 22910 12070 23000 12310
rect 23240 12070 23270 12310
rect 17840 12020 23270 12070
<< via4 >>
rect 11690 17560 11930 17610
rect 11690 17490 11760 17560
rect 11760 17490 11810 17560
rect 11810 17490 11880 17560
rect 11880 17490 11930 17560
rect 11690 17440 11930 17490
rect 11690 17370 11760 17440
rect 11760 17370 11810 17440
rect 11810 17370 11880 17440
rect 11880 17370 11930 17440
rect 12020 17560 12260 17610
rect 12020 17490 12090 17560
rect 12090 17490 12140 17560
rect 12140 17490 12210 17560
rect 12210 17490 12260 17560
rect 12020 17440 12260 17490
rect 12020 17370 12090 17440
rect 12090 17370 12140 17440
rect 12140 17370 12210 17440
rect 12210 17370 12260 17440
rect 12350 17560 12590 17610
rect 12350 17490 12420 17560
rect 12420 17490 12470 17560
rect 12470 17490 12540 17560
rect 12540 17490 12590 17560
rect 12350 17440 12590 17490
rect 12350 17370 12420 17440
rect 12420 17370 12470 17440
rect 12470 17370 12540 17440
rect 12540 17370 12590 17440
rect 12680 17560 12920 17610
rect 12680 17490 12750 17560
rect 12750 17490 12800 17560
rect 12800 17490 12870 17560
rect 12870 17490 12920 17560
rect 12680 17440 12920 17490
rect 12680 17370 12750 17440
rect 12750 17370 12800 17440
rect 12800 17370 12870 17440
rect 12870 17370 12920 17440
rect 13010 17560 13250 17610
rect 13010 17490 13080 17560
rect 13080 17490 13130 17560
rect 13130 17490 13200 17560
rect 13200 17490 13250 17560
rect 13010 17440 13250 17490
rect 13010 17370 13080 17440
rect 13080 17370 13130 17440
rect 13130 17370 13200 17440
rect 13200 17370 13250 17440
rect 13340 17560 13580 17610
rect 13340 17490 13410 17560
rect 13410 17490 13460 17560
rect 13460 17490 13530 17560
rect 13530 17490 13580 17560
rect 13340 17440 13580 17490
rect 13340 17370 13410 17440
rect 13410 17370 13460 17440
rect 13460 17370 13530 17440
rect 13530 17370 13580 17440
rect 13670 17560 13910 17610
rect 13670 17490 13740 17560
rect 13740 17490 13790 17560
rect 13790 17490 13860 17560
rect 13860 17490 13910 17560
rect 13670 17440 13910 17490
rect 13670 17370 13740 17440
rect 13740 17370 13790 17440
rect 13790 17370 13860 17440
rect 13860 17370 13910 17440
rect 14000 17560 14240 17610
rect 14000 17490 14070 17560
rect 14070 17490 14120 17560
rect 14120 17490 14190 17560
rect 14190 17490 14240 17560
rect 14000 17440 14240 17490
rect 14000 17370 14070 17440
rect 14070 17370 14120 17440
rect 14120 17370 14190 17440
rect 14190 17370 14240 17440
rect 14330 17560 14570 17610
rect 14330 17490 14400 17560
rect 14400 17490 14450 17560
rect 14450 17490 14520 17560
rect 14520 17490 14570 17560
rect 14330 17440 14570 17490
rect 14330 17370 14400 17440
rect 14400 17370 14450 17440
rect 14450 17370 14520 17440
rect 14520 17370 14570 17440
rect 14660 17570 14900 17610
rect 14660 17500 14730 17570
rect 14730 17500 14780 17570
rect 14780 17500 14850 17570
rect 14850 17500 14900 17570
rect 14660 17450 14900 17500
rect 14660 17380 14730 17450
rect 14730 17380 14780 17450
rect 14780 17380 14850 17450
rect 14850 17380 14900 17450
rect 14660 17370 14900 17380
rect 14990 17570 15230 17610
rect 14990 17500 15060 17570
rect 15060 17500 15110 17570
rect 15110 17500 15180 17570
rect 15180 17500 15230 17570
rect 14990 17450 15230 17500
rect 14990 17380 15060 17450
rect 15060 17380 15110 17450
rect 15110 17380 15180 17450
rect 15180 17380 15230 17450
rect 14990 17370 15230 17380
rect 15320 17570 15560 17610
rect 15320 17500 15390 17570
rect 15390 17500 15440 17570
rect 15440 17500 15510 17570
rect 15510 17500 15560 17570
rect 15320 17450 15560 17500
rect 15320 17380 15390 17450
rect 15390 17380 15440 17450
rect 15440 17380 15510 17450
rect 15510 17380 15560 17450
rect 15320 17370 15560 17380
rect 15650 17560 15890 17610
rect 15650 17490 15720 17560
rect 15720 17490 15770 17560
rect 15770 17490 15840 17560
rect 15840 17490 15890 17560
rect 15650 17440 15890 17490
rect 15650 17370 15720 17440
rect 15720 17370 15770 17440
rect 15770 17370 15840 17440
rect 15840 17370 15890 17440
rect 15980 17560 16220 17610
rect 15980 17490 16050 17560
rect 16050 17490 16100 17560
rect 16100 17490 16170 17560
rect 16170 17490 16220 17560
rect 15980 17440 16220 17490
rect 15980 17370 16050 17440
rect 16050 17370 16100 17440
rect 16100 17370 16170 17440
rect 16170 17370 16220 17440
rect 16310 17560 16550 17610
rect 16310 17490 16380 17560
rect 16380 17490 16430 17560
rect 16430 17490 16500 17560
rect 16500 17490 16550 17560
rect 16310 17440 16550 17490
rect 16310 17370 16380 17440
rect 16380 17370 16430 17440
rect 16430 17370 16500 17440
rect 16500 17370 16550 17440
rect 16640 17560 16880 17610
rect 16640 17490 16710 17560
rect 16710 17490 16760 17560
rect 16760 17490 16830 17560
rect 16830 17490 16880 17560
rect 16640 17440 16880 17490
rect 16640 17370 16710 17440
rect 16710 17370 16760 17440
rect 16760 17370 16830 17440
rect 16830 17370 16880 17440
rect 18050 17560 18290 17610
rect 18050 17490 18100 17560
rect 18100 17490 18170 17560
rect 18170 17490 18220 17560
rect 18220 17490 18290 17560
rect 18050 17440 18290 17490
rect 18050 17370 18100 17440
rect 18100 17370 18170 17440
rect 18170 17370 18220 17440
rect 18220 17370 18290 17440
rect 18380 17560 18620 17610
rect 18380 17490 18430 17560
rect 18430 17490 18500 17560
rect 18500 17490 18550 17560
rect 18550 17490 18620 17560
rect 18380 17440 18620 17490
rect 18380 17370 18430 17440
rect 18430 17370 18500 17440
rect 18500 17370 18550 17440
rect 18550 17370 18620 17440
rect 18710 17560 18950 17610
rect 18710 17490 18760 17560
rect 18760 17490 18830 17560
rect 18830 17490 18880 17560
rect 18880 17490 18950 17560
rect 18710 17440 18950 17490
rect 18710 17370 18760 17440
rect 18760 17370 18830 17440
rect 18830 17370 18880 17440
rect 18880 17370 18950 17440
rect 19040 17560 19280 17610
rect 19040 17490 19090 17560
rect 19090 17490 19160 17560
rect 19160 17490 19210 17560
rect 19210 17490 19280 17560
rect 19040 17440 19280 17490
rect 19040 17370 19090 17440
rect 19090 17370 19160 17440
rect 19160 17370 19210 17440
rect 19210 17370 19280 17440
rect 19370 17570 19610 17610
rect 19370 17500 19420 17570
rect 19420 17500 19490 17570
rect 19490 17500 19540 17570
rect 19540 17500 19610 17570
rect 19370 17450 19610 17500
rect 19370 17380 19420 17450
rect 19420 17380 19490 17450
rect 19490 17380 19540 17450
rect 19540 17380 19610 17450
rect 19370 17370 19610 17380
rect 19700 17570 19940 17610
rect 19700 17500 19750 17570
rect 19750 17500 19820 17570
rect 19820 17500 19870 17570
rect 19870 17500 19940 17570
rect 19700 17450 19940 17500
rect 19700 17380 19750 17450
rect 19750 17380 19820 17450
rect 19820 17380 19870 17450
rect 19870 17380 19940 17450
rect 19700 17370 19940 17380
rect 20030 17570 20270 17610
rect 20030 17500 20080 17570
rect 20080 17500 20150 17570
rect 20150 17500 20200 17570
rect 20200 17500 20270 17570
rect 20030 17450 20270 17500
rect 20030 17380 20080 17450
rect 20080 17380 20150 17450
rect 20150 17380 20200 17450
rect 20200 17380 20270 17450
rect 20030 17370 20270 17380
rect 20360 17560 20600 17610
rect 20360 17490 20410 17560
rect 20410 17490 20480 17560
rect 20480 17490 20530 17560
rect 20530 17490 20600 17560
rect 20360 17440 20600 17490
rect 20360 17370 20410 17440
rect 20410 17370 20480 17440
rect 20480 17370 20530 17440
rect 20530 17370 20600 17440
rect 20690 17560 20930 17610
rect 20690 17490 20740 17560
rect 20740 17490 20810 17560
rect 20810 17490 20860 17560
rect 20860 17490 20930 17560
rect 20690 17440 20930 17490
rect 20690 17370 20740 17440
rect 20740 17370 20810 17440
rect 20810 17370 20860 17440
rect 20860 17370 20930 17440
rect 21020 17560 21260 17610
rect 21020 17490 21070 17560
rect 21070 17490 21140 17560
rect 21140 17490 21190 17560
rect 21190 17490 21260 17560
rect 21020 17440 21260 17490
rect 21020 17370 21070 17440
rect 21070 17370 21140 17440
rect 21140 17370 21190 17440
rect 21190 17370 21260 17440
rect 21350 17560 21590 17610
rect 21350 17490 21400 17560
rect 21400 17490 21470 17560
rect 21470 17490 21520 17560
rect 21520 17490 21590 17560
rect 21350 17440 21590 17490
rect 21350 17370 21400 17440
rect 21400 17370 21470 17440
rect 21470 17370 21520 17440
rect 21520 17370 21590 17440
rect 21680 17560 21920 17610
rect 21680 17490 21730 17560
rect 21730 17490 21800 17560
rect 21800 17490 21850 17560
rect 21850 17490 21920 17560
rect 21680 17440 21920 17490
rect 21680 17370 21730 17440
rect 21730 17370 21800 17440
rect 21800 17370 21850 17440
rect 21850 17370 21920 17440
rect 22010 17560 22250 17610
rect 22010 17490 22060 17560
rect 22060 17490 22130 17560
rect 22130 17490 22180 17560
rect 22180 17490 22250 17560
rect 22010 17440 22250 17490
rect 22010 17370 22060 17440
rect 22060 17370 22130 17440
rect 22130 17370 22180 17440
rect 22180 17370 22250 17440
rect 22340 17560 22580 17610
rect 22340 17490 22390 17560
rect 22390 17490 22460 17560
rect 22460 17490 22510 17560
rect 22510 17490 22580 17560
rect 22340 17440 22580 17490
rect 22340 17370 22390 17440
rect 22390 17370 22460 17440
rect 22460 17370 22510 17440
rect 22510 17370 22580 17440
rect 22670 17560 22910 17610
rect 22670 17490 22720 17560
rect 22720 17490 22790 17560
rect 22790 17490 22840 17560
rect 22840 17490 22910 17560
rect 22670 17440 22910 17490
rect 22670 17370 22720 17440
rect 22720 17370 22790 17440
rect 22790 17370 22840 17440
rect 22840 17370 22910 17440
rect 23000 17560 23240 17610
rect 23000 17490 23050 17560
rect 23050 17490 23120 17560
rect 23120 17490 23170 17560
rect 23170 17490 23240 17560
rect 23000 17440 23240 17490
rect 23000 17370 23050 17440
rect 23050 17370 23120 17440
rect 23120 17370 23170 17440
rect 23170 17370 23240 17440
rect 11690 12240 11760 12310
rect 11760 12240 11810 12310
rect 11810 12240 11880 12310
rect 11880 12240 11930 12310
rect 11690 12190 11930 12240
rect 11690 12120 11760 12190
rect 11760 12120 11810 12190
rect 11810 12120 11880 12190
rect 11880 12120 11930 12190
rect 11690 12070 11930 12120
rect 12020 12240 12090 12310
rect 12090 12240 12140 12310
rect 12140 12240 12210 12310
rect 12210 12240 12260 12310
rect 12020 12190 12260 12240
rect 12020 12120 12090 12190
rect 12090 12120 12140 12190
rect 12140 12120 12210 12190
rect 12210 12120 12260 12190
rect 12020 12070 12260 12120
rect 12350 12240 12420 12310
rect 12420 12240 12470 12310
rect 12470 12240 12540 12310
rect 12540 12240 12590 12310
rect 12350 12190 12590 12240
rect 12350 12120 12420 12190
rect 12420 12120 12470 12190
rect 12470 12120 12540 12190
rect 12540 12120 12590 12190
rect 12350 12070 12590 12120
rect 12680 12240 12750 12310
rect 12750 12240 12800 12310
rect 12800 12240 12870 12310
rect 12870 12240 12920 12310
rect 12680 12190 12920 12240
rect 12680 12120 12750 12190
rect 12750 12120 12800 12190
rect 12800 12120 12870 12190
rect 12870 12120 12920 12190
rect 12680 12070 12920 12120
rect 13010 12240 13080 12310
rect 13080 12240 13130 12310
rect 13130 12240 13200 12310
rect 13200 12240 13250 12310
rect 13010 12190 13250 12240
rect 13010 12120 13080 12190
rect 13080 12120 13130 12190
rect 13130 12120 13200 12190
rect 13200 12120 13250 12190
rect 13010 12070 13250 12120
rect 13340 12240 13410 12310
rect 13410 12240 13460 12310
rect 13460 12240 13530 12310
rect 13530 12240 13580 12310
rect 13340 12190 13580 12240
rect 13340 12120 13410 12190
rect 13410 12120 13460 12190
rect 13460 12120 13530 12190
rect 13530 12120 13580 12190
rect 13340 12070 13580 12120
rect 13670 12240 13740 12310
rect 13740 12240 13790 12310
rect 13790 12240 13860 12310
rect 13860 12240 13910 12310
rect 13670 12190 13910 12240
rect 13670 12120 13740 12190
rect 13740 12120 13790 12190
rect 13790 12120 13860 12190
rect 13860 12120 13910 12190
rect 13670 12070 13910 12120
rect 14000 12240 14070 12310
rect 14070 12240 14120 12310
rect 14120 12240 14190 12310
rect 14190 12240 14240 12310
rect 14000 12190 14240 12240
rect 14000 12120 14070 12190
rect 14070 12120 14120 12190
rect 14120 12120 14190 12190
rect 14190 12120 14240 12190
rect 14000 12070 14240 12120
rect 14330 12240 14400 12310
rect 14400 12240 14450 12310
rect 14450 12240 14520 12310
rect 14520 12240 14570 12310
rect 14330 12190 14570 12240
rect 14330 12120 14400 12190
rect 14400 12120 14450 12190
rect 14450 12120 14520 12190
rect 14520 12120 14570 12190
rect 14330 12070 14570 12120
rect 14660 12300 14900 12310
rect 14660 12230 14730 12300
rect 14730 12230 14780 12300
rect 14780 12230 14850 12300
rect 14850 12230 14900 12300
rect 14660 12180 14900 12230
rect 14660 12110 14730 12180
rect 14730 12110 14780 12180
rect 14780 12110 14850 12180
rect 14850 12110 14900 12180
rect 14660 12070 14900 12110
rect 14990 12300 15230 12310
rect 14990 12230 15060 12300
rect 15060 12230 15110 12300
rect 15110 12230 15180 12300
rect 15180 12230 15230 12300
rect 14990 12180 15230 12230
rect 14990 12110 15060 12180
rect 15060 12110 15110 12180
rect 15110 12110 15180 12180
rect 15180 12110 15230 12180
rect 14990 12070 15230 12110
rect 15320 12300 15560 12310
rect 15320 12230 15390 12300
rect 15390 12230 15440 12300
rect 15440 12230 15510 12300
rect 15510 12230 15560 12300
rect 15320 12180 15560 12230
rect 15320 12110 15390 12180
rect 15390 12110 15440 12180
rect 15440 12110 15510 12180
rect 15510 12110 15560 12180
rect 15320 12070 15560 12110
rect 15650 12240 15720 12310
rect 15720 12240 15770 12310
rect 15770 12240 15840 12310
rect 15840 12240 15890 12310
rect 15650 12190 15890 12240
rect 15650 12120 15720 12190
rect 15720 12120 15770 12190
rect 15770 12120 15840 12190
rect 15840 12120 15890 12190
rect 15650 12070 15890 12120
rect 15980 12240 16050 12310
rect 16050 12240 16100 12310
rect 16100 12240 16170 12310
rect 16170 12240 16220 12310
rect 15980 12190 16220 12240
rect 15980 12120 16050 12190
rect 16050 12120 16100 12190
rect 16100 12120 16170 12190
rect 16170 12120 16220 12190
rect 15980 12070 16220 12120
rect 16310 12240 16380 12310
rect 16380 12240 16430 12310
rect 16430 12240 16500 12310
rect 16500 12240 16550 12310
rect 16310 12190 16550 12240
rect 16310 12120 16380 12190
rect 16380 12120 16430 12190
rect 16430 12120 16500 12190
rect 16500 12120 16550 12190
rect 16310 12070 16550 12120
rect 16640 12240 16710 12310
rect 16710 12240 16760 12310
rect 16760 12240 16830 12310
rect 16830 12240 16880 12310
rect 16640 12190 16880 12240
rect 16640 12120 16710 12190
rect 16710 12120 16760 12190
rect 16760 12120 16830 12190
rect 16830 12120 16880 12190
rect 16640 12070 16880 12120
rect 18050 12240 18100 12310
rect 18100 12240 18170 12310
rect 18170 12240 18220 12310
rect 18220 12240 18290 12310
rect 18050 12190 18290 12240
rect 18050 12120 18100 12190
rect 18100 12120 18170 12190
rect 18170 12120 18220 12190
rect 18220 12120 18290 12190
rect 18050 12070 18290 12120
rect 18380 12240 18430 12310
rect 18430 12240 18500 12310
rect 18500 12240 18550 12310
rect 18550 12240 18620 12310
rect 18380 12190 18620 12240
rect 18380 12120 18430 12190
rect 18430 12120 18500 12190
rect 18500 12120 18550 12190
rect 18550 12120 18620 12190
rect 18380 12070 18620 12120
rect 18710 12240 18760 12310
rect 18760 12240 18830 12310
rect 18830 12240 18880 12310
rect 18880 12240 18950 12310
rect 18710 12190 18950 12240
rect 18710 12120 18760 12190
rect 18760 12120 18830 12190
rect 18830 12120 18880 12190
rect 18880 12120 18950 12190
rect 18710 12070 18950 12120
rect 19040 12240 19090 12310
rect 19090 12240 19160 12310
rect 19160 12240 19210 12310
rect 19210 12240 19280 12310
rect 19040 12190 19280 12240
rect 19040 12120 19090 12190
rect 19090 12120 19160 12190
rect 19160 12120 19210 12190
rect 19210 12120 19280 12190
rect 19040 12070 19280 12120
rect 19370 12300 19610 12310
rect 19370 12230 19420 12300
rect 19420 12230 19490 12300
rect 19490 12230 19540 12300
rect 19540 12230 19610 12300
rect 19370 12180 19610 12230
rect 19370 12110 19420 12180
rect 19420 12110 19490 12180
rect 19490 12110 19540 12180
rect 19540 12110 19610 12180
rect 19370 12070 19610 12110
rect 19700 12300 19940 12310
rect 19700 12230 19750 12300
rect 19750 12230 19820 12300
rect 19820 12230 19870 12300
rect 19870 12230 19940 12300
rect 19700 12180 19940 12230
rect 19700 12110 19750 12180
rect 19750 12110 19820 12180
rect 19820 12110 19870 12180
rect 19870 12110 19940 12180
rect 19700 12070 19940 12110
rect 20030 12300 20270 12310
rect 20030 12230 20080 12300
rect 20080 12230 20150 12300
rect 20150 12230 20200 12300
rect 20200 12230 20270 12300
rect 20030 12180 20270 12230
rect 20030 12110 20080 12180
rect 20080 12110 20150 12180
rect 20150 12110 20200 12180
rect 20200 12110 20270 12180
rect 20030 12070 20270 12110
rect 20360 12240 20410 12310
rect 20410 12240 20480 12310
rect 20480 12240 20530 12310
rect 20530 12240 20600 12310
rect 20360 12190 20600 12240
rect 20360 12120 20410 12190
rect 20410 12120 20480 12190
rect 20480 12120 20530 12190
rect 20530 12120 20600 12190
rect 20360 12070 20600 12120
rect 20690 12240 20740 12310
rect 20740 12240 20810 12310
rect 20810 12240 20860 12310
rect 20860 12240 20930 12310
rect 20690 12190 20930 12240
rect 20690 12120 20740 12190
rect 20740 12120 20810 12190
rect 20810 12120 20860 12190
rect 20860 12120 20930 12190
rect 20690 12070 20930 12120
rect 21020 12240 21070 12310
rect 21070 12240 21140 12310
rect 21140 12240 21190 12310
rect 21190 12240 21260 12310
rect 21020 12190 21260 12240
rect 21020 12120 21070 12190
rect 21070 12120 21140 12190
rect 21140 12120 21190 12190
rect 21190 12120 21260 12190
rect 21020 12070 21260 12120
rect 21350 12240 21400 12310
rect 21400 12240 21470 12310
rect 21470 12240 21520 12310
rect 21520 12240 21590 12310
rect 21350 12190 21590 12240
rect 21350 12120 21400 12190
rect 21400 12120 21470 12190
rect 21470 12120 21520 12190
rect 21520 12120 21590 12190
rect 21350 12070 21590 12120
rect 21680 12240 21730 12310
rect 21730 12240 21800 12310
rect 21800 12240 21850 12310
rect 21850 12240 21920 12310
rect 21680 12190 21920 12240
rect 21680 12120 21730 12190
rect 21730 12120 21800 12190
rect 21800 12120 21850 12190
rect 21850 12120 21920 12190
rect 21680 12070 21920 12120
rect 22010 12240 22060 12310
rect 22060 12240 22130 12310
rect 22130 12240 22180 12310
rect 22180 12240 22250 12310
rect 22010 12190 22250 12240
rect 22010 12120 22060 12190
rect 22060 12120 22130 12190
rect 22130 12120 22180 12190
rect 22180 12120 22250 12190
rect 22010 12070 22250 12120
rect 22340 12240 22390 12310
rect 22390 12240 22460 12310
rect 22460 12240 22510 12310
rect 22510 12240 22580 12310
rect 22340 12190 22580 12240
rect 22340 12120 22390 12190
rect 22390 12120 22460 12190
rect 22460 12120 22510 12190
rect 22510 12120 22580 12190
rect 22340 12070 22580 12120
rect 22670 12240 22720 12310
rect 22720 12240 22790 12310
rect 22790 12240 22840 12310
rect 22840 12240 22910 12310
rect 22670 12190 22910 12240
rect 22670 12120 22720 12190
rect 22720 12120 22790 12190
rect 22790 12120 22840 12190
rect 22840 12120 22910 12190
rect 22670 12070 22910 12120
rect 23000 12240 23050 12310
rect 23050 12240 23120 12310
rect 23120 12240 23170 12310
rect 23170 12240 23240 12310
rect 23000 12190 23240 12240
rect 23000 12120 23050 12190
rect 23050 12120 23120 12190
rect 23120 12120 23170 12190
rect 23170 12120 23240 12190
rect 23000 12070 23240 12120
<< metal5 >>
rect 11660 17610 23270 17660
rect 11660 17370 11690 17610
rect 11930 17370 12020 17610
rect 12260 17370 12350 17610
rect 12590 17370 12680 17610
rect 12920 17370 13010 17610
rect 13250 17370 13340 17610
rect 13580 17370 13670 17610
rect 13910 17370 14000 17610
rect 14240 17370 14330 17610
rect 14570 17370 14660 17610
rect 14900 17370 14990 17610
rect 15230 17370 15320 17610
rect 15560 17370 15650 17610
rect 15890 17370 15980 17610
rect 16220 17370 16310 17610
rect 16550 17370 16640 17610
rect 16880 17370 18050 17610
rect 18290 17370 18380 17610
rect 18620 17370 18710 17610
rect 18950 17370 19040 17610
rect 19280 17370 19370 17610
rect 19610 17370 19700 17610
rect 19940 17370 20030 17610
rect 20270 17370 20360 17610
rect 20600 17370 20690 17610
rect 20930 17370 21020 17610
rect 21260 17370 21350 17610
rect 21590 17370 21680 17610
rect 21920 17370 22010 17610
rect 22250 17370 22340 17610
rect 22580 17370 22670 17610
rect 22910 17370 23000 17610
rect 23240 17370 23270 17610
rect 11660 17340 23270 17370
rect 11660 12310 23270 12340
rect 11660 12070 11690 12310
rect 11930 12070 12020 12310
rect 12260 12070 12350 12310
rect 12590 12070 12680 12310
rect 12920 12070 13010 12310
rect 13250 12070 13340 12310
rect 13580 12070 13670 12310
rect 13910 12070 14000 12310
rect 14240 12070 14330 12310
rect 14570 12070 14660 12310
rect 14900 12070 14990 12310
rect 15230 12070 15320 12310
rect 15560 12070 15650 12310
rect 15890 12070 15980 12310
rect 16220 12070 16310 12310
rect 16550 12070 16640 12310
rect 16880 12070 18050 12310
rect 18290 12070 18380 12310
rect 18620 12070 18710 12310
rect 18950 12070 19040 12310
rect 19280 12070 19370 12310
rect 19610 12070 19700 12310
rect 19940 12070 20030 12310
rect 20270 12070 20360 12310
rect 20600 12070 20690 12310
rect 20930 12070 21020 12310
rect 21260 12070 21350 12310
rect 21590 12070 21680 12310
rect 21920 12070 22010 12310
rect 22250 12070 22340 12310
rect 22580 12070 22670 12310
rect 22910 12070 23000 12310
rect 23240 12070 23270 12310
rect 11660 12020 23270 12070
<< comment >>
rect 11570 16320 11630 16350
rect 23300 16320 23360 16350
rect 11570 13350 11630 13380
rect 23300 13350 23360 13380
<< labels >>
rlabel metal4 17450 11600 17450 11600 1 out
port 1 n
rlabel metal4 17450 18150 17450 18150 1 in
port 2 n
rlabel metal5 16990 17630 16990 17630 1 VDD
port 3 n
rlabel metal5 17090 12040 17090 12040 1 GND
port 4 n
<< end >>
