magic
tech sky130A
magscale 1 2
timestamp 1637734600
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 703830 21194 704800
rect 16194 703760 18070 703830
rect 18140 703760 18160 703830
rect 18230 703760 18250 703830
rect 18320 703760 18340 703830
rect 18410 703760 18430 703830
rect 18500 703760 18520 703830
rect 18590 703760 18610 703830
rect 18680 703760 18700 703830
rect 18770 703760 18790 703830
rect 18860 703760 18880 703830
rect 18950 703760 18970 703830
rect 19040 703760 19060 703830
rect 19130 703760 19150 703830
rect 19220 703760 19240 703830
rect 19310 703760 19330 703830
rect 19400 703760 19420 703830
rect 19490 703760 19510 703830
rect 19580 703760 21194 703830
rect 16194 703740 21194 703760
rect 16194 703670 18070 703740
rect 18140 703670 18160 703740
rect 18230 703670 18250 703740
rect 18320 703670 18340 703740
rect 18410 703670 18430 703740
rect 18500 703670 18520 703740
rect 18590 703670 18610 703740
rect 18680 703670 18700 703740
rect 18770 703670 18790 703740
rect 18860 703670 18880 703740
rect 18950 703670 18970 703740
rect 19040 703670 19060 703740
rect 19130 703670 19150 703740
rect 19220 703670 19240 703740
rect 19310 703670 19330 703740
rect 19400 703670 19420 703740
rect 19490 703670 19510 703740
rect 19580 703670 21194 703740
rect 16194 703650 21194 703670
rect 16194 703580 18070 703650
rect 18140 703580 18160 703650
rect 18230 703580 18250 703650
rect 18320 703580 18340 703650
rect 18410 703580 18430 703650
rect 18500 703580 18520 703650
rect 18590 703580 18610 703650
rect 18680 703580 18700 703650
rect 18770 703580 18790 703650
rect 18860 703580 18880 703650
rect 18950 703580 18970 703650
rect 19040 703580 19060 703650
rect 19130 703580 19150 703650
rect 19220 703580 19240 703650
rect 19310 703580 19330 703650
rect 19400 703580 19420 703650
rect 19490 703580 19510 703650
rect 19580 703580 21194 703650
rect 16194 703560 21194 703580
rect 16194 703490 18070 703560
rect 18140 703490 18160 703560
rect 18230 703490 18250 703560
rect 18320 703490 18340 703560
rect 18410 703490 18430 703560
rect 18500 703490 18520 703560
rect 18590 703490 18610 703560
rect 18680 703490 18700 703560
rect 18770 703490 18790 703560
rect 18860 703490 18880 703560
rect 18950 703490 18970 703560
rect 19040 703490 19060 703560
rect 19130 703490 19150 703560
rect 19220 703490 19240 703560
rect 19310 703490 19330 703560
rect 19400 703490 19420 703560
rect 19490 703490 19510 703560
rect 19580 703490 21194 703560
rect 16194 703470 21194 703490
rect 16194 703400 18070 703470
rect 18140 703400 18160 703470
rect 18230 703400 18250 703470
rect 18320 703400 18340 703470
rect 18410 703400 18430 703470
rect 18500 703400 18520 703470
rect 18590 703400 18610 703470
rect 18680 703400 18700 703470
rect 18770 703400 18790 703470
rect 18860 703400 18880 703470
rect 18950 703400 18970 703470
rect 19040 703400 19060 703470
rect 19130 703400 19150 703470
rect 19220 703400 19240 703470
rect 19310 703400 19330 703470
rect 19400 703400 19420 703470
rect 19490 703400 19510 703470
rect 19580 703400 21194 703470
rect 16194 703380 21194 703400
rect 16194 703310 18070 703380
rect 18140 703310 18160 703380
rect 18230 703310 18250 703380
rect 18320 703310 18340 703380
rect 18410 703310 18430 703380
rect 18500 703310 18520 703380
rect 18590 703310 18610 703380
rect 18680 703310 18700 703380
rect 18770 703310 18790 703380
rect 18860 703310 18880 703380
rect 18950 703310 18970 703380
rect 19040 703310 19060 703380
rect 19130 703310 19150 703380
rect 19220 703310 19240 703380
rect 19310 703310 19330 703380
rect 19400 703310 19420 703380
rect 19490 703310 19510 703380
rect 19580 703310 21194 703380
rect 16194 703290 21194 703310
rect 16194 703220 18070 703290
rect 18140 703220 18160 703290
rect 18230 703220 18250 703290
rect 18320 703220 18340 703290
rect 18410 703220 18430 703290
rect 18500 703220 18520 703290
rect 18590 703220 18610 703290
rect 18680 703220 18700 703290
rect 18770 703220 18790 703290
rect 18860 703220 18880 703290
rect 18950 703220 18970 703290
rect 19040 703220 19060 703290
rect 19130 703220 19150 703290
rect 19220 703220 19240 703290
rect 19310 703220 19330 703290
rect 19400 703220 19420 703290
rect 19490 703220 19510 703290
rect 19580 703220 21194 703290
rect 16194 703200 21194 703220
rect 16194 703130 18070 703200
rect 18140 703130 18160 703200
rect 18230 703130 18250 703200
rect 18320 703130 18340 703200
rect 18410 703130 18430 703200
rect 18500 703130 18520 703200
rect 18590 703130 18610 703200
rect 18680 703130 18700 703200
rect 18770 703130 18790 703200
rect 18860 703130 18880 703200
rect 18950 703130 18970 703200
rect 19040 703130 19060 703200
rect 19130 703130 19150 703200
rect 19220 703130 19240 703200
rect 19310 703130 19330 703200
rect 19400 703130 19420 703200
rect 19490 703130 19510 703200
rect 19580 703130 21194 703200
rect 16194 703110 21194 703130
rect 16194 703040 18070 703110
rect 18140 703040 18160 703110
rect 18230 703040 18250 703110
rect 18320 703040 18340 703110
rect 18410 703040 18430 703110
rect 18500 703040 18520 703110
rect 18590 703040 18610 703110
rect 18680 703040 18700 703110
rect 18770 703040 18790 703110
rect 18860 703040 18880 703110
rect 18950 703040 18970 703110
rect 19040 703040 19060 703110
rect 19130 703040 19150 703110
rect 19220 703040 19240 703110
rect 19310 703040 19330 703110
rect 19400 703040 19420 703110
rect 19490 703040 19510 703110
rect 19580 703040 21194 703110
rect 16194 703020 21194 703040
rect 16194 702950 18070 703020
rect 18140 702950 18160 703020
rect 18230 702950 18250 703020
rect 18320 702950 18340 703020
rect 18410 702950 18430 703020
rect 18500 702950 18520 703020
rect 18590 702950 18610 703020
rect 18680 702950 18700 703020
rect 18770 702950 18790 703020
rect 18860 702950 18880 703020
rect 18950 702950 18970 703020
rect 19040 702950 19060 703020
rect 19130 702950 19150 703020
rect 19220 702950 19240 703020
rect 19310 702950 19330 703020
rect 19400 702950 19420 703020
rect 19490 702950 19510 703020
rect 19580 702950 21194 703020
rect 16194 702930 21194 702950
rect 16194 702860 18070 702930
rect 18140 702860 18160 702930
rect 18230 702860 18250 702930
rect 18320 702860 18340 702930
rect 18410 702860 18430 702930
rect 18500 702860 18520 702930
rect 18590 702860 18610 702930
rect 18680 702860 18700 702930
rect 18770 702860 18790 702930
rect 18860 702860 18880 702930
rect 18950 702860 18970 702930
rect 19040 702860 19060 702930
rect 19130 702860 19150 702930
rect 19220 702860 19240 702930
rect 19310 702860 19330 702930
rect 19400 702860 19420 702930
rect 19490 702860 19510 702930
rect 19580 702860 21194 702930
rect 16194 702840 21194 702860
rect 16194 702770 18070 702840
rect 18140 702770 18160 702840
rect 18230 702770 18250 702840
rect 18320 702770 18340 702840
rect 18410 702770 18430 702840
rect 18500 702770 18520 702840
rect 18590 702770 18610 702840
rect 18680 702770 18700 702840
rect 18770 702770 18790 702840
rect 18860 702770 18880 702840
rect 18950 702770 18970 702840
rect 19040 702770 19060 702840
rect 19130 702770 19150 702840
rect 19220 702770 19240 702840
rect 19310 702770 19330 702840
rect 19400 702770 19420 702840
rect 19490 702770 19510 702840
rect 19580 702770 21194 702840
rect 16194 702750 21194 702770
rect 16194 702680 18070 702750
rect 18140 702680 18160 702750
rect 18230 702680 18250 702750
rect 18320 702680 18340 702750
rect 18410 702680 18430 702750
rect 18500 702680 18520 702750
rect 18590 702680 18610 702750
rect 18680 702680 18700 702750
rect 18770 702680 18790 702750
rect 18860 702680 18880 702750
rect 18950 702680 18970 702750
rect 19040 702680 19060 702750
rect 19130 702680 19150 702750
rect 19220 702680 19240 702750
rect 19310 702680 19330 702750
rect 19400 702680 19420 702750
rect 19490 702680 19510 702750
rect 19580 702680 21194 702750
rect 16194 702660 21194 702680
rect 16194 702590 18070 702660
rect 18140 702590 18160 702660
rect 18230 702590 18250 702660
rect 18320 702590 18340 702660
rect 18410 702590 18430 702660
rect 18500 702590 18520 702660
rect 18590 702590 18610 702660
rect 18680 702590 18700 702660
rect 18770 702590 18790 702660
rect 18860 702590 18880 702660
rect 18950 702590 18970 702660
rect 19040 702590 19060 702660
rect 19130 702590 19150 702660
rect 19220 702590 19240 702660
rect 19310 702590 19330 702660
rect 19400 702590 19420 702660
rect 19490 702590 19510 702660
rect 19580 702590 21194 702660
rect 16194 702570 21194 702590
rect 16194 702500 18070 702570
rect 18140 702500 18160 702570
rect 18230 702500 18250 702570
rect 18320 702500 18340 702570
rect 18410 702500 18430 702570
rect 18500 702500 18520 702570
rect 18590 702500 18610 702570
rect 18680 702500 18700 702570
rect 18770 702500 18790 702570
rect 18860 702500 18880 702570
rect 18950 702500 18970 702570
rect 19040 702500 19060 702570
rect 19130 702500 19150 702570
rect 19220 702500 19240 702570
rect 19310 702500 19330 702570
rect 19400 702500 19420 702570
rect 19490 702500 19510 702570
rect 19580 702500 21194 702570
rect 16194 702480 21194 702500
rect 16194 702410 18070 702480
rect 18140 702410 18160 702480
rect 18230 702410 18250 702480
rect 18320 702410 18340 702480
rect 18410 702410 18430 702480
rect 18500 702410 18520 702480
rect 18590 702410 18610 702480
rect 18680 702410 18700 702480
rect 18770 702410 18790 702480
rect 18860 702410 18880 702480
rect 18950 702410 18970 702480
rect 19040 702410 19060 702480
rect 19130 702410 19150 702480
rect 19220 702410 19240 702480
rect 19310 702410 19330 702480
rect 19400 702410 19420 702480
rect 19490 702410 19510 702480
rect 19580 702410 21194 702480
rect 16194 702390 21194 702410
rect 16194 702320 18070 702390
rect 18140 702320 18160 702390
rect 18230 702320 18250 702390
rect 18320 702320 18340 702390
rect 18410 702320 18430 702390
rect 18500 702320 18520 702390
rect 18590 702320 18610 702390
rect 18680 702320 18700 702390
rect 18770 702320 18790 702390
rect 18860 702320 18880 702390
rect 18950 702320 18970 702390
rect 19040 702320 19060 702390
rect 19130 702320 19150 702390
rect 19220 702320 19240 702390
rect 19310 702320 19330 702390
rect 19400 702320 19420 702390
rect 19490 702320 19510 702390
rect 19580 702320 21194 702390
rect 16194 702300 21194 702320
rect 68194 703830 73194 704800
rect 68194 703760 70090 703830
rect 70160 703760 70180 703830
rect 70250 703760 70270 703830
rect 70340 703760 70360 703830
rect 70430 703760 70450 703830
rect 70520 703760 70540 703830
rect 70610 703760 70630 703830
rect 70700 703760 70720 703830
rect 70790 703760 70810 703830
rect 70880 703760 70900 703830
rect 70970 703760 70990 703830
rect 71060 703760 71080 703830
rect 71150 703760 71170 703830
rect 71240 703760 71260 703830
rect 71330 703760 71350 703830
rect 71420 703760 71440 703830
rect 71510 703760 71530 703830
rect 71600 703760 73194 703830
rect 68194 703740 73194 703760
rect 68194 703670 70090 703740
rect 70160 703670 70180 703740
rect 70250 703670 70270 703740
rect 70340 703670 70360 703740
rect 70430 703670 70450 703740
rect 70520 703670 70540 703740
rect 70610 703670 70630 703740
rect 70700 703670 70720 703740
rect 70790 703670 70810 703740
rect 70880 703670 70900 703740
rect 70970 703670 70990 703740
rect 71060 703670 71080 703740
rect 71150 703670 71170 703740
rect 71240 703670 71260 703740
rect 71330 703670 71350 703740
rect 71420 703670 71440 703740
rect 71510 703670 71530 703740
rect 71600 703670 73194 703740
rect 68194 703650 73194 703670
rect 68194 703580 70090 703650
rect 70160 703580 70180 703650
rect 70250 703580 70270 703650
rect 70340 703580 70360 703650
rect 70430 703580 70450 703650
rect 70520 703580 70540 703650
rect 70610 703580 70630 703650
rect 70700 703580 70720 703650
rect 70790 703580 70810 703650
rect 70880 703580 70900 703650
rect 70970 703580 70990 703650
rect 71060 703580 71080 703650
rect 71150 703580 71170 703650
rect 71240 703580 71260 703650
rect 71330 703580 71350 703650
rect 71420 703580 71440 703650
rect 71510 703580 71530 703650
rect 71600 703580 73194 703650
rect 68194 703560 73194 703580
rect 68194 703490 70090 703560
rect 70160 703490 70180 703560
rect 70250 703490 70270 703560
rect 70340 703490 70360 703560
rect 70430 703490 70450 703560
rect 70520 703490 70540 703560
rect 70610 703490 70630 703560
rect 70700 703490 70720 703560
rect 70790 703490 70810 703560
rect 70880 703490 70900 703560
rect 70970 703490 70990 703560
rect 71060 703490 71080 703560
rect 71150 703490 71170 703560
rect 71240 703490 71260 703560
rect 71330 703490 71350 703560
rect 71420 703490 71440 703560
rect 71510 703490 71530 703560
rect 71600 703490 73194 703560
rect 68194 703470 73194 703490
rect 68194 703400 70090 703470
rect 70160 703400 70180 703470
rect 70250 703400 70270 703470
rect 70340 703400 70360 703470
rect 70430 703400 70450 703470
rect 70520 703400 70540 703470
rect 70610 703400 70630 703470
rect 70700 703400 70720 703470
rect 70790 703400 70810 703470
rect 70880 703400 70900 703470
rect 70970 703400 70990 703470
rect 71060 703400 71080 703470
rect 71150 703400 71170 703470
rect 71240 703400 71260 703470
rect 71330 703400 71350 703470
rect 71420 703400 71440 703470
rect 71510 703400 71530 703470
rect 71600 703400 73194 703470
rect 68194 703380 73194 703400
rect 68194 703310 70090 703380
rect 70160 703310 70180 703380
rect 70250 703310 70270 703380
rect 70340 703310 70360 703380
rect 70430 703310 70450 703380
rect 70520 703310 70540 703380
rect 70610 703310 70630 703380
rect 70700 703310 70720 703380
rect 70790 703310 70810 703380
rect 70880 703310 70900 703380
rect 70970 703310 70990 703380
rect 71060 703310 71080 703380
rect 71150 703310 71170 703380
rect 71240 703310 71260 703380
rect 71330 703310 71350 703380
rect 71420 703310 71440 703380
rect 71510 703310 71530 703380
rect 71600 703310 73194 703380
rect 68194 703290 73194 703310
rect 68194 703220 70090 703290
rect 70160 703220 70180 703290
rect 70250 703220 70270 703290
rect 70340 703220 70360 703290
rect 70430 703220 70450 703290
rect 70520 703220 70540 703290
rect 70610 703220 70630 703290
rect 70700 703220 70720 703290
rect 70790 703220 70810 703290
rect 70880 703220 70900 703290
rect 70970 703220 70990 703290
rect 71060 703220 71080 703290
rect 71150 703220 71170 703290
rect 71240 703220 71260 703290
rect 71330 703220 71350 703290
rect 71420 703220 71440 703290
rect 71510 703220 71530 703290
rect 71600 703220 73194 703290
rect 68194 703200 73194 703220
rect 68194 703130 70090 703200
rect 70160 703130 70180 703200
rect 70250 703130 70270 703200
rect 70340 703130 70360 703200
rect 70430 703130 70450 703200
rect 70520 703130 70540 703200
rect 70610 703130 70630 703200
rect 70700 703130 70720 703200
rect 70790 703130 70810 703200
rect 70880 703130 70900 703200
rect 70970 703130 70990 703200
rect 71060 703130 71080 703200
rect 71150 703130 71170 703200
rect 71240 703130 71260 703200
rect 71330 703130 71350 703200
rect 71420 703130 71440 703200
rect 71510 703130 71530 703200
rect 71600 703130 73194 703200
rect 68194 703110 73194 703130
rect 68194 703040 70090 703110
rect 70160 703040 70180 703110
rect 70250 703040 70270 703110
rect 70340 703040 70360 703110
rect 70430 703040 70450 703110
rect 70520 703040 70540 703110
rect 70610 703040 70630 703110
rect 70700 703040 70720 703110
rect 70790 703040 70810 703110
rect 70880 703040 70900 703110
rect 70970 703040 70990 703110
rect 71060 703040 71080 703110
rect 71150 703040 71170 703110
rect 71240 703040 71260 703110
rect 71330 703040 71350 703110
rect 71420 703040 71440 703110
rect 71510 703040 71530 703110
rect 71600 703040 73194 703110
rect 68194 703020 73194 703040
rect 68194 702950 70090 703020
rect 70160 702950 70180 703020
rect 70250 702950 70270 703020
rect 70340 702950 70360 703020
rect 70430 702950 70450 703020
rect 70520 702950 70540 703020
rect 70610 702950 70630 703020
rect 70700 702950 70720 703020
rect 70790 702950 70810 703020
rect 70880 702950 70900 703020
rect 70970 702950 70990 703020
rect 71060 702950 71080 703020
rect 71150 702950 71170 703020
rect 71240 702950 71260 703020
rect 71330 702950 71350 703020
rect 71420 702950 71440 703020
rect 71510 702950 71530 703020
rect 71600 702950 73194 703020
rect 68194 702930 73194 702950
rect 68194 702860 70090 702930
rect 70160 702860 70180 702930
rect 70250 702860 70270 702930
rect 70340 702860 70360 702930
rect 70430 702860 70450 702930
rect 70520 702860 70540 702930
rect 70610 702860 70630 702930
rect 70700 702860 70720 702930
rect 70790 702860 70810 702930
rect 70880 702860 70900 702930
rect 70970 702860 70990 702930
rect 71060 702860 71080 702930
rect 71150 702860 71170 702930
rect 71240 702860 71260 702930
rect 71330 702860 71350 702930
rect 71420 702860 71440 702930
rect 71510 702860 71530 702930
rect 71600 702860 73194 702930
rect 68194 702840 73194 702860
rect 68194 702770 70090 702840
rect 70160 702770 70180 702840
rect 70250 702770 70270 702840
rect 70340 702770 70360 702840
rect 70430 702770 70450 702840
rect 70520 702770 70540 702840
rect 70610 702770 70630 702840
rect 70700 702770 70720 702840
rect 70790 702770 70810 702840
rect 70880 702770 70900 702840
rect 70970 702770 70990 702840
rect 71060 702770 71080 702840
rect 71150 702770 71170 702840
rect 71240 702770 71260 702840
rect 71330 702770 71350 702840
rect 71420 702770 71440 702840
rect 71510 702770 71530 702840
rect 71600 702770 73194 702840
rect 68194 702750 73194 702770
rect 68194 702680 70090 702750
rect 70160 702680 70180 702750
rect 70250 702680 70270 702750
rect 70340 702680 70360 702750
rect 70430 702680 70450 702750
rect 70520 702680 70540 702750
rect 70610 702680 70630 702750
rect 70700 702680 70720 702750
rect 70790 702680 70810 702750
rect 70880 702680 70900 702750
rect 70970 702680 70990 702750
rect 71060 702680 71080 702750
rect 71150 702680 71170 702750
rect 71240 702680 71260 702750
rect 71330 702680 71350 702750
rect 71420 702680 71440 702750
rect 71510 702680 71530 702750
rect 71600 702680 73194 702750
rect 68194 702660 73194 702680
rect 68194 702590 70090 702660
rect 70160 702590 70180 702660
rect 70250 702590 70270 702660
rect 70340 702590 70360 702660
rect 70430 702590 70450 702660
rect 70520 702590 70540 702660
rect 70610 702590 70630 702660
rect 70700 702590 70720 702660
rect 70790 702590 70810 702660
rect 70880 702590 70900 702660
rect 70970 702590 70990 702660
rect 71060 702590 71080 702660
rect 71150 702590 71170 702660
rect 71240 702590 71260 702660
rect 71330 702590 71350 702660
rect 71420 702590 71440 702660
rect 71510 702590 71530 702660
rect 71600 702590 73194 702660
rect 68194 702570 73194 702590
rect 68194 702500 70090 702570
rect 70160 702500 70180 702570
rect 70250 702500 70270 702570
rect 70340 702500 70360 702570
rect 70430 702500 70450 702570
rect 70520 702500 70540 702570
rect 70610 702500 70630 702570
rect 70700 702500 70720 702570
rect 70790 702500 70810 702570
rect 70880 702500 70900 702570
rect 70970 702500 70990 702570
rect 71060 702500 71080 702570
rect 71150 702500 71170 702570
rect 71240 702500 71260 702570
rect 71330 702500 71350 702570
rect 71420 702500 71440 702570
rect 71510 702500 71530 702570
rect 71600 702500 73194 702570
rect 68194 702480 73194 702500
rect 68194 702410 70090 702480
rect 70160 702410 70180 702480
rect 70250 702410 70270 702480
rect 70340 702410 70360 702480
rect 70430 702410 70450 702480
rect 70520 702410 70540 702480
rect 70610 702410 70630 702480
rect 70700 702410 70720 702480
rect 70790 702410 70810 702480
rect 70880 702410 70900 702480
rect 70970 702410 70990 702480
rect 71060 702410 71080 702480
rect 71150 702410 71170 702480
rect 71240 702410 71260 702480
rect 71330 702410 71350 702480
rect 71420 702410 71440 702480
rect 71510 702410 71530 702480
rect 71600 702410 73194 702480
rect 68194 702390 73194 702410
rect 68194 702320 70090 702390
rect 70160 702320 70180 702390
rect 70250 702320 70270 702390
rect 70340 702320 70360 702390
rect 70430 702320 70450 702390
rect 70520 702320 70540 702390
rect 70610 702320 70630 702390
rect 70700 702320 70720 702390
rect 70790 702320 70810 702390
rect 70880 702320 70900 702390
rect 70970 702320 70990 702390
rect 71060 702320 71080 702390
rect 71150 702320 71170 702390
rect 71240 702320 71260 702390
rect 71330 702320 71350 702390
rect 71420 702320 71440 702390
rect 71510 702320 71530 702390
rect 71600 702320 73194 702390
rect 68194 702300 73194 702320
rect 120194 703830 125194 704800
rect 120194 703760 121788 703830
rect 121858 703760 121878 703830
rect 121948 703760 121968 703830
rect 122038 703760 122058 703830
rect 122128 703760 122148 703830
rect 122218 703760 122238 703830
rect 122308 703760 122328 703830
rect 122398 703760 122418 703830
rect 122488 703760 122508 703830
rect 122578 703760 122598 703830
rect 122668 703760 122688 703830
rect 122758 703760 122778 703830
rect 122848 703760 122868 703830
rect 122938 703760 122958 703830
rect 123028 703760 123048 703830
rect 123118 703760 123138 703830
rect 123208 703760 123228 703830
rect 123298 703760 125194 703830
rect 120194 703740 125194 703760
rect 120194 703670 121788 703740
rect 121858 703670 121878 703740
rect 121948 703670 121968 703740
rect 122038 703670 122058 703740
rect 122128 703670 122148 703740
rect 122218 703670 122238 703740
rect 122308 703670 122328 703740
rect 122398 703670 122418 703740
rect 122488 703670 122508 703740
rect 122578 703670 122598 703740
rect 122668 703670 122688 703740
rect 122758 703670 122778 703740
rect 122848 703670 122868 703740
rect 122938 703670 122958 703740
rect 123028 703670 123048 703740
rect 123118 703670 123138 703740
rect 123208 703670 123228 703740
rect 123298 703670 125194 703740
rect 120194 703650 125194 703670
rect 120194 703580 121788 703650
rect 121858 703580 121878 703650
rect 121948 703580 121968 703650
rect 122038 703580 122058 703650
rect 122128 703580 122148 703650
rect 122218 703580 122238 703650
rect 122308 703580 122328 703650
rect 122398 703580 122418 703650
rect 122488 703580 122508 703650
rect 122578 703580 122598 703650
rect 122668 703580 122688 703650
rect 122758 703580 122778 703650
rect 122848 703580 122868 703650
rect 122938 703580 122958 703650
rect 123028 703580 123048 703650
rect 123118 703580 123138 703650
rect 123208 703580 123228 703650
rect 123298 703580 125194 703650
rect 120194 703560 125194 703580
rect 120194 703490 121788 703560
rect 121858 703490 121878 703560
rect 121948 703490 121968 703560
rect 122038 703490 122058 703560
rect 122128 703490 122148 703560
rect 122218 703490 122238 703560
rect 122308 703490 122328 703560
rect 122398 703490 122418 703560
rect 122488 703490 122508 703560
rect 122578 703490 122598 703560
rect 122668 703490 122688 703560
rect 122758 703490 122778 703560
rect 122848 703490 122868 703560
rect 122938 703490 122958 703560
rect 123028 703490 123048 703560
rect 123118 703490 123138 703560
rect 123208 703490 123228 703560
rect 123298 703490 125194 703560
rect 120194 703470 125194 703490
rect 120194 703400 121788 703470
rect 121858 703400 121878 703470
rect 121948 703400 121968 703470
rect 122038 703400 122058 703470
rect 122128 703400 122148 703470
rect 122218 703400 122238 703470
rect 122308 703400 122328 703470
rect 122398 703400 122418 703470
rect 122488 703400 122508 703470
rect 122578 703400 122598 703470
rect 122668 703400 122688 703470
rect 122758 703400 122778 703470
rect 122848 703400 122868 703470
rect 122938 703400 122958 703470
rect 123028 703400 123048 703470
rect 123118 703400 123138 703470
rect 123208 703400 123228 703470
rect 123298 703400 125194 703470
rect 120194 703380 125194 703400
rect 120194 703310 121788 703380
rect 121858 703310 121878 703380
rect 121948 703310 121968 703380
rect 122038 703310 122058 703380
rect 122128 703310 122148 703380
rect 122218 703310 122238 703380
rect 122308 703310 122328 703380
rect 122398 703310 122418 703380
rect 122488 703310 122508 703380
rect 122578 703310 122598 703380
rect 122668 703310 122688 703380
rect 122758 703310 122778 703380
rect 122848 703310 122868 703380
rect 122938 703310 122958 703380
rect 123028 703310 123048 703380
rect 123118 703310 123138 703380
rect 123208 703310 123228 703380
rect 123298 703310 125194 703380
rect 120194 703290 125194 703310
rect 120194 703220 121788 703290
rect 121858 703220 121878 703290
rect 121948 703220 121968 703290
rect 122038 703220 122058 703290
rect 122128 703220 122148 703290
rect 122218 703220 122238 703290
rect 122308 703220 122328 703290
rect 122398 703220 122418 703290
rect 122488 703220 122508 703290
rect 122578 703220 122598 703290
rect 122668 703220 122688 703290
rect 122758 703220 122778 703290
rect 122848 703220 122868 703290
rect 122938 703220 122958 703290
rect 123028 703220 123048 703290
rect 123118 703220 123138 703290
rect 123208 703220 123228 703290
rect 123298 703220 125194 703290
rect 120194 703200 125194 703220
rect 120194 703130 121788 703200
rect 121858 703130 121878 703200
rect 121948 703130 121968 703200
rect 122038 703130 122058 703200
rect 122128 703130 122148 703200
rect 122218 703130 122238 703200
rect 122308 703130 122328 703200
rect 122398 703130 122418 703200
rect 122488 703130 122508 703200
rect 122578 703130 122598 703200
rect 122668 703130 122688 703200
rect 122758 703130 122778 703200
rect 122848 703130 122868 703200
rect 122938 703130 122958 703200
rect 123028 703130 123048 703200
rect 123118 703130 123138 703200
rect 123208 703130 123228 703200
rect 123298 703130 125194 703200
rect 120194 703110 125194 703130
rect 120194 703040 121788 703110
rect 121858 703040 121878 703110
rect 121948 703040 121968 703110
rect 122038 703040 122058 703110
rect 122128 703040 122148 703110
rect 122218 703040 122238 703110
rect 122308 703040 122328 703110
rect 122398 703040 122418 703110
rect 122488 703040 122508 703110
rect 122578 703040 122598 703110
rect 122668 703040 122688 703110
rect 122758 703040 122778 703110
rect 122848 703040 122868 703110
rect 122938 703040 122958 703110
rect 123028 703040 123048 703110
rect 123118 703040 123138 703110
rect 123208 703040 123228 703110
rect 123298 703040 125194 703110
rect 120194 703020 125194 703040
rect 120194 702950 121788 703020
rect 121858 702950 121878 703020
rect 121948 702950 121968 703020
rect 122038 702950 122058 703020
rect 122128 702950 122148 703020
rect 122218 702950 122238 703020
rect 122308 702950 122328 703020
rect 122398 702950 122418 703020
rect 122488 702950 122508 703020
rect 122578 702950 122598 703020
rect 122668 702950 122688 703020
rect 122758 702950 122778 703020
rect 122848 702950 122868 703020
rect 122938 702950 122958 703020
rect 123028 702950 123048 703020
rect 123118 702950 123138 703020
rect 123208 702950 123228 703020
rect 123298 702950 125194 703020
rect 120194 702930 125194 702950
rect 120194 702860 121788 702930
rect 121858 702860 121878 702930
rect 121948 702860 121968 702930
rect 122038 702860 122058 702930
rect 122128 702860 122148 702930
rect 122218 702860 122238 702930
rect 122308 702860 122328 702930
rect 122398 702860 122418 702930
rect 122488 702860 122508 702930
rect 122578 702860 122598 702930
rect 122668 702860 122688 702930
rect 122758 702860 122778 702930
rect 122848 702860 122868 702930
rect 122938 702860 122958 702930
rect 123028 702860 123048 702930
rect 123118 702860 123138 702930
rect 123208 702860 123228 702930
rect 123298 702860 125194 702930
rect 120194 702840 125194 702860
rect 120194 702770 121788 702840
rect 121858 702770 121878 702840
rect 121948 702770 121968 702840
rect 122038 702770 122058 702840
rect 122128 702770 122148 702840
rect 122218 702770 122238 702840
rect 122308 702770 122328 702840
rect 122398 702770 122418 702840
rect 122488 702770 122508 702840
rect 122578 702770 122598 702840
rect 122668 702770 122688 702840
rect 122758 702770 122778 702840
rect 122848 702770 122868 702840
rect 122938 702770 122958 702840
rect 123028 702770 123048 702840
rect 123118 702770 123138 702840
rect 123208 702770 123228 702840
rect 123298 702770 125194 702840
rect 120194 702750 125194 702770
rect 120194 702680 121788 702750
rect 121858 702680 121878 702750
rect 121948 702680 121968 702750
rect 122038 702680 122058 702750
rect 122128 702680 122148 702750
rect 122218 702680 122238 702750
rect 122308 702680 122328 702750
rect 122398 702680 122418 702750
rect 122488 702680 122508 702750
rect 122578 702680 122598 702750
rect 122668 702680 122688 702750
rect 122758 702680 122778 702750
rect 122848 702680 122868 702750
rect 122938 702680 122958 702750
rect 123028 702680 123048 702750
rect 123118 702680 123138 702750
rect 123208 702680 123228 702750
rect 123298 702680 125194 702750
rect 120194 702660 125194 702680
rect 120194 702590 121788 702660
rect 121858 702590 121878 702660
rect 121948 702590 121968 702660
rect 122038 702590 122058 702660
rect 122128 702590 122148 702660
rect 122218 702590 122238 702660
rect 122308 702590 122328 702660
rect 122398 702590 122418 702660
rect 122488 702590 122508 702660
rect 122578 702590 122598 702660
rect 122668 702590 122688 702660
rect 122758 702590 122778 702660
rect 122848 702590 122868 702660
rect 122938 702590 122958 702660
rect 123028 702590 123048 702660
rect 123118 702590 123138 702660
rect 123208 702590 123228 702660
rect 123298 702590 125194 702660
rect 120194 702570 125194 702590
rect 120194 702500 121788 702570
rect 121858 702500 121878 702570
rect 121948 702500 121968 702570
rect 122038 702500 122058 702570
rect 122128 702500 122148 702570
rect 122218 702500 122238 702570
rect 122308 702500 122328 702570
rect 122398 702500 122418 702570
rect 122488 702500 122508 702570
rect 122578 702500 122598 702570
rect 122668 702500 122688 702570
rect 122758 702500 122778 702570
rect 122848 702500 122868 702570
rect 122938 702500 122958 702570
rect 123028 702500 123048 702570
rect 123118 702500 123138 702570
rect 123208 702500 123228 702570
rect 123298 702500 125194 702570
rect 120194 702480 125194 702500
rect 120194 702410 121788 702480
rect 121858 702410 121878 702480
rect 121948 702410 121968 702480
rect 122038 702410 122058 702480
rect 122128 702410 122148 702480
rect 122218 702410 122238 702480
rect 122308 702410 122328 702480
rect 122398 702410 122418 702480
rect 122488 702410 122508 702480
rect 122578 702410 122598 702480
rect 122668 702410 122688 702480
rect 122758 702410 122778 702480
rect 122848 702410 122868 702480
rect 122938 702410 122958 702480
rect 123028 702410 123048 702480
rect 123118 702410 123138 702480
rect 123208 702410 123228 702480
rect 123298 702410 125194 702480
rect 120194 702390 125194 702410
rect 120194 702320 121788 702390
rect 121858 702320 121878 702390
rect 121948 702320 121968 702390
rect 122038 702320 122058 702390
rect 122128 702320 122148 702390
rect 122218 702320 122238 702390
rect 122308 702320 122328 702390
rect 122398 702320 122418 702390
rect 122488 702320 122508 702390
rect 122578 702320 122598 702390
rect 122668 702320 122688 702390
rect 122758 702320 122778 702390
rect 122848 702320 122868 702390
rect 122938 702320 122958 702390
rect 123028 702320 123048 702390
rect 123118 702320 123138 702390
rect 123208 702320 123228 702390
rect 123298 702320 125194 702390
rect 120194 702300 125194 702320
rect 165594 702300 170594 704800
rect 170894 692930 173094 704800
rect 173394 704000 175594 704800
rect 175894 704000 180894 704800
rect 173394 702300 180894 704000
rect 217294 704000 222294 704800
rect 222594 704000 224794 704800
rect 217294 702300 224794 704000
rect 225094 700930 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702840 418394 704800
rect 413394 702770 415630 702840
rect 415700 702770 415720 702840
rect 415790 702770 415810 702840
rect 415880 702770 415900 702840
rect 415970 702770 415990 702840
rect 416060 702770 416080 702840
rect 416150 702770 418394 702840
rect 413394 702750 418394 702770
rect 413394 702680 415630 702750
rect 415700 702680 415720 702750
rect 415790 702680 415810 702750
rect 415880 702680 415900 702750
rect 415970 702680 415990 702750
rect 416060 702680 416080 702750
rect 416150 702680 418394 702750
rect 413394 702660 418394 702680
rect 413394 702590 415630 702660
rect 415700 702590 415720 702660
rect 415790 702590 415810 702660
rect 415880 702590 415900 702660
rect 415970 702590 415990 702660
rect 416060 702590 416080 702660
rect 416150 702590 418394 702660
rect 413394 702570 418394 702590
rect 413394 702500 415630 702570
rect 415700 702500 415720 702570
rect 415790 702500 415810 702570
rect 415880 702500 415900 702570
rect 415970 702500 415990 702570
rect 416060 702500 416080 702570
rect 416150 702500 418394 702570
rect 413394 702480 418394 702500
rect 413394 702410 415630 702480
rect 415700 702410 415720 702480
rect 415790 702410 415810 702480
rect 415880 702410 415900 702480
rect 415970 702410 415990 702480
rect 416060 702410 416080 702480
rect 416150 702410 418394 702480
rect 413394 702390 418394 702410
rect 413394 702320 415630 702390
rect 415700 702320 415720 702390
rect 415790 702320 415810 702390
rect 415880 702320 415900 702390
rect 415970 702320 415990 702390
rect 416060 702320 416080 702390
rect 416150 702320 418394 702390
rect 413394 702300 418394 702320
rect 465394 702840 470394 704800
rect 465394 702770 467630 702840
rect 467700 702770 467720 702840
rect 467790 702770 467810 702840
rect 467880 702770 467900 702840
rect 467970 702770 467990 702840
rect 468060 702770 468080 702840
rect 468150 702770 470394 702840
rect 465394 702750 470394 702770
rect 465394 702680 467630 702750
rect 467700 702680 467720 702750
rect 467790 702680 467810 702750
rect 467880 702680 467900 702750
rect 467970 702680 467990 702750
rect 468060 702680 468080 702750
rect 468150 702680 470394 702750
rect 465394 702660 470394 702680
rect 465394 702590 467630 702660
rect 467700 702590 467720 702660
rect 467790 702590 467810 702660
rect 467880 702590 467900 702660
rect 467970 702590 467990 702660
rect 468060 702590 468080 702660
rect 468150 702590 470394 702660
rect 465394 702570 470394 702590
rect 465394 702500 467630 702570
rect 467700 702500 467720 702570
rect 467790 702500 467810 702570
rect 467880 702500 467900 702570
rect 467970 702500 467990 702570
rect 468060 702500 468080 702570
rect 468150 702500 470394 702570
rect 465394 702480 470394 702500
rect 465394 702410 467630 702480
rect 467700 702410 467720 702480
rect 467790 702410 467810 702480
rect 467880 702410 467900 702480
rect 467970 702410 467990 702480
rect 468060 702410 468080 702480
rect 468150 702410 470394 702480
rect 465394 702390 470394 702410
rect 465394 702320 467630 702390
rect 467700 702320 467720 702390
rect 467790 702320 467810 702390
rect 467880 702320 467900 702390
rect 467970 702320 467990 702390
rect 468060 702320 468080 702390
rect 468150 702320 470394 702390
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702840 571594 704800
rect 566594 702770 566740 702840
rect 566810 702770 566830 702840
rect 566900 702770 566920 702840
rect 566990 702770 567010 702840
rect 567080 702770 567100 702840
rect 567170 702770 567190 702840
rect 567260 702770 571594 702840
rect 566594 702750 571594 702770
rect 566594 702680 566740 702750
rect 566810 702680 566830 702750
rect 566900 702680 566920 702750
rect 566990 702680 567010 702750
rect 567080 702680 567100 702750
rect 567170 702680 567190 702750
rect 567260 702680 571594 702750
rect 566594 702660 571594 702680
rect 566594 702590 566740 702660
rect 566810 702590 566830 702660
rect 566900 702590 566920 702660
rect 566990 702590 567010 702660
rect 567080 702590 567100 702660
rect 567170 702590 567190 702660
rect 567260 702590 571594 702660
rect 566594 702570 571594 702590
rect 566594 702500 566740 702570
rect 566810 702500 566830 702570
rect 566900 702500 566920 702570
rect 566990 702500 567010 702570
rect 567080 702500 567100 702570
rect 567170 702500 567190 702570
rect 567260 702500 571594 702570
rect 566594 702480 571594 702500
rect 566594 702410 566740 702480
rect 566810 702410 566830 702480
rect 566900 702410 566920 702480
rect 566990 702410 567010 702480
rect 567080 702410 567100 702480
rect 567170 702410 567190 702480
rect 567260 702410 571594 702480
rect 566594 702390 571594 702410
rect 465394 702300 470394 702320
rect 566594 702320 566740 702390
rect 566810 702320 566830 702390
rect 566900 702320 566920 702390
rect 566990 702320 567010 702390
rect 567080 702320 567100 702390
rect 567170 702320 567190 702390
rect 567260 702320 571594 702390
rect 566594 702300 571594 702320
rect 225094 700690 225164 700930
rect 225404 700690 225494 700930
rect 225734 700690 225824 700930
rect 226064 700690 226154 700930
rect 226394 700690 226484 700930
rect 226724 700690 226814 700930
rect 227054 700690 227294 700930
rect 225094 700600 227294 700690
rect 225094 700360 225164 700600
rect 225404 700360 225494 700600
rect 225734 700360 225824 700600
rect 226064 700360 226154 700600
rect 226394 700360 226484 700600
rect 226724 700360 226814 700600
rect 227054 700360 227294 700600
rect 225094 700270 227294 700360
rect 225094 700030 225164 700270
rect 225404 700030 225494 700270
rect 225734 700030 225824 700270
rect 226064 700030 226154 700270
rect 226394 700030 226484 700270
rect 226724 700030 226814 700270
rect 227054 700030 227294 700270
rect 225094 699940 227294 700030
rect 225094 699700 225164 699940
rect 225404 699700 225494 699940
rect 225734 699700 225824 699940
rect 226064 699700 226154 699940
rect 226394 699700 226484 699940
rect 226724 699700 226814 699940
rect 227054 699700 227294 699940
rect 225094 699610 227294 699700
rect 225094 699370 225164 699610
rect 225404 699370 225494 699610
rect 225734 699370 225824 699610
rect 226064 699370 226154 699610
rect 226394 699370 226484 699610
rect 226724 699370 226814 699610
rect 227054 699370 227294 699610
rect 225094 699280 227294 699370
rect 225094 699040 225164 699280
rect 225404 699040 225494 699280
rect 225734 699040 225824 699280
rect 226064 699040 226154 699280
rect 226394 699040 226484 699280
rect 226724 699040 226814 699280
rect 227054 699040 227294 699280
rect 225094 698950 227294 699040
rect 225094 698710 225164 698950
rect 225404 698710 225494 698950
rect 225734 698710 225824 698950
rect 226064 698710 226154 698950
rect 226394 698710 226484 698950
rect 226724 698710 226814 698950
rect 227054 698710 227294 698950
rect 225094 698620 227294 698710
rect 225094 698380 225164 698620
rect 225404 698380 225494 698620
rect 225734 698380 225824 698620
rect 226064 698380 226154 698620
rect 226394 698380 226484 698620
rect 226724 698380 226814 698620
rect 227054 698380 227294 698620
rect 225094 698290 227294 698380
rect 225094 698050 225164 698290
rect 225404 698050 225494 698290
rect 225734 698050 225824 698290
rect 226064 698050 226154 698290
rect 226394 698050 226484 698290
rect 226724 698050 226814 698290
rect 227054 698050 227294 698290
rect 225094 697960 227294 698050
rect 225094 697720 225164 697960
rect 225404 697720 225494 697960
rect 225734 697720 225824 697960
rect 226064 697720 226154 697960
rect 226394 697720 226484 697960
rect 226724 697720 226814 697960
rect 227054 697720 227294 697960
rect 225094 697630 227294 697720
rect 225094 697390 225164 697630
rect 225404 697390 225494 697630
rect 225734 697390 225824 697630
rect 226064 697390 226154 697630
rect 226394 697390 226484 697630
rect 226724 697390 226814 697630
rect 227054 697390 227294 697630
rect 225094 697300 227294 697390
rect 225094 697060 225164 697300
rect 225404 697060 225494 697300
rect 225734 697060 225824 697300
rect 226064 697060 226154 697300
rect 226394 697060 226484 697300
rect 226724 697060 226814 697300
rect 227054 697060 227294 697300
rect 225094 696970 227294 697060
rect 225094 696730 225164 696970
rect 225404 696730 225494 696970
rect 225734 696730 225824 696970
rect 226064 696730 226154 696970
rect 226394 696730 226484 696970
rect 226724 696730 226814 696970
rect 227054 696730 227294 696970
rect 225094 696640 227294 696730
rect 225094 696400 225164 696640
rect 225404 696400 225494 696640
rect 225734 696400 225824 696640
rect 226064 696400 226154 696640
rect 226394 696400 226484 696640
rect 226724 696400 226814 696640
rect 227054 696400 227294 696640
rect 225094 696310 227294 696400
rect 225094 696070 225164 696310
rect 225404 696070 225494 696310
rect 225734 696070 225824 696310
rect 226064 696070 226154 696310
rect 226394 696070 226484 696310
rect 226724 696070 226814 696310
rect 227054 696070 227294 696310
rect 225094 696000 227294 696070
rect 170894 692690 170964 692930
rect 171204 692690 171294 692930
rect 171534 692690 171624 692930
rect 171864 692690 171954 692930
rect 172194 692690 172284 692930
rect 172524 692690 172614 692930
rect 172854 692690 173094 692930
rect 170894 692600 173094 692690
rect 170894 692360 170964 692600
rect 171204 692360 171294 692600
rect 171534 692360 171624 692600
rect 171864 692360 171954 692600
rect 172194 692360 172284 692600
rect 172524 692360 172614 692600
rect 172854 692360 173094 692600
rect 170894 692270 173094 692360
rect 170894 692030 170964 692270
rect 171204 692030 171294 692270
rect 171534 692030 171624 692270
rect 171864 692030 171954 692270
rect 172194 692030 172284 692270
rect 172524 692030 172614 692270
rect 172854 692030 173094 692270
rect 170894 691940 173094 692030
rect 170894 691700 170964 691940
rect 171204 691700 171294 691940
rect 171534 691700 171624 691940
rect 171864 691700 171954 691940
rect 172194 691700 172284 691940
rect 172524 691700 172614 691940
rect 172854 691700 173094 691940
rect 170894 691610 173094 691700
rect 170894 691370 170964 691610
rect 171204 691370 171294 691610
rect 171534 691370 171624 691610
rect 171864 691370 171954 691610
rect 172194 691370 172284 691610
rect 172524 691370 172614 691610
rect 172854 691370 173094 691610
rect 170894 691280 173094 691370
rect 170894 691040 170964 691280
rect 171204 691040 171294 691280
rect 171534 691040 171624 691280
rect 171864 691040 171954 691280
rect 172194 691040 172284 691280
rect 172524 691040 172614 691280
rect 172854 691040 173094 691280
rect 170894 690950 173094 691040
rect 170894 690710 170964 690950
rect 171204 690710 171294 690950
rect 171534 690710 171624 690950
rect 171864 690710 171954 690950
rect 172194 690710 172284 690950
rect 172524 690710 172614 690950
rect 172854 690710 173094 690950
rect 170894 690620 173094 690710
rect 170894 690380 170964 690620
rect 171204 690380 171294 690620
rect 171534 690380 171624 690620
rect 171864 690380 171954 690620
rect 172194 690380 172284 690620
rect 172524 690380 172614 690620
rect 172854 690380 173094 690620
rect 170894 690290 173094 690380
rect 170894 690050 170964 690290
rect 171204 690050 171294 690290
rect 171534 690050 171624 690290
rect 171864 690050 171954 690290
rect 172194 690050 172284 690290
rect 172524 690050 172614 690290
rect 172854 690050 173094 690290
rect 170894 689960 173094 690050
rect 170894 689720 170964 689960
rect 171204 689720 171294 689960
rect 171534 689720 171624 689960
rect 171864 689720 171954 689960
rect 172194 689720 172284 689960
rect 172524 689720 172614 689960
rect 172854 689720 173094 689960
rect 170894 689630 173094 689720
rect 170894 689390 170964 689630
rect 171204 689390 171294 689630
rect 171534 689390 171624 689630
rect 171864 689390 171954 689630
rect 172194 689390 172284 689630
rect 172524 689390 172614 689630
rect 172854 689390 173094 689630
rect 170894 689300 173094 689390
rect 170894 689060 170964 689300
rect 171204 689060 171294 689300
rect 171534 689060 171624 689300
rect 171864 689060 171954 689300
rect 172194 689060 172284 689300
rect 172524 689060 172614 689300
rect 172854 689060 173094 689300
rect 170894 688970 173094 689060
rect 170894 688730 170964 688970
rect 171204 688730 171294 688970
rect 171534 688730 171624 688970
rect 171864 688730 171954 688970
rect 172194 688730 172284 688970
rect 172524 688730 172614 688970
rect 172854 688730 173094 688970
rect 170894 688640 173094 688730
rect 170894 688400 170964 688640
rect 171204 688400 171294 688640
rect 171534 688400 171624 688640
rect 171864 688400 171954 688640
rect 172194 688400 172284 688640
rect 172524 688400 172614 688640
rect 172854 688400 173094 688640
rect 170894 688310 173094 688400
rect 170894 688070 170964 688310
rect 171204 688070 171294 688310
rect 171534 688070 171624 688310
rect 171864 688070 171954 688310
rect 172194 688070 172284 688310
rect 172524 688070 172614 688310
rect 172854 688070 173094 688310
rect 170894 688000 173094 688070
rect 18050 687370 23946 687390
rect 18050 687300 18120 687370
rect 18190 687300 18210 687370
rect 18280 687300 18300 687370
rect 18370 687300 18390 687370
rect 18460 687300 18480 687370
rect 18550 687300 18570 687370
rect 18640 687300 18660 687370
rect 18730 687300 18750 687370
rect 18820 687300 18840 687370
rect 18910 687300 18930 687370
rect 19000 687300 19020 687370
rect 19090 687300 19110 687370
rect 19180 687300 19200 687370
rect 19270 687300 19290 687370
rect 19360 687300 19380 687370
rect 19450 687300 19470 687370
rect 19540 687300 19560 687370
rect 19630 687300 23946 687370
rect 18050 687280 23946 687300
rect 18050 687210 18120 687280
rect 18190 687210 18210 687280
rect 18280 687210 18300 687280
rect 18370 687210 18390 687280
rect 18460 687210 18480 687280
rect 18550 687210 18570 687280
rect 18640 687210 18660 687280
rect 18730 687210 18750 687280
rect 18820 687210 18840 687280
rect 18910 687210 18930 687280
rect 19000 687210 19020 687280
rect 19090 687210 19110 687280
rect 19180 687210 19200 687280
rect 19270 687210 19290 687280
rect 19360 687210 19380 687280
rect 19450 687210 19470 687280
rect 19540 687210 19560 687280
rect 19630 687210 23946 687280
rect 18050 687190 23946 687210
rect 18050 687120 18120 687190
rect 18190 687120 18210 687190
rect 18280 687120 18300 687190
rect 18370 687120 18390 687190
rect 18460 687120 18480 687190
rect 18550 687120 18570 687190
rect 18640 687120 18660 687190
rect 18730 687120 18750 687190
rect 18820 687120 18840 687190
rect 18910 687120 18930 687190
rect 19000 687120 19020 687190
rect 19090 687120 19110 687190
rect 19180 687120 19200 687190
rect 19270 687120 19290 687190
rect 19360 687120 19380 687190
rect 19450 687120 19470 687190
rect 19540 687120 19560 687190
rect 19630 687120 23946 687190
rect 18050 687100 23946 687120
rect 18050 687030 18120 687100
rect 18190 687030 18210 687100
rect 18280 687030 18300 687100
rect 18370 687030 18390 687100
rect 18460 687030 18480 687100
rect 18550 687030 18570 687100
rect 18640 687030 18660 687100
rect 18730 687030 18750 687100
rect 18820 687030 18840 687100
rect 18910 687030 18930 687100
rect 19000 687030 19020 687100
rect 19090 687030 19110 687100
rect 19180 687030 19200 687100
rect 19270 687030 19290 687100
rect 19360 687030 19380 687100
rect 19450 687030 19470 687100
rect 19540 687030 19560 687100
rect 19630 687030 23946 687100
rect 18050 687010 23946 687030
rect 18050 686940 18120 687010
rect 18190 686940 18210 687010
rect 18280 686940 18300 687010
rect 18370 686940 18390 687010
rect 18460 686940 18480 687010
rect 18550 686940 18570 687010
rect 18640 686940 18660 687010
rect 18730 686940 18750 687010
rect 18820 686940 18840 687010
rect 18910 686940 18930 687010
rect 19000 686940 19020 687010
rect 19090 686940 19110 687010
rect 19180 686940 19200 687010
rect 19270 686940 19290 687010
rect 19360 686940 19380 687010
rect 19450 686940 19470 687010
rect 19540 686940 19560 687010
rect 19630 686940 23946 687010
rect 18050 686920 23946 686940
rect 18050 686850 18120 686920
rect 18190 686850 18210 686920
rect 18280 686850 18300 686920
rect 18370 686850 18390 686920
rect 18460 686850 18480 686920
rect 18550 686850 18570 686920
rect 18640 686850 18660 686920
rect 18730 686850 18750 686920
rect 18820 686850 18840 686920
rect 18910 686850 18930 686920
rect 19000 686850 19020 686920
rect 19090 686850 19110 686920
rect 19180 686850 19200 686920
rect 19270 686850 19290 686920
rect 19360 686850 19380 686920
rect 19450 686850 19470 686920
rect 19540 686850 19560 686920
rect 19630 686850 23946 686920
rect 18050 686830 23946 686850
rect 18050 686760 18120 686830
rect 18190 686760 18210 686830
rect 18280 686760 18300 686830
rect 18370 686760 18390 686830
rect 18460 686760 18480 686830
rect 18550 686760 18570 686830
rect 18640 686760 18660 686830
rect 18730 686760 18750 686830
rect 18820 686760 18840 686830
rect 18910 686760 18930 686830
rect 19000 686760 19020 686830
rect 19090 686760 19110 686830
rect 19180 686760 19200 686830
rect 19270 686760 19290 686830
rect 19360 686760 19380 686830
rect 19450 686760 19470 686830
rect 19540 686760 19560 686830
rect 19630 686760 23946 686830
rect 18050 686740 23946 686760
rect 18050 686670 18120 686740
rect 18190 686670 18210 686740
rect 18280 686670 18300 686740
rect 18370 686670 18390 686740
rect 18460 686670 18480 686740
rect 18550 686670 18570 686740
rect 18640 686670 18660 686740
rect 18730 686670 18750 686740
rect 18820 686670 18840 686740
rect 18910 686670 18930 686740
rect 19000 686670 19020 686740
rect 19090 686670 19110 686740
rect 19180 686670 19200 686740
rect 19270 686670 19290 686740
rect 19360 686670 19380 686740
rect 19450 686670 19470 686740
rect 19540 686670 19560 686740
rect 19630 686670 23946 686740
rect 18050 686650 23946 686670
rect 18050 686580 18120 686650
rect 18190 686580 18210 686650
rect 18280 686580 18300 686650
rect 18370 686580 18390 686650
rect 18460 686580 18480 686650
rect 18550 686580 18570 686650
rect 18640 686580 18660 686650
rect 18730 686580 18750 686650
rect 18820 686580 18840 686650
rect 18910 686580 18930 686650
rect 19000 686580 19020 686650
rect 19090 686580 19110 686650
rect 19180 686580 19200 686650
rect 19270 686580 19290 686650
rect 19360 686580 19380 686650
rect 19450 686580 19470 686650
rect 19540 686580 19560 686650
rect 19630 686580 23946 686650
rect 18050 686560 23946 686580
rect 18050 686490 18120 686560
rect 18190 686490 18210 686560
rect 18280 686490 18300 686560
rect 18370 686490 18390 686560
rect 18460 686490 18480 686560
rect 18550 686490 18570 686560
rect 18640 686490 18660 686560
rect 18730 686490 18750 686560
rect 18820 686490 18840 686560
rect 18910 686490 18930 686560
rect 19000 686490 19020 686560
rect 19090 686490 19110 686560
rect 19180 686490 19200 686560
rect 19270 686490 19290 686560
rect 19360 686490 19380 686560
rect 19450 686490 19470 686560
rect 19540 686490 19560 686560
rect 19630 686490 23946 686560
rect 18050 686470 23946 686490
rect 18050 686400 18120 686470
rect 18190 686400 18210 686470
rect 18280 686400 18300 686470
rect 18370 686400 18390 686470
rect 18460 686400 18480 686470
rect 18550 686400 18570 686470
rect 18640 686400 18660 686470
rect 18730 686400 18750 686470
rect 18820 686400 18840 686470
rect 18910 686400 18930 686470
rect 19000 686400 19020 686470
rect 19090 686400 19110 686470
rect 19180 686400 19200 686470
rect 19270 686400 19290 686470
rect 19360 686400 19380 686470
rect 19450 686400 19470 686470
rect 19540 686400 19560 686470
rect 19630 686400 23946 686470
rect 18050 686380 23946 686400
rect 18050 686310 18120 686380
rect 18190 686310 18210 686380
rect 18280 686310 18300 686380
rect 18370 686310 18390 686380
rect 18460 686310 18480 686380
rect 18550 686310 18570 686380
rect 18640 686310 18660 686380
rect 18730 686310 18750 686380
rect 18820 686310 18840 686380
rect 18910 686310 18930 686380
rect 19000 686310 19020 686380
rect 19090 686310 19110 686380
rect 19180 686310 19200 686380
rect 19270 686310 19290 686380
rect 19360 686310 19380 686380
rect 19450 686310 19470 686380
rect 19540 686310 19560 686380
rect 19630 686310 23946 686380
rect 18050 686290 23946 686310
rect 18050 686220 18120 686290
rect 18190 686220 18210 686290
rect 18280 686220 18300 686290
rect 18370 686220 18390 686290
rect 18460 686220 18480 686290
rect 18550 686220 18570 686290
rect 18640 686220 18660 686290
rect 18730 686220 18750 686290
rect 18820 686220 18840 686290
rect 18910 686220 18930 686290
rect 19000 686220 19020 686290
rect 19090 686220 19110 686290
rect 19180 686220 19200 686290
rect 19270 686220 19290 686290
rect 19360 686220 19380 686290
rect 19450 686220 19470 686290
rect 19540 686220 19560 686290
rect 19630 686220 23946 686290
rect 18050 686200 23946 686220
rect 18050 686130 18120 686200
rect 18190 686130 18210 686200
rect 18280 686130 18300 686200
rect 18370 686130 18390 686200
rect 18460 686130 18480 686200
rect 18550 686130 18570 686200
rect 18640 686130 18660 686200
rect 18730 686130 18750 686200
rect 18820 686130 18840 686200
rect 18910 686130 18930 686200
rect 19000 686130 19020 686200
rect 19090 686130 19110 686200
rect 19180 686130 19200 686200
rect 19270 686130 19290 686200
rect 19360 686130 19380 686200
rect 19450 686130 19470 686200
rect 19540 686130 19560 686200
rect 19630 686130 23946 686200
rect 18050 686110 23946 686130
rect 18050 686040 18120 686110
rect 18190 686040 18210 686110
rect 18280 686040 18300 686110
rect 18370 686040 18390 686110
rect 18460 686040 18480 686110
rect 18550 686040 18570 686110
rect 18640 686040 18660 686110
rect 18730 686040 18750 686110
rect 18820 686040 18840 686110
rect 18910 686040 18930 686110
rect 19000 686040 19020 686110
rect 19090 686040 19110 686110
rect 19180 686040 19200 686110
rect 19270 686040 19290 686110
rect 19360 686040 19380 686110
rect 19450 686040 19470 686110
rect 19540 686040 19560 686110
rect 19630 686040 23946 686110
rect 18050 686020 23946 686040
rect 18050 685950 18120 686020
rect 18190 685950 18210 686020
rect 18280 685950 18300 686020
rect 18370 685950 18390 686020
rect 18460 685950 18480 686020
rect 18550 685950 18570 686020
rect 18640 685950 18660 686020
rect 18730 685950 18750 686020
rect 18820 685950 18840 686020
rect 18910 685950 18930 686020
rect 19000 685950 19020 686020
rect 19090 685950 19110 686020
rect 19180 685950 19200 686020
rect 19270 685950 19290 686020
rect 19360 685950 19380 686020
rect 19450 685950 19470 686020
rect 19540 685950 19560 686020
rect 19630 685950 23946 686020
rect 18050 685930 23946 685950
rect 18050 685860 18120 685930
rect 18190 685860 18210 685930
rect 18280 685860 18300 685930
rect 18370 685860 18390 685930
rect 18460 685860 18480 685930
rect 18550 685860 18570 685930
rect 18640 685860 18660 685930
rect 18730 685860 18750 685930
rect 18820 685860 18840 685930
rect 18910 685860 18930 685930
rect 19000 685860 19020 685930
rect 19090 685860 19110 685930
rect 19180 685860 19200 685930
rect 19270 685860 19290 685930
rect 19360 685860 19380 685930
rect 19450 685860 19470 685930
rect 19540 685860 19560 685930
rect 19630 685860 23946 685930
rect 18050 685840 23946 685860
rect 18050 685770 18120 685840
rect 18190 685770 18210 685840
rect 18280 685770 18300 685840
rect 18370 685770 18390 685840
rect 18460 685770 18480 685840
rect 18550 685770 18570 685840
rect 18640 685770 18660 685840
rect 18730 685770 18750 685840
rect 18820 685770 18840 685840
rect 18910 685770 18930 685840
rect 19000 685770 19020 685840
rect 19090 685770 19110 685840
rect 19180 685770 19200 685840
rect 19270 685770 19290 685840
rect 19360 685770 19380 685840
rect 19450 685770 19470 685840
rect 19540 685770 19560 685840
rect 19630 685770 23946 685840
rect 18050 685750 23946 685770
rect 18050 685680 18120 685750
rect 18190 685680 18210 685750
rect 18280 685680 18300 685750
rect 18370 685680 18390 685750
rect 18460 685680 18480 685750
rect 18550 685680 18570 685750
rect 18640 685680 18660 685750
rect 18730 685680 18750 685750
rect 18820 685680 18840 685750
rect 18910 685680 18930 685750
rect 19000 685680 19020 685750
rect 19090 685680 19110 685750
rect 19180 685680 19200 685750
rect 19270 685680 19290 685750
rect 19360 685680 19380 685750
rect 19450 685680 19470 685750
rect 19540 685680 19560 685750
rect 19630 685680 23946 685750
rect 18050 685660 23946 685680
rect 18050 685590 18120 685660
rect 18190 685590 18210 685660
rect 18280 685590 18300 685660
rect 18370 685590 18390 685660
rect 18460 685590 18480 685660
rect 18550 685590 18570 685660
rect 18640 685590 18660 685660
rect 18730 685590 18750 685660
rect 18820 685590 18840 685660
rect 18910 685590 18930 685660
rect 19000 685590 19020 685660
rect 19090 685590 19110 685660
rect 19180 685590 19200 685660
rect 19270 685590 19290 685660
rect 19360 685590 19380 685660
rect 19450 685590 19470 685660
rect 19540 685590 19560 685660
rect 19630 685590 23946 685660
rect 18050 685570 23946 685590
rect 18050 685500 18120 685570
rect 18190 685500 18210 685570
rect 18280 685500 18300 685570
rect 18370 685500 18390 685570
rect 18460 685500 18480 685570
rect 18550 685500 18570 685570
rect 18640 685500 18660 685570
rect 18730 685500 18750 685570
rect 18820 685500 18840 685570
rect 18910 685500 18930 685570
rect 19000 685500 19020 685570
rect 19090 685500 19110 685570
rect 19180 685500 19200 685570
rect 19270 685500 19290 685570
rect 19360 685500 19380 685570
rect 19450 685500 19470 685570
rect 19540 685500 19560 685570
rect 19630 685500 23946 685570
rect 18050 685480 23946 685500
rect 18050 685410 18120 685480
rect 18190 685410 18210 685480
rect 18280 685410 18300 685480
rect 18370 685410 18390 685480
rect 18460 685410 18480 685480
rect 18550 685410 18570 685480
rect 18640 685410 18660 685480
rect 18730 685410 18750 685480
rect 18820 685410 18840 685480
rect 18910 685410 18930 685480
rect 19000 685410 19020 685480
rect 19090 685410 19110 685480
rect 19180 685410 19200 685480
rect 19270 685410 19290 685480
rect 19360 685410 19380 685480
rect 19450 685410 19470 685480
rect 19540 685410 19560 685480
rect 19630 685410 23946 685480
rect 18050 685390 23946 685410
rect -800 683660 1700 685242
rect -800 683590 120 683660
rect 190 683590 210 683660
rect 280 683590 300 683660
rect 370 683590 390 683660
rect 460 683590 480 683660
rect 550 683590 570 683660
rect 640 683590 660 683660
rect 730 683590 750 683660
rect 820 683590 840 683660
rect 910 683590 930 683660
rect 1000 683590 1020 683660
rect 1090 683590 1110 683660
rect 1180 683590 1200 683660
rect 1270 683590 1290 683660
rect 1360 683590 1380 683660
rect 1450 683590 1470 683660
rect 1540 683590 1560 683660
rect 1630 683590 1700 683660
rect -800 683570 1700 683590
rect -800 683500 120 683570
rect 190 683500 210 683570
rect 280 683500 300 683570
rect 370 683500 390 683570
rect 460 683500 480 683570
rect 550 683500 570 683570
rect 640 683500 660 683570
rect 730 683500 750 683570
rect 820 683500 840 683570
rect 910 683500 930 683570
rect 1000 683500 1020 683570
rect 1090 683500 1110 683570
rect 1180 683500 1200 683570
rect 1270 683500 1290 683570
rect 1360 683500 1380 683570
rect 1450 683500 1470 683570
rect 1540 683500 1560 683570
rect 1630 683500 1700 683570
rect -800 683480 1700 683500
rect -800 683410 120 683480
rect 190 683410 210 683480
rect 280 683410 300 683480
rect 370 683410 390 683480
rect 460 683410 480 683480
rect 550 683410 570 683480
rect 640 683410 660 683480
rect 730 683410 750 683480
rect 820 683410 840 683480
rect 910 683410 930 683480
rect 1000 683410 1020 683480
rect 1090 683410 1110 683480
rect 1180 683410 1200 683480
rect 1270 683410 1290 683480
rect 1360 683410 1380 683480
rect 1450 683410 1470 683480
rect 1540 683410 1560 683480
rect 1630 683410 1700 683480
rect -800 683390 1700 683410
rect -800 683320 120 683390
rect 190 683320 210 683390
rect 280 683320 300 683390
rect 370 683320 390 683390
rect 460 683320 480 683390
rect 550 683320 570 683390
rect 640 683320 660 683390
rect 730 683320 750 683390
rect 820 683320 840 683390
rect 910 683320 930 683390
rect 1000 683320 1020 683390
rect 1090 683320 1110 683390
rect 1180 683320 1200 683390
rect 1270 683320 1290 683390
rect 1360 683320 1380 683390
rect 1450 683320 1470 683390
rect 1540 683320 1560 683390
rect 1630 683320 1700 683390
rect -800 683300 1700 683320
rect -800 683230 120 683300
rect 190 683230 210 683300
rect 280 683230 300 683300
rect 370 683230 390 683300
rect 460 683230 480 683300
rect 550 683230 570 683300
rect 640 683230 660 683300
rect 730 683230 750 683300
rect 820 683230 840 683300
rect 910 683230 930 683300
rect 1000 683230 1020 683300
rect 1090 683230 1110 683300
rect 1180 683230 1200 683300
rect 1270 683230 1290 683300
rect 1360 683230 1380 683300
rect 1450 683230 1470 683300
rect 1540 683230 1560 683300
rect 1630 683230 1700 683300
rect -800 683210 1700 683230
rect -800 683140 120 683210
rect 190 683140 210 683210
rect 280 683140 300 683210
rect 370 683140 390 683210
rect 460 683140 480 683210
rect 550 683140 570 683210
rect 640 683140 660 683210
rect 730 683140 750 683210
rect 820 683140 840 683210
rect 910 683140 930 683210
rect 1000 683140 1020 683210
rect 1090 683140 1110 683210
rect 1180 683140 1200 683210
rect 1270 683140 1290 683210
rect 1360 683140 1380 683210
rect 1450 683140 1470 683210
rect 1540 683140 1560 683210
rect 1630 683140 1700 683210
rect -800 683120 1700 683140
rect -800 683050 120 683120
rect 190 683050 210 683120
rect 280 683050 300 683120
rect 370 683050 390 683120
rect 460 683050 480 683120
rect 550 683050 570 683120
rect 640 683050 660 683120
rect 730 683050 750 683120
rect 820 683050 840 683120
rect 910 683050 930 683120
rect 1000 683050 1020 683120
rect 1090 683050 1110 683120
rect 1180 683050 1200 683120
rect 1270 683050 1290 683120
rect 1360 683050 1380 683120
rect 1450 683050 1470 683120
rect 1540 683050 1560 683120
rect 1630 683050 1700 683120
rect -800 683030 1700 683050
rect -800 682960 120 683030
rect 190 682960 210 683030
rect 280 682960 300 683030
rect 370 682960 390 683030
rect 460 682960 480 683030
rect 550 682960 570 683030
rect 640 682960 660 683030
rect 730 682960 750 683030
rect 820 682960 840 683030
rect 910 682960 930 683030
rect 1000 682960 1020 683030
rect 1090 682960 1110 683030
rect 1180 682960 1200 683030
rect 1270 682960 1290 683030
rect 1360 682960 1380 683030
rect 1450 682960 1470 683030
rect 1540 682960 1560 683030
rect 1630 682960 1700 683030
rect -800 682940 1700 682960
rect -800 682870 120 682940
rect 190 682870 210 682940
rect 280 682870 300 682940
rect 370 682870 390 682940
rect 460 682870 480 682940
rect 550 682870 570 682940
rect 640 682870 660 682940
rect 730 682870 750 682940
rect 820 682870 840 682940
rect 910 682870 930 682940
rect 1000 682870 1020 682940
rect 1090 682870 1110 682940
rect 1180 682870 1200 682940
rect 1270 682870 1290 682940
rect 1360 682870 1380 682940
rect 1450 682870 1470 682940
rect 1540 682870 1560 682940
rect 1630 682870 1700 682940
rect -800 682850 1700 682870
rect -800 682780 120 682850
rect 190 682780 210 682850
rect 280 682780 300 682850
rect 370 682780 390 682850
rect 460 682780 480 682850
rect 550 682780 570 682850
rect 640 682780 660 682850
rect 730 682780 750 682850
rect 820 682780 840 682850
rect 910 682780 930 682850
rect 1000 682780 1020 682850
rect 1090 682780 1110 682850
rect 1180 682780 1200 682850
rect 1270 682780 1290 682850
rect 1360 682780 1380 682850
rect 1450 682780 1470 682850
rect 1540 682780 1560 682850
rect 1630 682780 1700 682850
rect -800 682760 1700 682780
rect -800 682690 120 682760
rect 190 682690 210 682760
rect 280 682690 300 682760
rect 370 682690 390 682760
rect 460 682690 480 682760
rect 550 682690 570 682760
rect 640 682690 660 682760
rect 730 682690 750 682760
rect 820 682690 840 682760
rect 910 682690 930 682760
rect 1000 682690 1020 682760
rect 1090 682690 1110 682760
rect 1180 682690 1200 682760
rect 1270 682690 1290 682760
rect 1360 682690 1380 682760
rect 1450 682690 1470 682760
rect 1540 682690 1560 682760
rect 1630 682690 1700 682760
rect -800 682670 1700 682690
rect -800 682600 120 682670
rect 190 682600 210 682670
rect 280 682600 300 682670
rect 370 682600 390 682670
rect 460 682600 480 682670
rect 550 682600 570 682670
rect 640 682600 660 682670
rect 730 682600 750 682670
rect 820 682600 840 682670
rect 910 682600 930 682670
rect 1000 682600 1020 682670
rect 1090 682600 1110 682670
rect 1180 682600 1200 682670
rect 1270 682600 1290 682670
rect 1360 682600 1380 682670
rect 1450 682600 1470 682670
rect 1540 682600 1560 682670
rect 1630 682600 1700 682670
rect -800 682580 1700 682600
rect -800 682510 120 682580
rect 190 682510 210 682580
rect 280 682510 300 682580
rect 370 682510 390 682580
rect 460 682510 480 682580
rect 550 682510 570 682580
rect 640 682510 660 682580
rect 730 682510 750 682580
rect 820 682510 840 682580
rect 910 682510 930 682580
rect 1000 682510 1020 682580
rect 1090 682510 1110 682580
rect 1180 682510 1200 682580
rect 1270 682510 1290 682580
rect 1360 682510 1380 682580
rect 1450 682510 1470 682580
rect 1540 682510 1560 682580
rect 1630 682510 1700 682580
rect -800 682490 1700 682510
rect -800 682420 120 682490
rect 190 682420 210 682490
rect 280 682420 300 682490
rect 370 682420 390 682490
rect 460 682420 480 682490
rect 550 682420 570 682490
rect 640 682420 660 682490
rect 730 682420 750 682490
rect 820 682420 840 682490
rect 910 682420 930 682490
rect 1000 682420 1020 682490
rect 1090 682420 1110 682490
rect 1180 682420 1200 682490
rect 1270 682420 1290 682490
rect 1360 682420 1380 682490
rect 1450 682420 1470 682490
rect 1540 682420 1560 682490
rect 1630 682420 1700 682490
rect -800 682400 1700 682420
rect -800 682330 120 682400
rect 190 682330 210 682400
rect 280 682330 300 682400
rect 370 682330 390 682400
rect 460 682330 480 682400
rect 550 682330 570 682400
rect 640 682330 660 682400
rect 730 682330 750 682400
rect 820 682330 840 682400
rect 910 682330 930 682400
rect 1000 682330 1020 682400
rect 1090 682330 1110 682400
rect 1180 682330 1200 682400
rect 1270 682330 1290 682400
rect 1360 682330 1380 682400
rect 1450 682330 1470 682400
rect 1540 682330 1560 682400
rect 1630 682330 1700 682400
rect -800 682310 1700 682330
rect -800 682240 120 682310
rect 190 682240 210 682310
rect 280 682240 300 682310
rect 370 682240 390 682310
rect 460 682240 480 682310
rect 550 682240 570 682310
rect 640 682240 660 682310
rect 730 682240 750 682310
rect 820 682240 840 682310
rect 910 682240 930 682310
rect 1000 682240 1020 682310
rect 1090 682240 1110 682310
rect 1180 682240 1200 682310
rect 1270 682240 1290 682310
rect 1360 682240 1380 682310
rect 1450 682240 1470 682310
rect 1540 682240 1560 682310
rect 1630 682240 1700 682310
rect -800 682220 1700 682240
rect -800 682150 120 682220
rect 190 682150 210 682220
rect 280 682150 300 682220
rect 370 682150 390 682220
rect 460 682150 480 682220
rect 550 682150 570 682220
rect 640 682150 660 682220
rect 730 682150 750 682220
rect 820 682150 840 682220
rect 910 682150 930 682220
rect 1000 682150 1020 682220
rect 1090 682150 1110 682220
rect 1180 682150 1200 682220
rect 1270 682150 1290 682220
rect 1360 682150 1380 682220
rect 1450 682150 1470 682220
rect 1540 682150 1560 682220
rect 1630 682150 1700 682220
rect -800 680242 1700 682150
rect 17650 683660 19650 683730
rect 17650 683590 17670 683660
rect 17740 683590 17760 683660
rect 17830 683590 17850 683660
rect 17920 683590 17940 683660
rect 18010 683590 18030 683660
rect 18100 683590 18120 683660
rect 18190 683590 18210 683660
rect 18280 683590 18300 683660
rect 18370 683590 18390 683660
rect 18460 683590 18480 683660
rect 18550 683590 18570 683660
rect 18640 683590 18660 683660
rect 18730 683590 18750 683660
rect 18820 683590 18840 683660
rect 18910 683590 18930 683660
rect 19000 683590 19020 683660
rect 19090 683590 19110 683660
rect 19180 683590 19200 683660
rect 19270 683590 19290 683660
rect 19360 683590 19380 683660
rect 19450 683590 19470 683660
rect 19540 683590 19560 683660
rect 19630 683590 19650 683660
rect 17650 683570 19650 683590
rect 17650 683500 17670 683570
rect 17740 683500 17760 683570
rect 17830 683500 17850 683570
rect 17920 683500 17940 683570
rect 18010 683500 18030 683570
rect 18100 683500 18120 683570
rect 18190 683500 18210 683570
rect 18280 683500 18300 683570
rect 18370 683500 18390 683570
rect 18460 683500 18480 683570
rect 18550 683500 18570 683570
rect 18640 683500 18660 683570
rect 18730 683500 18750 683570
rect 18820 683500 18840 683570
rect 18910 683500 18930 683570
rect 19000 683500 19020 683570
rect 19090 683500 19110 683570
rect 19180 683500 19200 683570
rect 19270 683500 19290 683570
rect 19360 683500 19380 683570
rect 19450 683500 19470 683570
rect 19540 683500 19560 683570
rect 19630 683500 19650 683570
rect 17650 683480 19650 683500
rect 17650 683410 17670 683480
rect 17740 683410 17760 683480
rect 17830 683410 17850 683480
rect 17920 683410 17940 683480
rect 18010 683410 18030 683480
rect 18100 683410 18120 683480
rect 18190 683410 18210 683480
rect 18280 683410 18300 683480
rect 18370 683410 18390 683480
rect 18460 683410 18480 683480
rect 18550 683410 18570 683480
rect 18640 683410 18660 683480
rect 18730 683410 18750 683480
rect 18820 683410 18840 683480
rect 18910 683410 18930 683480
rect 19000 683410 19020 683480
rect 19090 683410 19110 683480
rect 19180 683410 19200 683480
rect 19270 683410 19290 683480
rect 19360 683410 19380 683480
rect 19450 683410 19470 683480
rect 19540 683410 19560 683480
rect 19630 683410 19650 683480
rect 17650 683390 19650 683410
rect 17650 683320 17670 683390
rect 17740 683320 17760 683390
rect 17830 683320 17850 683390
rect 17920 683320 17940 683390
rect 18010 683320 18030 683390
rect 18100 683320 18120 683390
rect 18190 683320 18210 683390
rect 18280 683320 18300 683390
rect 18370 683320 18390 683390
rect 18460 683320 18480 683390
rect 18550 683320 18570 683390
rect 18640 683320 18660 683390
rect 18730 683320 18750 683390
rect 18820 683320 18840 683390
rect 18910 683320 18930 683390
rect 19000 683320 19020 683390
rect 19090 683320 19110 683390
rect 19180 683320 19200 683390
rect 19270 683320 19290 683390
rect 19360 683320 19380 683390
rect 19450 683320 19470 683390
rect 19540 683320 19560 683390
rect 19630 683320 19650 683390
rect 17650 683300 19650 683320
rect 17650 683230 17670 683300
rect 17740 683230 17760 683300
rect 17830 683230 17850 683300
rect 17920 683230 17940 683300
rect 18010 683230 18030 683300
rect 18100 683230 18120 683300
rect 18190 683230 18210 683300
rect 18280 683230 18300 683300
rect 18370 683230 18390 683300
rect 18460 683230 18480 683300
rect 18550 683230 18570 683300
rect 18640 683230 18660 683300
rect 18730 683230 18750 683300
rect 18820 683230 18840 683300
rect 18910 683230 18930 683300
rect 19000 683230 19020 683300
rect 19090 683230 19110 683300
rect 19180 683230 19200 683300
rect 19270 683230 19290 683300
rect 19360 683230 19380 683300
rect 19450 683230 19470 683300
rect 19540 683230 19560 683300
rect 19630 683230 19650 683300
rect 17650 683210 19650 683230
rect 17650 683140 17670 683210
rect 17740 683140 17760 683210
rect 17830 683140 17850 683210
rect 17920 683140 17940 683210
rect 18010 683140 18030 683210
rect 18100 683140 18120 683210
rect 18190 683140 18210 683210
rect 18280 683140 18300 683210
rect 18370 683140 18390 683210
rect 18460 683140 18480 683210
rect 18550 683140 18570 683210
rect 18640 683140 18660 683210
rect 18730 683140 18750 683210
rect 18820 683140 18840 683210
rect 18910 683140 18930 683210
rect 19000 683140 19020 683210
rect 19090 683140 19110 683210
rect 19180 683140 19200 683210
rect 19270 683140 19290 683210
rect 19360 683140 19380 683210
rect 19450 683140 19470 683210
rect 19540 683140 19560 683210
rect 19630 683140 19650 683210
rect 17650 683120 19650 683140
rect 17650 683050 17670 683120
rect 17740 683050 17760 683120
rect 17830 683050 17850 683120
rect 17920 683050 17940 683120
rect 18010 683050 18030 683120
rect 18100 683050 18120 683120
rect 18190 683050 18210 683120
rect 18280 683050 18300 683120
rect 18370 683050 18390 683120
rect 18460 683050 18480 683120
rect 18550 683050 18570 683120
rect 18640 683050 18660 683120
rect 18730 683050 18750 683120
rect 18820 683050 18840 683120
rect 18910 683050 18930 683120
rect 19000 683050 19020 683120
rect 19090 683050 19110 683120
rect 19180 683050 19200 683120
rect 19270 683050 19290 683120
rect 19360 683050 19380 683120
rect 19450 683050 19470 683120
rect 19540 683050 19560 683120
rect 19630 683050 19650 683120
rect 17650 683030 19650 683050
rect 17650 682960 17670 683030
rect 17740 682960 17760 683030
rect 17830 682960 17850 683030
rect 17920 682960 17940 683030
rect 18010 682960 18030 683030
rect 18100 682960 18120 683030
rect 18190 682960 18210 683030
rect 18280 682960 18300 683030
rect 18370 682960 18390 683030
rect 18460 682960 18480 683030
rect 18550 682960 18570 683030
rect 18640 682960 18660 683030
rect 18730 682960 18750 683030
rect 18820 682960 18840 683030
rect 18910 682960 18930 683030
rect 19000 682960 19020 683030
rect 19090 682960 19110 683030
rect 19180 682960 19200 683030
rect 19270 682960 19290 683030
rect 19360 682960 19380 683030
rect 19450 682960 19470 683030
rect 19540 682960 19560 683030
rect 19630 682960 19650 683030
rect 17650 682940 19650 682960
rect 17650 682870 17670 682940
rect 17740 682870 17760 682940
rect 17830 682870 17850 682940
rect 17920 682870 17940 682940
rect 18010 682870 18030 682940
rect 18100 682870 18120 682940
rect 18190 682870 18210 682940
rect 18280 682870 18300 682940
rect 18370 682870 18390 682940
rect 18460 682870 18480 682940
rect 18550 682870 18570 682940
rect 18640 682870 18660 682940
rect 18730 682870 18750 682940
rect 18820 682870 18840 682940
rect 18910 682870 18930 682940
rect 19000 682870 19020 682940
rect 19090 682870 19110 682940
rect 19180 682870 19200 682940
rect 19270 682870 19290 682940
rect 19360 682870 19380 682940
rect 19450 682870 19470 682940
rect 19540 682870 19560 682940
rect 19630 682870 19650 682940
rect 17650 682850 19650 682870
rect 17650 682780 17670 682850
rect 17740 682780 17760 682850
rect 17830 682780 17850 682850
rect 17920 682780 17940 682850
rect 18010 682780 18030 682850
rect 18100 682780 18120 682850
rect 18190 682780 18210 682850
rect 18280 682780 18300 682850
rect 18370 682780 18390 682850
rect 18460 682780 18480 682850
rect 18550 682780 18570 682850
rect 18640 682780 18660 682850
rect 18730 682780 18750 682850
rect 18820 682780 18840 682850
rect 18910 682780 18930 682850
rect 19000 682780 19020 682850
rect 19090 682780 19110 682850
rect 19180 682780 19200 682850
rect 19270 682780 19290 682850
rect 19360 682780 19380 682850
rect 19450 682780 19470 682850
rect 19540 682780 19560 682850
rect 19630 682780 19650 682850
rect 17650 682760 19650 682780
rect 17650 682690 17670 682760
rect 17740 682690 17760 682760
rect 17830 682690 17850 682760
rect 17920 682690 17940 682760
rect 18010 682690 18030 682760
rect 18100 682690 18120 682760
rect 18190 682690 18210 682760
rect 18280 682690 18300 682760
rect 18370 682690 18390 682760
rect 18460 682690 18480 682760
rect 18550 682690 18570 682760
rect 18640 682690 18660 682760
rect 18730 682690 18750 682760
rect 18820 682690 18840 682760
rect 18910 682690 18930 682760
rect 19000 682690 19020 682760
rect 19090 682690 19110 682760
rect 19180 682690 19200 682760
rect 19270 682690 19290 682760
rect 19360 682690 19380 682760
rect 19450 682690 19470 682760
rect 19540 682690 19560 682760
rect 19630 682690 19650 682760
rect 17650 682670 19650 682690
rect 17650 682600 17670 682670
rect 17740 682600 17760 682670
rect 17830 682600 17850 682670
rect 17920 682600 17940 682670
rect 18010 682600 18030 682670
rect 18100 682600 18120 682670
rect 18190 682600 18210 682670
rect 18280 682600 18300 682670
rect 18370 682600 18390 682670
rect 18460 682600 18480 682670
rect 18550 682600 18570 682670
rect 18640 682600 18660 682670
rect 18730 682600 18750 682670
rect 18820 682600 18840 682670
rect 18910 682600 18930 682670
rect 19000 682600 19020 682670
rect 19090 682600 19110 682670
rect 19180 682600 19200 682670
rect 19270 682600 19290 682670
rect 19360 682600 19380 682670
rect 19450 682600 19470 682670
rect 19540 682600 19560 682670
rect 19630 682600 19650 682670
rect 17650 682580 19650 682600
rect 17650 682510 17670 682580
rect 17740 682510 17760 682580
rect 17830 682510 17850 682580
rect 17920 682510 17940 682580
rect 18010 682510 18030 682580
rect 18100 682510 18120 682580
rect 18190 682510 18210 682580
rect 18280 682510 18300 682580
rect 18370 682510 18390 682580
rect 18460 682510 18480 682580
rect 18550 682510 18570 682580
rect 18640 682510 18660 682580
rect 18730 682510 18750 682580
rect 18820 682510 18840 682580
rect 18910 682510 18930 682580
rect 19000 682510 19020 682580
rect 19090 682510 19110 682580
rect 19180 682510 19200 682580
rect 19270 682510 19290 682580
rect 19360 682510 19380 682580
rect 19450 682510 19470 682580
rect 19540 682510 19560 682580
rect 19630 682510 19650 682580
rect 17650 682490 19650 682510
rect 17650 682420 17670 682490
rect 17740 682420 17760 682490
rect 17830 682420 17850 682490
rect 17920 682420 17940 682490
rect 18010 682420 18030 682490
rect 18100 682420 18120 682490
rect 18190 682420 18210 682490
rect 18280 682420 18300 682490
rect 18370 682420 18390 682490
rect 18460 682420 18480 682490
rect 18550 682420 18570 682490
rect 18640 682420 18660 682490
rect 18730 682420 18750 682490
rect 18820 682420 18840 682490
rect 18910 682420 18930 682490
rect 19000 682420 19020 682490
rect 19090 682420 19110 682490
rect 19180 682420 19200 682490
rect 19270 682420 19290 682490
rect 19360 682420 19380 682490
rect 19450 682420 19470 682490
rect 19540 682420 19560 682490
rect 19630 682420 19650 682490
rect 17650 682400 19650 682420
rect 17650 682330 17670 682400
rect 17740 682330 17760 682400
rect 17830 682330 17850 682400
rect 17920 682330 17940 682400
rect 18010 682330 18030 682400
rect 18100 682330 18120 682400
rect 18190 682330 18210 682400
rect 18280 682330 18300 682400
rect 18370 682330 18390 682400
rect 18460 682330 18480 682400
rect 18550 682330 18570 682400
rect 18640 682330 18660 682400
rect 18730 682330 18750 682400
rect 18820 682330 18840 682400
rect 18910 682330 18930 682400
rect 19000 682330 19020 682400
rect 19090 682330 19110 682400
rect 19180 682330 19200 682400
rect 19270 682330 19290 682400
rect 19360 682330 19380 682400
rect 19450 682330 19470 682400
rect 19540 682330 19560 682400
rect 19630 682330 19650 682400
rect 17650 682310 19650 682330
rect 17650 682240 17670 682310
rect 17740 682240 17760 682310
rect 17830 682240 17850 682310
rect 17920 682240 17940 682310
rect 18010 682240 18030 682310
rect 18100 682240 18120 682310
rect 18190 682240 18210 682310
rect 18280 682240 18300 682310
rect 18370 682240 18390 682310
rect 18460 682240 18480 682310
rect 18550 682240 18570 682310
rect 18640 682240 18660 682310
rect 18730 682240 18750 682310
rect 18820 682240 18840 682310
rect 18910 682240 18930 682310
rect 19000 682240 19020 682310
rect 19090 682240 19110 682310
rect 19180 682240 19200 682310
rect 19270 682240 19290 682310
rect 19360 682240 19380 682310
rect 19450 682240 19470 682310
rect 19540 682240 19560 682310
rect 19630 682240 19650 682310
rect 17650 682220 19650 682240
rect 17650 682150 17670 682220
rect 17740 682150 17760 682220
rect 17830 682150 17850 682220
rect 17920 682150 17940 682220
rect 18010 682150 18030 682220
rect 18100 682150 18120 682220
rect 18190 682150 18210 682220
rect 18280 682150 18300 682220
rect 18370 682150 18390 682220
rect 18460 682150 18480 682220
rect 18550 682150 18570 682220
rect 18640 682150 18660 682220
rect 18730 682150 18750 682220
rect 18820 682150 18840 682220
rect 18910 682150 18930 682220
rect 19000 682150 19020 682220
rect 19090 682150 19110 682220
rect 19180 682150 19200 682220
rect 19270 682150 19290 682220
rect 19360 682150 19380 682220
rect 19450 682150 19470 682220
rect 19540 682150 19560 682220
rect 19630 682150 19650 682220
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 17650 619420 19650 682150
rect 21946 623528 23946 685390
rect 582300 679516 584800 682984
rect 582300 679446 582320 679516
rect 582390 679446 582410 679516
rect 582480 679446 582500 679516
rect 582570 679446 582590 679516
rect 582660 679446 582680 679516
rect 582750 679446 582770 679516
rect 582840 679446 584800 679516
rect 582300 679426 584800 679446
rect 582300 679356 582320 679426
rect 582390 679356 582410 679426
rect 582480 679356 582500 679426
rect 582570 679356 582590 679426
rect 582660 679356 582680 679426
rect 582750 679356 582770 679426
rect 582840 679356 584800 679426
rect 582300 679336 584800 679356
rect 582300 679266 582320 679336
rect 582390 679266 582410 679336
rect 582480 679266 582500 679336
rect 582570 679266 582590 679336
rect 582660 679266 582680 679336
rect 582750 679266 582770 679336
rect 582840 679266 584800 679336
rect 582300 679246 584800 679266
rect 582300 679176 582320 679246
rect 582390 679176 582410 679246
rect 582480 679176 582500 679246
rect 582570 679176 582590 679246
rect 582660 679176 582680 679246
rect 582750 679176 582770 679246
rect 582840 679176 584800 679246
rect 582300 679156 584800 679176
rect 582300 679086 582320 679156
rect 582390 679086 582410 679156
rect 582480 679086 582500 679156
rect 582570 679086 582590 679156
rect 582660 679086 582680 679156
rect 582750 679086 582770 679156
rect 582840 679086 584800 679156
rect 582300 679066 584800 679086
rect 582300 678996 582320 679066
rect 582390 678996 582410 679066
rect 582480 678996 582500 679066
rect 582570 678996 582590 679066
rect 582660 678996 582680 679066
rect 582750 678996 582770 679066
rect 582840 678996 584800 679066
rect 582300 677984 584800 678996
rect 582340 639784 584800 644584
rect 94254 638170 94574 638390
rect 94254 638100 94280 638170
rect 94350 638100 94380 638170
rect 94450 638100 94480 638170
rect 94550 638100 94574 638170
rect 94254 638080 94574 638100
rect 94254 638010 94280 638080
rect 94350 638010 94380 638080
rect 94450 638010 94480 638080
rect 94550 638010 94574 638080
rect 94254 637980 94574 638010
rect 98814 638170 99134 638390
rect 98814 638100 98838 638170
rect 98908 638100 98938 638170
rect 99008 638100 99038 638170
rect 99108 638100 99134 638170
rect 98814 638080 99134 638100
rect 98814 638010 98838 638080
rect 98908 638010 98938 638080
rect 99008 638010 99038 638080
rect 99108 638010 99134 638080
rect 98814 637980 99134 638010
rect 582340 629784 584800 634584
rect 21946 623458 21966 623528
rect 22036 623458 22056 623528
rect 22126 623458 22146 623528
rect 22216 623458 22236 623528
rect 22306 623458 22326 623528
rect 22396 623458 22416 623528
rect 22486 623458 22506 623528
rect 22576 623458 22596 623528
rect 22666 623458 22686 623528
rect 22756 623458 22776 623528
rect 22846 623458 22866 623528
rect 22936 623458 22956 623528
rect 23026 623458 23046 623528
rect 23116 623458 23136 623528
rect 23206 623458 23226 623528
rect 23296 623458 23316 623528
rect 23386 623458 23406 623528
rect 23476 623458 23496 623528
rect 23566 623458 23586 623528
rect 23656 623458 23676 623528
rect 23746 623458 23766 623528
rect 23836 623458 23856 623528
rect 23926 623458 23946 623528
rect 21946 623438 23946 623458
rect 21946 623368 21966 623438
rect 22036 623368 22056 623438
rect 22126 623368 22146 623438
rect 22216 623368 22236 623438
rect 22306 623368 22326 623438
rect 22396 623368 22416 623438
rect 22486 623368 22506 623438
rect 22576 623368 22596 623438
rect 22666 623368 22686 623438
rect 22756 623368 22776 623438
rect 22846 623368 22866 623438
rect 22936 623368 22956 623438
rect 23026 623368 23046 623438
rect 23116 623368 23136 623438
rect 23206 623368 23226 623438
rect 23296 623368 23316 623438
rect 23386 623368 23406 623438
rect 23476 623368 23496 623438
rect 23566 623368 23586 623438
rect 23656 623368 23676 623438
rect 23746 623368 23766 623438
rect 23836 623368 23856 623438
rect 23926 623368 23946 623438
rect 21946 623348 23946 623368
rect 21946 623278 21966 623348
rect 22036 623278 22056 623348
rect 22126 623278 22146 623348
rect 22216 623278 22236 623348
rect 22306 623278 22326 623348
rect 22396 623278 22416 623348
rect 22486 623278 22506 623348
rect 22576 623278 22596 623348
rect 22666 623278 22686 623348
rect 22756 623278 22776 623348
rect 22846 623278 22866 623348
rect 22936 623278 22956 623348
rect 23026 623278 23046 623348
rect 23116 623278 23136 623348
rect 23206 623278 23226 623348
rect 23296 623278 23316 623348
rect 23386 623278 23406 623348
rect 23476 623278 23496 623348
rect 23566 623278 23586 623348
rect 23656 623278 23676 623348
rect 23746 623278 23766 623348
rect 23836 623278 23856 623348
rect 23926 623278 23946 623348
rect 21946 623258 23946 623278
rect 21946 623188 21966 623258
rect 22036 623188 22056 623258
rect 22126 623188 22146 623258
rect 22216 623188 22236 623258
rect 22306 623188 22326 623258
rect 22396 623188 22416 623258
rect 22486 623188 22506 623258
rect 22576 623188 22596 623258
rect 22666 623188 22686 623258
rect 22756 623188 22776 623258
rect 22846 623188 22866 623258
rect 22936 623188 22956 623258
rect 23026 623188 23046 623258
rect 23116 623188 23136 623258
rect 23206 623188 23226 623258
rect 23296 623188 23316 623258
rect 23386 623188 23406 623258
rect 23476 623188 23496 623258
rect 23566 623188 23586 623258
rect 23656 623188 23676 623258
rect 23746 623188 23766 623258
rect 23836 623188 23856 623258
rect 23926 623188 23946 623258
rect 21946 623168 23946 623188
rect 21946 623098 21966 623168
rect 22036 623098 22056 623168
rect 22126 623098 22146 623168
rect 22216 623098 22236 623168
rect 22306 623098 22326 623168
rect 22396 623098 22416 623168
rect 22486 623098 22506 623168
rect 22576 623098 22596 623168
rect 22666 623098 22686 623168
rect 22756 623098 22776 623168
rect 22846 623098 22866 623168
rect 22936 623098 22956 623168
rect 23026 623098 23046 623168
rect 23116 623098 23136 623168
rect 23206 623098 23226 623168
rect 23296 623098 23316 623168
rect 23386 623098 23406 623168
rect 23476 623098 23496 623168
rect 23566 623098 23586 623168
rect 23656 623098 23676 623168
rect 23746 623098 23766 623168
rect 23836 623098 23856 623168
rect 23926 623098 23946 623168
rect 21946 623078 23946 623098
rect 21946 623008 21966 623078
rect 22036 623008 22056 623078
rect 22126 623008 22146 623078
rect 22216 623008 22236 623078
rect 22306 623008 22326 623078
rect 22396 623008 22416 623078
rect 22486 623008 22506 623078
rect 22576 623008 22596 623078
rect 22666 623008 22686 623078
rect 22756 623008 22776 623078
rect 22846 623008 22866 623078
rect 22936 623008 22956 623078
rect 23026 623008 23046 623078
rect 23116 623008 23136 623078
rect 23206 623008 23226 623078
rect 23296 623008 23316 623078
rect 23386 623008 23406 623078
rect 23476 623008 23496 623078
rect 23566 623008 23586 623078
rect 23656 623008 23676 623078
rect 23746 623008 23766 623078
rect 23836 623008 23856 623078
rect 23926 623008 23946 623078
rect 21946 622988 23946 623008
rect 21946 622918 21966 622988
rect 22036 622918 22056 622988
rect 22126 622918 22146 622988
rect 22216 622918 22236 622988
rect 22306 622918 22326 622988
rect 22396 622918 22416 622988
rect 22486 622918 22506 622988
rect 22576 622918 22596 622988
rect 22666 622918 22686 622988
rect 22756 622918 22776 622988
rect 22846 622918 22866 622988
rect 22936 622918 22956 622988
rect 23026 622918 23046 622988
rect 23116 622918 23136 622988
rect 23206 622918 23226 622988
rect 23296 622918 23316 622988
rect 23386 622918 23406 622988
rect 23476 622918 23496 622988
rect 23566 622918 23586 622988
rect 23656 622918 23676 622988
rect 23746 622918 23766 622988
rect 23836 622918 23856 622988
rect 23926 622918 23946 622988
rect 21946 622898 23946 622918
rect 21946 622828 21966 622898
rect 22036 622828 22056 622898
rect 22126 622828 22146 622898
rect 22216 622828 22236 622898
rect 22306 622828 22326 622898
rect 22396 622828 22416 622898
rect 22486 622828 22506 622898
rect 22576 622828 22596 622898
rect 22666 622828 22686 622898
rect 22756 622828 22776 622898
rect 22846 622828 22866 622898
rect 22936 622828 22956 622898
rect 23026 622828 23046 622898
rect 23116 622828 23136 622898
rect 23206 622828 23226 622898
rect 23296 622828 23316 622898
rect 23386 622828 23406 622898
rect 23476 622828 23496 622898
rect 23566 622828 23586 622898
rect 23656 622828 23676 622898
rect 23746 622828 23766 622898
rect 23836 622828 23856 622898
rect 23926 622828 23946 622898
rect 21946 622808 23946 622828
rect 21946 622738 21966 622808
rect 22036 622738 22056 622808
rect 22126 622738 22146 622808
rect 22216 622738 22236 622808
rect 22306 622738 22326 622808
rect 22396 622738 22416 622808
rect 22486 622738 22506 622808
rect 22576 622738 22596 622808
rect 22666 622738 22686 622808
rect 22756 622738 22776 622808
rect 22846 622738 22866 622808
rect 22936 622738 22956 622808
rect 23026 622738 23046 622808
rect 23116 622738 23136 622808
rect 23206 622738 23226 622808
rect 23296 622738 23316 622808
rect 23386 622738 23406 622808
rect 23476 622738 23496 622808
rect 23566 622738 23586 622808
rect 23656 622738 23676 622808
rect 23746 622738 23766 622808
rect 23836 622738 23856 622808
rect 23926 622738 23946 622808
rect 21946 622718 23946 622738
rect 21946 622648 21966 622718
rect 22036 622648 22056 622718
rect 22126 622648 22146 622718
rect 22216 622648 22236 622718
rect 22306 622648 22326 622718
rect 22396 622648 22416 622718
rect 22486 622648 22506 622718
rect 22576 622648 22596 622718
rect 22666 622648 22686 622718
rect 22756 622648 22776 622718
rect 22846 622648 22866 622718
rect 22936 622648 22956 622718
rect 23026 622648 23046 622718
rect 23116 622648 23136 622718
rect 23206 622648 23226 622718
rect 23296 622648 23316 622718
rect 23386 622648 23406 622718
rect 23476 622648 23496 622718
rect 23566 622648 23586 622718
rect 23656 622648 23676 622718
rect 23746 622648 23766 622718
rect 23836 622648 23856 622718
rect 23926 622648 23946 622718
rect 21946 622628 23946 622648
rect 21946 622558 21966 622628
rect 22036 622558 22056 622628
rect 22126 622558 22146 622628
rect 22216 622558 22236 622628
rect 22306 622558 22326 622628
rect 22396 622558 22416 622628
rect 22486 622558 22506 622628
rect 22576 622558 22596 622628
rect 22666 622558 22686 622628
rect 22756 622558 22776 622628
rect 22846 622558 22866 622628
rect 22936 622558 22956 622628
rect 23026 622558 23046 622628
rect 23116 622558 23136 622628
rect 23206 622558 23226 622628
rect 23296 622558 23316 622628
rect 23386 622558 23406 622628
rect 23476 622558 23496 622628
rect 23566 622558 23586 622628
rect 23656 622558 23676 622628
rect 23746 622558 23766 622628
rect 23836 622558 23856 622628
rect 23926 622558 23946 622628
rect 21946 622538 23946 622558
rect 21946 622468 21966 622538
rect 22036 622468 22056 622538
rect 22126 622468 22146 622538
rect 22216 622468 22236 622538
rect 22306 622468 22326 622538
rect 22396 622468 22416 622538
rect 22486 622468 22506 622538
rect 22576 622468 22596 622538
rect 22666 622468 22686 622538
rect 22756 622468 22776 622538
rect 22846 622468 22866 622538
rect 22936 622468 22956 622538
rect 23026 622468 23046 622538
rect 23116 622468 23136 622538
rect 23206 622468 23226 622538
rect 23296 622468 23316 622538
rect 23386 622468 23406 622538
rect 23476 622468 23496 622538
rect 23566 622468 23586 622538
rect 23656 622468 23676 622538
rect 23746 622468 23766 622538
rect 23836 622468 23856 622538
rect 23926 622468 23946 622538
rect 21946 622448 23946 622468
rect 21946 622378 21966 622448
rect 22036 622378 22056 622448
rect 22126 622378 22146 622448
rect 22216 622378 22236 622448
rect 22306 622378 22326 622448
rect 22396 622378 22416 622448
rect 22486 622378 22506 622448
rect 22576 622378 22596 622448
rect 22666 622378 22686 622448
rect 22756 622378 22776 622448
rect 22846 622378 22866 622448
rect 22936 622378 22956 622448
rect 23026 622378 23046 622448
rect 23116 622378 23136 622448
rect 23206 622378 23226 622448
rect 23296 622378 23316 622448
rect 23386 622378 23406 622448
rect 23476 622378 23496 622448
rect 23566 622378 23586 622448
rect 23656 622378 23676 622448
rect 23746 622378 23766 622448
rect 23836 622378 23856 622448
rect 23926 622378 23946 622448
rect 21946 622358 23946 622378
rect 21946 622288 21966 622358
rect 22036 622288 22056 622358
rect 22126 622288 22146 622358
rect 22216 622288 22236 622358
rect 22306 622288 22326 622358
rect 22396 622288 22416 622358
rect 22486 622288 22506 622358
rect 22576 622288 22596 622358
rect 22666 622288 22686 622358
rect 22756 622288 22776 622358
rect 22846 622288 22866 622358
rect 22936 622288 22956 622358
rect 23026 622288 23046 622358
rect 23116 622288 23136 622358
rect 23206 622288 23226 622358
rect 23296 622288 23316 622358
rect 23386 622288 23406 622358
rect 23476 622288 23496 622358
rect 23566 622288 23586 622358
rect 23656 622288 23676 622358
rect 23746 622288 23766 622358
rect 23836 622288 23856 622358
rect 23926 622288 23946 622358
rect 21946 622268 23946 622288
rect 21946 622198 21966 622268
rect 22036 622198 22056 622268
rect 22126 622198 22146 622268
rect 22216 622198 22236 622268
rect 22306 622198 22326 622268
rect 22396 622198 22416 622268
rect 22486 622198 22506 622268
rect 22576 622198 22596 622268
rect 22666 622198 22686 622268
rect 22756 622198 22776 622268
rect 22846 622198 22866 622268
rect 22936 622198 22956 622268
rect 23026 622198 23046 622268
rect 23116 622198 23136 622268
rect 23206 622198 23226 622268
rect 23296 622198 23316 622268
rect 23386 622198 23406 622268
rect 23476 622198 23496 622268
rect 23566 622198 23586 622268
rect 23656 622198 23676 622268
rect 23746 622198 23766 622268
rect 23836 622198 23856 622268
rect 23926 622198 23946 622268
rect 21946 622178 23946 622198
rect 21946 622108 21966 622178
rect 22036 622108 22056 622178
rect 22126 622108 22146 622178
rect 22216 622108 22236 622178
rect 22306 622108 22326 622178
rect 22396 622108 22416 622178
rect 22486 622108 22506 622178
rect 22576 622108 22596 622178
rect 22666 622108 22686 622178
rect 22756 622108 22776 622178
rect 22846 622108 22866 622178
rect 22936 622108 22956 622178
rect 23026 622108 23046 622178
rect 23116 622108 23136 622178
rect 23206 622108 23226 622178
rect 23296 622108 23316 622178
rect 23386 622108 23406 622178
rect 23476 622108 23496 622178
rect 23566 622108 23586 622178
rect 23656 622108 23676 622178
rect 23746 622108 23766 622178
rect 23836 622108 23856 622178
rect 23926 622108 23946 622178
rect 21946 622088 23946 622108
rect 21946 622018 21966 622088
rect 22036 622018 22056 622088
rect 22126 622018 22146 622088
rect 22216 622018 22236 622088
rect 22306 622018 22326 622088
rect 22396 622018 22416 622088
rect 22486 622018 22506 622088
rect 22576 622018 22596 622088
rect 22666 622018 22686 622088
rect 22756 622018 22776 622088
rect 22846 622018 22866 622088
rect 22936 622018 22956 622088
rect 23026 622018 23046 622088
rect 23116 622018 23136 622088
rect 23206 622018 23226 622088
rect 23296 622018 23316 622088
rect 23386 622018 23406 622088
rect 23476 622018 23496 622088
rect 23566 622018 23586 622088
rect 23656 622018 23676 622088
rect 23746 622018 23766 622088
rect 23836 622018 23856 622088
rect 23926 622018 23946 622088
rect 21946 621998 23946 622018
rect 21946 621928 21966 621998
rect 22036 621928 22056 621998
rect 22126 621928 22146 621998
rect 22216 621928 22236 621998
rect 22306 621928 22326 621998
rect 22396 621928 22416 621998
rect 22486 621928 22506 621998
rect 22576 621928 22596 621998
rect 22666 621928 22686 621998
rect 22756 621928 22776 621998
rect 22846 621928 22866 621998
rect 22936 621928 22956 621998
rect 23026 621928 23046 621998
rect 23116 621928 23136 621998
rect 23206 621928 23226 621998
rect 23296 621928 23316 621998
rect 23386 621928 23406 621998
rect 23476 621928 23496 621998
rect 23566 621928 23586 621998
rect 23656 621928 23676 621998
rect 23746 621928 23766 621998
rect 23836 621928 23856 621998
rect 23926 621928 23946 621998
rect 21946 621908 23946 621928
rect 21946 621838 21966 621908
rect 22036 621838 22056 621908
rect 22126 621838 22146 621908
rect 22216 621838 22236 621908
rect 22306 621838 22326 621908
rect 22396 621838 22416 621908
rect 22486 621838 22506 621908
rect 22576 621838 22596 621908
rect 22666 621838 22686 621908
rect 22756 621838 22776 621908
rect 22846 621838 22866 621908
rect 22936 621838 22956 621908
rect 23026 621838 23046 621908
rect 23116 621838 23136 621908
rect 23206 621838 23226 621908
rect 23296 621838 23316 621908
rect 23386 621838 23406 621908
rect 23476 621838 23496 621908
rect 23566 621838 23586 621908
rect 23656 621838 23676 621908
rect 23746 621838 23766 621908
rect 23836 621838 23856 621908
rect 23926 621838 23946 621908
rect 21946 621818 23946 621838
rect 21946 621748 21966 621818
rect 22036 621748 22056 621818
rect 22126 621748 22146 621818
rect 22216 621748 22236 621818
rect 22306 621748 22326 621818
rect 22396 621748 22416 621818
rect 22486 621748 22506 621818
rect 22576 621748 22596 621818
rect 22666 621748 22686 621818
rect 22756 621748 22776 621818
rect 22846 621748 22866 621818
rect 22936 621748 22956 621818
rect 23026 621748 23046 621818
rect 23116 621748 23136 621818
rect 23206 621748 23226 621818
rect 23296 621748 23316 621818
rect 23386 621748 23406 621818
rect 23476 621748 23496 621818
rect 23566 621748 23586 621818
rect 23656 621748 23676 621818
rect 23746 621748 23766 621818
rect 23836 621748 23856 621818
rect 23926 621748 23946 621818
rect 21946 621728 23946 621748
rect 21946 621658 21966 621728
rect 22036 621658 22056 621728
rect 22126 621658 22146 621728
rect 22216 621658 22236 621728
rect 22306 621658 22326 621728
rect 22396 621658 22416 621728
rect 22486 621658 22506 621728
rect 22576 621658 22596 621728
rect 22666 621658 22686 621728
rect 22756 621658 22776 621728
rect 22846 621658 22866 621728
rect 22936 621658 22956 621728
rect 23026 621658 23046 621728
rect 23116 621658 23136 621728
rect 23206 621658 23226 621728
rect 23296 621658 23316 621728
rect 23386 621658 23406 621728
rect 23476 621658 23496 621728
rect 23566 621658 23586 621728
rect 23656 621658 23676 621728
rect 23746 621658 23766 621728
rect 23836 621658 23856 621728
rect 23926 621658 23946 621728
rect 21946 621638 23946 621658
rect 21946 621568 21966 621638
rect 22036 621568 22056 621638
rect 22126 621568 22146 621638
rect 22216 621568 22236 621638
rect 22306 621568 22326 621638
rect 22396 621568 22416 621638
rect 22486 621568 22506 621638
rect 22576 621568 22596 621638
rect 22666 621568 22686 621638
rect 22756 621568 22776 621638
rect 22846 621568 22866 621638
rect 22936 621568 22956 621638
rect 23026 621568 23046 621638
rect 23116 621568 23136 621638
rect 23206 621568 23226 621638
rect 23296 621568 23316 621638
rect 23386 621568 23406 621638
rect 23476 621568 23496 621638
rect 23566 621568 23586 621638
rect 23656 621568 23676 621638
rect 23746 621568 23766 621638
rect 23836 621568 23856 621638
rect 23926 621568 23946 621638
rect 21946 621548 23946 621568
rect 17650 619350 17670 619420
rect 17740 619350 17760 619420
rect 17830 619350 17850 619420
rect 17920 619350 17940 619420
rect 18010 619350 18030 619420
rect 18100 619350 18120 619420
rect 18190 619350 18210 619420
rect 18280 619350 18300 619420
rect 18370 619350 18390 619420
rect 18460 619350 18480 619420
rect 18550 619350 18570 619420
rect 18640 619350 18660 619420
rect 18730 619350 18750 619420
rect 18820 619350 18840 619420
rect 18910 619350 18930 619420
rect 19000 619350 19020 619420
rect 19090 619350 19110 619420
rect 19180 619350 19200 619420
rect 19270 619350 19290 619420
rect 19360 619350 19380 619420
rect 19450 619350 19470 619420
rect 19540 619350 19560 619420
rect 19630 619350 19650 619420
rect 17650 619330 19650 619350
rect 17650 619260 17670 619330
rect 17740 619260 17760 619330
rect 17830 619260 17850 619330
rect 17920 619260 17940 619330
rect 18010 619260 18030 619330
rect 18100 619260 18120 619330
rect 18190 619260 18210 619330
rect 18280 619260 18300 619330
rect 18370 619260 18390 619330
rect 18460 619260 18480 619330
rect 18550 619260 18570 619330
rect 18640 619260 18660 619330
rect 18730 619260 18750 619330
rect 18820 619260 18840 619330
rect 18910 619260 18930 619330
rect 19000 619260 19020 619330
rect 19090 619260 19110 619330
rect 19180 619260 19200 619330
rect 19270 619260 19290 619330
rect 19360 619260 19380 619330
rect 19450 619260 19470 619330
rect 19540 619260 19560 619330
rect 19630 619260 19650 619330
rect 17650 619240 19650 619260
rect 17650 619170 17670 619240
rect 17740 619170 17760 619240
rect 17830 619170 17850 619240
rect 17920 619170 17940 619240
rect 18010 619170 18030 619240
rect 18100 619170 18120 619240
rect 18190 619170 18210 619240
rect 18280 619170 18300 619240
rect 18370 619170 18390 619240
rect 18460 619170 18480 619240
rect 18550 619170 18570 619240
rect 18640 619170 18660 619240
rect 18730 619170 18750 619240
rect 18820 619170 18840 619240
rect 18910 619170 18930 619240
rect 19000 619170 19020 619240
rect 19090 619170 19110 619240
rect 19180 619170 19200 619240
rect 19270 619170 19290 619240
rect 19360 619170 19380 619240
rect 19450 619170 19470 619240
rect 19540 619170 19560 619240
rect 19630 619170 19650 619240
rect 17650 619150 19650 619170
rect 17650 619080 17670 619150
rect 17740 619080 17760 619150
rect 17830 619080 17850 619150
rect 17920 619080 17940 619150
rect 18010 619080 18030 619150
rect 18100 619080 18120 619150
rect 18190 619080 18210 619150
rect 18280 619080 18300 619150
rect 18370 619080 18390 619150
rect 18460 619080 18480 619150
rect 18550 619080 18570 619150
rect 18640 619080 18660 619150
rect 18730 619080 18750 619150
rect 18820 619080 18840 619150
rect 18910 619080 18930 619150
rect 19000 619080 19020 619150
rect 19090 619080 19110 619150
rect 19180 619080 19200 619150
rect 19270 619080 19290 619150
rect 19360 619080 19380 619150
rect 19450 619080 19470 619150
rect 19540 619080 19560 619150
rect 19630 619080 19650 619150
rect 17650 619060 19650 619080
rect 17650 618990 17670 619060
rect 17740 618990 17760 619060
rect 17830 618990 17850 619060
rect 17920 618990 17940 619060
rect 18010 618990 18030 619060
rect 18100 618990 18120 619060
rect 18190 618990 18210 619060
rect 18280 618990 18300 619060
rect 18370 618990 18390 619060
rect 18460 618990 18480 619060
rect 18550 618990 18570 619060
rect 18640 618990 18660 619060
rect 18730 618990 18750 619060
rect 18820 618990 18840 619060
rect 18910 618990 18930 619060
rect 19000 618990 19020 619060
rect 19090 618990 19110 619060
rect 19180 618990 19200 619060
rect 19270 618990 19290 619060
rect 19360 618990 19380 619060
rect 19450 618990 19470 619060
rect 19540 618990 19560 619060
rect 19630 618990 19650 619060
rect 17650 618970 19650 618990
rect 17650 618900 17670 618970
rect 17740 618900 17760 618970
rect 17830 618900 17850 618970
rect 17920 618900 17940 618970
rect 18010 618900 18030 618970
rect 18100 618900 18120 618970
rect 18190 618900 18210 618970
rect 18280 618900 18300 618970
rect 18370 618900 18390 618970
rect 18460 618900 18480 618970
rect 18550 618900 18570 618970
rect 18640 618900 18660 618970
rect 18730 618900 18750 618970
rect 18820 618900 18840 618970
rect 18910 618900 18930 618970
rect 19000 618900 19020 618970
rect 19090 618900 19110 618970
rect 19180 618900 19200 618970
rect 19270 618900 19290 618970
rect 19360 618900 19380 618970
rect 19450 618900 19470 618970
rect 19540 618900 19560 618970
rect 19630 618900 19650 618970
rect 17650 618880 19650 618900
rect 17650 618810 17670 618880
rect 17740 618810 17760 618880
rect 17830 618810 17850 618880
rect 17920 618810 17940 618880
rect 18010 618810 18030 618880
rect 18100 618810 18120 618880
rect 18190 618810 18210 618880
rect 18280 618810 18300 618880
rect 18370 618810 18390 618880
rect 18460 618810 18480 618880
rect 18550 618810 18570 618880
rect 18640 618810 18660 618880
rect 18730 618810 18750 618880
rect 18820 618810 18840 618880
rect 18910 618810 18930 618880
rect 19000 618810 19020 618880
rect 19090 618810 19110 618880
rect 19180 618810 19200 618880
rect 19270 618810 19290 618880
rect 19360 618810 19380 618880
rect 19450 618810 19470 618880
rect 19540 618810 19560 618880
rect 19630 618810 19650 618880
rect 17650 618790 19650 618810
rect 17650 618720 17670 618790
rect 17740 618720 17760 618790
rect 17830 618720 17850 618790
rect 17920 618720 17940 618790
rect 18010 618720 18030 618790
rect 18100 618720 18120 618790
rect 18190 618720 18210 618790
rect 18280 618720 18300 618790
rect 18370 618720 18390 618790
rect 18460 618720 18480 618790
rect 18550 618720 18570 618790
rect 18640 618720 18660 618790
rect 18730 618720 18750 618790
rect 18820 618720 18840 618790
rect 18910 618720 18930 618790
rect 19000 618720 19020 618790
rect 19090 618720 19110 618790
rect 19180 618720 19200 618790
rect 19270 618720 19290 618790
rect 19360 618720 19380 618790
rect 19450 618720 19470 618790
rect 19540 618720 19560 618790
rect 19630 618720 19650 618790
rect 17650 618700 19650 618720
rect 17650 618630 17670 618700
rect 17740 618630 17760 618700
rect 17830 618630 17850 618700
rect 17920 618630 17940 618700
rect 18010 618630 18030 618700
rect 18100 618630 18120 618700
rect 18190 618630 18210 618700
rect 18280 618630 18300 618700
rect 18370 618630 18390 618700
rect 18460 618630 18480 618700
rect 18550 618630 18570 618700
rect 18640 618630 18660 618700
rect 18730 618630 18750 618700
rect 18820 618630 18840 618700
rect 18910 618630 18930 618700
rect 19000 618630 19020 618700
rect 19090 618630 19110 618700
rect 19180 618630 19200 618700
rect 19270 618630 19290 618700
rect 19360 618630 19380 618700
rect 19450 618630 19470 618700
rect 19540 618630 19560 618700
rect 19630 618630 19650 618700
rect 17650 618610 19650 618630
rect 17650 618540 17670 618610
rect 17740 618540 17760 618610
rect 17830 618540 17850 618610
rect 17920 618540 17940 618610
rect 18010 618540 18030 618610
rect 18100 618540 18120 618610
rect 18190 618540 18210 618610
rect 18280 618540 18300 618610
rect 18370 618540 18390 618610
rect 18460 618540 18480 618610
rect 18550 618540 18570 618610
rect 18640 618540 18660 618610
rect 18730 618540 18750 618610
rect 18820 618540 18840 618610
rect 18910 618540 18930 618610
rect 19000 618540 19020 618610
rect 19090 618540 19110 618610
rect 19180 618540 19200 618610
rect 19270 618540 19290 618610
rect 19360 618540 19380 618610
rect 19450 618540 19470 618610
rect 19540 618540 19560 618610
rect 19630 618540 19650 618610
rect 17650 618520 19650 618540
rect 17650 618450 17670 618520
rect 17740 618450 17760 618520
rect 17830 618450 17850 618520
rect 17920 618450 17940 618520
rect 18010 618450 18030 618520
rect 18100 618450 18120 618520
rect 18190 618450 18210 618520
rect 18280 618450 18300 618520
rect 18370 618450 18390 618520
rect 18460 618450 18480 618520
rect 18550 618450 18570 618520
rect 18640 618450 18660 618520
rect 18730 618450 18750 618520
rect 18820 618450 18840 618520
rect 18910 618450 18930 618520
rect 19000 618450 19020 618520
rect 19090 618450 19110 618520
rect 19180 618450 19200 618520
rect 19270 618450 19290 618520
rect 19360 618450 19380 618520
rect 19450 618450 19470 618520
rect 19540 618450 19560 618520
rect 19630 618450 19650 618520
rect 17650 618430 19650 618450
rect 17650 618360 17670 618430
rect 17740 618360 17760 618430
rect 17830 618360 17850 618430
rect 17920 618360 17940 618430
rect 18010 618360 18030 618430
rect 18100 618360 18120 618430
rect 18190 618360 18210 618430
rect 18280 618360 18300 618430
rect 18370 618360 18390 618430
rect 18460 618360 18480 618430
rect 18550 618360 18570 618430
rect 18640 618360 18660 618430
rect 18730 618360 18750 618430
rect 18820 618360 18840 618430
rect 18910 618360 18930 618430
rect 19000 618360 19020 618430
rect 19090 618360 19110 618430
rect 19180 618360 19200 618430
rect 19270 618360 19290 618430
rect 19360 618360 19380 618430
rect 19450 618360 19470 618430
rect 19540 618360 19560 618430
rect 19630 618360 19650 618430
rect 17650 618340 19650 618360
rect 17650 618270 17670 618340
rect 17740 618270 17760 618340
rect 17830 618270 17850 618340
rect 17920 618270 17940 618340
rect 18010 618270 18030 618340
rect 18100 618270 18120 618340
rect 18190 618270 18210 618340
rect 18280 618270 18300 618340
rect 18370 618270 18390 618340
rect 18460 618270 18480 618340
rect 18550 618270 18570 618340
rect 18640 618270 18660 618340
rect 18730 618270 18750 618340
rect 18820 618270 18840 618340
rect 18910 618270 18930 618340
rect 19000 618270 19020 618340
rect 19090 618270 19110 618340
rect 19180 618270 19200 618340
rect 19270 618270 19290 618340
rect 19360 618270 19380 618340
rect 19450 618270 19470 618340
rect 19540 618270 19560 618340
rect 19630 618270 19650 618340
rect 17650 618250 19650 618270
rect 17650 618180 17670 618250
rect 17740 618180 17760 618250
rect 17830 618180 17850 618250
rect 17920 618180 17940 618250
rect 18010 618180 18030 618250
rect 18100 618180 18120 618250
rect 18190 618180 18210 618250
rect 18280 618180 18300 618250
rect 18370 618180 18390 618250
rect 18460 618180 18480 618250
rect 18550 618180 18570 618250
rect 18640 618180 18660 618250
rect 18730 618180 18750 618250
rect 18820 618180 18840 618250
rect 18910 618180 18930 618250
rect 19000 618180 19020 618250
rect 19090 618180 19110 618250
rect 19180 618180 19200 618250
rect 19270 618180 19290 618250
rect 19360 618180 19380 618250
rect 19450 618180 19470 618250
rect 19540 618180 19560 618250
rect 19630 618180 19650 618250
rect 17650 618160 19650 618180
rect 17650 618090 17670 618160
rect 17740 618090 17760 618160
rect 17830 618090 17850 618160
rect 17920 618090 17940 618160
rect 18010 618090 18030 618160
rect 18100 618090 18120 618160
rect 18190 618090 18210 618160
rect 18280 618090 18300 618160
rect 18370 618090 18390 618160
rect 18460 618090 18480 618160
rect 18550 618090 18570 618160
rect 18640 618090 18660 618160
rect 18730 618090 18750 618160
rect 18820 618090 18840 618160
rect 18910 618090 18930 618160
rect 19000 618090 19020 618160
rect 19090 618090 19110 618160
rect 19180 618090 19200 618160
rect 19270 618090 19290 618160
rect 19360 618090 19380 618160
rect 19450 618090 19470 618160
rect 19540 618090 19560 618160
rect 19630 618090 19650 618160
rect 17650 618070 19650 618090
rect 17650 618000 17670 618070
rect 17740 618000 17760 618070
rect 17830 618000 17850 618070
rect 17920 618000 17940 618070
rect 18010 618000 18030 618070
rect 18100 618000 18120 618070
rect 18190 618000 18210 618070
rect 18280 618000 18300 618070
rect 18370 618000 18390 618070
rect 18460 618000 18480 618070
rect 18550 618000 18570 618070
rect 18640 618000 18660 618070
rect 18730 618000 18750 618070
rect 18820 618000 18840 618070
rect 18910 618000 18930 618070
rect 19000 618000 19020 618070
rect 19090 618000 19110 618070
rect 19180 618000 19200 618070
rect 19270 618000 19290 618070
rect 19360 618000 19380 618070
rect 19450 618000 19470 618070
rect 19540 618000 19560 618070
rect 19630 618000 19650 618070
rect 17650 617980 19650 618000
rect 17650 617910 17670 617980
rect 17740 617910 17760 617980
rect 17830 617910 17850 617980
rect 17920 617910 17940 617980
rect 18010 617910 18030 617980
rect 18100 617910 18120 617980
rect 18190 617910 18210 617980
rect 18280 617910 18300 617980
rect 18370 617910 18390 617980
rect 18460 617910 18480 617980
rect 18550 617910 18570 617980
rect 18640 617910 18660 617980
rect 18730 617910 18750 617980
rect 18820 617910 18840 617980
rect 18910 617910 18930 617980
rect 19000 617910 19020 617980
rect 19090 617910 19110 617980
rect 19180 617910 19200 617980
rect 19270 617910 19290 617980
rect 19360 617910 19380 617980
rect 19450 617910 19470 617980
rect 19540 617910 19560 617980
rect 19630 617910 19650 617980
rect 17650 617890 19650 617910
rect 17650 617820 17670 617890
rect 17740 617820 17760 617890
rect 17830 617820 17850 617890
rect 17920 617820 17940 617890
rect 18010 617820 18030 617890
rect 18100 617820 18120 617890
rect 18190 617820 18210 617890
rect 18280 617820 18300 617890
rect 18370 617820 18390 617890
rect 18460 617820 18480 617890
rect 18550 617820 18570 617890
rect 18640 617820 18660 617890
rect 18730 617820 18750 617890
rect 18820 617820 18840 617890
rect 18910 617820 18930 617890
rect 19000 617820 19020 617890
rect 19090 617820 19110 617890
rect 19180 617820 19200 617890
rect 19270 617820 19290 617890
rect 19360 617820 19380 617890
rect 19450 617820 19470 617890
rect 19540 617820 19560 617890
rect 19630 617820 19650 617890
rect 17650 617800 19650 617820
rect 17650 617730 17670 617800
rect 17740 617730 17760 617800
rect 17830 617730 17850 617800
rect 17920 617730 17940 617800
rect 18010 617730 18030 617800
rect 18100 617730 18120 617800
rect 18190 617730 18210 617800
rect 18280 617730 18300 617800
rect 18370 617730 18390 617800
rect 18460 617730 18480 617800
rect 18550 617730 18570 617800
rect 18640 617730 18660 617800
rect 18730 617730 18750 617800
rect 18820 617730 18840 617800
rect 18910 617730 18930 617800
rect 19000 617730 19020 617800
rect 19090 617730 19110 617800
rect 19180 617730 19200 617800
rect 19270 617730 19290 617800
rect 19360 617730 19380 617800
rect 19450 617730 19470 617800
rect 19540 617730 19560 617800
rect 19630 617730 19650 617800
rect 17650 617710 19650 617730
rect 17650 617640 17670 617710
rect 17740 617640 17760 617710
rect 17830 617640 17850 617710
rect 17920 617640 17940 617710
rect 18010 617640 18030 617710
rect 18100 617640 18120 617710
rect 18190 617640 18210 617710
rect 18280 617640 18300 617710
rect 18370 617640 18390 617710
rect 18460 617640 18480 617710
rect 18550 617640 18570 617710
rect 18640 617640 18660 617710
rect 18730 617640 18750 617710
rect 18820 617640 18840 617710
rect 18910 617640 18930 617710
rect 19000 617640 19020 617710
rect 19090 617640 19110 617710
rect 19180 617640 19200 617710
rect 19270 617640 19290 617710
rect 19360 617640 19380 617710
rect 19450 617640 19470 617710
rect 19540 617640 19560 617710
rect 19630 617640 19650 617710
rect 17650 617620 19650 617640
rect 17650 617550 17670 617620
rect 17740 617550 17760 617620
rect 17830 617550 17850 617620
rect 17920 617550 17940 617620
rect 18010 617550 18030 617620
rect 18100 617550 18120 617620
rect 18190 617550 18210 617620
rect 18280 617550 18300 617620
rect 18370 617550 18390 617620
rect 18460 617550 18480 617620
rect 18550 617550 18570 617620
rect 18640 617550 18660 617620
rect 18730 617550 18750 617620
rect 18820 617550 18840 617620
rect 18910 617550 18930 617620
rect 19000 617550 19020 617620
rect 19090 617550 19110 617620
rect 19180 617550 19200 617620
rect 19270 617550 19290 617620
rect 19360 617550 19380 617620
rect 19450 617550 19470 617620
rect 19540 617550 19560 617620
rect 19630 617550 19650 617620
rect 17650 617530 19650 617550
rect 17650 617460 17670 617530
rect 17740 617460 17760 617530
rect 17830 617460 17850 617530
rect 17920 617460 17940 617530
rect 18010 617460 18030 617530
rect 18100 617460 18120 617530
rect 18190 617460 18210 617530
rect 18280 617460 18300 617530
rect 18370 617460 18390 617530
rect 18460 617460 18480 617530
rect 18550 617460 18570 617530
rect 18640 617460 18660 617530
rect 18730 617460 18750 617530
rect 18820 617460 18840 617530
rect 18910 617460 18930 617530
rect 19000 617460 19020 617530
rect 19090 617460 19110 617530
rect 19180 617460 19200 617530
rect 19270 617460 19290 617530
rect 19360 617460 19380 617530
rect 19450 617460 19470 617530
rect 19540 617460 19560 617530
rect 19630 617460 19650 617530
rect 17650 617440 19650 617460
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 18070 703760 18140 703830
rect 18160 703760 18230 703830
rect 18250 703760 18320 703830
rect 18340 703760 18410 703830
rect 18430 703760 18500 703830
rect 18520 703760 18590 703830
rect 18610 703760 18680 703830
rect 18700 703760 18770 703830
rect 18790 703760 18860 703830
rect 18880 703760 18950 703830
rect 18970 703760 19040 703830
rect 19060 703760 19130 703830
rect 19150 703760 19220 703830
rect 19240 703760 19310 703830
rect 19330 703760 19400 703830
rect 19420 703760 19490 703830
rect 19510 703760 19580 703830
rect 18070 703670 18140 703740
rect 18160 703670 18230 703740
rect 18250 703670 18320 703740
rect 18340 703670 18410 703740
rect 18430 703670 18500 703740
rect 18520 703670 18590 703740
rect 18610 703670 18680 703740
rect 18700 703670 18770 703740
rect 18790 703670 18860 703740
rect 18880 703670 18950 703740
rect 18970 703670 19040 703740
rect 19060 703670 19130 703740
rect 19150 703670 19220 703740
rect 19240 703670 19310 703740
rect 19330 703670 19400 703740
rect 19420 703670 19490 703740
rect 19510 703670 19580 703740
rect 18070 703580 18140 703650
rect 18160 703580 18230 703650
rect 18250 703580 18320 703650
rect 18340 703580 18410 703650
rect 18430 703580 18500 703650
rect 18520 703580 18590 703650
rect 18610 703580 18680 703650
rect 18700 703580 18770 703650
rect 18790 703580 18860 703650
rect 18880 703580 18950 703650
rect 18970 703580 19040 703650
rect 19060 703580 19130 703650
rect 19150 703580 19220 703650
rect 19240 703580 19310 703650
rect 19330 703580 19400 703650
rect 19420 703580 19490 703650
rect 19510 703580 19580 703650
rect 18070 703490 18140 703560
rect 18160 703490 18230 703560
rect 18250 703490 18320 703560
rect 18340 703490 18410 703560
rect 18430 703490 18500 703560
rect 18520 703490 18590 703560
rect 18610 703490 18680 703560
rect 18700 703490 18770 703560
rect 18790 703490 18860 703560
rect 18880 703490 18950 703560
rect 18970 703490 19040 703560
rect 19060 703490 19130 703560
rect 19150 703490 19220 703560
rect 19240 703490 19310 703560
rect 19330 703490 19400 703560
rect 19420 703490 19490 703560
rect 19510 703490 19580 703560
rect 18070 703400 18140 703470
rect 18160 703400 18230 703470
rect 18250 703400 18320 703470
rect 18340 703400 18410 703470
rect 18430 703400 18500 703470
rect 18520 703400 18590 703470
rect 18610 703400 18680 703470
rect 18700 703400 18770 703470
rect 18790 703400 18860 703470
rect 18880 703400 18950 703470
rect 18970 703400 19040 703470
rect 19060 703400 19130 703470
rect 19150 703400 19220 703470
rect 19240 703400 19310 703470
rect 19330 703400 19400 703470
rect 19420 703400 19490 703470
rect 19510 703400 19580 703470
rect 18070 703310 18140 703380
rect 18160 703310 18230 703380
rect 18250 703310 18320 703380
rect 18340 703310 18410 703380
rect 18430 703310 18500 703380
rect 18520 703310 18590 703380
rect 18610 703310 18680 703380
rect 18700 703310 18770 703380
rect 18790 703310 18860 703380
rect 18880 703310 18950 703380
rect 18970 703310 19040 703380
rect 19060 703310 19130 703380
rect 19150 703310 19220 703380
rect 19240 703310 19310 703380
rect 19330 703310 19400 703380
rect 19420 703310 19490 703380
rect 19510 703310 19580 703380
rect 18070 703220 18140 703290
rect 18160 703220 18230 703290
rect 18250 703220 18320 703290
rect 18340 703220 18410 703290
rect 18430 703220 18500 703290
rect 18520 703220 18590 703290
rect 18610 703220 18680 703290
rect 18700 703220 18770 703290
rect 18790 703220 18860 703290
rect 18880 703220 18950 703290
rect 18970 703220 19040 703290
rect 19060 703220 19130 703290
rect 19150 703220 19220 703290
rect 19240 703220 19310 703290
rect 19330 703220 19400 703290
rect 19420 703220 19490 703290
rect 19510 703220 19580 703290
rect 18070 703130 18140 703200
rect 18160 703130 18230 703200
rect 18250 703130 18320 703200
rect 18340 703130 18410 703200
rect 18430 703130 18500 703200
rect 18520 703130 18590 703200
rect 18610 703130 18680 703200
rect 18700 703130 18770 703200
rect 18790 703130 18860 703200
rect 18880 703130 18950 703200
rect 18970 703130 19040 703200
rect 19060 703130 19130 703200
rect 19150 703130 19220 703200
rect 19240 703130 19310 703200
rect 19330 703130 19400 703200
rect 19420 703130 19490 703200
rect 19510 703130 19580 703200
rect 18070 703040 18140 703110
rect 18160 703040 18230 703110
rect 18250 703040 18320 703110
rect 18340 703040 18410 703110
rect 18430 703040 18500 703110
rect 18520 703040 18590 703110
rect 18610 703040 18680 703110
rect 18700 703040 18770 703110
rect 18790 703040 18860 703110
rect 18880 703040 18950 703110
rect 18970 703040 19040 703110
rect 19060 703040 19130 703110
rect 19150 703040 19220 703110
rect 19240 703040 19310 703110
rect 19330 703040 19400 703110
rect 19420 703040 19490 703110
rect 19510 703040 19580 703110
rect 18070 702950 18140 703020
rect 18160 702950 18230 703020
rect 18250 702950 18320 703020
rect 18340 702950 18410 703020
rect 18430 702950 18500 703020
rect 18520 702950 18590 703020
rect 18610 702950 18680 703020
rect 18700 702950 18770 703020
rect 18790 702950 18860 703020
rect 18880 702950 18950 703020
rect 18970 702950 19040 703020
rect 19060 702950 19130 703020
rect 19150 702950 19220 703020
rect 19240 702950 19310 703020
rect 19330 702950 19400 703020
rect 19420 702950 19490 703020
rect 19510 702950 19580 703020
rect 18070 702860 18140 702930
rect 18160 702860 18230 702930
rect 18250 702860 18320 702930
rect 18340 702860 18410 702930
rect 18430 702860 18500 702930
rect 18520 702860 18590 702930
rect 18610 702860 18680 702930
rect 18700 702860 18770 702930
rect 18790 702860 18860 702930
rect 18880 702860 18950 702930
rect 18970 702860 19040 702930
rect 19060 702860 19130 702930
rect 19150 702860 19220 702930
rect 19240 702860 19310 702930
rect 19330 702860 19400 702930
rect 19420 702860 19490 702930
rect 19510 702860 19580 702930
rect 18070 702770 18140 702840
rect 18160 702770 18230 702840
rect 18250 702770 18320 702840
rect 18340 702770 18410 702840
rect 18430 702770 18500 702840
rect 18520 702770 18590 702840
rect 18610 702770 18680 702840
rect 18700 702770 18770 702840
rect 18790 702770 18860 702840
rect 18880 702770 18950 702840
rect 18970 702770 19040 702840
rect 19060 702770 19130 702840
rect 19150 702770 19220 702840
rect 19240 702770 19310 702840
rect 19330 702770 19400 702840
rect 19420 702770 19490 702840
rect 19510 702770 19580 702840
rect 18070 702680 18140 702750
rect 18160 702680 18230 702750
rect 18250 702680 18320 702750
rect 18340 702680 18410 702750
rect 18430 702680 18500 702750
rect 18520 702680 18590 702750
rect 18610 702680 18680 702750
rect 18700 702680 18770 702750
rect 18790 702680 18860 702750
rect 18880 702680 18950 702750
rect 18970 702680 19040 702750
rect 19060 702680 19130 702750
rect 19150 702680 19220 702750
rect 19240 702680 19310 702750
rect 19330 702680 19400 702750
rect 19420 702680 19490 702750
rect 19510 702680 19580 702750
rect 18070 702590 18140 702660
rect 18160 702590 18230 702660
rect 18250 702590 18320 702660
rect 18340 702590 18410 702660
rect 18430 702590 18500 702660
rect 18520 702590 18590 702660
rect 18610 702590 18680 702660
rect 18700 702590 18770 702660
rect 18790 702590 18860 702660
rect 18880 702590 18950 702660
rect 18970 702590 19040 702660
rect 19060 702590 19130 702660
rect 19150 702590 19220 702660
rect 19240 702590 19310 702660
rect 19330 702590 19400 702660
rect 19420 702590 19490 702660
rect 19510 702590 19580 702660
rect 18070 702500 18140 702570
rect 18160 702500 18230 702570
rect 18250 702500 18320 702570
rect 18340 702500 18410 702570
rect 18430 702500 18500 702570
rect 18520 702500 18590 702570
rect 18610 702500 18680 702570
rect 18700 702500 18770 702570
rect 18790 702500 18860 702570
rect 18880 702500 18950 702570
rect 18970 702500 19040 702570
rect 19060 702500 19130 702570
rect 19150 702500 19220 702570
rect 19240 702500 19310 702570
rect 19330 702500 19400 702570
rect 19420 702500 19490 702570
rect 19510 702500 19580 702570
rect 18070 702410 18140 702480
rect 18160 702410 18230 702480
rect 18250 702410 18320 702480
rect 18340 702410 18410 702480
rect 18430 702410 18500 702480
rect 18520 702410 18590 702480
rect 18610 702410 18680 702480
rect 18700 702410 18770 702480
rect 18790 702410 18860 702480
rect 18880 702410 18950 702480
rect 18970 702410 19040 702480
rect 19060 702410 19130 702480
rect 19150 702410 19220 702480
rect 19240 702410 19310 702480
rect 19330 702410 19400 702480
rect 19420 702410 19490 702480
rect 19510 702410 19580 702480
rect 18070 702320 18140 702390
rect 18160 702320 18230 702390
rect 18250 702320 18320 702390
rect 18340 702320 18410 702390
rect 18430 702320 18500 702390
rect 18520 702320 18590 702390
rect 18610 702320 18680 702390
rect 18700 702320 18770 702390
rect 18790 702320 18860 702390
rect 18880 702320 18950 702390
rect 18970 702320 19040 702390
rect 19060 702320 19130 702390
rect 19150 702320 19220 702390
rect 19240 702320 19310 702390
rect 19330 702320 19400 702390
rect 19420 702320 19490 702390
rect 19510 702320 19580 702390
rect 70090 703760 70160 703830
rect 70180 703760 70250 703830
rect 70270 703760 70340 703830
rect 70360 703760 70430 703830
rect 70450 703760 70520 703830
rect 70540 703760 70610 703830
rect 70630 703760 70700 703830
rect 70720 703760 70790 703830
rect 70810 703760 70880 703830
rect 70900 703760 70970 703830
rect 70990 703760 71060 703830
rect 71080 703760 71150 703830
rect 71170 703760 71240 703830
rect 71260 703760 71330 703830
rect 71350 703760 71420 703830
rect 71440 703760 71510 703830
rect 71530 703760 71600 703830
rect 70090 703670 70160 703740
rect 70180 703670 70250 703740
rect 70270 703670 70340 703740
rect 70360 703670 70430 703740
rect 70450 703670 70520 703740
rect 70540 703670 70610 703740
rect 70630 703670 70700 703740
rect 70720 703670 70790 703740
rect 70810 703670 70880 703740
rect 70900 703670 70970 703740
rect 70990 703670 71060 703740
rect 71080 703670 71150 703740
rect 71170 703670 71240 703740
rect 71260 703670 71330 703740
rect 71350 703670 71420 703740
rect 71440 703670 71510 703740
rect 71530 703670 71600 703740
rect 70090 703580 70160 703650
rect 70180 703580 70250 703650
rect 70270 703580 70340 703650
rect 70360 703580 70430 703650
rect 70450 703580 70520 703650
rect 70540 703580 70610 703650
rect 70630 703580 70700 703650
rect 70720 703580 70790 703650
rect 70810 703580 70880 703650
rect 70900 703580 70970 703650
rect 70990 703580 71060 703650
rect 71080 703580 71150 703650
rect 71170 703580 71240 703650
rect 71260 703580 71330 703650
rect 71350 703580 71420 703650
rect 71440 703580 71510 703650
rect 71530 703580 71600 703650
rect 70090 703490 70160 703560
rect 70180 703490 70250 703560
rect 70270 703490 70340 703560
rect 70360 703490 70430 703560
rect 70450 703490 70520 703560
rect 70540 703490 70610 703560
rect 70630 703490 70700 703560
rect 70720 703490 70790 703560
rect 70810 703490 70880 703560
rect 70900 703490 70970 703560
rect 70990 703490 71060 703560
rect 71080 703490 71150 703560
rect 71170 703490 71240 703560
rect 71260 703490 71330 703560
rect 71350 703490 71420 703560
rect 71440 703490 71510 703560
rect 71530 703490 71600 703560
rect 70090 703400 70160 703470
rect 70180 703400 70250 703470
rect 70270 703400 70340 703470
rect 70360 703400 70430 703470
rect 70450 703400 70520 703470
rect 70540 703400 70610 703470
rect 70630 703400 70700 703470
rect 70720 703400 70790 703470
rect 70810 703400 70880 703470
rect 70900 703400 70970 703470
rect 70990 703400 71060 703470
rect 71080 703400 71150 703470
rect 71170 703400 71240 703470
rect 71260 703400 71330 703470
rect 71350 703400 71420 703470
rect 71440 703400 71510 703470
rect 71530 703400 71600 703470
rect 70090 703310 70160 703380
rect 70180 703310 70250 703380
rect 70270 703310 70340 703380
rect 70360 703310 70430 703380
rect 70450 703310 70520 703380
rect 70540 703310 70610 703380
rect 70630 703310 70700 703380
rect 70720 703310 70790 703380
rect 70810 703310 70880 703380
rect 70900 703310 70970 703380
rect 70990 703310 71060 703380
rect 71080 703310 71150 703380
rect 71170 703310 71240 703380
rect 71260 703310 71330 703380
rect 71350 703310 71420 703380
rect 71440 703310 71510 703380
rect 71530 703310 71600 703380
rect 70090 703220 70160 703290
rect 70180 703220 70250 703290
rect 70270 703220 70340 703290
rect 70360 703220 70430 703290
rect 70450 703220 70520 703290
rect 70540 703220 70610 703290
rect 70630 703220 70700 703290
rect 70720 703220 70790 703290
rect 70810 703220 70880 703290
rect 70900 703220 70970 703290
rect 70990 703220 71060 703290
rect 71080 703220 71150 703290
rect 71170 703220 71240 703290
rect 71260 703220 71330 703290
rect 71350 703220 71420 703290
rect 71440 703220 71510 703290
rect 71530 703220 71600 703290
rect 70090 703130 70160 703200
rect 70180 703130 70250 703200
rect 70270 703130 70340 703200
rect 70360 703130 70430 703200
rect 70450 703130 70520 703200
rect 70540 703130 70610 703200
rect 70630 703130 70700 703200
rect 70720 703130 70790 703200
rect 70810 703130 70880 703200
rect 70900 703130 70970 703200
rect 70990 703130 71060 703200
rect 71080 703130 71150 703200
rect 71170 703130 71240 703200
rect 71260 703130 71330 703200
rect 71350 703130 71420 703200
rect 71440 703130 71510 703200
rect 71530 703130 71600 703200
rect 70090 703040 70160 703110
rect 70180 703040 70250 703110
rect 70270 703040 70340 703110
rect 70360 703040 70430 703110
rect 70450 703040 70520 703110
rect 70540 703040 70610 703110
rect 70630 703040 70700 703110
rect 70720 703040 70790 703110
rect 70810 703040 70880 703110
rect 70900 703040 70970 703110
rect 70990 703040 71060 703110
rect 71080 703040 71150 703110
rect 71170 703040 71240 703110
rect 71260 703040 71330 703110
rect 71350 703040 71420 703110
rect 71440 703040 71510 703110
rect 71530 703040 71600 703110
rect 70090 702950 70160 703020
rect 70180 702950 70250 703020
rect 70270 702950 70340 703020
rect 70360 702950 70430 703020
rect 70450 702950 70520 703020
rect 70540 702950 70610 703020
rect 70630 702950 70700 703020
rect 70720 702950 70790 703020
rect 70810 702950 70880 703020
rect 70900 702950 70970 703020
rect 70990 702950 71060 703020
rect 71080 702950 71150 703020
rect 71170 702950 71240 703020
rect 71260 702950 71330 703020
rect 71350 702950 71420 703020
rect 71440 702950 71510 703020
rect 71530 702950 71600 703020
rect 70090 702860 70160 702930
rect 70180 702860 70250 702930
rect 70270 702860 70340 702930
rect 70360 702860 70430 702930
rect 70450 702860 70520 702930
rect 70540 702860 70610 702930
rect 70630 702860 70700 702930
rect 70720 702860 70790 702930
rect 70810 702860 70880 702930
rect 70900 702860 70970 702930
rect 70990 702860 71060 702930
rect 71080 702860 71150 702930
rect 71170 702860 71240 702930
rect 71260 702860 71330 702930
rect 71350 702860 71420 702930
rect 71440 702860 71510 702930
rect 71530 702860 71600 702930
rect 70090 702770 70160 702840
rect 70180 702770 70250 702840
rect 70270 702770 70340 702840
rect 70360 702770 70430 702840
rect 70450 702770 70520 702840
rect 70540 702770 70610 702840
rect 70630 702770 70700 702840
rect 70720 702770 70790 702840
rect 70810 702770 70880 702840
rect 70900 702770 70970 702840
rect 70990 702770 71060 702840
rect 71080 702770 71150 702840
rect 71170 702770 71240 702840
rect 71260 702770 71330 702840
rect 71350 702770 71420 702840
rect 71440 702770 71510 702840
rect 71530 702770 71600 702840
rect 70090 702680 70160 702750
rect 70180 702680 70250 702750
rect 70270 702680 70340 702750
rect 70360 702680 70430 702750
rect 70450 702680 70520 702750
rect 70540 702680 70610 702750
rect 70630 702680 70700 702750
rect 70720 702680 70790 702750
rect 70810 702680 70880 702750
rect 70900 702680 70970 702750
rect 70990 702680 71060 702750
rect 71080 702680 71150 702750
rect 71170 702680 71240 702750
rect 71260 702680 71330 702750
rect 71350 702680 71420 702750
rect 71440 702680 71510 702750
rect 71530 702680 71600 702750
rect 70090 702590 70160 702660
rect 70180 702590 70250 702660
rect 70270 702590 70340 702660
rect 70360 702590 70430 702660
rect 70450 702590 70520 702660
rect 70540 702590 70610 702660
rect 70630 702590 70700 702660
rect 70720 702590 70790 702660
rect 70810 702590 70880 702660
rect 70900 702590 70970 702660
rect 70990 702590 71060 702660
rect 71080 702590 71150 702660
rect 71170 702590 71240 702660
rect 71260 702590 71330 702660
rect 71350 702590 71420 702660
rect 71440 702590 71510 702660
rect 71530 702590 71600 702660
rect 70090 702500 70160 702570
rect 70180 702500 70250 702570
rect 70270 702500 70340 702570
rect 70360 702500 70430 702570
rect 70450 702500 70520 702570
rect 70540 702500 70610 702570
rect 70630 702500 70700 702570
rect 70720 702500 70790 702570
rect 70810 702500 70880 702570
rect 70900 702500 70970 702570
rect 70990 702500 71060 702570
rect 71080 702500 71150 702570
rect 71170 702500 71240 702570
rect 71260 702500 71330 702570
rect 71350 702500 71420 702570
rect 71440 702500 71510 702570
rect 71530 702500 71600 702570
rect 70090 702410 70160 702480
rect 70180 702410 70250 702480
rect 70270 702410 70340 702480
rect 70360 702410 70430 702480
rect 70450 702410 70520 702480
rect 70540 702410 70610 702480
rect 70630 702410 70700 702480
rect 70720 702410 70790 702480
rect 70810 702410 70880 702480
rect 70900 702410 70970 702480
rect 70990 702410 71060 702480
rect 71080 702410 71150 702480
rect 71170 702410 71240 702480
rect 71260 702410 71330 702480
rect 71350 702410 71420 702480
rect 71440 702410 71510 702480
rect 71530 702410 71600 702480
rect 70090 702320 70160 702390
rect 70180 702320 70250 702390
rect 70270 702320 70340 702390
rect 70360 702320 70430 702390
rect 70450 702320 70520 702390
rect 70540 702320 70610 702390
rect 70630 702320 70700 702390
rect 70720 702320 70790 702390
rect 70810 702320 70880 702390
rect 70900 702320 70970 702390
rect 70990 702320 71060 702390
rect 71080 702320 71150 702390
rect 71170 702320 71240 702390
rect 71260 702320 71330 702390
rect 71350 702320 71420 702390
rect 71440 702320 71510 702390
rect 71530 702320 71600 702390
rect 121788 703760 121858 703830
rect 121878 703760 121948 703830
rect 121968 703760 122038 703830
rect 122058 703760 122128 703830
rect 122148 703760 122218 703830
rect 122238 703760 122308 703830
rect 122328 703760 122398 703830
rect 122418 703760 122488 703830
rect 122508 703760 122578 703830
rect 122598 703760 122668 703830
rect 122688 703760 122758 703830
rect 122778 703760 122848 703830
rect 122868 703760 122938 703830
rect 122958 703760 123028 703830
rect 123048 703760 123118 703830
rect 123138 703760 123208 703830
rect 123228 703760 123298 703830
rect 121788 703670 121858 703740
rect 121878 703670 121948 703740
rect 121968 703670 122038 703740
rect 122058 703670 122128 703740
rect 122148 703670 122218 703740
rect 122238 703670 122308 703740
rect 122328 703670 122398 703740
rect 122418 703670 122488 703740
rect 122508 703670 122578 703740
rect 122598 703670 122668 703740
rect 122688 703670 122758 703740
rect 122778 703670 122848 703740
rect 122868 703670 122938 703740
rect 122958 703670 123028 703740
rect 123048 703670 123118 703740
rect 123138 703670 123208 703740
rect 123228 703670 123298 703740
rect 121788 703580 121858 703650
rect 121878 703580 121948 703650
rect 121968 703580 122038 703650
rect 122058 703580 122128 703650
rect 122148 703580 122218 703650
rect 122238 703580 122308 703650
rect 122328 703580 122398 703650
rect 122418 703580 122488 703650
rect 122508 703580 122578 703650
rect 122598 703580 122668 703650
rect 122688 703580 122758 703650
rect 122778 703580 122848 703650
rect 122868 703580 122938 703650
rect 122958 703580 123028 703650
rect 123048 703580 123118 703650
rect 123138 703580 123208 703650
rect 123228 703580 123298 703650
rect 121788 703490 121858 703560
rect 121878 703490 121948 703560
rect 121968 703490 122038 703560
rect 122058 703490 122128 703560
rect 122148 703490 122218 703560
rect 122238 703490 122308 703560
rect 122328 703490 122398 703560
rect 122418 703490 122488 703560
rect 122508 703490 122578 703560
rect 122598 703490 122668 703560
rect 122688 703490 122758 703560
rect 122778 703490 122848 703560
rect 122868 703490 122938 703560
rect 122958 703490 123028 703560
rect 123048 703490 123118 703560
rect 123138 703490 123208 703560
rect 123228 703490 123298 703560
rect 121788 703400 121858 703470
rect 121878 703400 121948 703470
rect 121968 703400 122038 703470
rect 122058 703400 122128 703470
rect 122148 703400 122218 703470
rect 122238 703400 122308 703470
rect 122328 703400 122398 703470
rect 122418 703400 122488 703470
rect 122508 703400 122578 703470
rect 122598 703400 122668 703470
rect 122688 703400 122758 703470
rect 122778 703400 122848 703470
rect 122868 703400 122938 703470
rect 122958 703400 123028 703470
rect 123048 703400 123118 703470
rect 123138 703400 123208 703470
rect 123228 703400 123298 703470
rect 121788 703310 121858 703380
rect 121878 703310 121948 703380
rect 121968 703310 122038 703380
rect 122058 703310 122128 703380
rect 122148 703310 122218 703380
rect 122238 703310 122308 703380
rect 122328 703310 122398 703380
rect 122418 703310 122488 703380
rect 122508 703310 122578 703380
rect 122598 703310 122668 703380
rect 122688 703310 122758 703380
rect 122778 703310 122848 703380
rect 122868 703310 122938 703380
rect 122958 703310 123028 703380
rect 123048 703310 123118 703380
rect 123138 703310 123208 703380
rect 123228 703310 123298 703380
rect 121788 703220 121858 703290
rect 121878 703220 121948 703290
rect 121968 703220 122038 703290
rect 122058 703220 122128 703290
rect 122148 703220 122218 703290
rect 122238 703220 122308 703290
rect 122328 703220 122398 703290
rect 122418 703220 122488 703290
rect 122508 703220 122578 703290
rect 122598 703220 122668 703290
rect 122688 703220 122758 703290
rect 122778 703220 122848 703290
rect 122868 703220 122938 703290
rect 122958 703220 123028 703290
rect 123048 703220 123118 703290
rect 123138 703220 123208 703290
rect 123228 703220 123298 703290
rect 121788 703130 121858 703200
rect 121878 703130 121948 703200
rect 121968 703130 122038 703200
rect 122058 703130 122128 703200
rect 122148 703130 122218 703200
rect 122238 703130 122308 703200
rect 122328 703130 122398 703200
rect 122418 703130 122488 703200
rect 122508 703130 122578 703200
rect 122598 703130 122668 703200
rect 122688 703130 122758 703200
rect 122778 703130 122848 703200
rect 122868 703130 122938 703200
rect 122958 703130 123028 703200
rect 123048 703130 123118 703200
rect 123138 703130 123208 703200
rect 123228 703130 123298 703200
rect 121788 703040 121858 703110
rect 121878 703040 121948 703110
rect 121968 703040 122038 703110
rect 122058 703040 122128 703110
rect 122148 703040 122218 703110
rect 122238 703040 122308 703110
rect 122328 703040 122398 703110
rect 122418 703040 122488 703110
rect 122508 703040 122578 703110
rect 122598 703040 122668 703110
rect 122688 703040 122758 703110
rect 122778 703040 122848 703110
rect 122868 703040 122938 703110
rect 122958 703040 123028 703110
rect 123048 703040 123118 703110
rect 123138 703040 123208 703110
rect 123228 703040 123298 703110
rect 121788 702950 121858 703020
rect 121878 702950 121948 703020
rect 121968 702950 122038 703020
rect 122058 702950 122128 703020
rect 122148 702950 122218 703020
rect 122238 702950 122308 703020
rect 122328 702950 122398 703020
rect 122418 702950 122488 703020
rect 122508 702950 122578 703020
rect 122598 702950 122668 703020
rect 122688 702950 122758 703020
rect 122778 702950 122848 703020
rect 122868 702950 122938 703020
rect 122958 702950 123028 703020
rect 123048 702950 123118 703020
rect 123138 702950 123208 703020
rect 123228 702950 123298 703020
rect 121788 702860 121858 702930
rect 121878 702860 121948 702930
rect 121968 702860 122038 702930
rect 122058 702860 122128 702930
rect 122148 702860 122218 702930
rect 122238 702860 122308 702930
rect 122328 702860 122398 702930
rect 122418 702860 122488 702930
rect 122508 702860 122578 702930
rect 122598 702860 122668 702930
rect 122688 702860 122758 702930
rect 122778 702860 122848 702930
rect 122868 702860 122938 702930
rect 122958 702860 123028 702930
rect 123048 702860 123118 702930
rect 123138 702860 123208 702930
rect 123228 702860 123298 702930
rect 121788 702770 121858 702840
rect 121878 702770 121948 702840
rect 121968 702770 122038 702840
rect 122058 702770 122128 702840
rect 122148 702770 122218 702840
rect 122238 702770 122308 702840
rect 122328 702770 122398 702840
rect 122418 702770 122488 702840
rect 122508 702770 122578 702840
rect 122598 702770 122668 702840
rect 122688 702770 122758 702840
rect 122778 702770 122848 702840
rect 122868 702770 122938 702840
rect 122958 702770 123028 702840
rect 123048 702770 123118 702840
rect 123138 702770 123208 702840
rect 123228 702770 123298 702840
rect 121788 702680 121858 702750
rect 121878 702680 121948 702750
rect 121968 702680 122038 702750
rect 122058 702680 122128 702750
rect 122148 702680 122218 702750
rect 122238 702680 122308 702750
rect 122328 702680 122398 702750
rect 122418 702680 122488 702750
rect 122508 702680 122578 702750
rect 122598 702680 122668 702750
rect 122688 702680 122758 702750
rect 122778 702680 122848 702750
rect 122868 702680 122938 702750
rect 122958 702680 123028 702750
rect 123048 702680 123118 702750
rect 123138 702680 123208 702750
rect 123228 702680 123298 702750
rect 121788 702590 121858 702660
rect 121878 702590 121948 702660
rect 121968 702590 122038 702660
rect 122058 702590 122128 702660
rect 122148 702590 122218 702660
rect 122238 702590 122308 702660
rect 122328 702590 122398 702660
rect 122418 702590 122488 702660
rect 122508 702590 122578 702660
rect 122598 702590 122668 702660
rect 122688 702590 122758 702660
rect 122778 702590 122848 702660
rect 122868 702590 122938 702660
rect 122958 702590 123028 702660
rect 123048 702590 123118 702660
rect 123138 702590 123208 702660
rect 123228 702590 123298 702660
rect 121788 702500 121858 702570
rect 121878 702500 121948 702570
rect 121968 702500 122038 702570
rect 122058 702500 122128 702570
rect 122148 702500 122218 702570
rect 122238 702500 122308 702570
rect 122328 702500 122398 702570
rect 122418 702500 122488 702570
rect 122508 702500 122578 702570
rect 122598 702500 122668 702570
rect 122688 702500 122758 702570
rect 122778 702500 122848 702570
rect 122868 702500 122938 702570
rect 122958 702500 123028 702570
rect 123048 702500 123118 702570
rect 123138 702500 123208 702570
rect 123228 702500 123298 702570
rect 121788 702410 121858 702480
rect 121878 702410 121948 702480
rect 121968 702410 122038 702480
rect 122058 702410 122128 702480
rect 122148 702410 122218 702480
rect 122238 702410 122308 702480
rect 122328 702410 122398 702480
rect 122418 702410 122488 702480
rect 122508 702410 122578 702480
rect 122598 702410 122668 702480
rect 122688 702410 122758 702480
rect 122778 702410 122848 702480
rect 122868 702410 122938 702480
rect 122958 702410 123028 702480
rect 123048 702410 123118 702480
rect 123138 702410 123208 702480
rect 123228 702410 123298 702480
rect 121788 702320 121858 702390
rect 121878 702320 121948 702390
rect 121968 702320 122038 702390
rect 122058 702320 122128 702390
rect 122148 702320 122218 702390
rect 122238 702320 122308 702390
rect 122328 702320 122398 702390
rect 122418 702320 122488 702390
rect 122508 702320 122578 702390
rect 122598 702320 122668 702390
rect 122688 702320 122758 702390
rect 122778 702320 122848 702390
rect 122868 702320 122938 702390
rect 122958 702320 123028 702390
rect 123048 702320 123118 702390
rect 123138 702320 123208 702390
rect 123228 702320 123298 702390
rect 415630 702770 415700 702840
rect 415720 702770 415790 702840
rect 415810 702770 415880 702840
rect 415900 702770 415970 702840
rect 415990 702770 416060 702840
rect 416080 702770 416150 702840
rect 415630 702680 415700 702750
rect 415720 702680 415790 702750
rect 415810 702680 415880 702750
rect 415900 702680 415970 702750
rect 415990 702680 416060 702750
rect 416080 702680 416150 702750
rect 415630 702590 415700 702660
rect 415720 702590 415790 702660
rect 415810 702590 415880 702660
rect 415900 702590 415970 702660
rect 415990 702590 416060 702660
rect 416080 702590 416150 702660
rect 415630 702500 415700 702570
rect 415720 702500 415790 702570
rect 415810 702500 415880 702570
rect 415900 702500 415970 702570
rect 415990 702500 416060 702570
rect 416080 702500 416150 702570
rect 415630 702410 415700 702480
rect 415720 702410 415790 702480
rect 415810 702410 415880 702480
rect 415900 702410 415970 702480
rect 415990 702410 416060 702480
rect 416080 702410 416150 702480
rect 415630 702320 415700 702390
rect 415720 702320 415790 702390
rect 415810 702320 415880 702390
rect 415900 702320 415970 702390
rect 415990 702320 416060 702390
rect 416080 702320 416150 702390
rect 467630 702770 467700 702840
rect 467720 702770 467790 702840
rect 467810 702770 467880 702840
rect 467900 702770 467970 702840
rect 467990 702770 468060 702840
rect 468080 702770 468150 702840
rect 467630 702680 467700 702750
rect 467720 702680 467790 702750
rect 467810 702680 467880 702750
rect 467900 702680 467970 702750
rect 467990 702680 468060 702750
rect 468080 702680 468150 702750
rect 467630 702590 467700 702660
rect 467720 702590 467790 702660
rect 467810 702590 467880 702660
rect 467900 702590 467970 702660
rect 467990 702590 468060 702660
rect 468080 702590 468150 702660
rect 467630 702500 467700 702570
rect 467720 702500 467790 702570
rect 467810 702500 467880 702570
rect 467900 702500 467970 702570
rect 467990 702500 468060 702570
rect 468080 702500 468150 702570
rect 467630 702410 467700 702480
rect 467720 702410 467790 702480
rect 467810 702410 467880 702480
rect 467900 702410 467970 702480
rect 467990 702410 468060 702480
rect 468080 702410 468150 702480
rect 467630 702320 467700 702390
rect 467720 702320 467790 702390
rect 467810 702320 467880 702390
rect 467900 702320 467970 702390
rect 467990 702320 468060 702390
rect 468080 702320 468150 702390
rect 566740 702770 566810 702840
rect 566830 702770 566900 702840
rect 566920 702770 566990 702840
rect 567010 702770 567080 702840
rect 567100 702770 567170 702840
rect 567190 702770 567260 702840
rect 566740 702680 566810 702750
rect 566830 702680 566900 702750
rect 566920 702680 566990 702750
rect 567010 702680 567080 702750
rect 567100 702680 567170 702750
rect 567190 702680 567260 702750
rect 566740 702590 566810 702660
rect 566830 702590 566900 702660
rect 566920 702590 566990 702660
rect 567010 702590 567080 702660
rect 567100 702590 567170 702660
rect 567190 702590 567260 702660
rect 566740 702500 566810 702570
rect 566830 702500 566900 702570
rect 566920 702500 566990 702570
rect 567010 702500 567080 702570
rect 567100 702500 567170 702570
rect 567190 702500 567260 702570
rect 566740 702410 566810 702480
rect 566830 702410 566900 702480
rect 566920 702410 566990 702480
rect 567010 702410 567080 702480
rect 567100 702410 567170 702480
rect 567190 702410 567260 702480
rect 566740 702320 566810 702390
rect 566830 702320 566900 702390
rect 566920 702320 566990 702390
rect 567010 702320 567080 702390
rect 567100 702320 567170 702390
rect 567190 702320 567260 702390
rect 225164 700690 225404 700930
rect 225494 700690 225734 700930
rect 225824 700690 226064 700930
rect 226154 700690 226394 700930
rect 226484 700690 226724 700930
rect 226814 700690 227054 700930
rect 225164 700360 225404 700600
rect 225494 700360 225734 700600
rect 225824 700360 226064 700600
rect 226154 700360 226394 700600
rect 226484 700360 226724 700600
rect 226814 700360 227054 700600
rect 225164 700030 225404 700270
rect 225494 700030 225734 700270
rect 225824 700030 226064 700270
rect 226154 700030 226394 700270
rect 226484 700030 226724 700270
rect 226814 700030 227054 700270
rect 225164 699700 225404 699940
rect 225494 699700 225734 699940
rect 225824 699700 226064 699940
rect 226154 699700 226394 699940
rect 226484 699700 226724 699940
rect 226814 699700 227054 699940
rect 225164 699370 225404 699610
rect 225494 699370 225734 699610
rect 225824 699370 226064 699610
rect 226154 699370 226394 699610
rect 226484 699370 226724 699610
rect 226814 699370 227054 699610
rect 225164 699040 225404 699280
rect 225494 699040 225734 699280
rect 225824 699040 226064 699280
rect 226154 699040 226394 699280
rect 226484 699040 226724 699280
rect 226814 699040 227054 699280
rect 225164 698710 225404 698950
rect 225494 698710 225734 698950
rect 225824 698710 226064 698950
rect 226154 698710 226394 698950
rect 226484 698710 226724 698950
rect 226814 698710 227054 698950
rect 225164 698380 225404 698620
rect 225494 698380 225734 698620
rect 225824 698380 226064 698620
rect 226154 698380 226394 698620
rect 226484 698380 226724 698620
rect 226814 698380 227054 698620
rect 225164 698050 225404 698290
rect 225494 698050 225734 698290
rect 225824 698050 226064 698290
rect 226154 698050 226394 698290
rect 226484 698050 226724 698290
rect 226814 698050 227054 698290
rect 225164 697720 225404 697960
rect 225494 697720 225734 697960
rect 225824 697720 226064 697960
rect 226154 697720 226394 697960
rect 226484 697720 226724 697960
rect 226814 697720 227054 697960
rect 225164 697390 225404 697630
rect 225494 697390 225734 697630
rect 225824 697390 226064 697630
rect 226154 697390 226394 697630
rect 226484 697390 226724 697630
rect 226814 697390 227054 697630
rect 225164 697060 225404 697300
rect 225494 697060 225734 697300
rect 225824 697060 226064 697300
rect 226154 697060 226394 697300
rect 226484 697060 226724 697300
rect 226814 697060 227054 697300
rect 225164 696730 225404 696970
rect 225494 696730 225734 696970
rect 225824 696730 226064 696970
rect 226154 696730 226394 696970
rect 226484 696730 226724 696970
rect 226814 696730 227054 696970
rect 225164 696400 225404 696640
rect 225494 696400 225734 696640
rect 225824 696400 226064 696640
rect 226154 696400 226394 696640
rect 226484 696400 226724 696640
rect 226814 696400 227054 696640
rect 225164 696070 225404 696310
rect 225494 696070 225734 696310
rect 225824 696070 226064 696310
rect 226154 696070 226394 696310
rect 226484 696070 226724 696310
rect 226814 696070 227054 696310
rect 170964 692690 171204 692930
rect 171294 692690 171534 692930
rect 171624 692690 171864 692930
rect 171954 692690 172194 692930
rect 172284 692690 172524 692930
rect 172614 692690 172854 692930
rect 170964 692360 171204 692600
rect 171294 692360 171534 692600
rect 171624 692360 171864 692600
rect 171954 692360 172194 692600
rect 172284 692360 172524 692600
rect 172614 692360 172854 692600
rect 170964 692030 171204 692270
rect 171294 692030 171534 692270
rect 171624 692030 171864 692270
rect 171954 692030 172194 692270
rect 172284 692030 172524 692270
rect 172614 692030 172854 692270
rect 170964 691700 171204 691940
rect 171294 691700 171534 691940
rect 171624 691700 171864 691940
rect 171954 691700 172194 691940
rect 172284 691700 172524 691940
rect 172614 691700 172854 691940
rect 170964 691370 171204 691610
rect 171294 691370 171534 691610
rect 171624 691370 171864 691610
rect 171954 691370 172194 691610
rect 172284 691370 172524 691610
rect 172614 691370 172854 691610
rect 170964 691040 171204 691280
rect 171294 691040 171534 691280
rect 171624 691040 171864 691280
rect 171954 691040 172194 691280
rect 172284 691040 172524 691280
rect 172614 691040 172854 691280
rect 170964 690710 171204 690950
rect 171294 690710 171534 690950
rect 171624 690710 171864 690950
rect 171954 690710 172194 690950
rect 172284 690710 172524 690950
rect 172614 690710 172854 690950
rect 170964 690380 171204 690620
rect 171294 690380 171534 690620
rect 171624 690380 171864 690620
rect 171954 690380 172194 690620
rect 172284 690380 172524 690620
rect 172614 690380 172854 690620
rect 170964 690050 171204 690290
rect 171294 690050 171534 690290
rect 171624 690050 171864 690290
rect 171954 690050 172194 690290
rect 172284 690050 172524 690290
rect 172614 690050 172854 690290
rect 170964 689720 171204 689960
rect 171294 689720 171534 689960
rect 171624 689720 171864 689960
rect 171954 689720 172194 689960
rect 172284 689720 172524 689960
rect 172614 689720 172854 689960
rect 170964 689390 171204 689630
rect 171294 689390 171534 689630
rect 171624 689390 171864 689630
rect 171954 689390 172194 689630
rect 172284 689390 172524 689630
rect 172614 689390 172854 689630
rect 170964 689060 171204 689300
rect 171294 689060 171534 689300
rect 171624 689060 171864 689300
rect 171954 689060 172194 689300
rect 172284 689060 172524 689300
rect 172614 689060 172854 689300
rect 170964 688730 171204 688970
rect 171294 688730 171534 688970
rect 171624 688730 171864 688970
rect 171954 688730 172194 688970
rect 172284 688730 172524 688970
rect 172614 688730 172854 688970
rect 170964 688400 171204 688640
rect 171294 688400 171534 688640
rect 171624 688400 171864 688640
rect 171954 688400 172194 688640
rect 172284 688400 172524 688640
rect 172614 688400 172854 688640
rect 170964 688070 171204 688310
rect 171294 688070 171534 688310
rect 171624 688070 171864 688310
rect 171954 688070 172194 688310
rect 172284 688070 172524 688310
rect 172614 688070 172854 688310
rect 18120 687300 18190 687370
rect 18210 687300 18280 687370
rect 18300 687300 18370 687370
rect 18390 687300 18460 687370
rect 18480 687300 18550 687370
rect 18570 687300 18640 687370
rect 18660 687300 18730 687370
rect 18750 687300 18820 687370
rect 18840 687300 18910 687370
rect 18930 687300 19000 687370
rect 19020 687300 19090 687370
rect 19110 687300 19180 687370
rect 19200 687300 19270 687370
rect 19290 687300 19360 687370
rect 19380 687300 19450 687370
rect 19470 687300 19540 687370
rect 19560 687300 19630 687370
rect 18120 687210 18190 687280
rect 18210 687210 18280 687280
rect 18300 687210 18370 687280
rect 18390 687210 18460 687280
rect 18480 687210 18550 687280
rect 18570 687210 18640 687280
rect 18660 687210 18730 687280
rect 18750 687210 18820 687280
rect 18840 687210 18910 687280
rect 18930 687210 19000 687280
rect 19020 687210 19090 687280
rect 19110 687210 19180 687280
rect 19200 687210 19270 687280
rect 19290 687210 19360 687280
rect 19380 687210 19450 687280
rect 19470 687210 19540 687280
rect 19560 687210 19630 687280
rect 18120 687120 18190 687190
rect 18210 687120 18280 687190
rect 18300 687120 18370 687190
rect 18390 687120 18460 687190
rect 18480 687120 18550 687190
rect 18570 687120 18640 687190
rect 18660 687120 18730 687190
rect 18750 687120 18820 687190
rect 18840 687120 18910 687190
rect 18930 687120 19000 687190
rect 19020 687120 19090 687190
rect 19110 687120 19180 687190
rect 19200 687120 19270 687190
rect 19290 687120 19360 687190
rect 19380 687120 19450 687190
rect 19470 687120 19540 687190
rect 19560 687120 19630 687190
rect 18120 687030 18190 687100
rect 18210 687030 18280 687100
rect 18300 687030 18370 687100
rect 18390 687030 18460 687100
rect 18480 687030 18550 687100
rect 18570 687030 18640 687100
rect 18660 687030 18730 687100
rect 18750 687030 18820 687100
rect 18840 687030 18910 687100
rect 18930 687030 19000 687100
rect 19020 687030 19090 687100
rect 19110 687030 19180 687100
rect 19200 687030 19270 687100
rect 19290 687030 19360 687100
rect 19380 687030 19450 687100
rect 19470 687030 19540 687100
rect 19560 687030 19630 687100
rect 18120 686940 18190 687010
rect 18210 686940 18280 687010
rect 18300 686940 18370 687010
rect 18390 686940 18460 687010
rect 18480 686940 18550 687010
rect 18570 686940 18640 687010
rect 18660 686940 18730 687010
rect 18750 686940 18820 687010
rect 18840 686940 18910 687010
rect 18930 686940 19000 687010
rect 19020 686940 19090 687010
rect 19110 686940 19180 687010
rect 19200 686940 19270 687010
rect 19290 686940 19360 687010
rect 19380 686940 19450 687010
rect 19470 686940 19540 687010
rect 19560 686940 19630 687010
rect 18120 686850 18190 686920
rect 18210 686850 18280 686920
rect 18300 686850 18370 686920
rect 18390 686850 18460 686920
rect 18480 686850 18550 686920
rect 18570 686850 18640 686920
rect 18660 686850 18730 686920
rect 18750 686850 18820 686920
rect 18840 686850 18910 686920
rect 18930 686850 19000 686920
rect 19020 686850 19090 686920
rect 19110 686850 19180 686920
rect 19200 686850 19270 686920
rect 19290 686850 19360 686920
rect 19380 686850 19450 686920
rect 19470 686850 19540 686920
rect 19560 686850 19630 686920
rect 18120 686760 18190 686830
rect 18210 686760 18280 686830
rect 18300 686760 18370 686830
rect 18390 686760 18460 686830
rect 18480 686760 18550 686830
rect 18570 686760 18640 686830
rect 18660 686760 18730 686830
rect 18750 686760 18820 686830
rect 18840 686760 18910 686830
rect 18930 686760 19000 686830
rect 19020 686760 19090 686830
rect 19110 686760 19180 686830
rect 19200 686760 19270 686830
rect 19290 686760 19360 686830
rect 19380 686760 19450 686830
rect 19470 686760 19540 686830
rect 19560 686760 19630 686830
rect 18120 686670 18190 686740
rect 18210 686670 18280 686740
rect 18300 686670 18370 686740
rect 18390 686670 18460 686740
rect 18480 686670 18550 686740
rect 18570 686670 18640 686740
rect 18660 686670 18730 686740
rect 18750 686670 18820 686740
rect 18840 686670 18910 686740
rect 18930 686670 19000 686740
rect 19020 686670 19090 686740
rect 19110 686670 19180 686740
rect 19200 686670 19270 686740
rect 19290 686670 19360 686740
rect 19380 686670 19450 686740
rect 19470 686670 19540 686740
rect 19560 686670 19630 686740
rect 18120 686580 18190 686650
rect 18210 686580 18280 686650
rect 18300 686580 18370 686650
rect 18390 686580 18460 686650
rect 18480 686580 18550 686650
rect 18570 686580 18640 686650
rect 18660 686580 18730 686650
rect 18750 686580 18820 686650
rect 18840 686580 18910 686650
rect 18930 686580 19000 686650
rect 19020 686580 19090 686650
rect 19110 686580 19180 686650
rect 19200 686580 19270 686650
rect 19290 686580 19360 686650
rect 19380 686580 19450 686650
rect 19470 686580 19540 686650
rect 19560 686580 19630 686650
rect 18120 686490 18190 686560
rect 18210 686490 18280 686560
rect 18300 686490 18370 686560
rect 18390 686490 18460 686560
rect 18480 686490 18550 686560
rect 18570 686490 18640 686560
rect 18660 686490 18730 686560
rect 18750 686490 18820 686560
rect 18840 686490 18910 686560
rect 18930 686490 19000 686560
rect 19020 686490 19090 686560
rect 19110 686490 19180 686560
rect 19200 686490 19270 686560
rect 19290 686490 19360 686560
rect 19380 686490 19450 686560
rect 19470 686490 19540 686560
rect 19560 686490 19630 686560
rect 18120 686400 18190 686470
rect 18210 686400 18280 686470
rect 18300 686400 18370 686470
rect 18390 686400 18460 686470
rect 18480 686400 18550 686470
rect 18570 686400 18640 686470
rect 18660 686400 18730 686470
rect 18750 686400 18820 686470
rect 18840 686400 18910 686470
rect 18930 686400 19000 686470
rect 19020 686400 19090 686470
rect 19110 686400 19180 686470
rect 19200 686400 19270 686470
rect 19290 686400 19360 686470
rect 19380 686400 19450 686470
rect 19470 686400 19540 686470
rect 19560 686400 19630 686470
rect 18120 686310 18190 686380
rect 18210 686310 18280 686380
rect 18300 686310 18370 686380
rect 18390 686310 18460 686380
rect 18480 686310 18550 686380
rect 18570 686310 18640 686380
rect 18660 686310 18730 686380
rect 18750 686310 18820 686380
rect 18840 686310 18910 686380
rect 18930 686310 19000 686380
rect 19020 686310 19090 686380
rect 19110 686310 19180 686380
rect 19200 686310 19270 686380
rect 19290 686310 19360 686380
rect 19380 686310 19450 686380
rect 19470 686310 19540 686380
rect 19560 686310 19630 686380
rect 18120 686220 18190 686290
rect 18210 686220 18280 686290
rect 18300 686220 18370 686290
rect 18390 686220 18460 686290
rect 18480 686220 18550 686290
rect 18570 686220 18640 686290
rect 18660 686220 18730 686290
rect 18750 686220 18820 686290
rect 18840 686220 18910 686290
rect 18930 686220 19000 686290
rect 19020 686220 19090 686290
rect 19110 686220 19180 686290
rect 19200 686220 19270 686290
rect 19290 686220 19360 686290
rect 19380 686220 19450 686290
rect 19470 686220 19540 686290
rect 19560 686220 19630 686290
rect 18120 686130 18190 686200
rect 18210 686130 18280 686200
rect 18300 686130 18370 686200
rect 18390 686130 18460 686200
rect 18480 686130 18550 686200
rect 18570 686130 18640 686200
rect 18660 686130 18730 686200
rect 18750 686130 18820 686200
rect 18840 686130 18910 686200
rect 18930 686130 19000 686200
rect 19020 686130 19090 686200
rect 19110 686130 19180 686200
rect 19200 686130 19270 686200
rect 19290 686130 19360 686200
rect 19380 686130 19450 686200
rect 19470 686130 19540 686200
rect 19560 686130 19630 686200
rect 18120 686040 18190 686110
rect 18210 686040 18280 686110
rect 18300 686040 18370 686110
rect 18390 686040 18460 686110
rect 18480 686040 18550 686110
rect 18570 686040 18640 686110
rect 18660 686040 18730 686110
rect 18750 686040 18820 686110
rect 18840 686040 18910 686110
rect 18930 686040 19000 686110
rect 19020 686040 19090 686110
rect 19110 686040 19180 686110
rect 19200 686040 19270 686110
rect 19290 686040 19360 686110
rect 19380 686040 19450 686110
rect 19470 686040 19540 686110
rect 19560 686040 19630 686110
rect 18120 685950 18190 686020
rect 18210 685950 18280 686020
rect 18300 685950 18370 686020
rect 18390 685950 18460 686020
rect 18480 685950 18550 686020
rect 18570 685950 18640 686020
rect 18660 685950 18730 686020
rect 18750 685950 18820 686020
rect 18840 685950 18910 686020
rect 18930 685950 19000 686020
rect 19020 685950 19090 686020
rect 19110 685950 19180 686020
rect 19200 685950 19270 686020
rect 19290 685950 19360 686020
rect 19380 685950 19450 686020
rect 19470 685950 19540 686020
rect 19560 685950 19630 686020
rect 18120 685860 18190 685930
rect 18210 685860 18280 685930
rect 18300 685860 18370 685930
rect 18390 685860 18460 685930
rect 18480 685860 18550 685930
rect 18570 685860 18640 685930
rect 18660 685860 18730 685930
rect 18750 685860 18820 685930
rect 18840 685860 18910 685930
rect 18930 685860 19000 685930
rect 19020 685860 19090 685930
rect 19110 685860 19180 685930
rect 19200 685860 19270 685930
rect 19290 685860 19360 685930
rect 19380 685860 19450 685930
rect 19470 685860 19540 685930
rect 19560 685860 19630 685930
rect 18120 685770 18190 685840
rect 18210 685770 18280 685840
rect 18300 685770 18370 685840
rect 18390 685770 18460 685840
rect 18480 685770 18550 685840
rect 18570 685770 18640 685840
rect 18660 685770 18730 685840
rect 18750 685770 18820 685840
rect 18840 685770 18910 685840
rect 18930 685770 19000 685840
rect 19020 685770 19090 685840
rect 19110 685770 19180 685840
rect 19200 685770 19270 685840
rect 19290 685770 19360 685840
rect 19380 685770 19450 685840
rect 19470 685770 19540 685840
rect 19560 685770 19630 685840
rect 18120 685680 18190 685750
rect 18210 685680 18280 685750
rect 18300 685680 18370 685750
rect 18390 685680 18460 685750
rect 18480 685680 18550 685750
rect 18570 685680 18640 685750
rect 18660 685680 18730 685750
rect 18750 685680 18820 685750
rect 18840 685680 18910 685750
rect 18930 685680 19000 685750
rect 19020 685680 19090 685750
rect 19110 685680 19180 685750
rect 19200 685680 19270 685750
rect 19290 685680 19360 685750
rect 19380 685680 19450 685750
rect 19470 685680 19540 685750
rect 19560 685680 19630 685750
rect 18120 685590 18190 685660
rect 18210 685590 18280 685660
rect 18300 685590 18370 685660
rect 18390 685590 18460 685660
rect 18480 685590 18550 685660
rect 18570 685590 18640 685660
rect 18660 685590 18730 685660
rect 18750 685590 18820 685660
rect 18840 685590 18910 685660
rect 18930 685590 19000 685660
rect 19020 685590 19090 685660
rect 19110 685590 19180 685660
rect 19200 685590 19270 685660
rect 19290 685590 19360 685660
rect 19380 685590 19450 685660
rect 19470 685590 19540 685660
rect 19560 685590 19630 685660
rect 18120 685500 18190 685570
rect 18210 685500 18280 685570
rect 18300 685500 18370 685570
rect 18390 685500 18460 685570
rect 18480 685500 18550 685570
rect 18570 685500 18640 685570
rect 18660 685500 18730 685570
rect 18750 685500 18820 685570
rect 18840 685500 18910 685570
rect 18930 685500 19000 685570
rect 19020 685500 19090 685570
rect 19110 685500 19180 685570
rect 19200 685500 19270 685570
rect 19290 685500 19360 685570
rect 19380 685500 19450 685570
rect 19470 685500 19540 685570
rect 19560 685500 19630 685570
rect 18120 685410 18190 685480
rect 18210 685410 18280 685480
rect 18300 685410 18370 685480
rect 18390 685410 18460 685480
rect 18480 685410 18550 685480
rect 18570 685410 18640 685480
rect 18660 685410 18730 685480
rect 18750 685410 18820 685480
rect 18840 685410 18910 685480
rect 18930 685410 19000 685480
rect 19020 685410 19090 685480
rect 19110 685410 19180 685480
rect 19200 685410 19270 685480
rect 19290 685410 19360 685480
rect 19380 685410 19450 685480
rect 19470 685410 19540 685480
rect 19560 685410 19630 685480
rect 120 683590 190 683660
rect 210 683590 280 683660
rect 300 683590 370 683660
rect 390 683590 460 683660
rect 480 683590 550 683660
rect 570 683590 640 683660
rect 660 683590 730 683660
rect 750 683590 820 683660
rect 840 683590 910 683660
rect 930 683590 1000 683660
rect 1020 683590 1090 683660
rect 1110 683590 1180 683660
rect 1200 683590 1270 683660
rect 1290 683590 1360 683660
rect 1380 683590 1450 683660
rect 1470 683590 1540 683660
rect 1560 683590 1630 683660
rect 120 683500 190 683570
rect 210 683500 280 683570
rect 300 683500 370 683570
rect 390 683500 460 683570
rect 480 683500 550 683570
rect 570 683500 640 683570
rect 660 683500 730 683570
rect 750 683500 820 683570
rect 840 683500 910 683570
rect 930 683500 1000 683570
rect 1020 683500 1090 683570
rect 1110 683500 1180 683570
rect 1200 683500 1270 683570
rect 1290 683500 1360 683570
rect 1380 683500 1450 683570
rect 1470 683500 1540 683570
rect 1560 683500 1630 683570
rect 120 683410 190 683480
rect 210 683410 280 683480
rect 300 683410 370 683480
rect 390 683410 460 683480
rect 480 683410 550 683480
rect 570 683410 640 683480
rect 660 683410 730 683480
rect 750 683410 820 683480
rect 840 683410 910 683480
rect 930 683410 1000 683480
rect 1020 683410 1090 683480
rect 1110 683410 1180 683480
rect 1200 683410 1270 683480
rect 1290 683410 1360 683480
rect 1380 683410 1450 683480
rect 1470 683410 1540 683480
rect 1560 683410 1630 683480
rect 120 683320 190 683390
rect 210 683320 280 683390
rect 300 683320 370 683390
rect 390 683320 460 683390
rect 480 683320 550 683390
rect 570 683320 640 683390
rect 660 683320 730 683390
rect 750 683320 820 683390
rect 840 683320 910 683390
rect 930 683320 1000 683390
rect 1020 683320 1090 683390
rect 1110 683320 1180 683390
rect 1200 683320 1270 683390
rect 1290 683320 1360 683390
rect 1380 683320 1450 683390
rect 1470 683320 1540 683390
rect 1560 683320 1630 683390
rect 120 683230 190 683300
rect 210 683230 280 683300
rect 300 683230 370 683300
rect 390 683230 460 683300
rect 480 683230 550 683300
rect 570 683230 640 683300
rect 660 683230 730 683300
rect 750 683230 820 683300
rect 840 683230 910 683300
rect 930 683230 1000 683300
rect 1020 683230 1090 683300
rect 1110 683230 1180 683300
rect 1200 683230 1270 683300
rect 1290 683230 1360 683300
rect 1380 683230 1450 683300
rect 1470 683230 1540 683300
rect 1560 683230 1630 683300
rect 120 683140 190 683210
rect 210 683140 280 683210
rect 300 683140 370 683210
rect 390 683140 460 683210
rect 480 683140 550 683210
rect 570 683140 640 683210
rect 660 683140 730 683210
rect 750 683140 820 683210
rect 840 683140 910 683210
rect 930 683140 1000 683210
rect 1020 683140 1090 683210
rect 1110 683140 1180 683210
rect 1200 683140 1270 683210
rect 1290 683140 1360 683210
rect 1380 683140 1450 683210
rect 1470 683140 1540 683210
rect 1560 683140 1630 683210
rect 120 683050 190 683120
rect 210 683050 280 683120
rect 300 683050 370 683120
rect 390 683050 460 683120
rect 480 683050 550 683120
rect 570 683050 640 683120
rect 660 683050 730 683120
rect 750 683050 820 683120
rect 840 683050 910 683120
rect 930 683050 1000 683120
rect 1020 683050 1090 683120
rect 1110 683050 1180 683120
rect 1200 683050 1270 683120
rect 1290 683050 1360 683120
rect 1380 683050 1450 683120
rect 1470 683050 1540 683120
rect 1560 683050 1630 683120
rect 120 682960 190 683030
rect 210 682960 280 683030
rect 300 682960 370 683030
rect 390 682960 460 683030
rect 480 682960 550 683030
rect 570 682960 640 683030
rect 660 682960 730 683030
rect 750 682960 820 683030
rect 840 682960 910 683030
rect 930 682960 1000 683030
rect 1020 682960 1090 683030
rect 1110 682960 1180 683030
rect 1200 682960 1270 683030
rect 1290 682960 1360 683030
rect 1380 682960 1450 683030
rect 1470 682960 1540 683030
rect 1560 682960 1630 683030
rect 120 682870 190 682940
rect 210 682870 280 682940
rect 300 682870 370 682940
rect 390 682870 460 682940
rect 480 682870 550 682940
rect 570 682870 640 682940
rect 660 682870 730 682940
rect 750 682870 820 682940
rect 840 682870 910 682940
rect 930 682870 1000 682940
rect 1020 682870 1090 682940
rect 1110 682870 1180 682940
rect 1200 682870 1270 682940
rect 1290 682870 1360 682940
rect 1380 682870 1450 682940
rect 1470 682870 1540 682940
rect 1560 682870 1630 682940
rect 120 682780 190 682850
rect 210 682780 280 682850
rect 300 682780 370 682850
rect 390 682780 460 682850
rect 480 682780 550 682850
rect 570 682780 640 682850
rect 660 682780 730 682850
rect 750 682780 820 682850
rect 840 682780 910 682850
rect 930 682780 1000 682850
rect 1020 682780 1090 682850
rect 1110 682780 1180 682850
rect 1200 682780 1270 682850
rect 1290 682780 1360 682850
rect 1380 682780 1450 682850
rect 1470 682780 1540 682850
rect 1560 682780 1630 682850
rect 120 682690 190 682760
rect 210 682690 280 682760
rect 300 682690 370 682760
rect 390 682690 460 682760
rect 480 682690 550 682760
rect 570 682690 640 682760
rect 660 682690 730 682760
rect 750 682690 820 682760
rect 840 682690 910 682760
rect 930 682690 1000 682760
rect 1020 682690 1090 682760
rect 1110 682690 1180 682760
rect 1200 682690 1270 682760
rect 1290 682690 1360 682760
rect 1380 682690 1450 682760
rect 1470 682690 1540 682760
rect 1560 682690 1630 682760
rect 120 682600 190 682670
rect 210 682600 280 682670
rect 300 682600 370 682670
rect 390 682600 460 682670
rect 480 682600 550 682670
rect 570 682600 640 682670
rect 660 682600 730 682670
rect 750 682600 820 682670
rect 840 682600 910 682670
rect 930 682600 1000 682670
rect 1020 682600 1090 682670
rect 1110 682600 1180 682670
rect 1200 682600 1270 682670
rect 1290 682600 1360 682670
rect 1380 682600 1450 682670
rect 1470 682600 1540 682670
rect 1560 682600 1630 682670
rect 120 682510 190 682580
rect 210 682510 280 682580
rect 300 682510 370 682580
rect 390 682510 460 682580
rect 480 682510 550 682580
rect 570 682510 640 682580
rect 660 682510 730 682580
rect 750 682510 820 682580
rect 840 682510 910 682580
rect 930 682510 1000 682580
rect 1020 682510 1090 682580
rect 1110 682510 1180 682580
rect 1200 682510 1270 682580
rect 1290 682510 1360 682580
rect 1380 682510 1450 682580
rect 1470 682510 1540 682580
rect 1560 682510 1630 682580
rect 120 682420 190 682490
rect 210 682420 280 682490
rect 300 682420 370 682490
rect 390 682420 460 682490
rect 480 682420 550 682490
rect 570 682420 640 682490
rect 660 682420 730 682490
rect 750 682420 820 682490
rect 840 682420 910 682490
rect 930 682420 1000 682490
rect 1020 682420 1090 682490
rect 1110 682420 1180 682490
rect 1200 682420 1270 682490
rect 1290 682420 1360 682490
rect 1380 682420 1450 682490
rect 1470 682420 1540 682490
rect 1560 682420 1630 682490
rect 120 682330 190 682400
rect 210 682330 280 682400
rect 300 682330 370 682400
rect 390 682330 460 682400
rect 480 682330 550 682400
rect 570 682330 640 682400
rect 660 682330 730 682400
rect 750 682330 820 682400
rect 840 682330 910 682400
rect 930 682330 1000 682400
rect 1020 682330 1090 682400
rect 1110 682330 1180 682400
rect 1200 682330 1270 682400
rect 1290 682330 1360 682400
rect 1380 682330 1450 682400
rect 1470 682330 1540 682400
rect 1560 682330 1630 682400
rect 120 682240 190 682310
rect 210 682240 280 682310
rect 300 682240 370 682310
rect 390 682240 460 682310
rect 480 682240 550 682310
rect 570 682240 640 682310
rect 660 682240 730 682310
rect 750 682240 820 682310
rect 840 682240 910 682310
rect 930 682240 1000 682310
rect 1020 682240 1090 682310
rect 1110 682240 1180 682310
rect 1200 682240 1270 682310
rect 1290 682240 1360 682310
rect 1380 682240 1450 682310
rect 1470 682240 1540 682310
rect 1560 682240 1630 682310
rect 120 682150 190 682220
rect 210 682150 280 682220
rect 300 682150 370 682220
rect 390 682150 460 682220
rect 480 682150 550 682220
rect 570 682150 640 682220
rect 660 682150 730 682220
rect 750 682150 820 682220
rect 840 682150 910 682220
rect 930 682150 1000 682220
rect 1020 682150 1090 682220
rect 1110 682150 1180 682220
rect 1200 682150 1270 682220
rect 1290 682150 1360 682220
rect 1380 682150 1450 682220
rect 1470 682150 1540 682220
rect 1560 682150 1630 682220
rect 17670 683590 17740 683660
rect 17760 683590 17830 683660
rect 17850 683590 17920 683660
rect 17940 683590 18010 683660
rect 18030 683590 18100 683660
rect 18120 683590 18190 683660
rect 18210 683590 18280 683660
rect 18300 683590 18370 683660
rect 18390 683590 18460 683660
rect 18480 683590 18550 683660
rect 18570 683590 18640 683660
rect 18660 683590 18730 683660
rect 18750 683590 18820 683660
rect 18840 683590 18910 683660
rect 18930 683590 19000 683660
rect 19020 683590 19090 683660
rect 19110 683590 19180 683660
rect 19200 683590 19270 683660
rect 19290 683590 19360 683660
rect 19380 683590 19450 683660
rect 19470 683590 19540 683660
rect 19560 683590 19630 683660
rect 17670 683500 17740 683570
rect 17760 683500 17830 683570
rect 17850 683500 17920 683570
rect 17940 683500 18010 683570
rect 18030 683500 18100 683570
rect 18120 683500 18190 683570
rect 18210 683500 18280 683570
rect 18300 683500 18370 683570
rect 18390 683500 18460 683570
rect 18480 683500 18550 683570
rect 18570 683500 18640 683570
rect 18660 683500 18730 683570
rect 18750 683500 18820 683570
rect 18840 683500 18910 683570
rect 18930 683500 19000 683570
rect 19020 683500 19090 683570
rect 19110 683500 19180 683570
rect 19200 683500 19270 683570
rect 19290 683500 19360 683570
rect 19380 683500 19450 683570
rect 19470 683500 19540 683570
rect 19560 683500 19630 683570
rect 17670 683410 17740 683480
rect 17760 683410 17830 683480
rect 17850 683410 17920 683480
rect 17940 683410 18010 683480
rect 18030 683410 18100 683480
rect 18120 683410 18190 683480
rect 18210 683410 18280 683480
rect 18300 683410 18370 683480
rect 18390 683410 18460 683480
rect 18480 683410 18550 683480
rect 18570 683410 18640 683480
rect 18660 683410 18730 683480
rect 18750 683410 18820 683480
rect 18840 683410 18910 683480
rect 18930 683410 19000 683480
rect 19020 683410 19090 683480
rect 19110 683410 19180 683480
rect 19200 683410 19270 683480
rect 19290 683410 19360 683480
rect 19380 683410 19450 683480
rect 19470 683410 19540 683480
rect 19560 683410 19630 683480
rect 17670 683320 17740 683390
rect 17760 683320 17830 683390
rect 17850 683320 17920 683390
rect 17940 683320 18010 683390
rect 18030 683320 18100 683390
rect 18120 683320 18190 683390
rect 18210 683320 18280 683390
rect 18300 683320 18370 683390
rect 18390 683320 18460 683390
rect 18480 683320 18550 683390
rect 18570 683320 18640 683390
rect 18660 683320 18730 683390
rect 18750 683320 18820 683390
rect 18840 683320 18910 683390
rect 18930 683320 19000 683390
rect 19020 683320 19090 683390
rect 19110 683320 19180 683390
rect 19200 683320 19270 683390
rect 19290 683320 19360 683390
rect 19380 683320 19450 683390
rect 19470 683320 19540 683390
rect 19560 683320 19630 683390
rect 17670 683230 17740 683300
rect 17760 683230 17830 683300
rect 17850 683230 17920 683300
rect 17940 683230 18010 683300
rect 18030 683230 18100 683300
rect 18120 683230 18190 683300
rect 18210 683230 18280 683300
rect 18300 683230 18370 683300
rect 18390 683230 18460 683300
rect 18480 683230 18550 683300
rect 18570 683230 18640 683300
rect 18660 683230 18730 683300
rect 18750 683230 18820 683300
rect 18840 683230 18910 683300
rect 18930 683230 19000 683300
rect 19020 683230 19090 683300
rect 19110 683230 19180 683300
rect 19200 683230 19270 683300
rect 19290 683230 19360 683300
rect 19380 683230 19450 683300
rect 19470 683230 19540 683300
rect 19560 683230 19630 683300
rect 17670 683140 17740 683210
rect 17760 683140 17830 683210
rect 17850 683140 17920 683210
rect 17940 683140 18010 683210
rect 18030 683140 18100 683210
rect 18120 683140 18190 683210
rect 18210 683140 18280 683210
rect 18300 683140 18370 683210
rect 18390 683140 18460 683210
rect 18480 683140 18550 683210
rect 18570 683140 18640 683210
rect 18660 683140 18730 683210
rect 18750 683140 18820 683210
rect 18840 683140 18910 683210
rect 18930 683140 19000 683210
rect 19020 683140 19090 683210
rect 19110 683140 19180 683210
rect 19200 683140 19270 683210
rect 19290 683140 19360 683210
rect 19380 683140 19450 683210
rect 19470 683140 19540 683210
rect 19560 683140 19630 683210
rect 17670 683050 17740 683120
rect 17760 683050 17830 683120
rect 17850 683050 17920 683120
rect 17940 683050 18010 683120
rect 18030 683050 18100 683120
rect 18120 683050 18190 683120
rect 18210 683050 18280 683120
rect 18300 683050 18370 683120
rect 18390 683050 18460 683120
rect 18480 683050 18550 683120
rect 18570 683050 18640 683120
rect 18660 683050 18730 683120
rect 18750 683050 18820 683120
rect 18840 683050 18910 683120
rect 18930 683050 19000 683120
rect 19020 683050 19090 683120
rect 19110 683050 19180 683120
rect 19200 683050 19270 683120
rect 19290 683050 19360 683120
rect 19380 683050 19450 683120
rect 19470 683050 19540 683120
rect 19560 683050 19630 683120
rect 17670 682960 17740 683030
rect 17760 682960 17830 683030
rect 17850 682960 17920 683030
rect 17940 682960 18010 683030
rect 18030 682960 18100 683030
rect 18120 682960 18190 683030
rect 18210 682960 18280 683030
rect 18300 682960 18370 683030
rect 18390 682960 18460 683030
rect 18480 682960 18550 683030
rect 18570 682960 18640 683030
rect 18660 682960 18730 683030
rect 18750 682960 18820 683030
rect 18840 682960 18910 683030
rect 18930 682960 19000 683030
rect 19020 682960 19090 683030
rect 19110 682960 19180 683030
rect 19200 682960 19270 683030
rect 19290 682960 19360 683030
rect 19380 682960 19450 683030
rect 19470 682960 19540 683030
rect 19560 682960 19630 683030
rect 17670 682870 17740 682940
rect 17760 682870 17830 682940
rect 17850 682870 17920 682940
rect 17940 682870 18010 682940
rect 18030 682870 18100 682940
rect 18120 682870 18190 682940
rect 18210 682870 18280 682940
rect 18300 682870 18370 682940
rect 18390 682870 18460 682940
rect 18480 682870 18550 682940
rect 18570 682870 18640 682940
rect 18660 682870 18730 682940
rect 18750 682870 18820 682940
rect 18840 682870 18910 682940
rect 18930 682870 19000 682940
rect 19020 682870 19090 682940
rect 19110 682870 19180 682940
rect 19200 682870 19270 682940
rect 19290 682870 19360 682940
rect 19380 682870 19450 682940
rect 19470 682870 19540 682940
rect 19560 682870 19630 682940
rect 17670 682780 17740 682850
rect 17760 682780 17830 682850
rect 17850 682780 17920 682850
rect 17940 682780 18010 682850
rect 18030 682780 18100 682850
rect 18120 682780 18190 682850
rect 18210 682780 18280 682850
rect 18300 682780 18370 682850
rect 18390 682780 18460 682850
rect 18480 682780 18550 682850
rect 18570 682780 18640 682850
rect 18660 682780 18730 682850
rect 18750 682780 18820 682850
rect 18840 682780 18910 682850
rect 18930 682780 19000 682850
rect 19020 682780 19090 682850
rect 19110 682780 19180 682850
rect 19200 682780 19270 682850
rect 19290 682780 19360 682850
rect 19380 682780 19450 682850
rect 19470 682780 19540 682850
rect 19560 682780 19630 682850
rect 17670 682690 17740 682760
rect 17760 682690 17830 682760
rect 17850 682690 17920 682760
rect 17940 682690 18010 682760
rect 18030 682690 18100 682760
rect 18120 682690 18190 682760
rect 18210 682690 18280 682760
rect 18300 682690 18370 682760
rect 18390 682690 18460 682760
rect 18480 682690 18550 682760
rect 18570 682690 18640 682760
rect 18660 682690 18730 682760
rect 18750 682690 18820 682760
rect 18840 682690 18910 682760
rect 18930 682690 19000 682760
rect 19020 682690 19090 682760
rect 19110 682690 19180 682760
rect 19200 682690 19270 682760
rect 19290 682690 19360 682760
rect 19380 682690 19450 682760
rect 19470 682690 19540 682760
rect 19560 682690 19630 682760
rect 17670 682600 17740 682670
rect 17760 682600 17830 682670
rect 17850 682600 17920 682670
rect 17940 682600 18010 682670
rect 18030 682600 18100 682670
rect 18120 682600 18190 682670
rect 18210 682600 18280 682670
rect 18300 682600 18370 682670
rect 18390 682600 18460 682670
rect 18480 682600 18550 682670
rect 18570 682600 18640 682670
rect 18660 682600 18730 682670
rect 18750 682600 18820 682670
rect 18840 682600 18910 682670
rect 18930 682600 19000 682670
rect 19020 682600 19090 682670
rect 19110 682600 19180 682670
rect 19200 682600 19270 682670
rect 19290 682600 19360 682670
rect 19380 682600 19450 682670
rect 19470 682600 19540 682670
rect 19560 682600 19630 682670
rect 17670 682510 17740 682580
rect 17760 682510 17830 682580
rect 17850 682510 17920 682580
rect 17940 682510 18010 682580
rect 18030 682510 18100 682580
rect 18120 682510 18190 682580
rect 18210 682510 18280 682580
rect 18300 682510 18370 682580
rect 18390 682510 18460 682580
rect 18480 682510 18550 682580
rect 18570 682510 18640 682580
rect 18660 682510 18730 682580
rect 18750 682510 18820 682580
rect 18840 682510 18910 682580
rect 18930 682510 19000 682580
rect 19020 682510 19090 682580
rect 19110 682510 19180 682580
rect 19200 682510 19270 682580
rect 19290 682510 19360 682580
rect 19380 682510 19450 682580
rect 19470 682510 19540 682580
rect 19560 682510 19630 682580
rect 17670 682420 17740 682490
rect 17760 682420 17830 682490
rect 17850 682420 17920 682490
rect 17940 682420 18010 682490
rect 18030 682420 18100 682490
rect 18120 682420 18190 682490
rect 18210 682420 18280 682490
rect 18300 682420 18370 682490
rect 18390 682420 18460 682490
rect 18480 682420 18550 682490
rect 18570 682420 18640 682490
rect 18660 682420 18730 682490
rect 18750 682420 18820 682490
rect 18840 682420 18910 682490
rect 18930 682420 19000 682490
rect 19020 682420 19090 682490
rect 19110 682420 19180 682490
rect 19200 682420 19270 682490
rect 19290 682420 19360 682490
rect 19380 682420 19450 682490
rect 19470 682420 19540 682490
rect 19560 682420 19630 682490
rect 17670 682330 17740 682400
rect 17760 682330 17830 682400
rect 17850 682330 17920 682400
rect 17940 682330 18010 682400
rect 18030 682330 18100 682400
rect 18120 682330 18190 682400
rect 18210 682330 18280 682400
rect 18300 682330 18370 682400
rect 18390 682330 18460 682400
rect 18480 682330 18550 682400
rect 18570 682330 18640 682400
rect 18660 682330 18730 682400
rect 18750 682330 18820 682400
rect 18840 682330 18910 682400
rect 18930 682330 19000 682400
rect 19020 682330 19090 682400
rect 19110 682330 19180 682400
rect 19200 682330 19270 682400
rect 19290 682330 19360 682400
rect 19380 682330 19450 682400
rect 19470 682330 19540 682400
rect 19560 682330 19630 682400
rect 17670 682240 17740 682310
rect 17760 682240 17830 682310
rect 17850 682240 17920 682310
rect 17940 682240 18010 682310
rect 18030 682240 18100 682310
rect 18120 682240 18190 682310
rect 18210 682240 18280 682310
rect 18300 682240 18370 682310
rect 18390 682240 18460 682310
rect 18480 682240 18550 682310
rect 18570 682240 18640 682310
rect 18660 682240 18730 682310
rect 18750 682240 18820 682310
rect 18840 682240 18910 682310
rect 18930 682240 19000 682310
rect 19020 682240 19090 682310
rect 19110 682240 19180 682310
rect 19200 682240 19270 682310
rect 19290 682240 19360 682310
rect 19380 682240 19450 682310
rect 19470 682240 19540 682310
rect 19560 682240 19630 682310
rect 17670 682150 17740 682220
rect 17760 682150 17830 682220
rect 17850 682150 17920 682220
rect 17940 682150 18010 682220
rect 18030 682150 18100 682220
rect 18120 682150 18190 682220
rect 18210 682150 18280 682220
rect 18300 682150 18370 682220
rect 18390 682150 18460 682220
rect 18480 682150 18550 682220
rect 18570 682150 18640 682220
rect 18660 682150 18730 682220
rect 18750 682150 18820 682220
rect 18840 682150 18910 682220
rect 18930 682150 19000 682220
rect 19020 682150 19090 682220
rect 19110 682150 19180 682220
rect 19200 682150 19270 682220
rect 19290 682150 19360 682220
rect 19380 682150 19450 682220
rect 19470 682150 19540 682220
rect 19560 682150 19630 682220
rect 582320 679446 582390 679516
rect 582410 679446 582480 679516
rect 582500 679446 582570 679516
rect 582590 679446 582660 679516
rect 582680 679446 582750 679516
rect 582770 679446 582840 679516
rect 582320 679356 582390 679426
rect 582410 679356 582480 679426
rect 582500 679356 582570 679426
rect 582590 679356 582660 679426
rect 582680 679356 582750 679426
rect 582770 679356 582840 679426
rect 582320 679266 582390 679336
rect 582410 679266 582480 679336
rect 582500 679266 582570 679336
rect 582590 679266 582660 679336
rect 582680 679266 582750 679336
rect 582770 679266 582840 679336
rect 582320 679176 582390 679246
rect 582410 679176 582480 679246
rect 582500 679176 582570 679246
rect 582590 679176 582660 679246
rect 582680 679176 582750 679246
rect 582770 679176 582840 679246
rect 582320 679086 582390 679156
rect 582410 679086 582480 679156
rect 582500 679086 582570 679156
rect 582590 679086 582660 679156
rect 582680 679086 582750 679156
rect 582770 679086 582840 679156
rect 582320 678996 582390 679066
rect 582410 678996 582480 679066
rect 582500 678996 582570 679066
rect 582590 678996 582660 679066
rect 582680 678996 582750 679066
rect 582770 678996 582840 679066
rect 94280 638100 94350 638170
rect 94380 638100 94450 638170
rect 94480 638100 94550 638170
rect 94280 638010 94350 638080
rect 94380 638010 94450 638080
rect 94480 638010 94550 638080
rect 98838 638100 98908 638170
rect 98938 638100 99008 638170
rect 99038 638100 99108 638170
rect 98838 638010 98908 638080
rect 98938 638010 99008 638080
rect 99038 638010 99108 638080
rect 21966 623458 22036 623528
rect 22056 623458 22126 623528
rect 22146 623458 22216 623528
rect 22236 623458 22306 623528
rect 22326 623458 22396 623528
rect 22416 623458 22486 623528
rect 22506 623458 22576 623528
rect 22596 623458 22666 623528
rect 22686 623458 22756 623528
rect 22776 623458 22846 623528
rect 22866 623458 22936 623528
rect 22956 623458 23026 623528
rect 23046 623458 23116 623528
rect 23136 623458 23206 623528
rect 23226 623458 23296 623528
rect 23316 623458 23386 623528
rect 23406 623458 23476 623528
rect 23496 623458 23566 623528
rect 23586 623458 23656 623528
rect 23676 623458 23746 623528
rect 23766 623458 23836 623528
rect 23856 623458 23926 623528
rect 21966 623368 22036 623438
rect 22056 623368 22126 623438
rect 22146 623368 22216 623438
rect 22236 623368 22306 623438
rect 22326 623368 22396 623438
rect 22416 623368 22486 623438
rect 22506 623368 22576 623438
rect 22596 623368 22666 623438
rect 22686 623368 22756 623438
rect 22776 623368 22846 623438
rect 22866 623368 22936 623438
rect 22956 623368 23026 623438
rect 23046 623368 23116 623438
rect 23136 623368 23206 623438
rect 23226 623368 23296 623438
rect 23316 623368 23386 623438
rect 23406 623368 23476 623438
rect 23496 623368 23566 623438
rect 23586 623368 23656 623438
rect 23676 623368 23746 623438
rect 23766 623368 23836 623438
rect 23856 623368 23926 623438
rect 21966 623278 22036 623348
rect 22056 623278 22126 623348
rect 22146 623278 22216 623348
rect 22236 623278 22306 623348
rect 22326 623278 22396 623348
rect 22416 623278 22486 623348
rect 22506 623278 22576 623348
rect 22596 623278 22666 623348
rect 22686 623278 22756 623348
rect 22776 623278 22846 623348
rect 22866 623278 22936 623348
rect 22956 623278 23026 623348
rect 23046 623278 23116 623348
rect 23136 623278 23206 623348
rect 23226 623278 23296 623348
rect 23316 623278 23386 623348
rect 23406 623278 23476 623348
rect 23496 623278 23566 623348
rect 23586 623278 23656 623348
rect 23676 623278 23746 623348
rect 23766 623278 23836 623348
rect 23856 623278 23926 623348
rect 21966 623188 22036 623258
rect 22056 623188 22126 623258
rect 22146 623188 22216 623258
rect 22236 623188 22306 623258
rect 22326 623188 22396 623258
rect 22416 623188 22486 623258
rect 22506 623188 22576 623258
rect 22596 623188 22666 623258
rect 22686 623188 22756 623258
rect 22776 623188 22846 623258
rect 22866 623188 22936 623258
rect 22956 623188 23026 623258
rect 23046 623188 23116 623258
rect 23136 623188 23206 623258
rect 23226 623188 23296 623258
rect 23316 623188 23386 623258
rect 23406 623188 23476 623258
rect 23496 623188 23566 623258
rect 23586 623188 23656 623258
rect 23676 623188 23746 623258
rect 23766 623188 23836 623258
rect 23856 623188 23926 623258
rect 21966 623098 22036 623168
rect 22056 623098 22126 623168
rect 22146 623098 22216 623168
rect 22236 623098 22306 623168
rect 22326 623098 22396 623168
rect 22416 623098 22486 623168
rect 22506 623098 22576 623168
rect 22596 623098 22666 623168
rect 22686 623098 22756 623168
rect 22776 623098 22846 623168
rect 22866 623098 22936 623168
rect 22956 623098 23026 623168
rect 23046 623098 23116 623168
rect 23136 623098 23206 623168
rect 23226 623098 23296 623168
rect 23316 623098 23386 623168
rect 23406 623098 23476 623168
rect 23496 623098 23566 623168
rect 23586 623098 23656 623168
rect 23676 623098 23746 623168
rect 23766 623098 23836 623168
rect 23856 623098 23926 623168
rect 21966 623008 22036 623078
rect 22056 623008 22126 623078
rect 22146 623008 22216 623078
rect 22236 623008 22306 623078
rect 22326 623008 22396 623078
rect 22416 623008 22486 623078
rect 22506 623008 22576 623078
rect 22596 623008 22666 623078
rect 22686 623008 22756 623078
rect 22776 623008 22846 623078
rect 22866 623008 22936 623078
rect 22956 623008 23026 623078
rect 23046 623008 23116 623078
rect 23136 623008 23206 623078
rect 23226 623008 23296 623078
rect 23316 623008 23386 623078
rect 23406 623008 23476 623078
rect 23496 623008 23566 623078
rect 23586 623008 23656 623078
rect 23676 623008 23746 623078
rect 23766 623008 23836 623078
rect 23856 623008 23926 623078
rect 21966 622918 22036 622988
rect 22056 622918 22126 622988
rect 22146 622918 22216 622988
rect 22236 622918 22306 622988
rect 22326 622918 22396 622988
rect 22416 622918 22486 622988
rect 22506 622918 22576 622988
rect 22596 622918 22666 622988
rect 22686 622918 22756 622988
rect 22776 622918 22846 622988
rect 22866 622918 22936 622988
rect 22956 622918 23026 622988
rect 23046 622918 23116 622988
rect 23136 622918 23206 622988
rect 23226 622918 23296 622988
rect 23316 622918 23386 622988
rect 23406 622918 23476 622988
rect 23496 622918 23566 622988
rect 23586 622918 23656 622988
rect 23676 622918 23746 622988
rect 23766 622918 23836 622988
rect 23856 622918 23926 622988
rect 21966 622828 22036 622898
rect 22056 622828 22126 622898
rect 22146 622828 22216 622898
rect 22236 622828 22306 622898
rect 22326 622828 22396 622898
rect 22416 622828 22486 622898
rect 22506 622828 22576 622898
rect 22596 622828 22666 622898
rect 22686 622828 22756 622898
rect 22776 622828 22846 622898
rect 22866 622828 22936 622898
rect 22956 622828 23026 622898
rect 23046 622828 23116 622898
rect 23136 622828 23206 622898
rect 23226 622828 23296 622898
rect 23316 622828 23386 622898
rect 23406 622828 23476 622898
rect 23496 622828 23566 622898
rect 23586 622828 23656 622898
rect 23676 622828 23746 622898
rect 23766 622828 23836 622898
rect 23856 622828 23926 622898
rect 21966 622738 22036 622808
rect 22056 622738 22126 622808
rect 22146 622738 22216 622808
rect 22236 622738 22306 622808
rect 22326 622738 22396 622808
rect 22416 622738 22486 622808
rect 22506 622738 22576 622808
rect 22596 622738 22666 622808
rect 22686 622738 22756 622808
rect 22776 622738 22846 622808
rect 22866 622738 22936 622808
rect 22956 622738 23026 622808
rect 23046 622738 23116 622808
rect 23136 622738 23206 622808
rect 23226 622738 23296 622808
rect 23316 622738 23386 622808
rect 23406 622738 23476 622808
rect 23496 622738 23566 622808
rect 23586 622738 23656 622808
rect 23676 622738 23746 622808
rect 23766 622738 23836 622808
rect 23856 622738 23926 622808
rect 21966 622648 22036 622718
rect 22056 622648 22126 622718
rect 22146 622648 22216 622718
rect 22236 622648 22306 622718
rect 22326 622648 22396 622718
rect 22416 622648 22486 622718
rect 22506 622648 22576 622718
rect 22596 622648 22666 622718
rect 22686 622648 22756 622718
rect 22776 622648 22846 622718
rect 22866 622648 22936 622718
rect 22956 622648 23026 622718
rect 23046 622648 23116 622718
rect 23136 622648 23206 622718
rect 23226 622648 23296 622718
rect 23316 622648 23386 622718
rect 23406 622648 23476 622718
rect 23496 622648 23566 622718
rect 23586 622648 23656 622718
rect 23676 622648 23746 622718
rect 23766 622648 23836 622718
rect 23856 622648 23926 622718
rect 21966 622558 22036 622628
rect 22056 622558 22126 622628
rect 22146 622558 22216 622628
rect 22236 622558 22306 622628
rect 22326 622558 22396 622628
rect 22416 622558 22486 622628
rect 22506 622558 22576 622628
rect 22596 622558 22666 622628
rect 22686 622558 22756 622628
rect 22776 622558 22846 622628
rect 22866 622558 22936 622628
rect 22956 622558 23026 622628
rect 23046 622558 23116 622628
rect 23136 622558 23206 622628
rect 23226 622558 23296 622628
rect 23316 622558 23386 622628
rect 23406 622558 23476 622628
rect 23496 622558 23566 622628
rect 23586 622558 23656 622628
rect 23676 622558 23746 622628
rect 23766 622558 23836 622628
rect 23856 622558 23926 622628
rect 21966 622468 22036 622538
rect 22056 622468 22126 622538
rect 22146 622468 22216 622538
rect 22236 622468 22306 622538
rect 22326 622468 22396 622538
rect 22416 622468 22486 622538
rect 22506 622468 22576 622538
rect 22596 622468 22666 622538
rect 22686 622468 22756 622538
rect 22776 622468 22846 622538
rect 22866 622468 22936 622538
rect 22956 622468 23026 622538
rect 23046 622468 23116 622538
rect 23136 622468 23206 622538
rect 23226 622468 23296 622538
rect 23316 622468 23386 622538
rect 23406 622468 23476 622538
rect 23496 622468 23566 622538
rect 23586 622468 23656 622538
rect 23676 622468 23746 622538
rect 23766 622468 23836 622538
rect 23856 622468 23926 622538
rect 21966 622378 22036 622448
rect 22056 622378 22126 622448
rect 22146 622378 22216 622448
rect 22236 622378 22306 622448
rect 22326 622378 22396 622448
rect 22416 622378 22486 622448
rect 22506 622378 22576 622448
rect 22596 622378 22666 622448
rect 22686 622378 22756 622448
rect 22776 622378 22846 622448
rect 22866 622378 22936 622448
rect 22956 622378 23026 622448
rect 23046 622378 23116 622448
rect 23136 622378 23206 622448
rect 23226 622378 23296 622448
rect 23316 622378 23386 622448
rect 23406 622378 23476 622448
rect 23496 622378 23566 622448
rect 23586 622378 23656 622448
rect 23676 622378 23746 622448
rect 23766 622378 23836 622448
rect 23856 622378 23926 622448
rect 21966 622288 22036 622358
rect 22056 622288 22126 622358
rect 22146 622288 22216 622358
rect 22236 622288 22306 622358
rect 22326 622288 22396 622358
rect 22416 622288 22486 622358
rect 22506 622288 22576 622358
rect 22596 622288 22666 622358
rect 22686 622288 22756 622358
rect 22776 622288 22846 622358
rect 22866 622288 22936 622358
rect 22956 622288 23026 622358
rect 23046 622288 23116 622358
rect 23136 622288 23206 622358
rect 23226 622288 23296 622358
rect 23316 622288 23386 622358
rect 23406 622288 23476 622358
rect 23496 622288 23566 622358
rect 23586 622288 23656 622358
rect 23676 622288 23746 622358
rect 23766 622288 23836 622358
rect 23856 622288 23926 622358
rect 21966 622198 22036 622268
rect 22056 622198 22126 622268
rect 22146 622198 22216 622268
rect 22236 622198 22306 622268
rect 22326 622198 22396 622268
rect 22416 622198 22486 622268
rect 22506 622198 22576 622268
rect 22596 622198 22666 622268
rect 22686 622198 22756 622268
rect 22776 622198 22846 622268
rect 22866 622198 22936 622268
rect 22956 622198 23026 622268
rect 23046 622198 23116 622268
rect 23136 622198 23206 622268
rect 23226 622198 23296 622268
rect 23316 622198 23386 622268
rect 23406 622198 23476 622268
rect 23496 622198 23566 622268
rect 23586 622198 23656 622268
rect 23676 622198 23746 622268
rect 23766 622198 23836 622268
rect 23856 622198 23926 622268
rect 21966 622108 22036 622178
rect 22056 622108 22126 622178
rect 22146 622108 22216 622178
rect 22236 622108 22306 622178
rect 22326 622108 22396 622178
rect 22416 622108 22486 622178
rect 22506 622108 22576 622178
rect 22596 622108 22666 622178
rect 22686 622108 22756 622178
rect 22776 622108 22846 622178
rect 22866 622108 22936 622178
rect 22956 622108 23026 622178
rect 23046 622108 23116 622178
rect 23136 622108 23206 622178
rect 23226 622108 23296 622178
rect 23316 622108 23386 622178
rect 23406 622108 23476 622178
rect 23496 622108 23566 622178
rect 23586 622108 23656 622178
rect 23676 622108 23746 622178
rect 23766 622108 23836 622178
rect 23856 622108 23926 622178
rect 21966 622018 22036 622088
rect 22056 622018 22126 622088
rect 22146 622018 22216 622088
rect 22236 622018 22306 622088
rect 22326 622018 22396 622088
rect 22416 622018 22486 622088
rect 22506 622018 22576 622088
rect 22596 622018 22666 622088
rect 22686 622018 22756 622088
rect 22776 622018 22846 622088
rect 22866 622018 22936 622088
rect 22956 622018 23026 622088
rect 23046 622018 23116 622088
rect 23136 622018 23206 622088
rect 23226 622018 23296 622088
rect 23316 622018 23386 622088
rect 23406 622018 23476 622088
rect 23496 622018 23566 622088
rect 23586 622018 23656 622088
rect 23676 622018 23746 622088
rect 23766 622018 23836 622088
rect 23856 622018 23926 622088
rect 21966 621928 22036 621998
rect 22056 621928 22126 621998
rect 22146 621928 22216 621998
rect 22236 621928 22306 621998
rect 22326 621928 22396 621998
rect 22416 621928 22486 621998
rect 22506 621928 22576 621998
rect 22596 621928 22666 621998
rect 22686 621928 22756 621998
rect 22776 621928 22846 621998
rect 22866 621928 22936 621998
rect 22956 621928 23026 621998
rect 23046 621928 23116 621998
rect 23136 621928 23206 621998
rect 23226 621928 23296 621998
rect 23316 621928 23386 621998
rect 23406 621928 23476 621998
rect 23496 621928 23566 621998
rect 23586 621928 23656 621998
rect 23676 621928 23746 621998
rect 23766 621928 23836 621998
rect 23856 621928 23926 621998
rect 21966 621838 22036 621908
rect 22056 621838 22126 621908
rect 22146 621838 22216 621908
rect 22236 621838 22306 621908
rect 22326 621838 22396 621908
rect 22416 621838 22486 621908
rect 22506 621838 22576 621908
rect 22596 621838 22666 621908
rect 22686 621838 22756 621908
rect 22776 621838 22846 621908
rect 22866 621838 22936 621908
rect 22956 621838 23026 621908
rect 23046 621838 23116 621908
rect 23136 621838 23206 621908
rect 23226 621838 23296 621908
rect 23316 621838 23386 621908
rect 23406 621838 23476 621908
rect 23496 621838 23566 621908
rect 23586 621838 23656 621908
rect 23676 621838 23746 621908
rect 23766 621838 23836 621908
rect 23856 621838 23926 621908
rect 21966 621748 22036 621818
rect 22056 621748 22126 621818
rect 22146 621748 22216 621818
rect 22236 621748 22306 621818
rect 22326 621748 22396 621818
rect 22416 621748 22486 621818
rect 22506 621748 22576 621818
rect 22596 621748 22666 621818
rect 22686 621748 22756 621818
rect 22776 621748 22846 621818
rect 22866 621748 22936 621818
rect 22956 621748 23026 621818
rect 23046 621748 23116 621818
rect 23136 621748 23206 621818
rect 23226 621748 23296 621818
rect 23316 621748 23386 621818
rect 23406 621748 23476 621818
rect 23496 621748 23566 621818
rect 23586 621748 23656 621818
rect 23676 621748 23746 621818
rect 23766 621748 23836 621818
rect 23856 621748 23926 621818
rect 21966 621658 22036 621728
rect 22056 621658 22126 621728
rect 22146 621658 22216 621728
rect 22236 621658 22306 621728
rect 22326 621658 22396 621728
rect 22416 621658 22486 621728
rect 22506 621658 22576 621728
rect 22596 621658 22666 621728
rect 22686 621658 22756 621728
rect 22776 621658 22846 621728
rect 22866 621658 22936 621728
rect 22956 621658 23026 621728
rect 23046 621658 23116 621728
rect 23136 621658 23206 621728
rect 23226 621658 23296 621728
rect 23316 621658 23386 621728
rect 23406 621658 23476 621728
rect 23496 621658 23566 621728
rect 23586 621658 23656 621728
rect 23676 621658 23746 621728
rect 23766 621658 23836 621728
rect 23856 621658 23926 621728
rect 21966 621568 22036 621638
rect 22056 621568 22126 621638
rect 22146 621568 22216 621638
rect 22236 621568 22306 621638
rect 22326 621568 22396 621638
rect 22416 621568 22486 621638
rect 22506 621568 22576 621638
rect 22596 621568 22666 621638
rect 22686 621568 22756 621638
rect 22776 621568 22846 621638
rect 22866 621568 22936 621638
rect 22956 621568 23026 621638
rect 23046 621568 23116 621638
rect 23136 621568 23206 621638
rect 23226 621568 23296 621638
rect 23316 621568 23386 621638
rect 23406 621568 23476 621638
rect 23496 621568 23566 621638
rect 23586 621568 23656 621638
rect 23676 621568 23746 621638
rect 23766 621568 23836 621638
rect 23856 621568 23926 621638
rect 17670 619350 17740 619420
rect 17760 619350 17830 619420
rect 17850 619350 17920 619420
rect 17940 619350 18010 619420
rect 18030 619350 18100 619420
rect 18120 619350 18190 619420
rect 18210 619350 18280 619420
rect 18300 619350 18370 619420
rect 18390 619350 18460 619420
rect 18480 619350 18550 619420
rect 18570 619350 18640 619420
rect 18660 619350 18730 619420
rect 18750 619350 18820 619420
rect 18840 619350 18910 619420
rect 18930 619350 19000 619420
rect 19020 619350 19090 619420
rect 19110 619350 19180 619420
rect 19200 619350 19270 619420
rect 19290 619350 19360 619420
rect 19380 619350 19450 619420
rect 19470 619350 19540 619420
rect 19560 619350 19630 619420
rect 17670 619260 17740 619330
rect 17760 619260 17830 619330
rect 17850 619260 17920 619330
rect 17940 619260 18010 619330
rect 18030 619260 18100 619330
rect 18120 619260 18190 619330
rect 18210 619260 18280 619330
rect 18300 619260 18370 619330
rect 18390 619260 18460 619330
rect 18480 619260 18550 619330
rect 18570 619260 18640 619330
rect 18660 619260 18730 619330
rect 18750 619260 18820 619330
rect 18840 619260 18910 619330
rect 18930 619260 19000 619330
rect 19020 619260 19090 619330
rect 19110 619260 19180 619330
rect 19200 619260 19270 619330
rect 19290 619260 19360 619330
rect 19380 619260 19450 619330
rect 19470 619260 19540 619330
rect 19560 619260 19630 619330
rect 17670 619170 17740 619240
rect 17760 619170 17830 619240
rect 17850 619170 17920 619240
rect 17940 619170 18010 619240
rect 18030 619170 18100 619240
rect 18120 619170 18190 619240
rect 18210 619170 18280 619240
rect 18300 619170 18370 619240
rect 18390 619170 18460 619240
rect 18480 619170 18550 619240
rect 18570 619170 18640 619240
rect 18660 619170 18730 619240
rect 18750 619170 18820 619240
rect 18840 619170 18910 619240
rect 18930 619170 19000 619240
rect 19020 619170 19090 619240
rect 19110 619170 19180 619240
rect 19200 619170 19270 619240
rect 19290 619170 19360 619240
rect 19380 619170 19450 619240
rect 19470 619170 19540 619240
rect 19560 619170 19630 619240
rect 17670 619080 17740 619150
rect 17760 619080 17830 619150
rect 17850 619080 17920 619150
rect 17940 619080 18010 619150
rect 18030 619080 18100 619150
rect 18120 619080 18190 619150
rect 18210 619080 18280 619150
rect 18300 619080 18370 619150
rect 18390 619080 18460 619150
rect 18480 619080 18550 619150
rect 18570 619080 18640 619150
rect 18660 619080 18730 619150
rect 18750 619080 18820 619150
rect 18840 619080 18910 619150
rect 18930 619080 19000 619150
rect 19020 619080 19090 619150
rect 19110 619080 19180 619150
rect 19200 619080 19270 619150
rect 19290 619080 19360 619150
rect 19380 619080 19450 619150
rect 19470 619080 19540 619150
rect 19560 619080 19630 619150
rect 17670 618990 17740 619060
rect 17760 618990 17830 619060
rect 17850 618990 17920 619060
rect 17940 618990 18010 619060
rect 18030 618990 18100 619060
rect 18120 618990 18190 619060
rect 18210 618990 18280 619060
rect 18300 618990 18370 619060
rect 18390 618990 18460 619060
rect 18480 618990 18550 619060
rect 18570 618990 18640 619060
rect 18660 618990 18730 619060
rect 18750 618990 18820 619060
rect 18840 618990 18910 619060
rect 18930 618990 19000 619060
rect 19020 618990 19090 619060
rect 19110 618990 19180 619060
rect 19200 618990 19270 619060
rect 19290 618990 19360 619060
rect 19380 618990 19450 619060
rect 19470 618990 19540 619060
rect 19560 618990 19630 619060
rect 17670 618900 17740 618970
rect 17760 618900 17830 618970
rect 17850 618900 17920 618970
rect 17940 618900 18010 618970
rect 18030 618900 18100 618970
rect 18120 618900 18190 618970
rect 18210 618900 18280 618970
rect 18300 618900 18370 618970
rect 18390 618900 18460 618970
rect 18480 618900 18550 618970
rect 18570 618900 18640 618970
rect 18660 618900 18730 618970
rect 18750 618900 18820 618970
rect 18840 618900 18910 618970
rect 18930 618900 19000 618970
rect 19020 618900 19090 618970
rect 19110 618900 19180 618970
rect 19200 618900 19270 618970
rect 19290 618900 19360 618970
rect 19380 618900 19450 618970
rect 19470 618900 19540 618970
rect 19560 618900 19630 618970
rect 17670 618810 17740 618880
rect 17760 618810 17830 618880
rect 17850 618810 17920 618880
rect 17940 618810 18010 618880
rect 18030 618810 18100 618880
rect 18120 618810 18190 618880
rect 18210 618810 18280 618880
rect 18300 618810 18370 618880
rect 18390 618810 18460 618880
rect 18480 618810 18550 618880
rect 18570 618810 18640 618880
rect 18660 618810 18730 618880
rect 18750 618810 18820 618880
rect 18840 618810 18910 618880
rect 18930 618810 19000 618880
rect 19020 618810 19090 618880
rect 19110 618810 19180 618880
rect 19200 618810 19270 618880
rect 19290 618810 19360 618880
rect 19380 618810 19450 618880
rect 19470 618810 19540 618880
rect 19560 618810 19630 618880
rect 17670 618720 17740 618790
rect 17760 618720 17830 618790
rect 17850 618720 17920 618790
rect 17940 618720 18010 618790
rect 18030 618720 18100 618790
rect 18120 618720 18190 618790
rect 18210 618720 18280 618790
rect 18300 618720 18370 618790
rect 18390 618720 18460 618790
rect 18480 618720 18550 618790
rect 18570 618720 18640 618790
rect 18660 618720 18730 618790
rect 18750 618720 18820 618790
rect 18840 618720 18910 618790
rect 18930 618720 19000 618790
rect 19020 618720 19090 618790
rect 19110 618720 19180 618790
rect 19200 618720 19270 618790
rect 19290 618720 19360 618790
rect 19380 618720 19450 618790
rect 19470 618720 19540 618790
rect 19560 618720 19630 618790
rect 17670 618630 17740 618700
rect 17760 618630 17830 618700
rect 17850 618630 17920 618700
rect 17940 618630 18010 618700
rect 18030 618630 18100 618700
rect 18120 618630 18190 618700
rect 18210 618630 18280 618700
rect 18300 618630 18370 618700
rect 18390 618630 18460 618700
rect 18480 618630 18550 618700
rect 18570 618630 18640 618700
rect 18660 618630 18730 618700
rect 18750 618630 18820 618700
rect 18840 618630 18910 618700
rect 18930 618630 19000 618700
rect 19020 618630 19090 618700
rect 19110 618630 19180 618700
rect 19200 618630 19270 618700
rect 19290 618630 19360 618700
rect 19380 618630 19450 618700
rect 19470 618630 19540 618700
rect 19560 618630 19630 618700
rect 17670 618540 17740 618610
rect 17760 618540 17830 618610
rect 17850 618540 17920 618610
rect 17940 618540 18010 618610
rect 18030 618540 18100 618610
rect 18120 618540 18190 618610
rect 18210 618540 18280 618610
rect 18300 618540 18370 618610
rect 18390 618540 18460 618610
rect 18480 618540 18550 618610
rect 18570 618540 18640 618610
rect 18660 618540 18730 618610
rect 18750 618540 18820 618610
rect 18840 618540 18910 618610
rect 18930 618540 19000 618610
rect 19020 618540 19090 618610
rect 19110 618540 19180 618610
rect 19200 618540 19270 618610
rect 19290 618540 19360 618610
rect 19380 618540 19450 618610
rect 19470 618540 19540 618610
rect 19560 618540 19630 618610
rect 17670 618450 17740 618520
rect 17760 618450 17830 618520
rect 17850 618450 17920 618520
rect 17940 618450 18010 618520
rect 18030 618450 18100 618520
rect 18120 618450 18190 618520
rect 18210 618450 18280 618520
rect 18300 618450 18370 618520
rect 18390 618450 18460 618520
rect 18480 618450 18550 618520
rect 18570 618450 18640 618520
rect 18660 618450 18730 618520
rect 18750 618450 18820 618520
rect 18840 618450 18910 618520
rect 18930 618450 19000 618520
rect 19020 618450 19090 618520
rect 19110 618450 19180 618520
rect 19200 618450 19270 618520
rect 19290 618450 19360 618520
rect 19380 618450 19450 618520
rect 19470 618450 19540 618520
rect 19560 618450 19630 618520
rect 17670 618360 17740 618430
rect 17760 618360 17830 618430
rect 17850 618360 17920 618430
rect 17940 618360 18010 618430
rect 18030 618360 18100 618430
rect 18120 618360 18190 618430
rect 18210 618360 18280 618430
rect 18300 618360 18370 618430
rect 18390 618360 18460 618430
rect 18480 618360 18550 618430
rect 18570 618360 18640 618430
rect 18660 618360 18730 618430
rect 18750 618360 18820 618430
rect 18840 618360 18910 618430
rect 18930 618360 19000 618430
rect 19020 618360 19090 618430
rect 19110 618360 19180 618430
rect 19200 618360 19270 618430
rect 19290 618360 19360 618430
rect 19380 618360 19450 618430
rect 19470 618360 19540 618430
rect 19560 618360 19630 618430
rect 17670 618270 17740 618340
rect 17760 618270 17830 618340
rect 17850 618270 17920 618340
rect 17940 618270 18010 618340
rect 18030 618270 18100 618340
rect 18120 618270 18190 618340
rect 18210 618270 18280 618340
rect 18300 618270 18370 618340
rect 18390 618270 18460 618340
rect 18480 618270 18550 618340
rect 18570 618270 18640 618340
rect 18660 618270 18730 618340
rect 18750 618270 18820 618340
rect 18840 618270 18910 618340
rect 18930 618270 19000 618340
rect 19020 618270 19090 618340
rect 19110 618270 19180 618340
rect 19200 618270 19270 618340
rect 19290 618270 19360 618340
rect 19380 618270 19450 618340
rect 19470 618270 19540 618340
rect 19560 618270 19630 618340
rect 17670 618180 17740 618250
rect 17760 618180 17830 618250
rect 17850 618180 17920 618250
rect 17940 618180 18010 618250
rect 18030 618180 18100 618250
rect 18120 618180 18190 618250
rect 18210 618180 18280 618250
rect 18300 618180 18370 618250
rect 18390 618180 18460 618250
rect 18480 618180 18550 618250
rect 18570 618180 18640 618250
rect 18660 618180 18730 618250
rect 18750 618180 18820 618250
rect 18840 618180 18910 618250
rect 18930 618180 19000 618250
rect 19020 618180 19090 618250
rect 19110 618180 19180 618250
rect 19200 618180 19270 618250
rect 19290 618180 19360 618250
rect 19380 618180 19450 618250
rect 19470 618180 19540 618250
rect 19560 618180 19630 618250
rect 17670 618090 17740 618160
rect 17760 618090 17830 618160
rect 17850 618090 17920 618160
rect 17940 618090 18010 618160
rect 18030 618090 18100 618160
rect 18120 618090 18190 618160
rect 18210 618090 18280 618160
rect 18300 618090 18370 618160
rect 18390 618090 18460 618160
rect 18480 618090 18550 618160
rect 18570 618090 18640 618160
rect 18660 618090 18730 618160
rect 18750 618090 18820 618160
rect 18840 618090 18910 618160
rect 18930 618090 19000 618160
rect 19020 618090 19090 618160
rect 19110 618090 19180 618160
rect 19200 618090 19270 618160
rect 19290 618090 19360 618160
rect 19380 618090 19450 618160
rect 19470 618090 19540 618160
rect 19560 618090 19630 618160
rect 17670 618000 17740 618070
rect 17760 618000 17830 618070
rect 17850 618000 17920 618070
rect 17940 618000 18010 618070
rect 18030 618000 18100 618070
rect 18120 618000 18190 618070
rect 18210 618000 18280 618070
rect 18300 618000 18370 618070
rect 18390 618000 18460 618070
rect 18480 618000 18550 618070
rect 18570 618000 18640 618070
rect 18660 618000 18730 618070
rect 18750 618000 18820 618070
rect 18840 618000 18910 618070
rect 18930 618000 19000 618070
rect 19020 618000 19090 618070
rect 19110 618000 19180 618070
rect 19200 618000 19270 618070
rect 19290 618000 19360 618070
rect 19380 618000 19450 618070
rect 19470 618000 19540 618070
rect 19560 618000 19630 618070
rect 17670 617910 17740 617980
rect 17760 617910 17830 617980
rect 17850 617910 17920 617980
rect 17940 617910 18010 617980
rect 18030 617910 18100 617980
rect 18120 617910 18190 617980
rect 18210 617910 18280 617980
rect 18300 617910 18370 617980
rect 18390 617910 18460 617980
rect 18480 617910 18550 617980
rect 18570 617910 18640 617980
rect 18660 617910 18730 617980
rect 18750 617910 18820 617980
rect 18840 617910 18910 617980
rect 18930 617910 19000 617980
rect 19020 617910 19090 617980
rect 19110 617910 19180 617980
rect 19200 617910 19270 617980
rect 19290 617910 19360 617980
rect 19380 617910 19450 617980
rect 19470 617910 19540 617980
rect 19560 617910 19630 617980
rect 17670 617820 17740 617890
rect 17760 617820 17830 617890
rect 17850 617820 17920 617890
rect 17940 617820 18010 617890
rect 18030 617820 18100 617890
rect 18120 617820 18190 617890
rect 18210 617820 18280 617890
rect 18300 617820 18370 617890
rect 18390 617820 18460 617890
rect 18480 617820 18550 617890
rect 18570 617820 18640 617890
rect 18660 617820 18730 617890
rect 18750 617820 18820 617890
rect 18840 617820 18910 617890
rect 18930 617820 19000 617890
rect 19020 617820 19090 617890
rect 19110 617820 19180 617890
rect 19200 617820 19270 617890
rect 19290 617820 19360 617890
rect 19380 617820 19450 617890
rect 19470 617820 19540 617890
rect 19560 617820 19630 617890
rect 17670 617730 17740 617800
rect 17760 617730 17830 617800
rect 17850 617730 17920 617800
rect 17940 617730 18010 617800
rect 18030 617730 18100 617800
rect 18120 617730 18190 617800
rect 18210 617730 18280 617800
rect 18300 617730 18370 617800
rect 18390 617730 18460 617800
rect 18480 617730 18550 617800
rect 18570 617730 18640 617800
rect 18660 617730 18730 617800
rect 18750 617730 18820 617800
rect 18840 617730 18910 617800
rect 18930 617730 19000 617800
rect 19020 617730 19090 617800
rect 19110 617730 19180 617800
rect 19200 617730 19270 617800
rect 19290 617730 19360 617800
rect 19380 617730 19450 617800
rect 19470 617730 19540 617800
rect 19560 617730 19630 617800
rect 17670 617640 17740 617710
rect 17760 617640 17830 617710
rect 17850 617640 17920 617710
rect 17940 617640 18010 617710
rect 18030 617640 18100 617710
rect 18120 617640 18190 617710
rect 18210 617640 18280 617710
rect 18300 617640 18370 617710
rect 18390 617640 18460 617710
rect 18480 617640 18550 617710
rect 18570 617640 18640 617710
rect 18660 617640 18730 617710
rect 18750 617640 18820 617710
rect 18840 617640 18910 617710
rect 18930 617640 19000 617710
rect 19020 617640 19090 617710
rect 19110 617640 19180 617710
rect 19200 617640 19270 617710
rect 19290 617640 19360 617710
rect 19380 617640 19450 617710
rect 19470 617640 19540 617710
rect 19560 617640 19630 617710
rect 17670 617550 17740 617620
rect 17760 617550 17830 617620
rect 17850 617550 17920 617620
rect 17940 617550 18010 617620
rect 18030 617550 18100 617620
rect 18120 617550 18190 617620
rect 18210 617550 18280 617620
rect 18300 617550 18370 617620
rect 18390 617550 18460 617620
rect 18480 617550 18550 617620
rect 18570 617550 18640 617620
rect 18660 617550 18730 617620
rect 18750 617550 18820 617620
rect 18840 617550 18910 617620
rect 18930 617550 19000 617620
rect 19020 617550 19090 617620
rect 19110 617550 19180 617620
rect 19200 617550 19270 617620
rect 19290 617550 19360 617620
rect 19380 617550 19450 617620
rect 19470 617550 19540 617620
rect 19560 617550 19630 617620
rect 17670 617460 17740 617530
rect 17760 617460 17830 617530
rect 17850 617460 17920 617530
rect 17940 617460 18010 617530
rect 18030 617460 18100 617530
rect 18120 617460 18190 617530
rect 18210 617460 18280 617530
rect 18300 617460 18370 617530
rect 18390 617460 18460 617530
rect 18480 617460 18550 617530
rect 18570 617460 18640 617530
rect 18660 617460 18730 617530
rect 18750 617460 18820 617530
rect 18840 617460 18910 617530
rect 18930 617460 19000 617530
rect 19020 617460 19090 617530
rect 19110 617460 19180 617530
rect 19200 617460 19270 617530
rect 19290 617460 19360 617530
rect 19380 617460 19450 617530
rect 19470 617460 19540 617530
rect 19560 617460 19630 617530
<< metal4 >>
rect 18050 703830 19650 703900
rect 18050 703760 18070 703830
rect 18140 703760 18160 703830
rect 18230 703760 18250 703830
rect 18320 703760 18340 703830
rect 18410 703760 18430 703830
rect 18500 703760 18520 703830
rect 18590 703760 18610 703830
rect 18680 703760 18700 703830
rect 18770 703760 18790 703830
rect 18860 703760 18880 703830
rect 18950 703760 18970 703830
rect 19040 703760 19060 703830
rect 19130 703760 19150 703830
rect 19220 703760 19240 703830
rect 19310 703760 19330 703830
rect 19400 703760 19420 703830
rect 19490 703760 19510 703830
rect 19580 703760 19650 703830
rect 18050 703740 19650 703760
rect 18050 703670 18070 703740
rect 18140 703670 18160 703740
rect 18230 703670 18250 703740
rect 18320 703670 18340 703740
rect 18410 703670 18430 703740
rect 18500 703670 18520 703740
rect 18590 703670 18610 703740
rect 18680 703670 18700 703740
rect 18770 703670 18790 703740
rect 18860 703670 18880 703740
rect 18950 703670 18970 703740
rect 19040 703670 19060 703740
rect 19130 703670 19150 703740
rect 19220 703670 19240 703740
rect 19310 703670 19330 703740
rect 19400 703670 19420 703740
rect 19490 703670 19510 703740
rect 19580 703670 19650 703740
rect 18050 703650 19650 703670
rect 18050 703580 18070 703650
rect 18140 703580 18160 703650
rect 18230 703580 18250 703650
rect 18320 703580 18340 703650
rect 18410 703580 18430 703650
rect 18500 703580 18520 703650
rect 18590 703580 18610 703650
rect 18680 703580 18700 703650
rect 18770 703580 18790 703650
rect 18860 703580 18880 703650
rect 18950 703580 18970 703650
rect 19040 703580 19060 703650
rect 19130 703580 19150 703650
rect 19220 703580 19240 703650
rect 19310 703580 19330 703650
rect 19400 703580 19420 703650
rect 19490 703580 19510 703650
rect 19580 703580 19650 703650
rect 18050 703560 19650 703580
rect 18050 703490 18070 703560
rect 18140 703490 18160 703560
rect 18230 703490 18250 703560
rect 18320 703490 18340 703560
rect 18410 703490 18430 703560
rect 18500 703490 18520 703560
rect 18590 703490 18610 703560
rect 18680 703490 18700 703560
rect 18770 703490 18790 703560
rect 18860 703490 18880 703560
rect 18950 703490 18970 703560
rect 19040 703490 19060 703560
rect 19130 703490 19150 703560
rect 19220 703490 19240 703560
rect 19310 703490 19330 703560
rect 19400 703490 19420 703560
rect 19490 703490 19510 703560
rect 19580 703490 19650 703560
rect 18050 703470 19650 703490
rect 18050 703400 18070 703470
rect 18140 703400 18160 703470
rect 18230 703400 18250 703470
rect 18320 703400 18340 703470
rect 18410 703400 18430 703470
rect 18500 703400 18520 703470
rect 18590 703400 18610 703470
rect 18680 703400 18700 703470
rect 18770 703400 18790 703470
rect 18860 703400 18880 703470
rect 18950 703400 18970 703470
rect 19040 703400 19060 703470
rect 19130 703400 19150 703470
rect 19220 703400 19240 703470
rect 19310 703400 19330 703470
rect 19400 703400 19420 703470
rect 19490 703400 19510 703470
rect 19580 703400 19650 703470
rect 18050 703380 19650 703400
rect 18050 703310 18070 703380
rect 18140 703310 18160 703380
rect 18230 703310 18250 703380
rect 18320 703310 18340 703380
rect 18410 703310 18430 703380
rect 18500 703310 18520 703380
rect 18590 703310 18610 703380
rect 18680 703310 18700 703380
rect 18770 703310 18790 703380
rect 18860 703310 18880 703380
rect 18950 703310 18970 703380
rect 19040 703310 19060 703380
rect 19130 703310 19150 703380
rect 19220 703310 19240 703380
rect 19310 703310 19330 703380
rect 19400 703310 19420 703380
rect 19490 703310 19510 703380
rect 19580 703310 19650 703380
rect 18050 703290 19650 703310
rect 18050 703220 18070 703290
rect 18140 703220 18160 703290
rect 18230 703220 18250 703290
rect 18320 703220 18340 703290
rect 18410 703220 18430 703290
rect 18500 703220 18520 703290
rect 18590 703220 18610 703290
rect 18680 703220 18700 703290
rect 18770 703220 18790 703290
rect 18860 703220 18880 703290
rect 18950 703220 18970 703290
rect 19040 703220 19060 703290
rect 19130 703220 19150 703290
rect 19220 703220 19240 703290
rect 19310 703220 19330 703290
rect 19400 703220 19420 703290
rect 19490 703220 19510 703290
rect 19580 703220 19650 703290
rect 18050 703200 19650 703220
rect 18050 703130 18070 703200
rect 18140 703130 18160 703200
rect 18230 703130 18250 703200
rect 18320 703130 18340 703200
rect 18410 703130 18430 703200
rect 18500 703130 18520 703200
rect 18590 703130 18610 703200
rect 18680 703130 18700 703200
rect 18770 703130 18790 703200
rect 18860 703130 18880 703200
rect 18950 703130 18970 703200
rect 19040 703130 19060 703200
rect 19130 703130 19150 703200
rect 19220 703130 19240 703200
rect 19310 703130 19330 703200
rect 19400 703130 19420 703200
rect 19490 703130 19510 703200
rect 19580 703130 19650 703200
rect 18050 703110 19650 703130
rect 18050 703040 18070 703110
rect 18140 703040 18160 703110
rect 18230 703040 18250 703110
rect 18320 703040 18340 703110
rect 18410 703040 18430 703110
rect 18500 703040 18520 703110
rect 18590 703040 18610 703110
rect 18680 703040 18700 703110
rect 18770 703040 18790 703110
rect 18860 703040 18880 703110
rect 18950 703040 18970 703110
rect 19040 703040 19060 703110
rect 19130 703040 19150 703110
rect 19220 703040 19240 703110
rect 19310 703040 19330 703110
rect 19400 703040 19420 703110
rect 19490 703040 19510 703110
rect 19580 703040 19650 703110
rect 18050 703020 19650 703040
rect 18050 702950 18070 703020
rect 18140 702950 18160 703020
rect 18230 702950 18250 703020
rect 18320 702950 18340 703020
rect 18410 702950 18430 703020
rect 18500 702950 18520 703020
rect 18590 702950 18610 703020
rect 18680 702950 18700 703020
rect 18770 702950 18790 703020
rect 18860 702950 18880 703020
rect 18950 702950 18970 703020
rect 19040 702950 19060 703020
rect 19130 702950 19150 703020
rect 19220 702950 19240 703020
rect 19310 702950 19330 703020
rect 19400 702950 19420 703020
rect 19490 702950 19510 703020
rect 19580 702950 19650 703020
rect 18050 702930 19650 702950
rect 18050 702860 18070 702930
rect 18140 702860 18160 702930
rect 18230 702860 18250 702930
rect 18320 702860 18340 702930
rect 18410 702860 18430 702930
rect 18500 702860 18520 702930
rect 18590 702860 18610 702930
rect 18680 702860 18700 702930
rect 18770 702860 18790 702930
rect 18860 702860 18880 702930
rect 18950 702860 18970 702930
rect 19040 702860 19060 702930
rect 19130 702860 19150 702930
rect 19220 702860 19240 702930
rect 19310 702860 19330 702930
rect 19400 702860 19420 702930
rect 19490 702860 19510 702930
rect 19580 702860 19650 702930
rect 18050 702840 19650 702860
rect 18050 702770 18070 702840
rect 18140 702770 18160 702840
rect 18230 702770 18250 702840
rect 18320 702770 18340 702840
rect 18410 702770 18430 702840
rect 18500 702770 18520 702840
rect 18590 702770 18610 702840
rect 18680 702770 18700 702840
rect 18770 702770 18790 702840
rect 18860 702770 18880 702840
rect 18950 702770 18970 702840
rect 19040 702770 19060 702840
rect 19130 702770 19150 702840
rect 19220 702770 19240 702840
rect 19310 702770 19330 702840
rect 19400 702770 19420 702840
rect 19490 702770 19510 702840
rect 19580 702770 19650 702840
rect 18050 702750 19650 702770
rect 18050 702680 18070 702750
rect 18140 702680 18160 702750
rect 18230 702680 18250 702750
rect 18320 702680 18340 702750
rect 18410 702680 18430 702750
rect 18500 702680 18520 702750
rect 18590 702680 18610 702750
rect 18680 702680 18700 702750
rect 18770 702680 18790 702750
rect 18860 702680 18880 702750
rect 18950 702680 18970 702750
rect 19040 702680 19060 702750
rect 19130 702680 19150 702750
rect 19220 702680 19240 702750
rect 19310 702680 19330 702750
rect 19400 702680 19420 702750
rect 19490 702680 19510 702750
rect 19580 702680 19650 702750
rect 18050 702660 19650 702680
rect 18050 702590 18070 702660
rect 18140 702590 18160 702660
rect 18230 702590 18250 702660
rect 18320 702590 18340 702660
rect 18410 702590 18430 702660
rect 18500 702590 18520 702660
rect 18590 702590 18610 702660
rect 18680 702590 18700 702660
rect 18770 702590 18790 702660
rect 18860 702590 18880 702660
rect 18950 702590 18970 702660
rect 19040 702590 19060 702660
rect 19130 702590 19150 702660
rect 19220 702590 19240 702660
rect 19310 702590 19330 702660
rect 19400 702590 19420 702660
rect 19490 702590 19510 702660
rect 19580 702590 19650 702660
rect 18050 702570 19650 702590
rect 18050 702500 18070 702570
rect 18140 702500 18160 702570
rect 18230 702500 18250 702570
rect 18320 702500 18340 702570
rect 18410 702500 18430 702570
rect 18500 702500 18520 702570
rect 18590 702500 18610 702570
rect 18680 702500 18700 702570
rect 18770 702500 18790 702570
rect 18860 702500 18880 702570
rect 18950 702500 18970 702570
rect 19040 702500 19060 702570
rect 19130 702500 19150 702570
rect 19220 702500 19240 702570
rect 19310 702500 19330 702570
rect 19400 702500 19420 702570
rect 19490 702500 19510 702570
rect 19580 702500 19650 702570
rect 18050 702480 19650 702500
rect 18050 702410 18070 702480
rect 18140 702410 18160 702480
rect 18230 702410 18250 702480
rect 18320 702410 18340 702480
rect 18410 702410 18430 702480
rect 18500 702410 18520 702480
rect 18590 702410 18610 702480
rect 18680 702410 18700 702480
rect 18770 702410 18790 702480
rect 18860 702410 18880 702480
rect 18950 702410 18970 702480
rect 19040 702410 19060 702480
rect 19130 702410 19150 702480
rect 19220 702410 19240 702480
rect 19310 702410 19330 702480
rect 19400 702410 19420 702480
rect 19490 702410 19510 702480
rect 19580 702410 19650 702480
rect 18050 702390 19650 702410
rect 18050 702320 18070 702390
rect 18140 702320 18160 702390
rect 18230 702320 18250 702390
rect 18320 702320 18340 702390
rect 18410 702320 18430 702390
rect 18500 702320 18520 702390
rect 18590 702320 18610 702390
rect 18680 702320 18700 702390
rect 18770 702320 18790 702390
rect 18860 702320 18880 702390
rect 18950 702320 18970 702390
rect 19040 702320 19060 702390
rect 19130 702320 19150 702390
rect 19220 702320 19240 702390
rect 19310 702320 19330 702390
rect 19400 702320 19420 702390
rect 19490 702320 19510 702390
rect 19580 702320 19650 702390
rect 18050 695790 19650 702320
rect 70070 703830 71670 703900
rect 70070 703760 70090 703830
rect 70160 703760 70180 703830
rect 70250 703760 70270 703830
rect 70340 703760 70360 703830
rect 70430 703760 70450 703830
rect 70520 703760 70540 703830
rect 70610 703760 70630 703830
rect 70700 703760 70720 703830
rect 70790 703760 70810 703830
rect 70880 703760 70900 703830
rect 70970 703760 70990 703830
rect 71060 703760 71080 703830
rect 71150 703760 71170 703830
rect 71240 703760 71260 703830
rect 71330 703760 71350 703830
rect 71420 703760 71440 703830
rect 71510 703760 71530 703830
rect 71600 703760 71670 703830
rect 70070 703740 71670 703760
rect 70070 703670 70090 703740
rect 70160 703670 70180 703740
rect 70250 703670 70270 703740
rect 70340 703670 70360 703740
rect 70430 703670 70450 703740
rect 70520 703670 70540 703740
rect 70610 703670 70630 703740
rect 70700 703670 70720 703740
rect 70790 703670 70810 703740
rect 70880 703670 70900 703740
rect 70970 703670 70990 703740
rect 71060 703670 71080 703740
rect 71150 703670 71170 703740
rect 71240 703670 71260 703740
rect 71330 703670 71350 703740
rect 71420 703670 71440 703740
rect 71510 703670 71530 703740
rect 71600 703670 71670 703740
rect 70070 703650 71670 703670
rect 70070 703580 70090 703650
rect 70160 703580 70180 703650
rect 70250 703580 70270 703650
rect 70340 703580 70360 703650
rect 70430 703580 70450 703650
rect 70520 703580 70540 703650
rect 70610 703580 70630 703650
rect 70700 703580 70720 703650
rect 70790 703580 70810 703650
rect 70880 703580 70900 703650
rect 70970 703580 70990 703650
rect 71060 703580 71080 703650
rect 71150 703580 71170 703650
rect 71240 703580 71260 703650
rect 71330 703580 71350 703650
rect 71420 703580 71440 703650
rect 71510 703580 71530 703650
rect 71600 703580 71670 703650
rect 70070 703560 71670 703580
rect 70070 703490 70090 703560
rect 70160 703490 70180 703560
rect 70250 703490 70270 703560
rect 70340 703490 70360 703560
rect 70430 703490 70450 703560
rect 70520 703490 70540 703560
rect 70610 703490 70630 703560
rect 70700 703490 70720 703560
rect 70790 703490 70810 703560
rect 70880 703490 70900 703560
rect 70970 703490 70990 703560
rect 71060 703490 71080 703560
rect 71150 703490 71170 703560
rect 71240 703490 71260 703560
rect 71330 703490 71350 703560
rect 71420 703490 71440 703560
rect 71510 703490 71530 703560
rect 71600 703490 71670 703560
rect 70070 703470 71670 703490
rect 70070 703400 70090 703470
rect 70160 703400 70180 703470
rect 70250 703400 70270 703470
rect 70340 703400 70360 703470
rect 70430 703400 70450 703470
rect 70520 703400 70540 703470
rect 70610 703400 70630 703470
rect 70700 703400 70720 703470
rect 70790 703400 70810 703470
rect 70880 703400 70900 703470
rect 70970 703400 70990 703470
rect 71060 703400 71080 703470
rect 71150 703400 71170 703470
rect 71240 703400 71260 703470
rect 71330 703400 71350 703470
rect 71420 703400 71440 703470
rect 71510 703400 71530 703470
rect 71600 703400 71670 703470
rect 70070 703380 71670 703400
rect 70070 703310 70090 703380
rect 70160 703310 70180 703380
rect 70250 703310 70270 703380
rect 70340 703310 70360 703380
rect 70430 703310 70450 703380
rect 70520 703310 70540 703380
rect 70610 703310 70630 703380
rect 70700 703310 70720 703380
rect 70790 703310 70810 703380
rect 70880 703310 70900 703380
rect 70970 703310 70990 703380
rect 71060 703310 71080 703380
rect 71150 703310 71170 703380
rect 71240 703310 71260 703380
rect 71330 703310 71350 703380
rect 71420 703310 71440 703380
rect 71510 703310 71530 703380
rect 71600 703310 71670 703380
rect 70070 703290 71670 703310
rect 70070 703220 70090 703290
rect 70160 703220 70180 703290
rect 70250 703220 70270 703290
rect 70340 703220 70360 703290
rect 70430 703220 70450 703290
rect 70520 703220 70540 703290
rect 70610 703220 70630 703290
rect 70700 703220 70720 703290
rect 70790 703220 70810 703290
rect 70880 703220 70900 703290
rect 70970 703220 70990 703290
rect 71060 703220 71080 703290
rect 71150 703220 71170 703290
rect 71240 703220 71260 703290
rect 71330 703220 71350 703290
rect 71420 703220 71440 703290
rect 71510 703220 71530 703290
rect 71600 703220 71670 703290
rect 70070 703200 71670 703220
rect 70070 703130 70090 703200
rect 70160 703130 70180 703200
rect 70250 703130 70270 703200
rect 70340 703130 70360 703200
rect 70430 703130 70450 703200
rect 70520 703130 70540 703200
rect 70610 703130 70630 703200
rect 70700 703130 70720 703200
rect 70790 703130 70810 703200
rect 70880 703130 70900 703200
rect 70970 703130 70990 703200
rect 71060 703130 71080 703200
rect 71150 703130 71170 703200
rect 71240 703130 71260 703200
rect 71330 703130 71350 703200
rect 71420 703130 71440 703200
rect 71510 703130 71530 703200
rect 71600 703130 71670 703200
rect 70070 703110 71670 703130
rect 70070 703040 70090 703110
rect 70160 703040 70180 703110
rect 70250 703040 70270 703110
rect 70340 703040 70360 703110
rect 70430 703040 70450 703110
rect 70520 703040 70540 703110
rect 70610 703040 70630 703110
rect 70700 703040 70720 703110
rect 70790 703040 70810 703110
rect 70880 703040 70900 703110
rect 70970 703040 70990 703110
rect 71060 703040 71080 703110
rect 71150 703040 71170 703110
rect 71240 703040 71260 703110
rect 71330 703040 71350 703110
rect 71420 703040 71440 703110
rect 71510 703040 71530 703110
rect 71600 703040 71670 703110
rect 70070 703020 71670 703040
rect 70070 702950 70090 703020
rect 70160 702950 70180 703020
rect 70250 702950 70270 703020
rect 70340 702950 70360 703020
rect 70430 702950 70450 703020
rect 70520 702950 70540 703020
rect 70610 702950 70630 703020
rect 70700 702950 70720 703020
rect 70790 702950 70810 703020
rect 70880 702950 70900 703020
rect 70970 702950 70990 703020
rect 71060 702950 71080 703020
rect 71150 702950 71170 703020
rect 71240 702950 71260 703020
rect 71330 702950 71350 703020
rect 71420 702950 71440 703020
rect 71510 702950 71530 703020
rect 71600 702950 71670 703020
rect 70070 702930 71670 702950
rect 70070 702860 70090 702930
rect 70160 702860 70180 702930
rect 70250 702860 70270 702930
rect 70340 702860 70360 702930
rect 70430 702860 70450 702930
rect 70520 702860 70540 702930
rect 70610 702860 70630 702930
rect 70700 702860 70720 702930
rect 70790 702860 70810 702930
rect 70880 702860 70900 702930
rect 70970 702860 70990 702930
rect 71060 702860 71080 702930
rect 71150 702860 71170 702930
rect 71240 702860 71260 702930
rect 71330 702860 71350 702930
rect 71420 702860 71440 702930
rect 71510 702860 71530 702930
rect 71600 702860 71670 702930
rect 70070 702840 71670 702860
rect 70070 702770 70090 702840
rect 70160 702770 70180 702840
rect 70250 702770 70270 702840
rect 70340 702770 70360 702840
rect 70430 702770 70450 702840
rect 70520 702770 70540 702840
rect 70610 702770 70630 702840
rect 70700 702770 70720 702840
rect 70790 702770 70810 702840
rect 70880 702770 70900 702840
rect 70970 702770 70990 702840
rect 71060 702770 71080 702840
rect 71150 702770 71170 702840
rect 71240 702770 71260 702840
rect 71330 702770 71350 702840
rect 71420 702770 71440 702840
rect 71510 702770 71530 702840
rect 71600 702770 71670 702840
rect 70070 702750 71670 702770
rect 70070 702680 70090 702750
rect 70160 702680 70180 702750
rect 70250 702680 70270 702750
rect 70340 702680 70360 702750
rect 70430 702680 70450 702750
rect 70520 702680 70540 702750
rect 70610 702680 70630 702750
rect 70700 702680 70720 702750
rect 70790 702680 70810 702750
rect 70880 702680 70900 702750
rect 70970 702680 70990 702750
rect 71060 702680 71080 702750
rect 71150 702680 71170 702750
rect 71240 702680 71260 702750
rect 71330 702680 71350 702750
rect 71420 702680 71440 702750
rect 71510 702680 71530 702750
rect 71600 702680 71670 702750
rect 70070 702660 71670 702680
rect 70070 702590 70090 702660
rect 70160 702590 70180 702660
rect 70250 702590 70270 702660
rect 70340 702590 70360 702660
rect 70430 702590 70450 702660
rect 70520 702590 70540 702660
rect 70610 702590 70630 702660
rect 70700 702590 70720 702660
rect 70790 702590 70810 702660
rect 70880 702590 70900 702660
rect 70970 702590 70990 702660
rect 71060 702590 71080 702660
rect 71150 702590 71170 702660
rect 71240 702590 71260 702660
rect 71330 702590 71350 702660
rect 71420 702590 71440 702660
rect 71510 702590 71530 702660
rect 71600 702590 71670 702660
rect 70070 702570 71670 702590
rect 70070 702500 70090 702570
rect 70160 702500 70180 702570
rect 70250 702500 70270 702570
rect 70340 702500 70360 702570
rect 70430 702500 70450 702570
rect 70520 702500 70540 702570
rect 70610 702500 70630 702570
rect 70700 702500 70720 702570
rect 70790 702500 70810 702570
rect 70880 702500 70900 702570
rect 70970 702500 70990 702570
rect 71060 702500 71080 702570
rect 71150 702500 71170 702570
rect 71240 702500 71260 702570
rect 71330 702500 71350 702570
rect 71420 702500 71440 702570
rect 71510 702500 71530 702570
rect 71600 702500 71670 702570
rect 70070 702480 71670 702500
rect 70070 702410 70090 702480
rect 70160 702410 70180 702480
rect 70250 702410 70270 702480
rect 70340 702410 70360 702480
rect 70430 702410 70450 702480
rect 70520 702410 70540 702480
rect 70610 702410 70630 702480
rect 70700 702410 70720 702480
rect 70790 702410 70810 702480
rect 70880 702410 70900 702480
rect 70970 702410 70990 702480
rect 71060 702410 71080 702480
rect 71150 702410 71170 702480
rect 71240 702410 71260 702480
rect 71330 702410 71350 702480
rect 71420 702410 71440 702480
rect 71510 702410 71530 702480
rect 71600 702410 71670 702480
rect 70070 702390 71670 702410
rect 70070 702320 70090 702390
rect 70160 702320 70180 702390
rect 70250 702320 70270 702390
rect 70340 702320 70360 702390
rect 70430 702320 70450 702390
rect 70520 702320 70540 702390
rect 70610 702320 70630 702390
rect 70700 702320 70720 702390
rect 70790 702320 70810 702390
rect 70880 702320 70900 702390
rect 70970 702320 70990 702390
rect 71060 702320 71080 702390
rect 71150 702320 71170 702390
rect 71240 702320 71260 702390
rect 71330 702320 71350 702390
rect 71420 702320 71440 702390
rect 71510 702320 71530 702390
rect 71600 702320 71670 702390
rect 18050 687370 19650 693230
rect 18050 687300 18120 687370
rect 18190 687300 18210 687370
rect 18280 687300 18300 687370
rect 18370 687300 18390 687370
rect 18460 687300 18480 687370
rect 18550 687300 18570 687370
rect 18640 687300 18660 687370
rect 18730 687300 18750 687370
rect 18820 687300 18840 687370
rect 18910 687300 18930 687370
rect 19000 687300 19020 687370
rect 19090 687300 19110 687370
rect 19180 687300 19200 687370
rect 19270 687300 19290 687370
rect 19360 687300 19380 687370
rect 19450 687300 19470 687370
rect 19540 687300 19560 687370
rect 19630 687300 19650 687370
rect 18050 687280 19650 687300
rect 18050 687210 18120 687280
rect 18190 687210 18210 687280
rect 18280 687210 18300 687280
rect 18370 687210 18390 687280
rect 18460 687210 18480 687280
rect 18550 687210 18570 687280
rect 18640 687210 18660 687280
rect 18730 687210 18750 687280
rect 18820 687210 18840 687280
rect 18910 687210 18930 687280
rect 19000 687210 19020 687280
rect 19090 687210 19110 687280
rect 19180 687210 19200 687280
rect 19270 687210 19290 687280
rect 19360 687210 19380 687280
rect 19450 687210 19470 687280
rect 19540 687210 19560 687280
rect 19630 687210 19650 687280
rect 18050 687190 19650 687210
rect 18050 687120 18120 687190
rect 18190 687120 18210 687190
rect 18280 687120 18300 687190
rect 18370 687120 18390 687190
rect 18460 687120 18480 687190
rect 18550 687120 18570 687190
rect 18640 687120 18660 687190
rect 18730 687120 18750 687190
rect 18820 687120 18840 687190
rect 18910 687120 18930 687190
rect 19000 687120 19020 687190
rect 19090 687120 19110 687190
rect 19180 687120 19200 687190
rect 19270 687120 19290 687190
rect 19360 687120 19380 687190
rect 19450 687120 19470 687190
rect 19540 687120 19560 687190
rect 19630 687120 19650 687190
rect 18050 687100 19650 687120
rect 18050 687030 18120 687100
rect 18190 687030 18210 687100
rect 18280 687030 18300 687100
rect 18370 687030 18390 687100
rect 18460 687030 18480 687100
rect 18550 687030 18570 687100
rect 18640 687030 18660 687100
rect 18730 687030 18750 687100
rect 18820 687030 18840 687100
rect 18910 687030 18930 687100
rect 19000 687030 19020 687100
rect 19090 687030 19110 687100
rect 19180 687030 19200 687100
rect 19270 687030 19290 687100
rect 19360 687030 19380 687100
rect 19450 687030 19470 687100
rect 19540 687030 19560 687100
rect 19630 687030 19650 687100
rect 18050 687010 19650 687030
rect 18050 686940 18120 687010
rect 18190 686940 18210 687010
rect 18280 686940 18300 687010
rect 18370 686940 18390 687010
rect 18460 686940 18480 687010
rect 18550 686940 18570 687010
rect 18640 686940 18660 687010
rect 18730 686940 18750 687010
rect 18820 686940 18840 687010
rect 18910 686940 18930 687010
rect 19000 686940 19020 687010
rect 19090 686940 19110 687010
rect 19180 686940 19200 687010
rect 19270 686940 19290 687010
rect 19360 686940 19380 687010
rect 19450 686940 19470 687010
rect 19540 686940 19560 687010
rect 19630 686940 19650 687010
rect 18050 686920 19650 686940
rect 18050 686850 18120 686920
rect 18190 686850 18210 686920
rect 18280 686850 18300 686920
rect 18370 686850 18390 686920
rect 18460 686850 18480 686920
rect 18550 686850 18570 686920
rect 18640 686850 18660 686920
rect 18730 686850 18750 686920
rect 18820 686850 18840 686920
rect 18910 686850 18930 686920
rect 19000 686850 19020 686920
rect 19090 686850 19110 686920
rect 19180 686850 19200 686920
rect 19270 686850 19290 686920
rect 19360 686850 19380 686920
rect 19450 686850 19470 686920
rect 19540 686850 19560 686920
rect 19630 686850 19650 686920
rect 18050 686830 19650 686850
rect 18050 686760 18120 686830
rect 18190 686760 18210 686830
rect 18280 686760 18300 686830
rect 18370 686760 18390 686830
rect 18460 686760 18480 686830
rect 18550 686760 18570 686830
rect 18640 686760 18660 686830
rect 18730 686760 18750 686830
rect 18820 686760 18840 686830
rect 18910 686760 18930 686830
rect 19000 686760 19020 686830
rect 19090 686760 19110 686830
rect 19180 686760 19200 686830
rect 19270 686760 19290 686830
rect 19360 686760 19380 686830
rect 19450 686760 19470 686830
rect 19540 686760 19560 686830
rect 19630 686760 19650 686830
rect 18050 686740 19650 686760
rect 18050 686670 18120 686740
rect 18190 686670 18210 686740
rect 18280 686670 18300 686740
rect 18370 686670 18390 686740
rect 18460 686670 18480 686740
rect 18550 686670 18570 686740
rect 18640 686670 18660 686740
rect 18730 686670 18750 686740
rect 18820 686670 18840 686740
rect 18910 686670 18930 686740
rect 19000 686670 19020 686740
rect 19090 686670 19110 686740
rect 19180 686670 19200 686740
rect 19270 686670 19290 686740
rect 19360 686670 19380 686740
rect 19450 686670 19470 686740
rect 19540 686670 19560 686740
rect 19630 686670 19650 686740
rect 18050 686650 19650 686670
rect 18050 686580 18120 686650
rect 18190 686580 18210 686650
rect 18280 686580 18300 686650
rect 18370 686580 18390 686650
rect 18460 686580 18480 686650
rect 18550 686580 18570 686650
rect 18640 686580 18660 686650
rect 18730 686580 18750 686650
rect 18820 686580 18840 686650
rect 18910 686580 18930 686650
rect 19000 686580 19020 686650
rect 19090 686580 19110 686650
rect 19180 686580 19200 686650
rect 19270 686580 19290 686650
rect 19360 686580 19380 686650
rect 19450 686580 19470 686650
rect 19540 686580 19560 686650
rect 19630 686580 19650 686650
rect 18050 686560 19650 686580
rect 18050 686490 18120 686560
rect 18190 686490 18210 686560
rect 18280 686490 18300 686560
rect 18370 686490 18390 686560
rect 18460 686490 18480 686560
rect 18550 686490 18570 686560
rect 18640 686490 18660 686560
rect 18730 686490 18750 686560
rect 18820 686490 18840 686560
rect 18910 686490 18930 686560
rect 19000 686490 19020 686560
rect 19090 686490 19110 686560
rect 19180 686490 19200 686560
rect 19270 686490 19290 686560
rect 19360 686490 19380 686560
rect 19450 686490 19470 686560
rect 19540 686490 19560 686560
rect 19630 686490 19650 686560
rect 18050 686470 19650 686490
rect 18050 686400 18120 686470
rect 18190 686400 18210 686470
rect 18280 686400 18300 686470
rect 18370 686400 18390 686470
rect 18460 686400 18480 686470
rect 18550 686400 18570 686470
rect 18640 686400 18660 686470
rect 18730 686400 18750 686470
rect 18820 686400 18840 686470
rect 18910 686400 18930 686470
rect 19000 686400 19020 686470
rect 19090 686400 19110 686470
rect 19180 686400 19200 686470
rect 19270 686400 19290 686470
rect 19360 686400 19380 686470
rect 19450 686400 19470 686470
rect 19540 686400 19560 686470
rect 19630 686400 19650 686470
rect 18050 686380 19650 686400
rect 18050 686310 18120 686380
rect 18190 686310 18210 686380
rect 18280 686310 18300 686380
rect 18370 686310 18390 686380
rect 18460 686310 18480 686380
rect 18550 686310 18570 686380
rect 18640 686310 18660 686380
rect 18730 686310 18750 686380
rect 18820 686310 18840 686380
rect 18910 686310 18930 686380
rect 19000 686310 19020 686380
rect 19090 686310 19110 686380
rect 19180 686310 19200 686380
rect 19270 686310 19290 686380
rect 19360 686310 19380 686380
rect 19450 686310 19470 686380
rect 19540 686310 19560 686380
rect 19630 686310 19650 686380
rect 18050 686290 19650 686310
rect 18050 686220 18120 686290
rect 18190 686220 18210 686290
rect 18280 686220 18300 686290
rect 18370 686220 18390 686290
rect 18460 686220 18480 686290
rect 18550 686220 18570 686290
rect 18640 686220 18660 686290
rect 18730 686220 18750 686290
rect 18820 686220 18840 686290
rect 18910 686220 18930 686290
rect 19000 686220 19020 686290
rect 19090 686220 19110 686290
rect 19180 686220 19200 686290
rect 19270 686220 19290 686290
rect 19360 686220 19380 686290
rect 19450 686220 19470 686290
rect 19540 686220 19560 686290
rect 19630 686220 19650 686290
rect 18050 686200 19650 686220
rect 18050 686130 18120 686200
rect 18190 686130 18210 686200
rect 18280 686130 18300 686200
rect 18370 686130 18390 686200
rect 18460 686130 18480 686200
rect 18550 686130 18570 686200
rect 18640 686130 18660 686200
rect 18730 686130 18750 686200
rect 18820 686130 18840 686200
rect 18910 686130 18930 686200
rect 19000 686130 19020 686200
rect 19090 686130 19110 686200
rect 19180 686130 19200 686200
rect 19270 686130 19290 686200
rect 19360 686130 19380 686200
rect 19450 686130 19470 686200
rect 19540 686130 19560 686200
rect 19630 686130 19650 686200
rect 18050 686110 19650 686130
rect 18050 686040 18120 686110
rect 18190 686040 18210 686110
rect 18280 686040 18300 686110
rect 18370 686040 18390 686110
rect 18460 686040 18480 686110
rect 18550 686040 18570 686110
rect 18640 686040 18660 686110
rect 18730 686040 18750 686110
rect 18820 686040 18840 686110
rect 18910 686040 18930 686110
rect 19000 686040 19020 686110
rect 19090 686040 19110 686110
rect 19180 686040 19200 686110
rect 19270 686040 19290 686110
rect 19360 686040 19380 686110
rect 19450 686040 19470 686110
rect 19540 686040 19560 686110
rect 19630 686040 19650 686110
rect 18050 686020 19650 686040
rect 18050 685950 18120 686020
rect 18190 685950 18210 686020
rect 18280 685950 18300 686020
rect 18370 685950 18390 686020
rect 18460 685950 18480 686020
rect 18550 685950 18570 686020
rect 18640 685950 18660 686020
rect 18730 685950 18750 686020
rect 18820 685950 18840 686020
rect 18910 685950 18930 686020
rect 19000 685950 19020 686020
rect 19090 685950 19110 686020
rect 19180 685950 19200 686020
rect 19270 685950 19290 686020
rect 19360 685950 19380 686020
rect 19450 685950 19470 686020
rect 19540 685950 19560 686020
rect 19630 685950 19650 686020
rect 18050 685930 19650 685950
rect 18050 685860 18120 685930
rect 18190 685860 18210 685930
rect 18280 685860 18300 685930
rect 18370 685860 18390 685930
rect 18460 685860 18480 685930
rect 18550 685860 18570 685930
rect 18640 685860 18660 685930
rect 18730 685860 18750 685930
rect 18820 685860 18840 685930
rect 18910 685860 18930 685930
rect 19000 685860 19020 685930
rect 19090 685860 19110 685930
rect 19180 685860 19200 685930
rect 19270 685860 19290 685930
rect 19360 685860 19380 685930
rect 19450 685860 19470 685930
rect 19540 685860 19560 685930
rect 19630 685860 19650 685930
rect 18050 685840 19650 685860
rect 18050 685770 18120 685840
rect 18190 685770 18210 685840
rect 18280 685770 18300 685840
rect 18370 685770 18390 685840
rect 18460 685770 18480 685840
rect 18550 685770 18570 685840
rect 18640 685770 18660 685840
rect 18730 685770 18750 685840
rect 18820 685770 18840 685840
rect 18910 685770 18930 685840
rect 19000 685770 19020 685840
rect 19090 685770 19110 685840
rect 19180 685770 19200 685840
rect 19270 685770 19290 685840
rect 19360 685770 19380 685840
rect 19450 685770 19470 685840
rect 19540 685770 19560 685840
rect 19630 685770 19650 685840
rect 18050 685750 19650 685770
rect 18050 685680 18120 685750
rect 18190 685680 18210 685750
rect 18280 685680 18300 685750
rect 18370 685680 18390 685750
rect 18460 685680 18480 685750
rect 18550 685680 18570 685750
rect 18640 685680 18660 685750
rect 18730 685680 18750 685750
rect 18820 685680 18840 685750
rect 18910 685680 18930 685750
rect 19000 685680 19020 685750
rect 19090 685680 19110 685750
rect 19180 685680 19200 685750
rect 19270 685680 19290 685750
rect 19360 685680 19380 685750
rect 19450 685680 19470 685750
rect 19540 685680 19560 685750
rect 19630 685680 19650 685750
rect 18050 685660 19650 685680
rect 18050 685590 18120 685660
rect 18190 685590 18210 685660
rect 18280 685590 18300 685660
rect 18370 685590 18390 685660
rect 18460 685590 18480 685660
rect 18550 685590 18570 685660
rect 18640 685590 18660 685660
rect 18730 685590 18750 685660
rect 18820 685590 18840 685660
rect 18910 685590 18930 685660
rect 19000 685590 19020 685660
rect 19090 685590 19110 685660
rect 19180 685590 19200 685660
rect 19270 685590 19290 685660
rect 19360 685590 19380 685660
rect 19450 685590 19470 685660
rect 19540 685590 19560 685660
rect 19630 685590 19650 685660
rect 18050 685570 19650 685590
rect 18050 685500 18120 685570
rect 18190 685500 18210 685570
rect 18280 685500 18300 685570
rect 18370 685500 18390 685570
rect 18460 685500 18480 685570
rect 18550 685500 18570 685570
rect 18640 685500 18660 685570
rect 18730 685500 18750 685570
rect 18820 685500 18840 685570
rect 18910 685500 18930 685570
rect 19000 685500 19020 685570
rect 19090 685500 19110 685570
rect 19180 685500 19200 685570
rect 19270 685500 19290 685570
rect 19360 685500 19380 685570
rect 19450 685500 19470 685570
rect 19540 685500 19560 685570
rect 19630 685500 19650 685570
rect 18050 685480 19650 685500
rect 18050 685410 18120 685480
rect 18190 685410 18210 685480
rect 18280 685410 18300 685480
rect 18370 685410 18390 685480
rect 18460 685410 18480 685480
rect 18550 685410 18570 685480
rect 18640 685410 18660 685480
rect 18730 685410 18750 685480
rect 18820 685410 18840 685480
rect 18910 685410 18930 685480
rect 19000 685410 19020 685480
rect 19090 685410 19110 685480
rect 19180 685410 19200 685480
rect 19270 685410 19290 685480
rect 19360 685410 19380 685480
rect 19450 685410 19470 685480
rect 19540 685410 19560 685480
rect 19630 685410 19650 685480
rect 18050 685390 19650 685410
rect 70070 685370 71670 702320
rect 70068 685070 71670 685370
rect 121718 703830 123318 703900
rect 121718 703760 121788 703830
rect 121858 703760 121878 703830
rect 121948 703760 121968 703830
rect 122038 703760 122058 703830
rect 122128 703760 122148 703830
rect 122218 703760 122238 703830
rect 122308 703760 122328 703830
rect 122398 703760 122418 703830
rect 122488 703760 122508 703830
rect 122578 703760 122598 703830
rect 122668 703760 122688 703830
rect 122758 703760 122778 703830
rect 122848 703760 122868 703830
rect 122938 703760 122958 703830
rect 123028 703760 123048 703830
rect 123118 703760 123138 703830
rect 123208 703760 123228 703830
rect 123298 703760 123318 703830
rect 121718 703740 123318 703760
rect 121718 703670 121788 703740
rect 121858 703670 121878 703740
rect 121948 703670 121968 703740
rect 122038 703670 122058 703740
rect 122128 703670 122148 703740
rect 122218 703670 122238 703740
rect 122308 703670 122328 703740
rect 122398 703670 122418 703740
rect 122488 703670 122508 703740
rect 122578 703670 122598 703740
rect 122668 703670 122688 703740
rect 122758 703670 122778 703740
rect 122848 703670 122868 703740
rect 122938 703670 122958 703740
rect 123028 703670 123048 703740
rect 123118 703670 123138 703740
rect 123208 703670 123228 703740
rect 123298 703670 123318 703740
rect 121718 703650 123318 703670
rect 121718 703580 121788 703650
rect 121858 703580 121878 703650
rect 121948 703580 121968 703650
rect 122038 703580 122058 703650
rect 122128 703580 122148 703650
rect 122218 703580 122238 703650
rect 122308 703580 122328 703650
rect 122398 703580 122418 703650
rect 122488 703580 122508 703650
rect 122578 703580 122598 703650
rect 122668 703580 122688 703650
rect 122758 703580 122778 703650
rect 122848 703580 122868 703650
rect 122938 703580 122958 703650
rect 123028 703580 123048 703650
rect 123118 703580 123138 703650
rect 123208 703580 123228 703650
rect 123298 703580 123318 703650
rect 121718 703560 123318 703580
rect 121718 703490 121788 703560
rect 121858 703490 121878 703560
rect 121948 703490 121968 703560
rect 122038 703490 122058 703560
rect 122128 703490 122148 703560
rect 122218 703490 122238 703560
rect 122308 703490 122328 703560
rect 122398 703490 122418 703560
rect 122488 703490 122508 703560
rect 122578 703490 122598 703560
rect 122668 703490 122688 703560
rect 122758 703490 122778 703560
rect 122848 703490 122868 703560
rect 122938 703490 122958 703560
rect 123028 703490 123048 703560
rect 123118 703490 123138 703560
rect 123208 703490 123228 703560
rect 123298 703490 123318 703560
rect 121718 703470 123318 703490
rect 121718 703400 121788 703470
rect 121858 703400 121878 703470
rect 121948 703400 121968 703470
rect 122038 703400 122058 703470
rect 122128 703400 122148 703470
rect 122218 703400 122238 703470
rect 122308 703400 122328 703470
rect 122398 703400 122418 703470
rect 122488 703400 122508 703470
rect 122578 703400 122598 703470
rect 122668 703400 122688 703470
rect 122758 703400 122778 703470
rect 122848 703400 122868 703470
rect 122938 703400 122958 703470
rect 123028 703400 123048 703470
rect 123118 703400 123138 703470
rect 123208 703400 123228 703470
rect 123298 703400 123318 703470
rect 121718 703380 123318 703400
rect 121718 703310 121788 703380
rect 121858 703310 121878 703380
rect 121948 703310 121968 703380
rect 122038 703310 122058 703380
rect 122128 703310 122148 703380
rect 122218 703310 122238 703380
rect 122308 703310 122328 703380
rect 122398 703310 122418 703380
rect 122488 703310 122508 703380
rect 122578 703310 122598 703380
rect 122668 703310 122688 703380
rect 122758 703310 122778 703380
rect 122848 703310 122868 703380
rect 122938 703310 122958 703380
rect 123028 703310 123048 703380
rect 123118 703310 123138 703380
rect 123208 703310 123228 703380
rect 123298 703310 123318 703380
rect 121718 703290 123318 703310
rect 121718 703220 121788 703290
rect 121858 703220 121878 703290
rect 121948 703220 121968 703290
rect 122038 703220 122058 703290
rect 122128 703220 122148 703290
rect 122218 703220 122238 703290
rect 122308 703220 122328 703290
rect 122398 703220 122418 703290
rect 122488 703220 122508 703290
rect 122578 703220 122598 703290
rect 122668 703220 122688 703290
rect 122758 703220 122778 703290
rect 122848 703220 122868 703290
rect 122938 703220 122958 703290
rect 123028 703220 123048 703290
rect 123118 703220 123138 703290
rect 123208 703220 123228 703290
rect 123298 703220 123318 703290
rect 121718 703200 123318 703220
rect 121718 703130 121788 703200
rect 121858 703130 121878 703200
rect 121948 703130 121968 703200
rect 122038 703130 122058 703200
rect 122128 703130 122148 703200
rect 122218 703130 122238 703200
rect 122308 703130 122328 703200
rect 122398 703130 122418 703200
rect 122488 703130 122508 703200
rect 122578 703130 122598 703200
rect 122668 703130 122688 703200
rect 122758 703130 122778 703200
rect 122848 703130 122868 703200
rect 122938 703130 122958 703200
rect 123028 703130 123048 703200
rect 123118 703130 123138 703200
rect 123208 703130 123228 703200
rect 123298 703130 123318 703200
rect 121718 703110 123318 703130
rect 121718 703040 121788 703110
rect 121858 703040 121878 703110
rect 121948 703040 121968 703110
rect 122038 703040 122058 703110
rect 122128 703040 122148 703110
rect 122218 703040 122238 703110
rect 122308 703040 122328 703110
rect 122398 703040 122418 703110
rect 122488 703040 122508 703110
rect 122578 703040 122598 703110
rect 122668 703040 122688 703110
rect 122758 703040 122778 703110
rect 122848 703040 122868 703110
rect 122938 703040 122958 703110
rect 123028 703040 123048 703110
rect 123118 703040 123138 703110
rect 123208 703040 123228 703110
rect 123298 703040 123318 703110
rect 121718 703020 123318 703040
rect 121718 702950 121788 703020
rect 121858 702950 121878 703020
rect 121948 702950 121968 703020
rect 122038 702950 122058 703020
rect 122128 702950 122148 703020
rect 122218 702950 122238 703020
rect 122308 702950 122328 703020
rect 122398 702950 122418 703020
rect 122488 702950 122508 703020
rect 122578 702950 122598 703020
rect 122668 702950 122688 703020
rect 122758 702950 122778 703020
rect 122848 702950 122868 703020
rect 122938 702950 122958 703020
rect 123028 702950 123048 703020
rect 123118 702950 123138 703020
rect 123208 702950 123228 703020
rect 123298 702950 123318 703020
rect 121718 702930 123318 702950
rect 121718 702860 121788 702930
rect 121858 702860 121878 702930
rect 121948 702860 121968 702930
rect 122038 702860 122058 702930
rect 122128 702860 122148 702930
rect 122218 702860 122238 702930
rect 122308 702860 122328 702930
rect 122398 702860 122418 702930
rect 122488 702860 122508 702930
rect 122578 702860 122598 702930
rect 122668 702860 122688 702930
rect 122758 702860 122778 702930
rect 122848 702860 122868 702930
rect 122938 702860 122958 702930
rect 123028 702860 123048 702930
rect 123118 702860 123138 702930
rect 123208 702860 123228 702930
rect 123298 702860 123318 702930
rect 121718 702840 123318 702860
rect 121718 702770 121788 702840
rect 121858 702770 121878 702840
rect 121948 702770 121968 702840
rect 122038 702770 122058 702840
rect 122128 702770 122148 702840
rect 122218 702770 122238 702840
rect 122308 702770 122328 702840
rect 122398 702770 122418 702840
rect 122488 702770 122508 702840
rect 122578 702770 122598 702840
rect 122668 702770 122688 702840
rect 122758 702770 122778 702840
rect 122848 702770 122868 702840
rect 122938 702770 122958 702840
rect 123028 702770 123048 702840
rect 123118 702770 123138 702840
rect 123208 702770 123228 702840
rect 123298 702770 123318 702840
rect 121718 702750 123318 702770
rect 121718 702680 121788 702750
rect 121858 702680 121878 702750
rect 121948 702680 121968 702750
rect 122038 702680 122058 702750
rect 122128 702680 122148 702750
rect 122218 702680 122238 702750
rect 122308 702680 122328 702750
rect 122398 702680 122418 702750
rect 122488 702680 122508 702750
rect 122578 702680 122598 702750
rect 122668 702680 122688 702750
rect 122758 702680 122778 702750
rect 122848 702680 122868 702750
rect 122938 702680 122958 702750
rect 123028 702680 123048 702750
rect 123118 702680 123138 702750
rect 123208 702680 123228 702750
rect 123298 702680 123318 702750
rect 121718 702660 123318 702680
rect 121718 702590 121788 702660
rect 121858 702590 121878 702660
rect 121948 702590 121968 702660
rect 122038 702590 122058 702660
rect 122128 702590 122148 702660
rect 122218 702590 122238 702660
rect 122308 702590 122328 702660
rect 122398 702590 122418 702660
rect 122488 702590 122508 702660
rect 122578 702590 122598 702660
rect 122668 702590 122688 702660
rect 122758 702590 122778 702660
rect 122848 702590 122868 702660
rect 122938 702590 122958 702660
rect 123028 702590 123048 702660
rect 123118 702590 123138 702660
rect 123208 702590 123228 702660
rect 123298 702590 123318 702660
rect 121718 702570 123318 702590
rect 121718 702500 121788 702570
rect 121858 702500 121878 702570
rect 121948 702500 121968 702570
rect 122038 702500 122058 702570
rect 122128 702500 122148 702570
rect 122218 702500 122238 702570
rect 122308 702500 122328 702570
rect 122398 702500 122418 702570
rect 122488 702500 122508 702570
rect 122578 702500 122598 702570
rect 122668 702500 122688 702570
rect 122758 702500 122778 702570
rect 122848 702500 122868 702570
rect 122938 702500 122958 702570
rect 123028 702500 123048 702570
rect 123118 702500 123138 702570
rect 123208 702500 123228 702570
rect 123298 702500 123318 702570
rect 121718 702480 123318 702500
rect 121718 702410 121788 702480
rect 121858 702410 121878 702480
rect 121948 702410 121968 702480
rect 122038 702410 122058 702480
rect 122128 702410 122148 702480
rect 122218 702410 122238 702480
rect 122308 702410 122328 702480
rect 122398 702410 122418 702480
rect 122488 702410 122508 702480
rect 122578 702410 122598 702480
rect 122668 702410 122688 702480
rect 122758 702410 122778 702480
rect 122848 702410 122868 702480
rect 122938 702410 122958 702480
rect 123028 702410 123048 702480
rect 123118 702410 123138 702480
rect 123208 702410 123228 702480
rect 123298 702410 123318 702480
rect 121718 702390 123318 702410
rect 121718 702320 121788 702390
rect 121858 702320 121878 702390
rect 121948 702320 121968 702390
rect 122038 702320 122058 702390
rect 122128 702320 122148 702390
rect 122218 702320 122238 702390
rect 122308 702320 122328 702390
rect 122398 702320 122418 702390
rect 122488 702320 122508 702390
rect 122578 702320 122598 702390
rect 122668 702320 122688 702390
rect 122758 702320 122778 702390
rect 122848 702320 122868 702390
rect 122938 702320 122958 702390
rect 123028 702320 123048 702390
rect 123118 702320 123138 702390
rect 123208 702320 123228 702390
rect 123298 702320 123318 702390
rect 121718 685070 123318 702320
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 170894 692930 173094 693000
rect 170894 692690 170964 692930
rect 171204 692690 171294 692930
rect 171534 692690 171624 692930
rect 171864 692690 171954 692930
rect 172194 692690 172284 692930
rect 172524 692690 172614 692930
rect 172854 692690 173094 692930
rect 170894 692600 173094 692690
rect 170894 692360 170964 692600
rect 171204 692360 171294 692600
rect 171534 692360 171624 692600
rect 171864 692360 171954 692600
rect 172194 692360 172284 692600
rect 172524 692360 172614 692600
rect 172854 692360 173094 692600
rect 170894 692270 173094 692360
rect 170894 692030 170964 692270
rect 171204 692030 171294 692270
rect 171534 692030 171624 692270
rect 171864 692030 171954 692270
rect 172194 692030 172284 692270
rect 172524 692030 172614 692270
rect 172854 692030 173094 692270
rect 170894 691940 173094 692030
rect 170894 691700 170964 691940
rect 171204 691700 171294 691940
rect 171534 691700 171624 691940
rect 171864 691700 171954 691940
rect 172194 691700 172284 691940
rect 172524 691700 172614 691940
rect 172854 691700 173094 691940
rect 170894 691610 173094 691700
rect 170894 691370 170964 691610
rect 171204 691370 171294 691610
rect 171534 691370 171624 691610
rect 171864 691370 171954 691610
rect 172194 691370 172284 691610
rect 172524 691370 172614 691610
rect 172854 691370 173094 691610
rect 170894 691280 173094 691370
rect 170894 691040 170964 691280
rect 171204 691040 171294 691280
rect 171534 691040 171624 691280
rect 171864 691040 171954 691280
rect 172194 691040 172284 691280
rect 172524 691040 172614 691280
rect 172854 691040 173094 691280
rect 170894 690950 173094 691040
rect 170894 690710 170964 690950
rect 171204 690710 171294 690950
rect 171534 690710 171624 690950
rect 171864 690710 171954 690950
rect 172194 690710 172284 690950
rect 172524 690710 172614 690950
rect 172854 690710 173094 690950
rect 170894 690620 173094 690710
rect 170894 690380 170964 690620
rect 171204 690380 171294 690620
rect 171534 690380 171624 690620
rect 171864 690380 171954 690620
rect 172194 690380 172284 690620
rect 172524 690380 172614 690620
rect 172854 690380 173094 690620
rect 170894 690290 173094 690380
rect 170894 690050 170964 690290
rect 171204 690050 171294 690290
rect 171534 690050 171624 690290
rect 171864 690050 171954 690290
rect 172194 690050 172284 690290
rect 172524 690050 172614 690290
rect 172854 690050 173094 690290
rect 170894 689960 173094 690050
rect 170894 689720 170964 689960
rect 171204 689720 171294 689960
rect 171534 689720 171624 689960
rect 171864 689720 171954 689960
rect 172194 689720 172284 689960
rect 172524 689720 172614 689960
rect 172854 689720 173094 689960
rect 170894 689630 173094 689720
rect 170894 689390 170964 689630
rect 171204 689390 171294 689630
rect 171534 689390 171624 689630
rect 171864 689390 171954 689630
rect 172194 689390 172284 689630
rect 172524 689390 172614 689630
rect 172854 689390 173094 689630
rect 170894 689300 173094 689390
rect 170894 689060 170964 689300
rect 171204 689060 171294 689300
rect 171534 689060 171624 689300
rect 171864 689060 171954 689300
rect 172194 689060 172284 689300
rect 172524 689060 172614 689300
rect 172854 689060 173094 689300
rect 170894 688970 173094 689060
rect 170894 688730 170964 688970
rect 171204 688730 171294 688970
rect 171534 688730 171624 688970
rect 171864 688730 171954 688970
rect 172194 688730 172284 688970
rect 172524 688730 172614 688970
rect 172854 688730 173094 688970
rect 170894 688640 173094 688730
rect 170894 688400 170964 688640
rect 171204 688400 171294 688640
rect 171534 688400 171624 688640
rect 171864 688400 171954 688640
rect 172194 688400 172284 688640
rect 172524 688400 172614 688640
rect 172854 688400 173094 688640
rect 170894 688310 173094 688400
rect 170894 688070 170964 688310
rect 171204 688070 171294 688310
rect 171534 688070 171624 688310
rect 171864 688070 171954 688310
rect 172194 688070 172284 688310
rect 172524 688070 172614 688310
rect 172854 688070 173094 688310
rect 170894 688000 173094 688070
rect 217294 692930 222294 704800
rect 225094 700930 227294 701000
rect 225094 700690 225164 700930
rect 225404 700690 225494 700930
rect 225734 700690 225824 700930
rect 226064 700690 226154 700930
rect 226394 700690 226484 700930
rect 226724 700690 226814 700930
rect 227054 700690 227294 700930
rect 225094 700600 227294 700690
rect 225094 700360 225164 700600
rect 225404 700360 225494 700600
rect 225734 700360 225824 700600
rect 226064 700360 226154 700600
rect 226394 700360 226484 700600
rect 226724 700360 226814 700600
rect 227054 700360 227294 700600
rect 225094 700270 227294 700360
rect 225094 700030 225164 700270
rect 225404 700030 225494 700270
rect 225734 700030 225824 700270
rect 226064 700030 226154 700270
rect 226394 700030 226484 700270
rect 226724 700030 226814 700270
rect 227054 700030 227294 700270
rect 225094 699940 227294 700030
rect 225094 699700 225164 699940
rect 225404 699700 225494 699940
rect 225734 699700 225824 699940
rect 226064 699700 226154 699940
rect 226394 699700 226484 699940
rect 226724 699700 226814 699940
rect 227054 699700 227294 699940
rect 225094 699610 227294 699700
rect 225094 699370 225164 699610
rect 225404 699370 225494 699610
rect 225734 699370 225824 699610
rect 226064 699370 226154 699610
rect 226394 699370 226484 699610
rect 226724 699370 226814 699610
rect 227054 699370 227294 699610
rect 225094 699280 227294 699370
rect 225094 699040 225164 699280
rect 225404 699040 225494 699280
rect 225734 699040 225824 699280
rect 226064 699040 226154 699280
rect 226394 699040 226484 699280
rect 226724 699040 226814 699280
rect 227054 699040 227294 699280
rect 225094 698950 227294 699040
rect 225094 698710 225164 698950
rect 225404 698710 225494 698950
rect 225734 698710 225824 698950
rect 226064 698710 226154 698950
rect 226394 698710 226484 698950
rect 226724 698710 226814 698950
rect 227054 698710 227294 698950
rect 225094 698620 227294 698710
rect 225094 698380 225164 698620
rect 225404 698380 225494 698620
rect 225734 698380 225824 698620
rect 226064 698380 226154 698620
rect 226394 698380 226484 698620
rect 226724 698380 226814 698620
rect 227054 698380 227294 698620
rect 225094 698290 227294 698380
rect 225094 698050 225164 698290
rect 225404 698050 225494 698290
rect 225734 698050 225824 698290
rect 226064 698050 226154 698290
rect 226394 698050 226484 698290
rect 226724 698050 226814 698290
rect 227054 698050 227294 698290
rect 225094 697960 227294 698050
rect 225094 697720 225164 697960
rect 225404 697720 225494 697960
rect 225734 697720 225824 697960
rect 226064 697720 226154 697960
rect 226394 697720 226484 697960
rect 226724 697720 226814 697960
rect 227054 697720 227294 697960
rect 225094 697630 227294 697720
rect 225094 697390 225164 697630
rect 225404 697390 225494 697630
rect 225734 697390 225824 697630
rect 226064 697390 226154 697630
rect 226394 697390 226484 697630
rect 226724 697390 226814 697630
rect 227054 697390 227294 697630
rect 225094 697300 227294 697390
rect 225094 697060 225164 697300
rect 225404 697060 225494 697300
rect 225734 697060 225824 697300
rect 226064 697060 226154 697300
rect 226394 697060 226484 697300
rect 226724 697060 226814 697300
rect 227054 697060 227294 697300
rect 225094 696970 227294 697060
rect 225094 696730 225164 696970
rect 225404 696730 225494 696970
rect 225734 696730 225824 696970
rect 226064 696730 226154 696970
rect 226394 696730 226484 696970
rect 226724 696730 226814 696970
rect 227054 696730 227294 696970
rect 225094 696640 227294 696730
rect 225094 696400 225164 696640
rect 225404 696400 225494 696640
rect 225734 696400 225824 696640
rect 226064 696400 226154 696640
rect 226394 696400 226484 696640
rect 226724 696400 226814 696640
rect 227054 696400 227294 696640
rect 225094 696310 227294 696400
rect 225094 696070 225164 696310
rect 225404 696070 225494 696310
rect 225734 696070 225824 696310
rect 226064 696070 226154 696310
rect 226394 696070 226484 696310
rect 226724 696070 226814 696310
rect 227054 696070 227294 696310
rect 225094 696000 227294 696070
rect 217294 692690 217364 692930
rect 217604 692690 217694 692930
rect 217934 692690 218024 692930
rect 218264 692690 218354 692930
rect 218594 692690 218684 692930
rect 218924 692690 219014 692930
rect 219254 692690 219344 692930
rect 219584 692690 219674 692930
rect 219914 692690 220004 692930
rect 220244 692690 220334 692930
rect 220574 692690 220664 692930
rect 220904 692690 220994 692930
rect 221234 692690 221324 692930
rect 221564 692690 221654 692930
rect 221894 692690 221984 692930
rect 222224 692690 222294 692930
rect 217294 692600 222294 692690
rect 217294 692360 217364 692600
rect 217604 692360 217694 692600
rect 217934 692360 218024 692600
rect 218264 692360 218354 692600
rect 218594 692360 218684 692600
rect 218924 692360 219014 692600
rect 219254 692360 219344 692600
rect 219584 692360 219674 692600
rect 219914 692360 220004 692600
rect 220244 692360 220334 692600
rect 220574 692360 220664 692600
rect 220904 692360 220994 692600
rect 221234 692360 221324 692600
rect 221564 692360 221654 692600
rect 221894 692360 221984 692600
rect 222224 692360 222294 692600
rect 217294 692270 222294 692360
rect 217294 692030 217364 692270
rect 217604 692030 217694 692270
rect 217934 692030 218024 692270
rect 218264 692030 218354 692270
rect 218594 692030 218684 692270
rect 218924 692030 219014 692270
rect 219254 692030 219344 692270
rect 219584 692030 219674 692270
rect 219914 692030 220004 692270
rect 220244 692030 220334 692270
rect 220574 692030 220664 692270
rect 220904 692030 220994 692270
rect 221234 692030 221324 692270
rect 221564 692030 221654 692270
rect 221894 692030 221984 692270
rect 222224 692030 222294 692270
rect 217294 691940 222294 692030
rect 217294 691700 217364 691940
rect 217604 691700 217694 691940
rect 217934 691700 218024 691940
rect 218264 691700 218354 691940
rect 218594 691700 218684 691940
rect 218924 691700 219014 691940
rect 219254 691700 219344 691940
rect 219584 691700 219674 691940
rect 219914 691700 220004 691940
rect 220244 691700 220334 691940
rect 220574 691700 220664 691940
rect 220904 691700 220994 691940
rect 221234 691700 221324 691940
rect 221564 691700 221654 691940
rect 221894 691700 221984 691940
rect 222224 691700 222294 691940
rect 217294 691610 222294 691700
rect 217294 691370 217364 691610
rect 217604 691370 217694 691610
rect 217934 691370 218024 691610
rect 218264 691370 218354 691610
rect 218594 691370 218684 691610
rect 218924 691370 219014 691610
rect 219254 691370 219344 691610
rect 219584 691370 219674 691610
rect 219914 691370 220004 691610
rect 220244 691370 220334 691610
rect 220574 691370 220664 691610
rect 220904 691370 220994 691610
rect 221234 691370 221324 691610
rect 221564 691370 221654 691610
rect 221894 691370 221984 691610
rect 222224 691370 222294 691610
rect 217294 691280 222294 691370
rect 217294 691040 217364 691280
rect 217604 691040 217694 691280
rect 217934 691040 218024 691280
rect 218264 691040 218354 691280
rect 218594 691040 218684 691280
rect 218924 691040 219014 691280
rect 219254 691040 219344 691280
rect 219584 691040 219674 691280
rect 219914 691040 220004 691280
rect 220244 691040 220334 691280
rect 220574 691040 220664 691280
rect 220904 691040 220994 691280
rect 221234 691040 221324 691280
rect 221564 691040 221654 691280
rect 221894 691040 221984 691280
rect 222224 691040 222294 691280
rect 217294 690950 222294 691040
rect 217294 690710 217364 690950
rect 217604 690710 217694 690950
rect 217934 690710 218024 690950
rect 218264 690710 218354 690950
rect 218594 690710 218684 690950
rect 218924 690710 219014 690950
rect 219254 690710 219344 690950
rect 219584 690710 219674 690950
rect 219914 690710 220004 690950
rect 220244 690710 220334 690950
rect 220574 690710 220664 690950
rect 220904 690710 220994 690950
rect 221234 690710 221324 690950
rect 221564 690710 221654 690950
rect 221894 690710 221984 690950
rect 222224 690710 222294 690950
rect 217294 690620 222294 690710
rect 217294 690380 217364 690620
rect 217604 690380 217694 690620
rect 217934 690380 218024 690620
rect 218264 690380 218354 690620
rect 218594 690380 218684 690620
rect 218924 690380 219014 690620
rect 219254 690380 219344 690620
rect 219584 690380 219674 690620
rect 219914 690380 220004 690620
rect 220244 690380 220334 690620
rect 220574 690380 220664 690620
rect 220904 690380 220994 690620
rect 221234 690380 221324 690620
rect 221564 690380 221654 690620
rect 221894 690380 221984 690620
rect 222224 690380 222294 690620
rect 217294 690290 222294 690380
rect 217294 690050 217364 690290
rect 217604 690050 217694 690290
rect 217934 690050 218024 690290
rect 218264 690050 218354 690290
rect 218594 690050 218684 690290
rect 218924 690050 219014 690290
rect 219254 690050 219344 690290
rect 219584 690050 219674 690290
rect 219914 690050 220004 690290
rect 220244 690050 220334 690290
rect 220574 690050 220664 690290
rect 220904 690050 220994 690290
rect 221234 690050 221324 690290
rect 221564 690050 221654 690290
rect 221894 690050 221984 690290
rect 222224 690050 222294 690290
rect 217294 689960 222294 690050
rect 217294 689720 217364 689960
rect 217604 689720 217694 689960
rect 217934 689720 218024 689960
rect 218264 689720 218354 689960
rect 218594 689720 218684 689960
rect 218924 689720 219014 689960
rect 219254 689720 219344 689960
rect 219584 689720 219674 689960
rect 219914 689720 220004 689960
rect 220244 689720 220334 689960
rect 220574 689720 220664 689960
rect 220904 689720 220994 689960
rect 221234 689720 221324 689960
rect 221564 689720 221654 689960
rect 221894 689720 221984 689960
rect 222224 689720 222294 689960
rect 217294 689630 222294 689720
rect 217294 689390 217364 689630
rect 217604 689390 217694 689630
rect 217934 689390 218024 689630
rect 218264 689390 218354 689630
rect 218594 689390 218684 689630
rect 218924 689390 219014 689630
rect 219254 689390 219344 689630
rect 219584 689390 219674 689630
rect 219914 689390 220004 689630
rect 220244 689390 220334 689630
rect 220574 689390 220664 689630
rect 220904 689390 220994 689630
rect 221234 689390 221324 689630
rect 221564 689390 221654 689630
rect 221894 689390 221984 689630
rect 222224 689390 222294 689630
rect 217294 689300 222294 689390
rect 217294 689060 217364 689300
rect 217604 689060 217694 689300
rect 217934 689060 218024 689300
rect 218264 689060 218354 689300
rect 218594 689060 218684 689300
rect 218924 689060 219014 689300
rect 219254 689060 219344 689300
rect 219584 689060 219674 689300
rect 219914 689060 220004 689300
rect 220244 689060 220334 689300
rect 220574 689060 220664 689300
rect 220904 689060 220994 689300
rect 221234 689060 221324 689300
rect 221564 689060 221654 689300
rect 221894 689060 221984 689300
rect 222224 689060 222294 689300
rect 217294 688970 222294 689060
rect 217294 688730 217364 688970
rect 217604 688730 217694 688970
rect 217934 688730 218024 688970
rect 218264 688730 218354 688970
rect 218594 688730 218684 688970
rect 218924 688730 219014 688970
rect 219254 688730 219344 688970
rect 219584 688730 219674 688970
rect 219914 688730 220004 688970
rect 220244 688730 220334 688970
rect 220574 688730 220664 688970
rect 220904 688730 220994 688970
rect 221234 688730 221324 688970
rect 221564 688730 221654 688970
rect 221894 688730 221984 688970
rect 222224 688730 222294 688970
rect 217294 688640 222294 688730
rect 217294 688400 217364 688640
rect 217604 688400 217694 688640
rect 217934 688400 218024 688640
rect 218264 688400 218354 688640
rect 218594 688400 218684 688640
rect 218924 688400 219014 688640
rect 219254 688400 219344 688640
rect 219584 688400 219674 688640
rect 219914 688400 220004 688640
rect 220244 688400 220334 688640
rect 220574 688400 220664 688640
rect 220904 688400 220994 688640
rect 221234 688400 221324 688640
rect 221564 688400 221654 688640
rect 221894 688400 221984 688640
rect 222224 688400 222294 688640
rect 217294 688310 222294 688400
rect 217294 688070 217364 688310
rect 217604 688070 217694 688310
rect 217934 688070 218024 688310
rect 218264 688070 218354 688310
rect 218594 688070 218684 688310
rect 218924 688070 219014 688310
rect 219254 688070 219344 688310
rect 219584 688070 219674 688310
rect 219914 688070 220004 688310
rect 220244 688070 220334 688310
rect 220574 688070 220664 688310
rect 220904 688070 220994 688310
rect 221234 688070 221324 688310
rect 221564 688070 221654 688310
rect 221894 688070 221984 688310
rect 222224 688070 222294 688310
rect 217294 688000 222294 688070
rect 227594 692930 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 415610 702840 416180 702870
rect 415610 702770 415630 702840
rect 415700 702770 415720 702840
rect 415790 702770 415810 702840
rect 415880 702770 415900 702840
rect 415970 702770 415990 702840
rect 416060 702770 416080 702840
rect 416150 702770 416180 702840
rect 415610 702750 416180 702770
rect 415610 702680 415630 702750
rect 415700 702680 415720 702750
rect 415790 702680 415810 702750
rect 415880 702680 415900 702750
rect 415970 702680 415990 702750
rect 416060 702680 416080 702750
rect 416150 702680 416180 702750
rect 415610 702660 416180 702680
rect 415610 702590 415630 702660
rect 415700 702590 415720 702660
rect 415790 702590 415810 702660
rect 415880 702590 415900 702660
rect 415970 702590 415990 702660
rect 416060 702590 416080 702660
rect 416150 702590 416180 702660
rect 415610 702570 416180 702590
rect 415610 702500 415630 702570
rect 415700 702500 415720 702570
rect 415790 702500 415810 702570
rect 415880 702500 415900 702570
rect 415970 702500 415990 702570
rect 416060 702500 416080 702570
rect 416150 702500 416180 702570
rect 415610 702480 416180 702500
rect 415610 702410 415630 702480
rect 415700 702410 415720 702480
rect 415790 702410 415810 702480
rect 415880 702410 415900 702480
rect 415970 702410 415990 702480
rect 416060 702410 416080 702480
rect 416150 702410 416180 702480
rect 415610 702390 416180 702410
rect 415610 702320 415630 702390
rect 415700 702320 415720 702390
rect 415790 702320 415810 702390
rect 415880 702320 415900 702390
rect 415970 702320 415990 702390
rect 416060 702320 416080 702390
rect 416150 702320 416180 702390
rect 321210 697305 321780 702300
rect 415610 697305 416180 702320
rect 467610 702840 468180 702870
rect 467610 702770 467630 702840
rect 467700 702770 467720 702840
rect 467790 702770 467810 702840
rect 467880 702770 467900 702840
rect 467970 702770 467990 702840
rect 468060 702770 468080 702840
rect 468150 702770 468180 702840
rect 467610 702750 468180 702770
rect 467610 702680 467630 702750
rect 467700 702680 467720 702750
rect 467790 702680 467810 702750
rect 467880 702680 467900 702750
rect 467970 702680 467990 702750
rect 468060 702680 468080 702750
rect 468150 702680 468180 702750
rect 467610 702660 468180 702680
rect 467610 702590 467630 702660
rect 467700 702590 467720 702660
rect 467790 702590 467810 702660
rect 467880 702590 467900 702660
rect 467970 702590 467990 702660
rect 468060 702590 468080 702660
rect 468150 702590 468180 702660
rect 467610 702570 468180 702590
rect 467610 702500 467630 702570
rect 467700 702500 467720 702570
rect 467790 702500 467810 702570
rect 467880 702500 467900 702570
rect 467970 702500 467990 702570
rect 468060 702500 468080 702570
rect 468150 702500 468180 702570
rect 467610 702480 468180 702500
rect 467610 702410 467630 702480
rect 467700 702410 467720 702480
rect 467790 702410 467810 702480
rect 467880 702410 467900 702480
rect 467970 702410 467990 702480
rect 468060 702410 468080 702480
rect 468150 702410 468180 702480
rect 467610 702390 468180 702410
rect 467610 702320 467630 702390
rect 467700 702320 467720 702390
rect 467790 702320 467810 702390
rect 467880 702320 467900 702390
rect 467970 702320 467990 702390
rect 468060 702320 468080 702390
rect 468150 702320 468180 702390
rect 467610 697305 468180 702320
rect 566720 702840 567290 702870
rect 566720 702770 566740 702840
rect 566810 702770 566830 702840
rect 566900 702770 566920 702840
rect 566990 702770 567010 702840
rect 567080 702770 567100 702840
rect 567170 702770 567190 702840
rect 567260 702770 567290 702840
rect 566720 702750 567290 702770
rect 566720 702680 566740 702750
rect 566810 702680 566830 702750
rect 566900 702680 566920 702750
rect 566990 702680 567010 702750
rect 567080 702680 567100 702750
rect 567170 702680 567190 702750
rect 567260 702680 567290 702750
rect 566720 702660 567290 702680
rect 566720 702590 566740 702660
rect 566810 702590 566830 702660
rect 566900 702590 566920 702660
rect 566990 702590 567010 702660
rect 567080 702590 567100 702660
rect 567170 702590 567190 702660
rect 567260 702590 567290 702660
rect 566720 702570 567290 702590
rect 566720 702500 566740 702570
rect 566810 702500 566830 702570
rect 566900 702500 566920 702570
rect 566990 702500 567010 702570
rect 567080 702500 567100 702570
rect 567170 702500 567190 702570
rect 567260 702500 567290 702570
rect 566720 702480 567290 702500
rect 566720 702410 566740 702480
rect 566810 702410 566830 702480
rect 566900 702410 566920 702480
rect 566990 702410 567010 702480
rect 567080 702410 567100 702480
rect 567170 702410 567190 702480
rect 567260 702410 567290 702480
rect 566720 702390 567290 702410
rect 566720 702320 566740 702390
rect 566810 702320 566830 702390
rect 566900 702320 566920 702390
rect 566990 702320 567010 702390
rect 567080 702320 567100 702390
rect 567170 702320 567190 702390
rect 567260 702320 567290 702390
rect 566720 697305 567290 702320
rect 227594 692690 227664 692930
rect 227904 692690 227994 692930
rect 228234 692690 228324 692930
rect 228564 692690 228654 692930
rect 228894 692690 228984 692930
rect 229224 692690 229314 692930
rect 229554 692690 229644 692930
rect 229884 692690 229974 692930
rect 230214 692690 230304 692930
rect 230544 692690 230634 692930
rect 230874 692690 230964 692930
rect 231204 692690 231294 692930
rect 231534 692690 231624 692930
rect 231864 692690 231954 692930
rect 232194 692690 232284 692930
rect 232524 692690 232594 692930
rect 227594 692600 232594 692690
rect 227594 692360 227664 692600
rect 227904 692360 227994 692600
rect 228234 692360 228324 692600
rect 228564 692360 228654 692600
rect 228894 692360 228984 692600
rect 229224 692360 229314 692600
rect 229554 692360 229644 692600
rect 229884 692360 229974 692600
rect 230214 692360 230304 692600
rect 230544 692360 230634 692600
rect 230874 692360 230964 692600
rect 231204 692360 231294 692600
rect 231534 692360 231624 692600
rect 231864 692360 231954 692600
rect 232194 692360 232284 692600
rect 232524 692360 232594 692600
rect 227594 692270 232594 692360
rect 227594 692030 227664 692270
rect 227904 692030 227994 692270
rect 228234 692030 228324 692270
rect 228564 692030 228654 692270
rect 228894 692030 228984 692270
rect 229224 692030 229314 692270
rect 229554 692030 229644 692270
rect 229884 692030 229974 692270
rect 230214 692030 230304 692270
rect 230544 692030 230634 692270
rect 230874 692030 230964 692270
rect 231204 692030 231294 692270
rect 231534 692030 231624 692270
rect 231864 692030 231954 692270
rect 232194 692030 232284 692270
rect 232524 692030 232594 692270
rect 227594 691940 232594 692030
rect 227594 691700 227664 691940
rect 227904 691700 227994 691940
rect 228234 691700 228324 691940
rect 228564 691700 228654 691940
rect 228894 691700 228984 691940
rect 229224 691700 229314 691940
rect 229554 691700 229644 691940
rect 229884 691700 229974 691940
rect 230214 691700 230304 691940
rect 230544 691700 230634 691940
rect 230874 691700 230964 691940
rect 231204 691700 231294 691940
rect 231534 691700 231624 691940
rect 231864 691700 231954 691940
rect 232194 691700 232284 691940
rect 232524 691700 232594 691940
rect 227594 691610 232594 691700
rect 227594 691370 227664 691610
rect 227904 691370 227994 691610
rect 228234 691370 228324 691610
rect 228564 691370 228654 691610
rect 228894 691370 228984 691610
rect 229224 691370 229314 691610
rect 229554 691370 229644 691610
rect 229884 691370 229974 691610
rect 230214 691370 230304 691610
rect 230544 691370 230634 691610
rect 230874 691370 230964 691610
rect 231204 691370 231294 691610
rect 231534 691370 231624 691610
rect 231864 691370 231954 691610
rect 232194 691370 232284 691610
rect 232524 691370 232594 691610
rect 227594 691280 232594 691370
rect 227594 691040 227664 691280
rect 227904 691040 227994 691280
rect 228234 691040 228324 691280
rect 228564 691040 228654 691280
rect 228894 691040 228984 691280
rect 229224 691040 229314 691280
rect 229554 691040 229644 691280
rect 229884 691040 229974 691280
rect 230214 691040 230304 691280
rect 230544 691040 230634 691280
rect 230874 691040 230964 691280
rect 231204 691040 231294 691280
rect 231534 691040 231624 691280
rect 231864 691040 231954 691280
rect 232194 691040 232284 691280
rect 232524 691040 232594 691280
rect 227594 690950 232594 691040
rect 227594 690710 227664 690950
rect 227904 690710 227994 690950
rect 228234 690710 228324 690950
rect 228564 690710 228654 690950
rect 228894 690710 228984 690950
rect 229224 690710 229314 690950
rect 229554 690710 229644 690950
rect 229884 690710 229974 690950
rect 230214 690710 230304 690950
rect 230544 690710 230634 690950
rect 230874 690710 230964 690950
rect 231204 690710 231294 690950
rect 231534 690710 231624 690950
rect 231864 690710 231954 690950
rect 232194 690710 232284 690950
rect 232524 690710 232594 690950
rect 227594 690620 232594 690710
rect 227594 690380 227664 690620
rect 227904 690380 227994 690620
rect 228234 690380 228324 690620
rect 228564 690380 228654 690620
rect 228894 690380 228984 690620
rect 229224 690380 229314 690620
rect 229554 690380 229644 690620
rect 229884 690380 229974 690620
rect 230214 690380 230304 690620
rect 230544 690380 230634 690620
rect 230874 690380 230964 690620
rect 231204 690380 231294 690620
rect 231534 690380 231624 690620
rect 231864 690380 231954 690620
rect 232194 690380 232284 690620
rect 232524 690380 232594 690620
rect 227594 690290 232594 690380
rect 227594 690050 227664 690290
rect 227904 690050 227994 690290
rect 228234 690050 228324 690290
rect 228564 690050 228654 690290
rect 228894 690050 228984 690290
rect 229224 690050 229314 690290
rect 229554 690050 229644 690290
rect 229884 690050 229974 690290
rect 230214 690050 230304 690290
rect 230544 690050 230634 690290
rect 230874 690050 230964 690290
rect 231204 690050 231294 690290
rect 231534 690050 231624 690290
rect 231864 690050 231954 690290
rect 232194 690050 232284 690290
rect 232524 690050 232594 690290
rect 227594 689960 232594 690050
rect 227594 689720 227664 689960
rect 227904 689720 227994 689960
rect 228234 689720 228324 689960
rect 228564 689720 228654 689960
rect 228894 689720 228984 689960
rect 229224 689720 229314 689960
rect 229554 689720 229644 689960
rect 229884 689720 229974 689960
rect 230214 689720 230304 689960
rect 230544 689720 230634 689960
rect 230874 689720 230964 689960
rect 231204 689720 231294 689960
rect 231534 689720 231624 689960
rect 231864 689720 231954 689960
rect 232194 689720 232284 689960
rect 232524 689720 232594 689960
rect 227594 689630 232594 689720
rect 227594 689390 227664 689630
rect 227904 689390 227994 689630
rect 228234 689390 228324 689630
rect 228564 689390 228654 689630
rect 228894 689390 228984 689630
rect 229224 689390 229314 689630
rect 229554 689390 229644 689630
rect 229884 689390 229974 689630
rect 230214 689390 230304 689630
rect 230544 689390 230634 689630
rect 230874 689390 230964 689630
rect 231204 689390 231294 689630
rect 231534 689390 231624 689630
rect 231864 689390 231954 689630
rect 232194 689390 232284 689630
rect 232524 689390 232594 689630
rect 227594 689300 232594 689390
rect 227594 689060 227664 689300
rect 227904 689060 227994 689300
rect 228234 689060 228324 689300
rect 228564 689060 228654 689300
rect 228894 689060 228984 689300
rect 229224 689060 229314 689300
rect 229554 689060 229644 689300
rect 229884 689060 229974 689300
rect 230214 689060 230304 689300
rect 230544 689060 230634 689300
rect 230874 689060 230964 689300
rect 231204 689060 231294 689300
rect 231534 689060 231624 689300
rect 231864 689060 231954 689300
rect 232194 689060 232284 689300
rect 232524 689060 232594 689300
rect 227594 688970 232594 689060
rect 227594 688730 227664 688970
rect 227904 688730 227994 688970
rect 228234 688730 228324 688970
rect 228564 688730 228654 688970
rect 228894 688730 228984 688970
rect 229224 688730 229314 688970
rect 229554 688730 229644 688970
rect 229884 688730 229974 688970
rect 230214 688730 230304 688970
rect 230544 688730 230634 688970
rect 230874 688730 230964 688970
rect 231204 688730 231294 688970
rect 231534 688730 231624 688970
rect 231864 688730 231954 688970
rect 232194 688730 232284 688970
rect 232524 688730 232594 688970
rect 227594 688640 232594 688730
rect 227594 688400 227664 688640
rect 227904 688400 227994 688640
rect 228234 688400 228324 688640
rect 228564 688400 228654 688640
rect 228894 688400 228984 688640
rect 229224 688400 229314 688640
rect 229554 688400 229644 688640
rect 229884 688400 229974 688640
rect 230214 688400 230304 688640
rect 230544 688400 230634 688640
rect 230874 688400 230964 688640
rect 231204 688400 231294 688640
rect 231534 688400 231624 688640
rect 231864 688400 231954 688640
rect 232194 688400 232284 688640
rect 232524 688400 232594 688640
rect 227594 688310 232594 688400
rect 227594 688070 227664 688310
rect 227904 688070 227994 688310
rect 228234 688070 228324 688310
rect 228564 688070 228654 688310
rect 228894 688070 228984 688310
rect 229224 688070 229314 688310
rect 229554 688070 229644 688310
rect 229884 688070 229974 688310
rect 230214 688070 230304 688310
rect 230544 688070 230634 688310
rect 230874 688070 230964 688310
rect 231204 688070 231294 688310
rect 231534 688070 231624 688310
rect 231864 688070 231954 688310
rect 232194 688070 232284 688310
rect 232524 688070 232594 688310
rect 227594 688000 232594 688070
rect 321210 685238 321780 691785
rect 100 683660 8100 683730
rect 100 683590 120 683660
rect 190 683590 210 683660
rect 280 683590 300 683660
rect 370 683590 390 683660
rect 460 683590 480 683660
rect 550 683590 570 683660
rect 640 683590 660 683660
rect 730 683590 750 683660
rect 820 683590 840 683660
rect 910 683590 930 683660
rect 1000 683590 1020 683660
rect 1090 683590 1110 683660
rect 1180 683590 1200 683660
rect 1270 683590 1290 683660
rect 1360 683590 1380 683660
rect 1450 683590 1470 683660
rect 1540 683590 1560 683660
rect 1630 683590 8100 683660
rect 100 683570 8100 683590
rect 100 683500 120 683570
rect 190 683500 210 683570
rect 280 683500 300 683570
rect 370 683500 390 683570
rect 460 683500 480 683570
rect 550 683500 570 683570
rect 640 683500 660 683570
rect 730 683500 750 683570
rect 820 683500 840 683570
rect 910 683500 930 683570
rect 1000 683500 1020 683570
rect 1090 683500 1110 683570
rect 1180 683500 1200 683570
rect 1270 683500 1290 683570
rect 1360 683500 1380 683570
rect 1450 683500 1470 683570
rect 1540 683500 1560 683570
rect 1630 683500 8100 683570
rect 100 683480 8100 683500
rect 100 683410 120 683480
rect 190 683410 210 683480
rect 280 683410 300 683480
rect 370 683410 390 683480
rect 460 683410 480 683480
rect 550 683410 570 683480
rect 640 683410 660 683480
rect 730 683410 750 683480
rect 820 683410 840 683480
rect 910 683410 930 683480
rect 1000 683410 1020 683480
rect 1090 683410 1110 683480
rect 1180 683410 1200 683480
rect 1270 683410 1290 683480
rect 1360 683410 1380 683480
rect 1450 683410 1470 683480
rect 1540 683410 1560 683480
rect 1630 683410 8100 683480
rect 100 683390 8100 683410
rect 100 683320 120 683390
rect 190 683320 210 683390
rect 280 683320 300 683390
rect 370 683320 390 683390
rect 460 683320 480 683390
rect 550 683320 570 683390
rect 640 683320 660 683390
rect 730 683320 750 683390
rect 820 683320 840 683390
rect 910 683320 930 683390
rect 1000 683320 1020 683390
rect 1090 683320 1110 683390
rect 1180 683320 1200 683390
rect 1270 683320 1290 683390
rect 1360 683320 1380 683390
rect 1450 683320 1470 683390
rect 1540 683320 1560 683390
rect 1630 683320 8100 683390
rect 100 683300 8100 683320
rect 100 683230 120 683300
rect 190 683230 210 683300
rect 280 683230 300 683300
rect 370 683230 390 683300
rect 460 683230 480 683300
rect 550 683230 570 683300
rect 640 683230 660 683300
rect 730 683230 750 683300
rect 820 683230 840 683300
rect 910 683230 930 683300
rect 1000 683230 1020 683300
rect 1090 683230 1110 683300
rect 1180 683230 1200 683300
rect 1270 683230 1290 683300
rect 1360 683230 1380 683300
rect 1450 683230 1470 683300
rect 1540 683230 1560 683300
rect 1630 683230 8100 683300
rect 100 683210 8100 683230
rect 100 683140 120 683210
rect 190 683140 210 683210
rect 280 683140 300 683210
rect 370 683140 390 683210
rect 460 683140 480 683210
rect 550 683140 570 683210
rect 640 683140 660 683210
rect 730 683140 750 683210
rect 820 683140 840 683210
rect 910 683140 930 683210
rect 1000 683140 1020 683210
rect 1090 683140 1110 683210
rect 1180 683140 1200 683210
rect 1270 683140 1290 683210
rect 1360 683140 1380 683210
rect 1450 683140 1470 683210
rect 1540 683140 1560 683210
rect 1630 683140 8100 683210
rect 100 683120 8100 683140
rect 100 683050 120 683120
rect 190 683050 210 683120
rect 280 683050 300 683120
rect 370 683050 390 683120
rect 460 683050 480 683120
rect 550 683050 570 683120
rect 640 683050 660 683120
rect 730 683050 750 683120
rect 820 683050 840 683120
rect 910 683050 930 683120
rect 1000 683050 1020 683120
rect 1090 683050 1110 683120
rect 1180 683050 1200 683120
rect 1270 683050 1290 683120
rect 1360 683050 1380 683120
rect 1450 683050 1470 683120
rect 1540 683050 1560 683120
rect 1630 683050 8100 683120
rect 100 683030 8100 683050
rect 100 682960 120 683030
rect 190 682960 210 683030
rect 280 682960 300 683030
rect 370 682960 390 683030
rect 460 682960 480 683030
rect 550 682960 570 683030
rect 640 682960 660 683030
rect 730 682960 750 683030
rect 820 682960 840 683030
rect 910 682960 930 683030
rect 1000 682960 1020 683030
rect 1090 682960 1110 683030
rect 1180 682960 1200 683030
rect 1270 682960 1290 683030
rect 1360 682960 1380 683030
rect 1450 682960 1470 683030
rect 1540 682960 1560 683030
rect 1630 682960 8100 683030
rect 100 682940 8100 682960
rect 100 682870 120 682940
rect 190 682870 210 682940
rect 280 682870 300 682940
rect 370 682870 390 682940
rect 460 682870 480 682940
rect 550 682870 570 682940
rect 640 682870 660 682940
rect 730 682870 750 682940
rect 820 682870 840 682940
rect 910 682870 930 682940
rect 1000 682870 1020 682940
rect 1090 682870 1110 682940
rect 1180 682870 1200 682940
rect 1270 682870 1290 682940
rect 1360 682870 1380 682940
rect 1450 682870 1470 682940
rect 1540 682870 1560 682940
rect 1630 682870 8100 682940
rect 100 682850 8100 682870
rect 100 682780 120 682850
rect 190 682780 210 682850
rect 280 682780 300 682850
rect 370 682780 390 682850
rect 460 682780 480 682850
rect 550 682780 570 682850
rect 640 682780 660 682850
rect 730 682780 750 682850
rect 820 682780 840 682850
rect 910 682780 930 682850
rect 1000 682780 1020 682850
rect 1090 682780 1110 682850
rect 1180 682780 1200 682850
rect 1270 682780 1290 682850
rect 1360 682780 1380 682850
rect 1450 682780 1470 682850
rect 1540 682780 1560 682850
rect 1630 682780 8100 682850
rect 100 682760 8100 682780
rect 100 682690 120 682760
rect 190 682690 210 682760
rect 280 682690 300 682760
rect 370 682690 390 682760
rect 460 682690 480 682760
rect 550 682690 570 682760
rect 640 682690 660 682760
rect 730 682690 750 682760
rect 820 682690 840 682760
rect 910 682690 930 682760
rect 1000 682690 1020 682760
rect 1090 682690 1110 682760
rect 1180 682690 1200 682760
rect 1270 682690 1290 682760
rect 1360 682690 1380 682760
rect 1450 682690 1470 682760
rect 1540 682690 1560 682760
rect 1630 682690 8100 682760
rect 100 682670 8100 682690
rect 100 682600 120 682670
rect 190 682600 210 682670
rect 280 682600 300 682670
rect 370 682600 390 682670
rect 460 682600 480 682670
rect 550 682600 570 682670
rect 640 682600 660 682670
rect 730 682600 750 682670
rect 820 682600 840 682670
rect 910 682600 930 682670
rect 1000 682600 1020 682670
rect 1090 682600 1110 682670
rect 1180 682600 1200 682670
rect 1270 682600 1290 682670
rect 1360 682600 1380 682670
rect 1450 682600 1470 682670
rect 1540 682600 1560 682670
rect 1630 682600 8100 682670
rect 100 682580 8100 682600
rect 100 682510 120 682580
rect 190 682510 210 682580
rect 280 682510 300 682580
rect 370 682510 390 682580
rect 460 682510 480 682580
rect 550 682510 570 682580
rect 640 682510 660 682580
rect 730 682510 750 682580
rect 820 682510 840 682580
rect 910 682510 930 682580
rect 1000 682510 1020 682580
rect 1090 682510 1110 682580
rect 1180 682510 1200 682580
rect 1270 682510 1290 682580
rect 1360 682510 1380 682580
rect 1450 682510 1470 682580
rect 1540 682510 1560 682580
rect 1630 682510 8100 682580
rect 100 682490 8100 682510
rect 100 682420 120 682490
rect 190 682420 210 682490
rect 280 682420 300 682490
rect 370 682420 390 682490
rect 460 682420 480 682490
rect 550 682420 570 682490
rect 640 682420 660 682490
rect 730 682420 750 682490
rect 820 682420 840 682490
rect 910 682420 930 682490
rect 1000 682420 1020 682490
rect 1090 682420 1110 682490
rect 1180 682420 1200 682490
rect 1270 682420 1290 682490
rect 1360 682420 1380 682490
rect 1450 682420 1470 682490
rect 1540 682420 1560 682490
rect 1630 682420 8100 682490
rect 100 682400 8100 682420
rect 100 682330 120 682400
rect 190 682330 210 682400
rect 280 682330 300 682400
rect 370 682330 390 682400
rect 460 682330 480 682400
rect 550 682330 570 682400
rect 640 682330 660 682400
rect 730 682330 750 682400
rect 820 682330 840 682400
rect 910 682330 930 682400
rect 1000 682330 1020 682400
rect 1090 682330 1110 682400
rect 1180 682330 1200 682400
rect 1270 682330 1290 682400
rect 1360 682330 1380 682400
rect 1450 682330 1470 682400
rect 1540 682330 1560 682400
rect 1630 682330 8100 682400
rect 100 682310 8100 682330
rect 100 682240 120 682310
rect 190 682240 210 682310
rect 280 682240 300 682310
rect 370 682240 390 682310
rect 460 682240 480 682310
rect 550 682240 570 682310
rect 640 682240 660 682310
rect 730 682240 750 682310
rect 820 682240 840 682310
rect 910 682240 930 682310
rect 1000 682240 1020 682310
rect 1090 682240 1110 682310
rect 1180 682240 1200 682310
rect 1270 682240 1290 682310
rect 1360 682240 1380 682310
rect 1450 682240 1470 682310
rect 1540 682240 1560 682310
rect 1630 682240 8100 682310
rect 100 682220 8100 682240
rect 100 682150 120 682220
rect 190 682150 210 682220
rect 280 682150 300 682220
rect 370 682150 390 682220
rect 460 682150 480 682220
rect 550 682150 570 682220
rect 640 682150 660 682220
rect 730 682150 750 682220
rect 820 682150 840 682220
rect 910 682150 930 682220
rect 1000 682150 1020 682220
rect 1090 682150 1110 682220
rect 1180 682150 1200 682220
rect 1270 682150 1290 682220
rect 1360 682150 1380 682220
rect 1450 682150 1470 682220
rect 1540 682150 1560 682220
rect 1630 682150 8100 682220
rect 100 682130 8100 682150
rect 10770 683660 19650 683730
rect 10770 683590 17670 683660
rect 17740 683590 17760 683660
rect 17830 683590 17850 683660
rect 17920 683590 17940 683660
rect 18010 683590 18030 683660
rect 18100 683590 18120 683660
rect 18190 683590 18210 683660
rect 18280 683590 18300 683660
rect 18370 683590 18390 683660
rect 18460 683590 18480 683660
rect 18550 683590 18570 683660
rect 18640 683590 18660 683660
rect 18730 683590 18750 683660
rect 18820 683590 18840 683660
rect 18910 683590 18930 683660
rect 19000 683590 19020 683660
rect 19090 683590 19110 683660
rect 19180 683590 19200 683660
rect 19270 683590 19290 683660
rect 19360 683590 19380 683660
rect 19450 683590 19470 683660
rect 19540 683590 19560 683660
rect 19630 683590 19650 683660
rect 10770 683570 19650 683590
rect 10770 683500 17670 683570
rect 17740 683500 17760 683570
rect 17830 683500 17850 683570
rect 17920 683500 17940 683570
rect 18010 683500 18030 683570
rect 18100 683500 18120 683570
rect 18190 683500 18210 683570
rect 18280 683500 18300 683570
rect 18370 683500 18390 683570
rect 18460 683500 18480 683570
rect 18550 683500 18570 683570
rect 18640 683500 18660 683570
rect 18730 683500 18750 683570
rect 18820 683500 18840 683570
rect 18910 683500 18930 683570
rect 19000 683500 19020 683570
rect 19090 683500 19110 683570
rect 19180 683500 19200 683570
rect 19270 683500 19290 683570
rect 19360 683500 19380 683570
rect 19450 683500 19470 683570
rect 19540 683500 19560 683570
rect 19630 683500 19650 683570
rect 10770 683480 19650 683500
rect 10770 683410 17670 683480
rect 17740 683410 17760 683480
rect 17830 683410 17850 683480
rect 17920 683410 17940 683480
rect 18010 683410 18030 683480
rect 18100 683410 18120 683480
rect 18190 683410 18210 683480
rect 18280 683410 18300 683480
rect 18370 683410 18390 683480
rect 18460 683410 18480 683480
rect 18550 683410 18570 683480
rect 18640 683410 18660 683480
rect 18730 683410 18750 683480
rect 18820 683410 18840 683480
rect 18910 683410 18930 683480
rect 19000 683410 19020 683480
rect 19090 683410 19110 683480
rect 19180 683410 19200 683480
rect 19270 683410 19290 683480
rect 19360 683410 19380 683480
rect 19450 683410 19470 683480
rect 19540 683410 19560 683480
rect 19630 683410 19650 683480
rect 70068 683470 96534 685070
rect 96854 683470 123320 685070
rect 131494 684668 321780 685238
rect 10770 683390 19650 683410
rect 10770 683320 17670 683390
rect 17740 683320 17760 683390
rect 17830 683320 17850 683390
rect 17920 683320 17940 683390
rect 18010 683320 18030 683390
rect 18100 683320 18120 683390
rect 18190 683320 18210 683390
rect 18280 683320 18300 683390
rect 18370 683320 18390 683390
rect 18460 683320 18480 683390
rect 18550 683320 18570 683390
rect 18640 683320 18660 683390
rect 18730 683320 18750 683390
rect 18820 683320 18840 683390
rect 18910 683320 18930 683390
rect 19000 683320 19020 683390
rect 19090 683320 19110 683390
rect 19180 683320 19200 683390
rect 19270 683320 19290 683390
rect 19360 683320 19380 683390
rect 19450 683320 19470 683390
rect 19540 683320 19560 683390
rect 19630 683320 19650 683390
rect 10770 683300 19650 683320
rect 10770 683230 17670 683300
rect 17740 683230 17760 683300
rect 17830 683230 17850 683300
rect 17920 683230 17940 683300
rect 18010 683230 18030 683300
rect 18100 683230 18120 683300
rect 18190 683230 18210 683300
rect 18280 683230 18300 683300
rect 18370 683230 18390 683300
rect 18460 683230 18480 683300
rect 18550 683230 18570 683300
rect 18640 683230 18660 683300
rect 18730 683230 18750 683300
rect 18820 683230 18840 683300
rect 18910 683230 18930 683300
rect 19000 683230 19020 683300
rect 19090 683230 19110 683300
rect 19180 683230 19200 683300
rect 19270 683230 19290 683300
rect 19360 683230 19380 683300
rect 19450 683230 19470 683300
rect 19540 683230 19560 683300
rect 19630 683230 19650 683300
rect 10770 683210 19650 683230
rect 10770 683140 17670 683210
rect 17740 683140 17760 683210
rect 17830 683140 17850 683210
rect 17920 683140 17940 683210
rect 18010 683140 18030 683210
rect 18100 683140 18120 683210
rect 18190 683140 18210 683210
rect 18280 683140 18300 683210
rect 18370 683140 18390 683210
rect 18460 683140 18480 683210
rect 18550 683140 18570 683210
rect 18640 683140 18660 683210
rect 18730 683140 18750 683210
rect 18820 683140 18840 683210
rect 18910 683140 18930 683210
rect 19000 683140 19020 683210
rect 19090 683140 19110 683210
rect 19180 683140 19200 683210
rect 19270 683140 19290 683210
rect 19360 683140 19380 683210
rect 19450 683140 19470 683210
rect 19540 683140 19560 683210
rect 19630 683140 19650 683210
rect 10770 683120 19650 683140
rect 10770 683050 17670 683120
rect 17740 683050 17760 683120
rect 17830 683050 17850 683120
rect 17920 683050 17940 683120
rect 18010 683050 18030 683120
rect 18100 683050 18120 683120
rect 18190 683050 18210 683120
rect 18280 683050 18300 683120
rect 18370 683050 18390 683120
rect 18460 683050 18480 683120
rect 18550 683050 18570 683120
rect 18640 683050 18660 683120
rect 18730 683050 18750 683120
rect 18820 683050 18840 683120
rect 18910 683050 18930 683120
rect 19000 683050 19020 683120
rect 19090 683050 19110 683120
rect 19180 683050 19200 683120
rect 19270 683050 19290 683120
rect 19360 683050 19380 683120
rect 19450 683050 19470 683120
rect 19540 683050 19560 683120
rect 19630 683050 19650 683120
rect 10770 683030 19650 683050
rect 10770 682960 17670 683030
rect 17740 682960 17760 683030
rect 17830 682960 17850 683030
rect 17920 682960 17940 683030
rect 18010 682960 18030 683030
rect 18100 682960 18120 683030
rect 18190 682960 18210 683030
rect 18280 682960 18300 683030
rect 18370 682960 18390 683030
rect 18460 682960 18480 683030
rect 18550 682960 18570 683030
rect 18640 682960 18660 683030
rect 18730 682960 18750 683030
rect 18820 682960 18840 683030
rect 18910 682960 18930 683030
rect 19000 682960 19020 683030
rect 19090 682960 19110 683030
rect 19180 682960 19200 683030
rect 19270 682960 19290 683030
rect 19360 682960 19380 683030
rect 19450 682960 19470 683030
rect 19540 682960 19560 683030
rect 19630 682960 19650 683030
rect 10770 682940 19650 682960
rect 10770 682870 17670 682940
rect 17740 682870 17760 682940
rect 17830 682870 17850 682940
rect 17920 682870 17940 682940
rect 18010 682870 18030 682940
rect 18100 682870 18120 682940
rect 18190 682870 18210 682940
rect 18280 682870 18300 682940
rect 18370 682870 18390 682940
rect 18460 682870 18480 682940
rect 18550 682870 18570 682940
rect 18640 682870 18660 682940
rect 18730 682870 18750 682940
rect 18820 682870 18840 682940
rect 18910 682870 18930 682940
rect 19000 682870 19020 682940
rect 19090 682870 19110 682940
rect 19180 682870 19200 682940
rect 19270 682870 19290 682940
rect 19360 682870 19380 682940
rect 19450 682870 19470 682940
rect 19540 682870 19560 682940
rect 19630 682870 19650 682940
rect 10770 682850 19650 682870
rect 10770 682780 17670 682850
rect 17740 682780 17760 682850
rect 17830 682780 17850 682850
rect 17920 682780 17940 682850
rect 18010 682780 18030 682850
rect 18100 682780 18120 682850
rect 18190 682780 18210 682850
rect 18280 682780 18300 682850
rect 18370 682780 18390 682850
rect 18460 682780 18480 682850
rect 18550 682780 18570 682850
rect 18640 682780 18660 682850
rect 18730 682780 18750 682850
rect 18820 682780 18840 682850
rect 18910 682780 18930 682850
rect 19000 682780 19020 682850
rect 19090 682780 19110 682850
rect 19180 682780 19200 682850
rect 19270 682780 19290 682850
rect 19360 682780 19380 682850
rect 19450 682780 19470 682850
rect 19540 682780 19560 682850
rect 19630 682780 19650 682850
rect 10770 682760 19650 682780
rect 10770 682690 17670 682760
rect 17740 682690 17760 682760
rect 17830 682690 17850 682760
rect 17920 682690 17940 682760
rect 18010 682690 18030 682760
rect 18100 682690 18120 682760
rect 18190 682690 18210 682760
rect 18280 682690 18300 682760
rect 18370 682690 18390 682760
rect 18460 682690 18480 682760
rect 18550 682690 18570 682760
rect 18640 682690 18660 682760
rect 18730 682690 18750 682760
rect 18820 682690 18840 682760
rect 18910 682690 18930 682760
rect 19000 682690 19020 682760
rect 19090 682690 19110 682760
rect 19180 682690 19200 682760
rect 19270 682690 19290 682760
rect 19360 682690 19380 682760
rect 19450 682690 19470 682760
rect 19540 682690 19560 682760
rect 19630 682690 19650 682760
rect 10770 682670 19650 682690
rect 10770 682600 17670 682670
rect 17740 682600 17760 682670
rect 17830 682600 17850 682670
rect 17920 682600 17940 682670
rect 18010 682600 18030 682670
rect 18100 682600 18120 682670
rect 18190 682600 18210 682670
rect 18280 682600 18300 682670
rect 18370 682600 18390 682670
rect 18460 682600 18480 682670
rect 18550 682600 18570 682670
rect 18640 682600 18660 682670
rect 18730 682600 18750 682670
rect 18820 682600 18840 682670
rect 18910 682600 18930 682670
rect 19000 682600 19020 682670
rect 19090 682600 19110 682670
rect 19180 682600 19200 682670
rect 19270 682600 19290 682670
rect 19360 682600 19380 682670
rect 19450 682600 19470 682670
rect 19540 682600 19560 682670
rect 19630 682600 19650 682670
rect 10770 682580 19650 682600
rect 10770 682510 17670 682580
rect 17740 682510 17760 682580
rect 17830 682510 17850 682580
rect 17920 682510 17940 682580
rect 18010 682510 18030 682580
rect 18100 682510 18120 682580
rect 18190 682510 18210 682580
rect 18280 682510 18300 682580
rect 18370 682510 18390 682580
rect 18460 682510 18480 682580
rect 18550 682510 18570 682580
rect 18640 682510 18660 682580
rect 18730 682510 18750 682580
rect 18820 682510 18840 682580
rect 18910 682510 18930 682580
rect 19000 682510 19020 682580
rect 19090 682510 19110 682580
rect 19180 682510 19200 682580
rect 19270 682510 19290 682580
rect 19360 682510 19380 682580
rect 19450 682510 19470 682580
rect 19540 682510 19560 682580
rect 19630 682510 19650 682580
rect 10770 682490 19650 682510
rect 10770 682420 17670 682490
rect 17740 682420 17760 682490
rect 17830 682420 17850 682490
rect 17920 682420 17940 682490
rect 18010 682420 18030 682490
rect 18100 682420 18120 682490
rect 18190 682420 18210 682490
rect 18280 682420 18300 682490
rect 18370 682420 18390 682490
rect 18460 682420 18480 682490
rect 18550 682420 18570 682490
rect 18640 682420 18660 682490
rect 18730 682420 18750 682490
rect 18820 682420 18840 682490
rect 18910 682420 18930 682490
rect 19000 682420 19020 682490
rect 19090 682420 19110 682490
rect 19180 682420 19200 682490
rect 19270 682420 19290 682490
rect 19360 682420 19380 682490
rect 19450 682420 19470 682490
rect 19540 682420 19560 682490
rect 19630 682420 19650 682490
rect 10770 682400 19650 682420
rect 10770 682330 17670 682400
rect 17740 682330 17760 682400
rect 17830 682330 17850 682400
rect 17920 682330 17940 682400
rect 18010 682330 18030 682400
rect 18100 682330 18120 682400
rect 18190 682330 18210 682400
rect 18280 682330 18300 682400
rect 18370 682330 18390 682400
rect 18460 682330 18480 682400
rect 18550 682330 18570 682400
rect 18640 682330 18660 682400
rect 18730 682330 18750 682400
rect 18820 682330 18840 682400
rect 18910 682330 18930 682400
rect 19000 682330 19020 682400
rect 19090 682330 19110 682400
rect 19180 682330 19200 682400
rect 19270 682330 19290 682400
rect 19360 682330 19380 682400
rect 19450 682330 19470 682400
rect 19540 682330 19560 682400
rect 19630 682330 19650 682400
rect 10770 682310 19650 682330
rect 10770 682240 17670 682310
rect 17740 682240 17760 682310
rect 17830 682240 17850 682310
rect 17920 682240 17940 682310
rect 18010 682240 18030 682310
rect 18100 682240 18120 682310
rect 18190 682240 18210 682310
rect 18280 682240 18300 682310
rect 18370 682240 18390 682310
rect 18460 682240 18480 682310
rect 18550 682240 18570 682310
rect 18640 682240 18660 682310
rect 18730 682240 18750 682310
rect 18820 682240 18840 682310
rect 18910 682240 18930 682310
rect 19000 682240 19020 682310
rect 19090 682240 19110 682310
rect 19180 682240 19200 682310
rect 19270 682240 19290 682310
rect 19360 682240 19380 682310
rect 19450 682240 19470 682310
rect 19540 682240 19560 682310
rect 19630 682240 19650 682310
rect 10770 682220 19650 682240
rect 10770 682150 17670 682220
rect 17740 682150 17760 682220
rect 17830 682150 17850 682220
rect 17920 682150 17940 682220
rect 18010 682150 18030 682220
rect 18100 682150 18120 682220
rect 18190 682150 18210 682220
rect 18280 682150 18300 682220
rect 18370 682150 18390 682220
rect 18460 682150 18480 682220
rect 18550 682150 18570 682220
rect 18640 682150 18660 682220
rect 18730 682150 18750 682220
rect 18820 682150 18840 682220
rect 18910 682150 18930 682220
rect 19000 682150 19020 682220
rect 19090 682150 19110 682220
rect 19180 682150 19200 682220
rect 19270 682150 19290 682220
rect 19360 682150 19380 682220
rect 19450 682150 19470 682220
rect 19540 682150 19560 682220
rect 19630 682150 19650 682220
rect 10770 682130 19650 682150
rect 131494 672440 132064 684668
rect 415610 684024 416180 691785
rect 110364 671870 132064 672440
rect 132936 683454 416180 684024
rect 110364 670830 110524 671870
rect 132936 670950 133506 683454
rect 467610 682866 468180 691785
rect 111044 670380 133506 670950
rect 134191 682296 468180 682866
rect 27350 668910 85310 669188
rect 27350 668670 82750 668910
rect 82990 668670 83080 668910
rect 83320 668670 83410 668910
rect 83650 668670 83770 668910
rect 84010 668670 84100 668910
rect 84340 668670 84460 668910
rect 84700 668670 84790 668910
rect 85030 668670 85310 668910
rect 27350 668580 85310 668670
rect 27350 668340 82750 668580
rect 82990 668340 83080 668580
rect 83320 668340 83410 668580
rect 83650 668340 83770 668580
rect 84010 668340 84100 668580
rect 84340 668340 84460 668580
rect 84700 668340 84790 668580
rect 85030 668340 85310 668580
rect 27350 668250 85310 668340
rect 27350 668010 82750 668250
rect 82990 668010 83080 668250
rect 83320 668010 83410 668250
rect 83650 668010 83770 668250
rect 84010 668010 84100 668250
rect 84340 668010 84460 668250
rect 84700 668010 84790 668250
rect 85030 668010 85310 668250
rect 27350 667890 85310 668010
rect 27350 667650 82750 667890
rect 82990 667650 83080 667890
rect 83320 667650 83410 667890
rect 83650 667650 83770 667890
rect 84010 667650 84100 667890
rect 84340 667650 84460 667890
rect 84700 667650 84790 667890
rect 85030 667650 85310 667890
rect 27350 667560 85310 667650
rect 27350 667320 82750 667560
rect 82990 667320 83080 667560
rect 83320 667320 83410 667560
rect 83650 667320 83770 667560
rect 84010 667320 84100 667560
rect 84340 667320 84460 667560
rect 84700 667320 84790 667560
rect 85030 667320 85310 667560
rect 27350 667200 85310 667320
rect 27350 666960 82750 667200
rect 82990 666960 83080 667200
rect 83320 666960 83410 667200
rect 83650 666960 83770 667200
rect 84010 666960 84100 667200
rect 84340 666960 84460 667200
rect 84700 666960 84790 667200
rect 85030 666960 85310 667200
rect 27350 666870 85310 666960
rect 27350 666630 82750 666870
rect 82990 666630 83080 666870
rect 83320 666630 83410 666870
rect 83650 666630 83770 666870
rect 84010 666630 84100 666870
rect 84340 666630 84460 666870
rect 84700 666630 84790 666870
rect 85030 666630 85310 666870
rect 27350 666510 85310 666630
rect 27350 666270 82750 666510
rect 82990 666270 83080 666510
rect 83320 666270 83410 666510
rect 83650 666270 83770 666510
rect 84010 666270 84100 666510
rect 84340 666270 84460 666510
rect 84700 666270 84790 666510
rect 85030 666270 85310 666510
rect 27350 666180 85310 666270
rect 27350 665940 82750 666180
rect 82990 665940 83080 666180
rect 83320 665940 83410 666180
rect 83650 665940 83770 666180
rect 84010 665940 84100 666180
rect 84340 665940 84460 666180
rect 84700 665940 84790 666180
rect 85030 665940 85310 666180
rect 27350 665820 85310 665940
rect 27350 665580 82750 665820
rect 82990 665580 83080 665820
rect 83320 665580 83410 665820
rect 83650 665580 83770 665820
rect 84010 665580 84100 665820
rect 84340 665580 84460 665820
rect 84700 665580 84790 665820
rect 85030 665580 85310 665820
rect 27350 665490 85310 665580
rect 27350 665250 82750 665490
rect 82990 665250 83080 665490
rect 83320 665250 83410 665490
rect 83650 665250 83770 665490
rect 84010 665250 84100 665490
rect 84340 665250 84460 665490
rect 84700 665250 84790 665490
rect 85030 665250 85310 665490
rect 27350 665130 85310 665250
rect 27350 664890 82750 665130
rect 82990 664890 83080 665130
rect 83320 664890 83410 665130
rect 83650 664890 83770 665130
rect 84010 664890 84100 665130
rect 84340 664890 84460 665130
rect 84700 664890 84790 665130
rect 85030 664890 85310 665130
rect 27350 664800 85310 664890
rect 27350 664560 82750 664800
rect 82990 664560 83080 664800
rect 83320 664560 83410 664800
rect 83650 664560 83770 664800
rect 84010 664560 84100 664800
rect 84340 664560 84460 664800
rect 84700 664560 84790 664800
rect 85030 664560 85310 664800
rect 27350 664470 85310 664560
rect 27350 664230 82750 664470
rect 82990 664230 83080 664470
rect 83320 664230 83410 664470
rect 83650 664230 83770 664470
rect 84010 664230 84100 664470
rect 84340 664230 84460 664470
rect 84700 664230 84790 664470
rect 85030 664230 85310 664470
rect 27350 664192 85310 664230
rect 27350 657307 32350 664192
rect 34110 657307 85310 657308
rect 27350 657030 85310 657307
rect 27350 656790 82750 657030
rect 82990 656790 83080 657030
rect 83320 656790 83410 657030
rect 83650 656790 83770 657030
rect 84010 656790 84100 657030
rect 84340 656790 84460 657030
rect 84700 656790 84790 657030
rect 85030 656790 85310 657030
rect 27350 656700 85310 656790
rect 27350 656460 82750 656700
rect 82990 656460 83080 656700
rect 83320 656460 83410 656700
rect 83650 656460 83770 656700
rect 84010 656460 84100 656700
rect 84340 656460 84460 656700
rect 84700 656460 84790 656700
rect 85030 656460 85310 656700
rect 27350 656370 85310 656460
rect 27350 656130 82750 656370
rect 82990 656130 83080 656370
rect 83320 656130 83410 656370
rect 83650 656130 83770 656370
rect 84010 656130 84100 656370
rect 84340 656130 84460 656370
rect 84700 656130 84790 656370
rect 85030 656130 85310 656370
rect 27350 656010 85310 656130
rect 27350 656000 82750 656010
rect 3000 655930 82750 656000
rect 3000 655690 3070 655930
rect 3310 655690 3400 655930
rect 3640 655690 3730 655930
rect 3970 655690 4060 655930
rect 4300 655690 4390 655930
rect 4630 655690 4720 655930
rect 4960 655690 5050 655930
rect 5290 655690 5380 655930
rect 5620 655690 5710 655930
rect 5950 655690 6040 655930
rect 6280 655690 6370 655930
rect 6610 655690 6700 655930
rect 6940 655690 7030 655930
rect 7270 655690 7360 655930
rect 7600 655690 7690 655930
rect 7930 655770 82750 655930
rect 82990 655770 83080 656010
rect 83320 655770 83410 656010
rect 83650 655770 83770 656010
rect 84010 655770 84100 656010
rect 84340 655770 84460 656010
rect 84700 655770 84790 656010
rect 85030 655770 85310 656010
rect 7930 655690 85310 655770
rect 3000 655680 85310 655690
rect 3000 655600 82750 655680
rect 3000 655360 3070 655600
rect 3310 655360 3400 655600
rect 3640 655360 3730 655600
rect 3970 655360 4060 655600
rect 4300 655360 4390 655600
rect 4630 655360 4720 655600
rect 4960 655360 5050 655600
rect 5290 655360 5380 655600
rect 5620 655360 5710 655600
rect 5950 655360 6040 655600
rect 6280 655360 6370 655600
rect 6610 655360 6700 655600
rect 6940 655360 7030 655600
rect 7270 655360 7360 655600
rect 7600 655360 7690 655600
rect 7930 655440 82750 655600
rect 82990 655440 83080 655680
rect 83320 655440 83410 655680
rect 83650 655440 83770 655680
rect 84010 655440 84100 655680
rect 84340 655440 84460 655680
rect 84700 655440 84790 655680
rect 85030 655440 85310 655680
rect 7930 655360 85310 655440
rect 3000 655320 85310 655360
rect 3000 655270 82750 655320
rect 3000 655030 3070 655270
rect 3310 655030 3400 655270
rect 3640 655030 3730 655270
rect 3970 655030 4060 655270
rect 4300 655030 4390 655270
rect 4630 655030 4720 655270
rect 4960 655030 5050 655270
rect 5290 655030 5380 655270
rect 5620 655030 5710 655270
rect 5950 655030 6040 655270
rect 6280 655030 6370 655270
rect 6610 655030 6700 655270
rect 6940 655030 7030 655270
rect 7270 655030 7360 655270
rect 7600 655030 7690 655270
rect 7930 655080 82750 655270
rect 82990 655080 83080 655320
rect 83320 655080 83410 655320
rect 83650 655080 83770 655320
rect 84010 655080 84100 655320
rect 84340 655080 84460 655320
rect 84700 655080 84790 655320
rect 85030 655080 85310 655320
rect 7930 655030 85310 655080
rect 3000 654990 85310 655030
rect 3000 654940 82750 654990
rect 3000 654700 3070 654940
rect 3310 654700 3400 654940
rect 3640 654700 3730 654940
rect 3970 654700 4060 654940
rect 4300 654700 4390 654940
rect 4630 654700 4720 654940
rect 4960 654700 5050 654940
rect 5290 654700 5380 654940
rect 5620 654700 5710 654940
rect 5950 654700 6040 654940
rect 6280 654700 6370 654940
rect 6610 654700 6700 654940
rect 6940 654700 7030 654940
rect 7270 654700 7360 654940
rect 7600 654700 7690 654940
rect 7930 654750 82750 654940
rect 82990 654750 83080 654990
rect 83320 654750 83410 654990
rect 83650 654750 83770 654990
rect 84010 654750 84100 654990
rect 84340 654750 84460 654990
rect 84700 654750 84790 654990
rect 85030 654750 85310 654990
rect 7930 654700 85310 654750
rect 3000 654630 85310 654700
rect 3000 654610 82750 654630
rect 3000 654370 3070 654610
rect 3310 654370 3400 654610
rect 3640 654370 3730 654610
rect 3970 654370 4060 654610
rect 4300 654370 4390 654610
rect 4630 654370 4720 654610
rect 4960 654370 5050 654610
rect 5290 654370 5380 654610
rect 5620 654370 5710 654610
rect 5950 654370 6040 654610
rect 6280 654370 6370 654610
rect 6610 654370 6700 654610
rect 6940 654370 7030 654610
rect 7270 654370 7360 654610
rect 7600 654370 7690 654610
rect 7930 654390 82750 654610
rect 82990 654390 83080 654630
rect 83320 654390 83410 654630
rect 83650 654390 83770 654630
rect 84010 654390 84100 654630
rect 84340 654390 84460 654630
rect 84700 654390 84790 654630
rect 85030 654390 85310 654630
rect 7930 654370 85310 654390
rect 3000 654300 85310 654370
rect 3000 654280 82750 654300
rect 3000 654040 3070 654280
rect 3310 654040 3400 654280
rect 3640 654040 3730 654280
rect 3970 654040 4060 654280
rect 4300 654040 4390 654280
rect 4630 654040 4720 654280
rect 4960 654040 5050 654280
rect 5290 654040 5380 654280
rect 5620 654040 5710 654280
rect 5950 654040 6040 654280
rect 6280 654040 6370 654280
rect 6610 654040 6700 654280
rect 6940 654040 7030 654280
rect 7270 654040 7360 654280
rect 7600 654040 7690 654280
rect 7930 654060 82750 654280
rect 82990 654060 83080 654300
rect 83320 654060 83410 654300
rect 83650 654060 83770 654300
rect 84010 654060 84100 654300
rect 84340 654060 84460 654300
rect 84700 654060 84790 654300
rect 85030 654060 85310 654300
rect 7930 654040 85310 654060
rect 3000 653950 85310 654040
rect 3000 653710 3070 653950
rect 3310 653710 3400 653950
rect 3640 653710 3730 653950
rect 3970 653710 4060 653950
rect 4300 653710 4390 653950
rect 4630 653710 4720 653950
rect 4960 653710 5050 653950
rect 5290 653710 5380 653950
rect 5620 653710 5710 653950
rect 5950 653710 6040 653950
rect 6280 653710 6370 653950
rect 6610 653710 6700 653950
rect 6940 653710 7030 653950
rect 7270 653710 7360 653950
rect 7600 653710 7690 653950
rect 7930 653940 85310 653950
rect 7930 653710 82750 653940
rect 3000 653700 82750 653710
rect 82990 653700 83080 653940
rect 83320 653700 83410 653940
rect 83650 653700 83770 653940
rect 84010 653700 84100 653940
rect 84340 653700 84460 653940
rect 84700 653700 84790 653940
rect 85030 653700 85310 653940
rect 3000 653620 85310 653700
rect 3000 653380 3070 653620
rect 3310 653380 3400 653620
rect 3640 653380 3730 653620
rect 3970 653380 4060 653620
rect 4300 653380 4390 653620
rect 4630 653380 4720 653620
rect 4960 653380 5050 653620
rect 5290 653380 5380 653620
rect 5620 653380 5710 653620
rect 5950 653380 6040 653620
rect 6280 653380 6370 653620
rect 6610 653380 6700 653620
rect 6940 653380 7030 653620
rect 7270 653380 7360 653620
rect 7600 653380 7690 653620
rect 7930 653610 85310 653620
rect 7930 653380 82750 653610
rect 3000 653370 82750 653380
rect 82990 653370 83080 653610
rect 83320 653370 83410 653610
rect 83650 653370 83770 653610
rect 84010 653370 84100 653610
rect 84340 653370 84460 653610
rect 84700 653370 84790 653610
rect 85030 653370 85310 653610
rect 3000 653290 85310 653370
rect 3000 653050 3070 653290
rect 3310 653050 3400 653290
rect 3640 653050 3730 653290
rect 3970 653050 4060 653290
rect 4300 653050 4390 653290
rect 4630 653050 4720 653290
rect 4960 653050 5050 653290
rect 5290 653050 5380 653290
rect 5620 653050 5710 653290
rect 5950 653050 6040 653290
rect 6280 653050 6370 653290
rect 6610 653050 6700 653290
rect 6940 653050 7030 653290
rect 7270 653050 7360 653290
rect 7600 653050 7690 653290
rect 7930 653250 85310 653290
rect 7930 653050 82750 653250
rect 3000 653010 82750 653050
rect 82990 653010 83080 653250
rect 83320 653010 83410 653250
rect 83650 653010 83770 653250
rect 84010 653010 84100 653250
rect 84340 653010 84460 653250
rect 84700 653010 84790 653250
rect 85030 653010 85310 653250
rect 3000 652960 85310 653010
rect 3000 652720 3070 652960
rect 3310 652720 3400 652960
rect 3640 652720 3730 652960
rect 3970 652720 4060 652960
rect 4300 652720 4390 652960
rect 4630 652720 4720 652960
rect 4960 652720 5050 652960
rect 5290 652720 5380 652960
rect 5620 652720 5710 652960
rect 5950 652720 6040 652960
rect 6280 652720 6370 652960
rect 6610 652720 6700 652960
rect 6940 652720 7030 652960
rect 7270 652720 7360 652960
rect 7600 652720 7690 652960
rect 7930 652920 85310 652960
rect 7930 652720 82750 652920
rect 3000 652680 82750 652720
rect 82990 652680 83080 652920
rect 83320 652680 83410 652920
rect 83650 652680 83770 652920
rect 84010 652680 84100 652920
rect 84340 652680 84460 652920
rect 84700 652680 84790 652920
rect 85030 652680 85310 652920
rect 3000 652630 85310 652680
rect 3000 652390 3070 652630
rect 3310 652390 3400 652630
rect 3640 652390 3730 652630
rect 3970 652390 4060 652630
rect 4300 652390 4390 652630
rect 4630 652390 4720 652630
rect 4960 652390 5050 652630
rect 5290 652390 5380 652630
rect 5620 652390 5710 652630
rect 5950 652390 6040 652630
rect 6280 652390 6370 652630
rect 6610 652390 6700 652630
rect 6940 652390 7030 652630
rect 7270 652390 7360 652630
rect 7600 652390 7690 652630
rect 7930 652590 85310 652630
rect 7930 652390 82750 652590
rect 3000 652350 82750 652390
rect 82990 652350 83080 652590
rect 83320 652350 83410 652590
rect 83650 652350 83770 652590
rect 84010 652350 84100 652590
rect 84340 652350 84460 652590
rect 84700 652350 84790 652590
rect 85030 652350 85310 652590
rect 3000 652312 85310 652350
rect 3000 652300 32350 652312
rect 3000 652060 3070 652300
rect 3310 652060 3400 652300
rect 3640 652060 3730 652300
rect 3970 652060 4060 652300
rect 4300 652060 4390 652300
rect 4630 652060 4720 652300
rect 4960 652060 5050 652300
rect 5290 652060 5380 652300
rect 5620 652060 5710 652300
rect 5950 652060 6040 652300
rect 6280 652060 6370 652300
rect 6610 652060 6700 652300
rect 6940 652060 7030 652300
rect 7270 652060 7360 652300
rect 7600 652060 7690 652300
rect 7930 652060 32350 652300
rect 3000 651970 32350 652060
rect 3000 651730 3070 651970
rect 3310 651730 3400 651970
rect 3640 651730 3730 651970
rect 3970 651730 4060 651970
rect 4300 651730 4390 651970
rect 4630 651730 4720 651970
rect 4960 651730 5050 651970
rect 5290 651730 5380 651970
rect 5620 651730 5710 651970
rect 5950 651730 6040 651970
rect 6280 651730 6370 651970
rect 6610 651730 6700 651970
rect 6940 651730 7030 651970
rect 7270 651730 7360 651970
rect 7600 651730 7690 651970
rect 7930 651730 32350 651970
rect 3000 651640 32350 651730
rect 134191 651640 134761 682296
rect 566720 681240 567290 691785
rect 566270 681239 567290 681240
rect 3000 651400 3070 651640
rect 3310 651400 3400 651640
rect 3640 651400 3730 651640
rect 3970 651400 4060 651640
rect 4300 651400 4390 651640
rect 4630 651400 4720 651640
rect 4960 651400 5050 651640
rect 5290 651400 5380 651640
rect 5620 651400 5710 651640
rect 5950 651400 6040 651640
rect 6280 651400 6370 651640
rect 6610 651400 6700 651640
rect 6940 651400 7030 651640
rect 7270 651400 7360 651640
rect 7600 651400 7690 651640
rect 7930 651400 32350 651640
rect 3000 651310 32350 651400
rect 120014 651320 134761 651640
rect 135741 680670 567290 681239
rect 135741 680669 566840 680670
rect 3000 651070 3070 651310
rect 3310 651070 3400 651310
rect 3640 651070 3730 651310
rect 3970 651070 4060 651310
rect 4300 651070 4390 651310
rect 4630 651070 4720 651310
rect 4960 651070 5050 651310
rect 5290 651070 5380 651310
rect 5620 651070 5710 651310
rect 5950 651070 6040 651310
rect 6280 651070 6370 651310
rect 6610 651070 6700 651310
rect 6940 651070 7030 651310
rect 7270 651070 7360 651310
rect 7600 651070 7690 651310
rect 7930 651070 32350 651310
rect 3000 651000 32350 651070
rect 27350 648719 32350 651000
rect 27350 643722 79310 648719
rect 135741 645780 136311 680669
rect 112144 645210 136311 645780
rect 137524 678966 571785 679536
rect 577305 679516 582870 679536
rect 577305 679446 582320 679516
rect 582390 679446 582410 679516
rect 582480 679446 582500 679516
rect 582570 679446 582590 679516
rect 582660 679446 582680 679516
rect 582750 679446 582770 679516
rect 582840 679446 582870 679516
rect 577305 679426 582870 679446
rect 577305 679356 582320 679426
rect 582390 679356 582410 679426
rect 582480 679356 582500 679426
rect 582570 679356 582590 679426
rect 582660 679356 582680 679426
rect 582750 679356 582770 679426
rect 582840 679356 582870 679426
rect 577305 679336 582870 679356
rect 577305 679266 582320 679336
rect 582390 679266 582410 679336
rect 582480 679266 582500 679336
rect 582570 679266 582590 679336
rect 582660 679266 582680 679336
rect 582750 679266 582770 679336
rect 582840 679266 582870 679336
rect 577305 679246 582870 679266
rect 577305 679176 582320 679246
rect 582390 679176 582410 679246
rect 582480 679176 582500 679246
rect 582570 679176 582590 679246
rect 582660 679176 582680 679246
rect 582750 679176 582770 679246
rect 582840 679176 582870 679246
rect 577305 679156 582870 679176
rect 577305 679086 582320 679156
rect 582390 679086 582410 679156
rect 582480 679086 582500 679156
rect 582570 679086 582590 679156
rect 582660 679086 582680 679156
rect 582750 679086 582770 679156
rect 582840 679086 582870 679156
rect 577305 679066 582870 679086
rect 577305 678996 582320 679066
rect 582390 678996 582410 679066
rect 582480 678996 582500 679066
rect 582570 678996 582590 679066
rect 582660 678996 582680 679066
rect 582750 678996 582770 679066
rect 582840 678996 582870 679066
rect 577305 678966 582870 678996
rect 27350 632894 32350 643722
rect 137524 639921 138094 678966
rect 111924 639351 138094 639921
rect 111924 639350 112363 639351
rect 93369 638170 95369 638207
rect 93369 638100 94280 638170
rect 94350 638100 94380 638170
rect 94450 638100 94480 638170
rect 94550 638100 95369 638170
rect 93369 638080 95369 638100
rect 93369 638010 94280 638080
rect 94350 638010 94380 638080
rect 94450 638010 94480 638080
rect 94550 638010 95369 638080
rect 27350 627894 79310 632894
rect 93369 623548 95369 638010
rect 21946 623528 95369 623548
rect 21946 623458 21966 623528
rect 22036 623458 22056 623528
rect 22126 623458 22146 623528
rect 22216 623458 22236 623528
rect 22306 623458 22326 623528
rect 22396 623458 22416 623528
rect 22486 623458 22506 623528
rect 22576 623458 22596 623528
rect 22666 623458 22686 623528
rect 22756 623458 22776 623528
rect 22846 623458 22866 623528
rect 22936 623458 22956 623528
rect 23026 623458 23046 623528
rect 23116 623458 23136 623528
rect 23206 623458 23226 623528
rect 23296 623458 23316 623528
rect 23386 623458 23406 623528
rect 23476 623458 23496 623528
rect 23566 623458 23586 623528
rect 23656 623458 23676 623528
rect 23746 623458 23766 623528
rect 23836 623458 23856 623528
rect 23926 623458 95369 623528
rect 21946 623438 95369 623458
rect 21946 623368 21966 623438
rect 22036 623368 22056 623438
rect 22126 623368 22146 623438
rect 22216 623368 22236 623438
rect 22306 623368 22326 623438
rect 22396 623368 22416 623438
rect 22486 623368 22506 623438
rect 22576 623368 22596 623438
rect 22666 623368 22686 623438
rect 22756 623368 22776 623438
rect 22846 623368 22866 623438
rect 22936 623368 22956 623438
rect 23026 623368 23046 623438
rect 23116 623368 23136 623438
rect 23206 623368 23226 623438
rect 23296 623368 23316 623438
rect 23386 623368 23406 623438
rect 23476 623368 23496 623438
rect 23566 623368 23586 623438
rect 23656 623368 23676 623438
rect 23746 623368 23766 623438
rect 23836 623368 23856 623438
rect 23926 623368 95369 623438
rect 21946 623348 95369 623368
rect 21946 623278 21966 623348
rect 22036 623278 22056 623348
rect 22126 623278 22146 623348
rect 22216 623278 22236 623348
rect 22306 623278 22326 623348
rect 22396 623278 22416 623348
rect 22486 623278 22506 623348
rect 22576 623278 22596 623348
rect 22666 623278 22686 623348
rect 22756 623278 22776 623348
rect 22846 623278 22866 623348
rect 22936 623278 22956 623348
rect 23026 623278 23046 623348
rect 23116 623278 23136 623348
rect 23206 623278 23226 623348
rect 23296 623278 23316 623348
rect 23386 623278 23406 623348
rect 23476 623278 23496 623348
rect 23566 623278 23586 623348
rect 23656 623278 23676 623348
rect 23746 623278 23766 623348
rect 23836 623278 23856 623348
rect 23926 623278 95369 623348
rect 21946 623258 95369 623278
rect 21946 623188 21966 623258
rect 22036 623188 22056 623258
rect 22126 623188 22146 623258
rect 22216 623188 22236 623258
rect 22306 623188 22326 623258
rect 22396 623188 22416 623258
rect 22486 623188 22506 623258
rect 22576 623188 22596 623258
rect 22666 623188 22686 623258
rect 22756 623188 22776 623258
rect 22846 623188 22866 623258
rect 22936 623188 22956 623258
rect 23026 623188 23046 623258
rect 23116 623188 23136 623258
rect 23206 623188 23226 623258
rect 23296 623188 23316 623258
rect 23386 623188 23406 623258
rect 23476 623188 23496 623258
rect 23566 623188 23586 623258
rect 23656 623188 23676 623258
rect 23746 623188 23766 623258
rect 23836 623188 23856 623258
rect 23926 623188 95369 623258
rect 21946 623168 95369 623188
rect 21946 623098 21966 623168
rect 22036 623098 22056 623168
rect 22126 623098 22146 623168
rect 22216 623098 22236 623168
rect 22306 623098 22326 623168
rect 22396 623098 22416 623168
rect 22486 623098 22506 623168
rect 22576 623098 22596 623168
rect 22666 623098 22686 623168
rect 22756 623098 22776 623168
rect 22846 623098 22866 623168
rect 22936 623098 22956 623168
rect 23026 623098 23046 623168
rect 23116 623098 23136 623168
rect 23206 623098 23226 623168
rect 23296 623098 23316 623168
rect 23386 623098 23406 623168
rect 23476 623098 23496 623168
rect 23566 623098 23586 623168
rect 23656 623098 23676 623168
rect 23746 623098 23766 623168
rect 23836 623098 23856 623168
rect 23926 623098 95369 623168
rect 21946 623078 95369 623098
rect 21946 623008 21966 623078
rect 22036 623008 22056 623078
rect 22126 623008 22146 623078
rect 22216 623008 22236 623078
rect 22306 623008 22326 623078
rect 22396 623008 22416 623078
rect 22486 623008 22506 623078
rect 22576 623008 22596 623078
rect 22666 623008 22686 623078
rect 22756 623008 22776 623078
rect 22846 623008 22866 623078
rect 22936 623008 22956 623078
rect 23026 623008 23046 623078
rect 23116 623008 23136 623078
rect 23206 623008 23226 623078
rect 23296 623008 23316 623078
rect 23386 623008 23406 623078
rect 23476 623008 23496 623078
rect 23566 623008 23586 623078
rect 23656 623008 23676 623078
rect 23746 623008 23766 623078
rect 23836 623008 23856 623078
rect 23926 623008 95369 623078
rect 21946 622988 95369 623008
rect 21946 622918 21966 622988
rect 22036 622918 22056 622988
rect 22126 622918 22146 622988
rect 22216 622918 22236 622988
rect 22306 622918 22326 622988
rect 22396 622918 22416 622988
rect 22486 622918 22506 622988
rect 22576 622918 22596 622988
rect 22666 622918 22686 622988
rect 22756 622918 22776 622988
rect 22846 622918 22866 622988
rect 22936 622918 22956 622988
rect 23026 622918 23046 622988
rect 23116 622918 23136 622988
rect 23206 622918 23226 622988
rect 23296 622918 23316 622988
rect 23386 622918 23406 622988
rect 23476 622918 23496 622988
rect 23566 622918 23586 622988
rect 23656 622918 23676 622988
rect 23746 622918 23766 622988
rect 23836 622918 23856 622988
rect 23926 622918 95369 622988
rect 21946 622898 95369 622918
rect 21946 622828 21966 622898
rect 22036 622828 22056 622898
rect 22126 622828 22146 622898
rect 22216 622828 22236 622898
rect 22306 622828 22326 622898
rect 22396 622828 22416 622898
rect 22486 622828 22506 622898
rect 22576 622828 22596 622898
rect 22666 622828 22686 622898
rect 22756 622828 22776 622898
rect 22846 622828 22866 622898
rect 22936 622828 22956 622898
rect 23026 622828 23046 622898
rect 23116 622828 23136 622898
rect 23206 622828 23226 622898
rect 23296 622828 23316 622898
rect 23386 622828 23406 622898
rect 23476 622828 23496 622898
rect 23566 622828 23586 622898
rect 23656 622828 23676 622898
rect 23746 622828 23766 622898
rect 23836 622828 23856 622898
rect 23926 622828 95369 622898
rect 21946 622808 95369 622828
rect 21946 622738 21966 622808
rect 22036 622738 22056 622808
rect 22126 622738 22146 622808
rect 22216 622738 22236 622808
rect 22306 622738 22326 622808
rect 22396 622738 22416 622808
rect 22486 622738 22506 622808
rect 22576 622738 22596 622808
rect 22666 622738 22686 622808
rect 22756 622738 22776 622808
rect 22846 622738 22866 622808
rect 22936 622738 22956 622808
rect 23026 622738 23046 622808
rect 23116 622738 23136 622808
rect 23206 622738 23226 622808
rect 23296 622738 23316 622808
rect 23386 622738 23406 622808
rect 23476 622738 23496 622808
rect 23566 622738 23586 622808
rect 23656 622738 23676 622808
rect 23746 622738 23766 622808
rect 23836 622738 23856 622808
rect 23926 622738 95369 622808
rect 21946 622718 95369 622738
rect 21946 622648 21966 622718
rect 22036 622648 22056 622718
rect 22126 622648 22146 622718
rect 22216 622648 22236 622718
rect 22306 622648 22326 622718
rect 22396 622648 22416 622718
rect 22486 622648 22506 622718
rect 22576 622648 22596 622718
rect 22666 622648 22686 622718
rect 22756 622648 22776 622718
rect 22846 622648 22866 622718
rect 22936 622648 22956 622718
rect 23026 622648 23046 622718
rect 23116 622648 23136 622718
rect 23206 622648 23226 622718
rect 23296 622648 23316 622718
rect 23386 622648 23406 622718
rect 23476 622648 23496 622718
rect 23566 622648 23586 622718
rect 23656 622648 23676 622718
rect 23746 622648 23766 622718
rect 23836 622648 23856 622718
rect 23926 622648 95369 622718
rect 21946 622628 95369 622648
rect 21946 622558 21966 622628
rect 22036 622558 22056 622628
rect 22126 622558 22146 622628
rect 22216 622558 22236 622628
rect 22306 622558 22326 622628
rect 22396 622558 22416 622628
rect 22486 622558 22506 622628
rect 22576 622558 22596 622628
rect 22666 622558 22686 622628
rect 22756 622558 22776 622628
rect 22846 622558 22866 622628
rect 22936 622558 22956 622628
rect 23026 622558 23046 622628
rect 23116 622558 23136 622628
rect 23206 622558 23226 622628
rect 23296 622558 23316 622628
rect 23386 622558 23406 622628
rect 23476 622558 23496 622628
rect 23566 622558 23586 622628
rect 23656 622558 23676 622628
rect 23746 622558 23766 622628
rect 23836 622558 23856 622628
rect 23926 622558 95369 622628
rect 21946 622538 95369 622558
rect 21946 622468 21966 622538
rect 22036 622468 22056 622538
rect 22126 622468 22146 622538
rect 22216 622468 22236 622538
rect 22306 622468 22326 622538
rect 22396 622468 22416 622538
rect 22486 622468 22506 622538
rect 22576 622468 22596 622538
rect 22666 622468 22686 622538
rect 22756 622468 22776 622538
rect 22846 622468 22866 622538
rect 22936 622468 22956 622538
rect 23026 622468 23046 622538
rect 23116 622468 23136 622538
rect 23206 622468 23226 622538
rect 23296 622468 23316 622538
rect 23386 622468 23406 622538
rect 23476 622468 23496 622538
rect 23566 622468 23586 622538
rect 23656 622468 23676 622538
rect 23746 622468 23766 622538
rect 23836 622468 23856 622538
rect 23926 622468 95369 622538
rect 21946 622448 95369 622468
rect 21946 622378 21966 622448
rect 22036 622378 22056 622448
rect 22126 622378 22146 622448
rect 22216 622378 22236 622448
rect 22306 622378 22326 622448
rect 22396 622378 22416 622448
rect 22486 622378 22506 622448
rect 22576 622378 22596 622448
rect 22666 622378 22686 622448
rect 22756 622378 22776 622448
rect 22846 622378 22866 622448
rect 22936 622378 22956 622448
rect 23026 622378 23046 622448
rect 23116 622378 23136 622448
rect 23206 622378 23226 622448
rect 23296 622378 23316 622448
rect 23386 622378 23406 622448
rect 23476 622378 23496 622448
rect 23566 622378 23586 622448
rect 23656 622378 23676 622448
rect 23746 622378 23766 622448
rect 23836 622378 23856 622448
rect 23926 622378 95369 622448
rect 21946 622358 95369 622378
rect 21946 622288 21966 622358
rect 22036 622288 22056 622358
rect 22126 622288 22146 622358
rect 22216 622288 22236 622358
rect 22306 622288 22326 622358
rect 22396 622288 22416 622358
rect 22486 622288 22506 622358
rect 22576 622288 22596 622358
rect 22666 622288 22686 622358
rect 22756 622288 22776 622358
rect 22846 622288 22866 622358
rect 22936 622288 22956 622358
rect 23026 622288 23046 622358
rect 23116 622288 23136 622358
rect 23206 622288 23226 622358
rect 23296 622288 23316 622358
rect 23386 622288 23406 622358
rect 23476 622288 23496 622358
rect 23566 622288 23586 622358
rect 23656 622288 23676 622358
rect 23746 622288 23766 622358
rect 23836 622288 23856 622358
rect 23926 622288 95369 622358
rect 21946 622268 95369 622288
rect 21946 622198 21966 622268
rect 22036 622198 22056 622268
rect 22126 622198 22146 622268
rect 22216 622198 22236 622268
rect 22306 622198 22326 622268
rect 22396 622198 22416 622268
rect 22486 622198 22506 622268
rect 22576 622198 22596 622268
rect 22666 622198 22686 622268
rect 22756 622198 22776 622268
rect 22846 622198 22866 622268
rect 22936 622198 22956 622268
rect 23026 622198 23046 622268
rect 23116 622198 23136 622268
rect 23206 622198 23226 622268
rect 23296 622198 23316 622268
rect 23386 622198 23406 622268
rect 23476 622198 23496 622268
rect 23566 622198 23586 622268
rect 23656 622198 23676 622268
rect 23746 622198 23766 622268
rect 23836 622198 23856 622268
rect 23926 622198 95369 622268
rect 21946 622178 95369 622198
rect 21946 622108 21966 622178
rect 22036 622108 22056 622178
rect 22126 622108 22146 622178
rect 22216 622108 22236 622178
rect 22306 622108 22326 622178
rect 22396 622108 22416 622178
rect 22486 622108 22506 622178
rect 22576 622108 22596 622178
rect 22666 622108 22686 622178
rect 22756 622108 22776 622178
rect 22846 622108 22866 622178
rect 22936 622108 22956 622178
rect 23026 622108 23046 622178
rect 23116 622108 23136 622178
rect 23206 622108 23226 622178
rect 23296 622108 23316 622178
rect 23386 622108 23406 622178
rect 23476 622108 23496 622178
rect 23566 622108 23586 622178
rect 23656 622108 23676 622178
rect 23746 622108 23766 622178
rect 23836 622108 23856 622178
rect 23926 622108 95369 622178
rect 21946 622088 95369 622108
rect 21946 622018 21966 622088
rect 22036 622018 22056 622088
rect 22126 622018 22146 622088
rect 22216 622018 22236 622088
rect 22306 622018 22326 622088
rect 22396 622018 22416 622088
rect 22486 622018 22506 622088
rect 22576 622018 22596 622088
rect 22666 622018 22686 622088
rect 22756 622018 22776 622088
rect 22846 622018 22866 622088
rect 22936 622018 22956 622088
rect 23026 622018 23046 622088
rect 23116 622018 23136 622088
rect 23206 622018 23226 622088
rect 23296 622018 23316 622088
rect 23386 622018 23406 622088
rect 23476 622018 23496 622088
rect 23566 622018 23586 622088
rect 23656 622018 23676 622088
rect 23746 622018 23766 622088
rect 23836 622018 23856 622088
rect 23926 622018 95369 622088
rect 21946 621998 95369 622018
rect 21946 621928 21966 621998
rect 22036 621928 22056 621998
rect 22126 621928 22146 621998
rect 22216 621928 22236 621998
rect 22306 621928 22326 621998
rect 22396 621928 22416 621998
rect 22486 621928 22506 621998
rect 22576 621928 22596 621998
rect 22666 621928 22686 621998
rect 22756 621928 22776 621998
rect 22846 621928 22866 621998
rect 22936 621928 22956 621998
rect 23026 621928 23046 621998
rect 23116 621928 23136 621998
rect 23206 621928 23226 621998
rect 23296 621928 23316 621998
rect 23386 621928 23406 621998
rect 23476 621928 23496 621998
rect 23566 621928 23586 621998
rect 23656 621928 23676 621998
rect 23746 621928 23766 621998
rect 23836 621928 23856 621998
rect 23926 621928 95369 621998
rect 21946 621908 95369 621928
rect 21946 621838 21966 621908
rect 22036 621838 22056 621908
rect 22126 621838 22146 621908
rect 22216 621838 22236 621908
rect 22306 621838 22326 621908
rect 22396 621838 22416 621908
rect 22486 621838 22506 621908
rect 22576 621838 22596 621908
rect 22666 621838 22686 621908
rect 22756 621838 22776 621908
rect 22846 621838 22866 621908
rect 22936 621838 22956 621908
rect 23026 621838 23046 621908
rect 23116 621838 23136 621908
rect 23206 621838 23226 621908
rect 23296 621838 23316 621908
rect 23386 621838 23406 621908
rect 23476 621838 23496 621908
rect 23566 621838 23586 621908
rect 23656 621838 23676 621908
rect 23746 621838 23766 621908
rect 23836 621838 23856 621908
rect 23926 621838 95369 621908
rect 21946 621818 95369 621838
rect 21946 621748 21966 621818
rect 22036 621748 22056 621818
rect 22126 621748 22146 621818
rect 22216 621748 22236 621818
rect 22306 621748 22326 621818
rect 22396 621748 22416 621818
rect 22486 621748 22506 621818
rect 22576 621748 22596 621818
rect 22666 621748 22686 621818
rect 22756 621748 22776 621818
rect 22846 621748 22866 621818
rect 22936 621748 22956 621818
rect 23026 621748 23046 621818
rect 23116 621748 23136 621818
rect 23206 621748 23226 621818
rect 23296 621748 23316 621818
rect 23386 621748 23406 621818
rect 23476 621748 23496 621818
rect 23566 621748 23586 621818
rect 23656 621748 23676 621818
rect 23746 621748 23766 621818
rect 23836 621748 23856 621818
rect 23926 621748 95369 621818
rect 21946 621728 95369 621748
rect 21946 621658 21966 621728
rect 22036 621658 22056 621728
rect 22126 621658 22146 621728
rect 22216 621658 22236 621728
rect 22306 621658 22326 621728
rect 22396 621658 22416 621728
rect 22486 621658 22506 621728
rect 22576 621658 22596 621728
rect 22666 621658 22686 621728
rect 22756 621658 22776 621728
rect 22846 621658 22866 621728
rect 22936 621658 22956 621728
rect 23026 621658 23046 621728
rect 23116 621658 23136 621728
rect 23206 621658 23226 621728
rect 23296 621658 23316 621728
rect 23386 621658 23406 621728
rect 23476 621658 23496 621728
rect 23566 621658 23586 621728
rect 23656 621658 23676 621728
rect 23746 621658 23766 621728
rect 23836 621658 23856 621728
rect 23926 621658 95369 621728
rect 21946 621638 95369 621658
rect 21946 621568 21966 621638
rect 22036 621568 22056 621638
rect 22126 621568 22146 621638
rect 22216 621568 22236 621638
rect 22306 621568 22326 621638
rect 22396 621568 22416 621638
rect 22486 621568 22506 621638
rect 22576 621568 22596 621638
rect 22666 621568 22686 621638
rect 22756 621568 22776 621638
rect 22846 621568 22866 621638
rect 22936 621568 22956 621638
rect 23026 621568 23046 621638
rect 23116 621568 23136 621638
rect 23206 621568 23226 621638
rect 23296 621568 23316 621638
rect 23386 621568 23406 621638
rect 23476 621568 23496 621638
rect 23566 621568 23586 621638
rect 23656 621568 23676 621638
rect 23746 621568 23766 621638
rect 23836 621568 23856 621638
rect 23926 621568 95369 621638
rect 21946 621548 95369 621568
rect 97956 638170 99956 638193
rect 97956 638100 98838 638170
rect 98908 638100 98938 638170
rect 99008 638100 99038 638170
rect 99108 638100 99956 638170
rect 97956 638080 99956 638100
rect 97956 638010 98838 638080
rect 98908 638010 98938 638080
rect 99008 638010 99038 638080
rect 99108 638010 99956 638080
rect 97956 619440 99956 638010
rect 17650 619420 99956 619440
rect 17650 619350 17670 619420
rect 17740 619350 17760 619420
rect 17830 619350 17850 619420
rect 17920 619350 17940 619420
rect 18010 619350 18030 619420
rect 18100 619350 18120 619420
rect 18190 619350 18210 619420
rect 18280 619350 18300 619420
rect 18370 619350 18390 619420
rect 18460 619350 18480 619420
rect 18550 619350 18570 619420
rect 18640 619350 18660 619420
rect 18730 619350 18750 619420
rect 18820 619350 18840 619420
rect 18910 619350 18930 619420
rect 19000 619350 19020 619420
rect 19090 619350 19110 619420
rect 19180 619350 19200 619420
rect 19270 619350 19290 619420
rect 19360 619350 19380 619420
rect 19450 619350 19470 619420
rect 19540 619350 19560 619420
rect 19630 619350 99956 619420
rect 17650 619330 99956 619350
rect 17650 619260 17670 619330
rect 17740 619260 17760 619330
rect 17830 619260 17850 619330
rect 17920 619260 17940 619330
rect 18010 619260 18030 619330
rect 18100 619260 18120 619330
rect 18190 619260 18210 619330
rect 18280 619260 18300 619330
rect 18370 619260 18390 619330
rect 18460 619260 18480 619330
rect 18550 619260 18570 619330
rect 18640 619260 18660 619330
rect 18730 619260 18750 619330
rect 18820 619260 18840 619330
rect 18910 619260 18930 619330
rect 19000 619260 19020 619330
rect 19090 619260 19110 619330
rect 19180 619260 19200 619330
rect 19270 619260 19290 619330
rect 19360 619260 19380 619330
rect 19450 619260 19470 619330
rect 19540 619260 19560 619330
rect 19630 619260 99956 619330
rect 17650 619240 99956 619260
rect 17650 619170 17670 619240
rect 17740 619170 17760 619240
rect 17830 619170 17850 619240
rect 17920 619170 17940 619240
rect 18010 619170 18030 619240
rect 18100 619170 18120 619240
rect 18190 619170 18210 619240
rect 18280 619170 18300 619240
rect 18370 619170 18390 619240
rect 18460 619170 18480 619240
rect 18550 619170 18570 619240
rect 18640 619170 18660 619240
rect 18730 619170 18750 619240
rect 18820 619170 18840 619240
rect 18910 619170 18930 619240
rect 19000 619170 19020 619240
rect 19090 619170 19110 619240
rect 19180 619170 19200 619240
rect 19270 619170 19290 619240
rect 19360 619170 19380 619240
rect 19450 619170 19470 619240
rect 19540 619170 19560 619240
rect 19630 619170 99956 619240
rect 17650 619150 99956 619170
rect 17650 619080 17670 619150
rect 17740 619080 17760 619150
rect 17830 619080 17850 619150
rect 17920 619080 17940 619150
rect 18010 619080 18030 619150
rect 18100 619080 18120 619150
rect 18190 619080 18210 619150
rect 18280 619080 18300 619150
rect 18370 619080 18390 619150
rect 18460 619080 18480 619150
rect 18550 619080 18570 619150
rect 18640 619080 18660 619150
rect 18730 619080 18750 619150
rect 18820 619080 18840 619150
rect 18910 619080 18930 619150
rect 19000 619080 19020 619150
rect 19090 619080 19110 619150
rect 19180 619080 19200 619150
rect 19270 619080 19290 619150
rect 19360 619080 19380 619150
rect 19450 619080 19470 619150
rect 19540 619080 19560 619150
rect 19630 619080 99956 619150
rect 17650 619060 99956 619080
rect 17650 618990 17670 619060
rect 17740 618990 17760 619060
rect 17830 618990 17850 619060
rect 17920 618990 17940 619060
rect 18010 618990 18030 619060
rect 18100 618990 18120 619060
rect 18190 618990 18210 619060
rect 18280 618990 18300 619060
rect 18370 618990 18390 619060
rect 18460 618990 18480 619060
rect 18550 618990 18570 619060
rect 18640 618990 18660 619060
rect 18730 618990 18750 619060
rect 18820 618990 18840 619060
rect 18910 618990 18930 619060
rect 19000 618990 19020 619060
rect 19090 618990 19110 619060
rect 19180 618990 19200 619060
rect 19270 618990 19290 619060
rect 19360 618990 19380 619060
rect 19450 618990 19470 619060
rect 19540 618990 19560 619060
rect 19630 618990 99956 619060
rect 17650 618970 99956 618990
rect 17650 618900 17670 618970
rect 17740 618900 17760 618970
rect 17830 618900 17850 618970
rect 17920 618900 17940 618970
rect 18010 618900 18030 618970
rect 18100 618900 18120 618970
rect 18190 618900 18210 618970
rect 18280 618900 18300 618970
rect 18370 618900 18390 618970
rect 18460 618900 18480 618970
rect 18550 618900 18570 618970
rect 18640 618900 18660 618970
rect 18730 618900 18750 618970
rect 18820 618900 18840 618970
rect 18910 618900 18930 618970
rect 19000 618900 19020 618970
rect 19090 618900 19110 618970
rect 19180 618900 19200 618970
rect 19270 618900 19290 618970
rect 19360 618900 19380 618970
rect 19450 618900 19470 618970
rect 19540 618900 19560 618970
rect 19630 618900 99956 618970
rect 17650 618880 99956 618900
rect 17650 618810 17670 618880
rect 17740 618810 17760 618880
rect 17830 618810 17850 618880
rect 17920 618810 17940 618880
rect 18010 618810 18030 618880
rect 18100 618810 18120 618880
rect 18190 618810 18210 618880
rect 18280 618810 18300 618880
rect 18370 618810 18390 618880
rect 18460 618810 18480 618880
rect 18550 618810 18570 618880
rect 18640 618810 18660 618880
rect 18730 618810 18750 618880
rect 18820 618810 18840 618880
rect 18910 618810 18930 618880
rect 19000 618810 19020 618880
rect 19090 618810 19110 618880
rect 19180 618810 19200 618880
rect 19270 618810 19290 618880
rect 19360 618810 19380 618880
rect 19450 618810 19470 618880
rect 19540 618810 19560 618880
rect 19630 618810 99956 618880
rect 17650 618790 99956 618810
rect 17650 618720 17670 618790
rect 17740 618720 17760 618790
rect 17830 618720 17850 618790
rect 17920 618720 17940 618790
rect 18010 618720 18030 618790
rect 18100 618720 18120 618790
rect 18190 618720 18210 618790
rect 18280 618720 18300 618790
rect 18370 618720 18390 618790
rect 18460 618720 18480 618790
rect 18550 618720 18570 618790
rect 18640 618720 18660 618790
rect 18730 618720 18750 618790
rect 18820 618720 18840 618790
rect 18910 618720 18930 618790
rect 19000 618720 19020 618790
rect 19090 618720 19110 618790
rect 19180 618720 19200 618790
rect 19270 618720 19290 618790
rect 19360 618720 19380 618790
rect 19450 618720 19470 618790
rect 19540 618720 19560 618790
rect 19630 618720 99956 618790
rect 17650 618700 99956 618720
rect 17650 618630 17670 618700
rect 17740 618630 17760 618700
rect 17830 618630 17850 618700
rect 17920 618630 17940 618700
rect 18010 618630 18030 618700
rect 18100 618630 18120 618700
rect 18190 618630 18210 618700
rect 18280 618630 18300 618700
rect 18370 618630 18390 618700
rect 18460 618630 18480 618700
rect 18550 618630 18570 618700
rect 18640 618630 18660 618700
rect 18730 618630 18750 618700
rect 18820 618630 18840 618700
rect 18910 618630 18930 618700
rect 19000 618630 19020 618700
rect 19090 618630 19110 618700
rect 19180 618630 19200 618700
rect 19270 618630 19290 618700
rect 19360 618630 19380 618700
rect 19450 618630 19470 618700
rect 19540 618630 19560 618700
rect 19630 618630 99956 618700
rect 17650 618610 99956 618630
rect 17650 618540 17670 618610
rect 17740 618540 17760 618610
rect 17830 618540 17850 618610
rect 17920 618540 17940 618610
rect 18010 618540 18030 618610
rect 18100 618540 18120 618610
rect 18190 618540 18210 618610
rect 18280 618540 18300 618610
rect 18370 618540 18390 618610
rect 18460 618540 18480 618610
rect 18550 618540 18570 618610
rect 18640 618540 18660 618610
rect 18730 618540 18750 618610
rect 18820 618540 18840 618610
rect 18910 618540 18930 618610
rect 19000 618540 19020 618610
rect 19090 618540 19110 618610
rect 19180 618540 19200 618610
rect 19270 618540 19290 618610
rect 19360 618540 19380 618610
rect 19450 618540 19470 618610
rect 19540 618540 19560 618610
rect 19630 618540 99956 618610
rect 17650 618520 99956 618540
rect 17650 618450 17670 618520
rect 17740 618450 17760 618520
rect 17830 618450 17850 618520
rect 17920 618450 17940 618520
rect 18010 618450 18030 618520
rect 18100 618450 18120 618520
rect 18190 618450 18210 618520
rect 18280 618450 18300 618520
rect 18370 618450 18390 618520
rect 18460 618450 18480 618520
rect 18550 618450 18570 618520
rect 18640 618450 18660 618520
rect 18730 618450 18750 618520
rect 18820 618450 18840 618520
rect 18910 618450 18930 618520
rect 19000 618450 19020 618520
rect 19090 618450 19110 618520
rect 19180 618450 19200 618520
rect 19270 618450 19290 618520
rect 19360 618450 19380 618520
rect 19450 618450 19470 618520
rect 19540 618450 19560 618520
rect 19630 618450 99956 618520
rect 17650 618430 99956 618450
rect 17650 618360 17670 618430
rect 17740 618360 17760 618430
rect 17830 618360 17850 618430
rect 17920 618360 17940 618430
rect 18010 618360 18030 618430
rect 18100 618360 18120 618430
rect 18190 618360 18210 618430
rect 18280 618360 18300 618430
rect 18370 618360 18390 618430
rect 18460 618360 18480 618430
rect 18550 618360 18570 618430
rect 18640 618360 18660 618430
rect 18730 618360 18750 618430
rect 18820 618360 18840 618430
rect 18910 618360 18930 618430
rect 19000 618360 19020 618430
rect 19090 618360 19110 618430
rect 19180 618360 19200 618430
rect 19270 618360 19290 618430
rect 19360 618360 19380 618430
rect 19450 618360 19470 618430
rect 19540 618360 19560 618430
rect 19630 618360 99956 618430
rect 17650 618340 99956 618360
rect 17650 618270 17670 618340
rect 17740 618270 17760 618340
rect 17830 618270 17850 618340
rect 17920 618270 17940 618340
rect 18010 618270 18030 618340
rect 18100 618270 18120 618340
rect 18190 618270 18210 618340
rect 18280 618270 18300 618340
rect 18370 618270 18390 618340
rect 18460 618270 18480 618340
rect 18550 618270 18570 618340
rect 18640 618270 18660 618340
rect 18730 618270 18750 618340
rect 18820 618270 18840 618340
rect 18910 618270 18930 618340
rect 19000 618270 19020 618340
rect 19090 618270 19110 618340
rect 19180 618270 19200 618340
rect 19270 618270 19290 618340
rect 19360 618270 19380 618340
rect 19450 618270 19470 618340
rect 19540 618270 19560 618340
rect 19630 618270 99956 618340
rect 17650 618250 99956 618270
rect 17650 618180 17670 618250
rect 17740 618180 17760 618250
rect 17830 618180 17850 618250
rect 17920 618180 17940 618250
rect 18010 618180 18030 618250
rect 18100 618180 18120 618250
rect 18190 618180 18210 618250
rect 18280 618180 18300 618250
rect 18370 618180 18390 618250
rect 18460 618180 18480 618250
rect 18550 618180 18570 618250
rect 18640 618180 18660 618250
rect 18730 618180 18750 618250
rect 18820 618180 18840 618250
rect 18910 618180 18930 618250
rect 19000 618180 19020 618250
rect 19090 618180 19110 618250
rect 19180 618180 19200 618250
rect 19270 618180 19290 618250
rect 19360 618180 19380 618250
rect 19450 618180 19470 618250
rect 19540 618180 19560 618250
rect 19630 618180 99956 618250
rect 17650 618160 99956 618180
rect 17650 618090 17670 618160
rect 17740 618090 17760 618160
rect 17830 618090 17850 618160
rect 17920 618090 17940 618160
rect 18010 618090 18030 618160
rect 18100 618090 18120 618160
rect 18190 618090 18210 618160
rect 18280 618090 18300 618160
rect 18370 618090 18390 618160
rect 18460 618090 18480 618160
rect 18550 618090 18570 618160
rect 18640 618090 18660 618160
rect 18730 618090 18750 618160
rect 18820 618090 18840 618160
rect 18910 618090 18930 618160
rect 19000 618090 19020 618160
rect 19090 618090 19110 618160
rect 19180 618090 19200 618160
rect 19270 618090 19290 618160
rect 19360 618090 19380 618160
rect 19450 618090 19470 618160
rect 19540 618090 19560 618160
rect 19630 618090 99956 618160
rect 17650 618070 99956 618090
rect 17650 618000 17670 618070
rect 17740 618000 17760 618070
rect 17830 618000 17850 618070
rect 17920 618000 17940 618070
rect 18010 618000 18030 618070
rect 18100 618000 18120 618070
rect 18190 618000 18210 618070
rect 18280 618000 18300 618070
rect 18370 618000 18390 618070
rect 18460 618000 18480 618070
rect 18550 618000 18570 618070
rect 18640 618000 18660 618070
rect 18730 618000 18750 618070
rect 18820 618000 18840 618070
rect 18910 618000 18930 618070
rect 19000 618000 19020 618070
rect 19090 618000 19110 618070
rect 19180 618000 19200 618070
rect 19270 618000 19290 618070
rect 19360 618000 19380 618070
rect 19450 618000 19470 618070
rect 19540 618000 19560 618070
rect 19630 618000 99956 618070
rect 17650 617980 99956 618000
rect 17650 617910 17670 617980
rect 17740 617910 17760 617980
rect 17830 617910 17850 617980
rect 17920 617910 17940 617980
rect 18010 617910 18030 617980
rect 18100 617910 18120 617980
rect 18190 617910 18210 617980
rect 18280 617910 18300 617980
rect 18370 617910 18390 617980
rect 18460 617910 18480 617980
rect 18550 617910 18570 617980
rect 18640 617910 18660 617980
rect 18730 617910 18750 617980
rect 18820 617910 18840 617980
rect 18910 617910 18930 617980
rect 19000 617910 19020 617980
rect 19090 617910 19110 617980
rect 19180 617910 19200 617980
rect 19270 617910 19290 617980
rect 19360 617910 19380 617980
rect 19450 617910 19470 617980
rect 19540 617910 19560 617980
rect 19630 617910 99956 617980
rect 17650 617890 99956 617910
rect 17650 617820 17670 617890
rect 17740 617820 17760 617890
rect 17830 617820 17850 617890
rect 17920 617820 17940 617890
rect 18010 617820 18030 617890
rect 18100 617820 18120 617890
rect 18190 617820 18210 617890
rect 18280 617820 18300 617890
rect 18370 617820 18390 617890
rect 18460 617820 18480 617890
rect 18550 617820 18570 617890
rect 18640 617820 18660 617890
rect 18730 617820 18750 617890
rect 18820 617820 18840 617890
rect 18910 617820 18930 617890
rect 19000 617820 19020 617890
rect 19090 617820 19110 617890
rect 19180 617820 19200 617890
rect 19270 617820 19290 617890
rect 19360 617820 19380 617890
rect 19450 617820 19470 617890
rect 19540 617820 19560 617890
rect 19630 617820 99956 617890
rect 17650 617800 99956 617820
rect 17650 617730 17670 617800
rect 17740 617730 17760 617800
rect 17830 617730 17850 617800
rect 17920 617730 17940 617800
rect 18010 617730 18030 617800
rect 18100 617730 18120 617800
rect 18190 617730 18210 617800
rect 18280 617730 18300 617800
rect 18370 617730 18390 617800
rect 18460 617730 18480 617800
rect 18550 617730 18570 617800
rect 18640 617730 18660 617800
rect 18730 617730 18750 617800
rect 18820 617730 18840 617800
rect 18910 617730 18930 617800
rect 19000 617730 19020 617800
rect 19090 617730 19110 617800
rect 19180 617730 19200 617800
rect 19270 617730 19290 617800
rect 19360 617730 19380 617800
rect 19450 617730 19470 617800
rect 19540 617730 19560 617800
rect 19630 617730 99956 617800
rect 17650 617710 99956 617730
rect 17650 617640 17670 617710
rect 17740 617640 17760 617710
rect 17830 617640 17850 617710
rect 17920 617640 17940 617710
rect 18010 617640 18030 617710
rect 18100 617640 18120 617710
rect 18190 617640 18210 617710
rect 18280 617640 18300 617710
rect 18370 617640 18390 617710
rect 18460 617640 18480 617710
rect 18550 617640 18570 617710
rect 18640 617640 18660 617710
rect 18730 617640 18750 617710
rect 18820 617640 18840 617710
rect 18910 617640 18930 617710
rect 19000 617640 19020 617710
rect 19090 617640 19110 617710
rect 19180 617640 19200 617710
rect 19270 617640 19290 617710
rect 19360 617640 19380 617710
rect 19450 617640 19470 617710
rect 19540 617640 19560 617710
rect 19630 617640 99956 617710
rect 17650 617620 99956 617640
rect 17650 617550 17670 617620
rect 17740 617550 17760 617620
rect 17830 617550 17850 617620
rect 17920 617550 17940 617620
rect 18010 617550 18030 617620
rect 18100 617550 18120 617620
rect 18190 617550 18210 617620
rect 18280 617550 18300 617620
rect 18370 617550 18390 617620
rect 18460 617550 18480 617620
rect 18550 617550 18570 617620
rect 18640 617550 18660 617620
rect 18730 617550 18750 617620
rect 18820 617550 18840 617620
rect 18910 617550 18930 617620
rect 19000 617550 19020 617620
rect 19090 617550 19110 617620
rect 19180 617550 19200 617620
rect 19270 617550 19290 617620
rect 19360 617550 19380 617620
rect 19450 617550 19470 617620
rect 19540 617550 19560 617620
rect 19630 617550 99956 617620
rect 17650 617530 99956 617550
rect 17650 617460 17670 617530
rect 17740 617460 17760 617530
rect 17830 617460 17850 617530
rect 17920 617460 17940 617530
rect 18010 617460 18030 617530
rect 18100 617460 18120 617530
rect 18190 617460 18210 617530
rect 18280 617460 18300 617530
rect 18370 617460 18390 617530
rect 18460 617460 18480 617530
rect 18550 617460 18570 617530
rect 18640 617460 18660 617530
rect 18730 617460 18750 617530
rect 18820 617460 18840 617530
rect 18910 617460 18930 617530
rect 19000 617460 19020 617530
rect 19090 617460 19110 617530
rect 19180 617460 19200 617530
rect 19270 617460 19290 617530
rect 19360 617460 19380 617530
rect 19450 617460 19470 617530
rect 19540 617460 19560 617530
rect 19630 617460 99956 617530
rect 17650 617440 99956 617460
<< via4 >>
rect 170964 692690 171204 692930
rect 171294 692690 171534 692930
rect 171624 692690 171864 692930
rect 171954 692690 172194 692930
rect 172284 692690 172524 692930
rect 172614 692690 172854 692930
rect 170964 692360 171204 692600
rect 171294 692360 171534 692600
rect 171624 692360 171864 692600
rect 171954 692360 172194 692600
rect 172284 692360 172524 692600
rect 172614 692360 172854 692600
rect 170964 692030 171204 692270
rect 171294 692030 171534 692270
rect 171624 692030 171864 692270
rect 171954 692030 172194 692270
rect 172284 692030 172524 692270
rect 172614 692030 172854 692270
rect 170964 691700 171204 691940
rect 171294 691700 171534 691940
rect 171624 691700 171864 691940
rect 171954 691700 172194 691940
rect 172284 691700 172524 691940
rect 172614 691700 172854 691940
rect 170964 691370 171204 691610
rect 171294 691370 171534 691610
rect 171624 691370 171864 691610
rect 171954 691370 172194 691610
rect 172284 691370 172524 691610
rect 172614 691370 172854 691610
rect 170964 691040 171204 691280
rect 171294 691040 171534 691280
rect 171624 691040 171864 691280
rect 171954 691040 172194 691280
rect 172284 691040 172524 691280
rect 172614 691040 172854 691280
rect 170964 690710 171204 690950
rect 171294 690710 171534 690950
rect 171624 690710 171864 690950
rect 171954 690710 172194 690950
rect 172284 690710 172524 690950
rect 172614 690710 172854 690950
rect 170964 690380 171204 690620
rect 171294 690380 171534 690620
rect 171624 690380 171864 690620
rect 171954 690380 172194 690620
rect 172284 690380 172524 690620
rect 172614 690380 172854 690620
rect 170964 690050 171204 690290
rect 171294 690050 171534 690290
rect 171624 690050 171864 690290
rect 171954 690050 172194 690290
rect 172284 690050 172524 690290
rect 172614 690050 172854 690290
rect 170964 689720 171204 689960
rect 171294 689720 171534 689960
rect 171624 689720 171864 689960
rect 171954 689720 172194 689960
rect 172284 689720 172524 689960
rect 172614 689720 172854 689960
rect 170964 689390 171204 689630
rect 171294 689390 171534 689630
rect 171624 689390 171864 689630
rect 171954 689390 172194 689630
rect 172284 689390 172524 689630
rect 172614 689390 172854 689630
rect 170964 689060 171204 689300
rect 171294 689060 171534 689300
rect 171624 689060 171864 689300
rect 171954 689060 172194 689300
rect 172284 689060 172524 689300
rect 172614 689060 172854 689300
rect 170964 688730 171204 688970
rect 171294 688730 171534 688970
rect 171624 688730 171864 688970
rect 171954 688730 172194 688970
rect 172284 688730 172524 688970
rect 172614 688730 172854 688970
rect 170964 688400 171204 688640
rect 171294 688400 171534 688640
rect 171624 688400 171864 688640
rect 171954 688400 172194 688640
rect 172284 688400 172524 688640
rect 172614 688400 172854 688640
rect 170964 688070 171204 688310
rect 171294 688070 171534 688310
rect 171624 688070 171864 688310
rect 171954 688070 172194 688310
rect 172284 688070 172524 688310
rect 172614 688070 172854 688310
rect 225164 700690 225404 700930
rect 225494 700690 225734 700930
rect 225824 700690 226064 700930
rect 226154 700690 226394 700930
rect 226484 700690 226724 700930
rect 226814 700690 227054 700930
rect 225164 700360 225404 700600
rect 225494 700360 225734 700600
rect 225824 700360 226064 700600
rect 226154 700360 226394 700600
rect 226484 700360 226724 700600
rect 226814 700360 227054 700600
rect 225164 700030 225404 700270
rect 225494 700030 225734 700270
rect 225824 700030 226064 700270
rect 226154 700030 226394 700270
rect 226484 700030 226724 700270
rect 226814 700030 227054 700270
rect 225164 699700 225404 699940
rect 225494 699700 225734 699940
rect 225824 699700 226064 699940
rect 226154 699700 226394 699940
rect 226484 699700 226724 699940
rect 226814 699700 227054 699940
rect 225164 699370 225404 699610
rect 225494 699370 225734 699610
rect 225824 699370 226064 699610
rect 226154 699370 226394 699610
rect 226484 699370 226724 699610
rect 226814 699370 227054 699610
rect 225164 699040 225404 699280
rect 225494 699040 225734 699280
rect 225824 699040 226064 699280
rect 226154 699040 226394 699280
rect 226484 699040 226724 699280
rect 226814 699040 227054 699280
rect 225164 698710 225404 698950
rect 225494 698710 225734 698950
rect 225824 698710 226064 698950
rect 226154 698710 226394 698950
rect 226484 698710 226724 698950
rect 226814 698710 227054 698950
rect 225164 698380 225404 698620
rect 225494 698380 225734 698620
rect 225824 698380 226064 698620
rect 226154 698380 226394 698620
rect 226484 698380 226724 698620
rect 226814 698380 227054 698620
rect 225164 698050 225404 698290
rect 225494 698050 225734 698290
rect 225824 698050 226064 698290
rect 226154 698050 226394 698290
rect 226484 698050 226724 698290
rect 226814 698050 227054 698290
rect 225164 697720 225404 697960
rect 225494 697720 225734 697960
rect 225824 697720 226064 697960
rect 226154 697720 226394 697960
rect 226484 697720 226724 697960
rect 226814 697720 227054 697960
rect 225164 697390 225404 697630
rect 225494 697390 225734 697630
rect 225824 697390 226064 697630
rect 226154 697390 226394 697630
rect 226484 697390 226724 697630
rect 226814 697390 227054 697630
rect 225164 697060 225404 697300
rect 225494 697060 225734 697300
rect 225824 697060 226064 697300
rect 226154 697060 226394 697300
rect 226484 697060 226724 697300
rect 226814 697060 227054 697300
rect 225164 696730 225404 696970
rect 225494 696730 225734 696970
rect 225824 696730 226064 696970
rect 226154 696730 226394 696970
rect 226484 696730 226724 696970
rect 226814 696730 227054 696970
rect 225164 696400 225404 696640
rect 225494 696400 225734 696640
rect 225824 696400 226064 696640
rect 226154 696400 226394 696640
rect 226484 696400 226724 696640
rect 226814 696400 227054 696640
rect 225164 696070 225404 696310
rect 225494 696070 225734 696310
rect 225824 696070 226064 696310
rect 226154 696070 226394 696310
rect 226484 696070 226724 696310
rect 226814 696070 227054 696310
rect 217364 692690 217604 692930
rect 217694 692690 217934 692930
rect 218024 692690 218264 692930
rect 218354 692690 218594 692930
rect 218684 692690 218924 692930
rect 219014 692690 219254 692930
rect 219344 692690 219584 692930
rect 219674 692690 219914 692930
rect 220004 692690 220244 692930
rect 220334 692690 220574 692930
rect 220664 692690 220904 692930
rect 220994 692690 221234 692930
rect 221324 692690 221564 692930
rect 221654 692690 221894 692930
rect 221984 692690 222224 692930
rect 217364 692360 217604 692600
rect 217694 692360 217934 692600
rect 218024 692360 218264 692600
rect 218354 692360 218594 692600
rect 218684 692360 218924 692600
rect 219014 692360 219254 692600
rect 219344 692360 219584 692600
rect 219674 692360 219914 692600
rect 220004 692360 220244 692600
rect 220334 692360 220574 692600
rect 220664 692360 220904 692600
rect 220994 692360 221234 692600
rect 221324 692360 221564 692600
rect 221654 692360 221894 692600
rect 221984 692360 222224 692600
rect 217364 692030 217604 692270
rect 217694 692030 217934 692270
rect 218024 692030 218264 692270
rect 218354 692030 218594 692270
rect 218684 692030 218924 692270
rect 219014 692030 219254 692270
rect 219344 692030 219584 692270
rect 219674 692030 219914 692270
rect 220004 692030 220244 692270
rect 220334 692030 220574 692270
rect 220664 692030 220904 692270
rect 220994 692030 221234 692270
rect 221324 692030 221564 692270
rect 221654 692030 221894 692270
rect 221984 692030 222224 692270
rect 217364 691700 217604 691940
rect 217694 691700 217934 691940
rect 218024 691700 218264 691940
rect 218354 691700 218594 691940
rect 218684 691700 218924 691940
rect 219014 691700 219254 691940
rect 219344 691700 219584 691940
rect 219674 691700 219914 691940
rect 220004 691700 220244 691940
rect 220334 691700 220574 691940
rect 220664 691700 220904 691940
rect 220994 691700 221234 691940
rect 221324 691700 221564 691940
rect 221654 691700 221894 691940
rect 221984 691700 222224 691940
rect 217364 691370 217604 691610
rect 217694 691370 217934 691610
rect 218024 691370 218264 691610
rect 218354 691370 218594 691610
rect 218684 691370 218924 691610
rect 219014 691370 219254 691610
rect 219344 691370 219584 691610
rect 219674 691370 219914 691610
rect 220004 691370 220244 691610
rect 220334 691370 220574 691610
rect 220664 691370 220904 691610
rect 220994 691370 221234 691610
rect 221324 691370 221564 691610
rect 221654 691370 221894 691610
rect 221984 691370 222224 691610
rect 217364 691040 217604 691280
rect 217694 691040 217934 691280
rect 218024 691040 218264 691280
rect 218354 691040 218594 691280
rect 218684 691040 218924 691280
rect 219014 691040 219254 691280
rect 219344 691040 219584 691280
rect 219674 691040 219914 691280
rect 220004 691040 220244 691280
rect 220334 691040 220574 691280
rect 220664 691040 220904 691280
rect 220994 691040 221234 691280
rect 221324 691040 221564 691280
rect 221654 691040 221894 691280
rect 221984 691040 222224 691280
rect 217364 690710 217604 690950
rect 217694 690710 217934 690950
rect 218024 690710 218264 690950
rect 218354 690710 218594 690950
rect 218684 690710 218924 690950
rect 219014 690710 219254 690950
rect 219344 690710 219584 690950
rect 219674 690710 219914 690950
rect 220004 690710 220244 690950
rect 220334 690710 220574 690950
rect 220664 690710 220904 690950
rect 220994 690710 221234 690950
rect 221324 690710 221564 690950
rect 221654 690710 221894 690950
rect 221984 690710 222224 690950
rect 217364 690380 217604 690620
rect 217694 690380 217934 690620
rect 218024 690380 218264 690620
rect 218354 690380 218594 690620
rect 218684 690380 218924 690620
rect 219014 690380 219254 690620
rect 219344 690380 219584 690620
rect 219674 690380 219914 690620
rect 220004 690380 220244 690620
rect 220334 690380 220574 690620
rect 220664 690380 220904 690620
rect 220994 690380 221234 690620
rect 221324 690380 221564 690620
rect 221654 690380 221894 690620
rect 221984 690380 222224 690620
rect 217364 690050 217604 690290
rect 217694 690050 217934 690290
rect 218024 690050 218264 690290
rect 218354 690050 218594 690290
rect 218684 690050 218924 690290
rect 219014 690050 219254 690290
rect 219344 690050 219584 690290
rect 219674 690050 219914 690290
rect 220004 690050 220244 690290
rect 220334 690050 220574 690290
rect 220664 690050 220904 690290
rect 220994 690050 221234 690290
rect 221324 690050 221564 690290
rect 221654 690050 221894 690290
rect 221984 690050 222224 690290
rect 217364 689720 217604 689960
rect 217694 689720 217934 689960
rect 218024 689720 218264 689960
rect 218354 689720 218594 689960
rect 218684 689720 218924 689960
rect 219014 689720 219254 689960
rect 219344 689720 219584 689960
rect 219674 689720 219914 689960
rect 220004 689720 220244 689960
rect 220334 689720 220574 689960
rect 220664 689720 220904 689960
rect 220994 689720 221234 689960
rect 221324 689720 221564 689960
rect 221654 689720 221894 689960
rect 221984 689720 222224 689960
rect 217364 689390 217604 689630
rect 217694 689390 217934 689630
rect 218024 689390 218264 689630
rect 218354 689390 218594 689630
rect 218684 689390 218924 689630
rect 219014 689390 219254 689630
rect 219344 689390 219584 689630
rect 219674 689390 219914 689630
rect 220004 689390 220244 689630
rect 220334 689390 220574 689630
rect 220664 689390 220904 689630
rect 220994 689390 221234 689630
rect 221324 689390 221564 689630
rect 221654 689390 221894 689630
rect 221984 689390 222224 689630
rect 217364 689060 217604 689300
rect 217694 689060 217934 689300
rect 218024 689060 218264 689300
rect 218354 689060 218594 689300
rect 218684 689060 218924 689300
rect 219014 689060 219254 689300
rect 219344 689060 219584 689300
rect 219674 689060 219914 689300
rect 220004 689060 220244 689300
rect 220334 689060 220574 689300
rect 220664 689060 220904 689300
rect 220994 689060 221234 689300
rect 221324 689060 221564 689300
rect 221654 689060 221894 689300
rect 221984 689060 222224 689300
rect 217364 688730 217604 688970
rect 217694 688730 217934 688970
rect 218024 688730 218264 688970
rect 218354 688730 218594 688970
rect 218684 688730 218924 688970
rect 219014 688730 219254 688970
rect 219344 688730 219584 688970
rect 219674 688730 219914 688970
rect 220004 688730 220244 688970
rect 220334 688730 220574 688970
rect 220664 688730 220904 688970
rect 220994 688730 221234 688970
rect 221324 688730 221564 688970
rect 221654 688730 221894 688970
rect 221984 688730 222224 688970
rect 217364 688400 217604 688640
rect 217694 688400 217934 688640
rect 218024 688400 218264 688640
rect 218354 688400 218594 688640
rect 218684 688400 218924 688640
rect 219014 688400 219254 688640
rect 219344 688400 219584 688640
rect 219674 688400 219914 688640
rect 220004 688400 220244 688640
rect 220334 688400 220574 688640
rect 220664 688400 220904 688640
rect 220994 688400 221234 688640
rect 221324 688400 221564 688640
rect 221654 688400 221894 688640
rect 221984 688400 222224 688640
rect 217364 688070 217604 688310
rect 217694 688070 217934 688310
rect 218024 688070 218264 688310
rect 218354 688070 218594 688310
rect 218684 688070 218924 688310
rect 219014 688070 219254 688310
rect 219344 688070 219584 688310
rect 219674 688070 219914 688310
rect 220004 688070 220244 688310
rect 220334 688070 220574 688310
rect 220664 688070 220904 688310
rect 220994 688070 221234 688310
rect 221324 688070 221564 688310
rect 221654 688070 221894 688310
rect 221984 688070 222224 688310
rect 227664 692690 227904 692930
rect 227994 692690 228234 692930
rect 228324 692690 228564 692930
rect 228654 692690 228894 692930
rect 228984 692690 229224 692930
rect 229314 692690 229554 692930
rect 229644 692690 229884 692930
rect 229974 692690 230214 692930
rect 230304 692690 230544 692930
rect 230634 692690 230874 692930
rect 230964 692690 231204 692930
rect 231294 692690 231534 692930
rect 231624 692690 231864 692930
rect 231954 692690 232194 692930
rect 232284 692690 232524 692930
rect 227664 692360 227904 692600
rect 227994 692360 228234 692600
rect 228324 692360 228564 692600
rect 228654 692360 228894 692600
rect 228984 692360 229224 692600
rect 229314 692360 229554 692600
rect 229644 692360 229884 692600
rect 229974 692360 230214 692600
rect 230304 692360 230544 692600
rect 230634 692360 230874 692600
rect 230964 692360 231204 692600
rect 231294 692360 231534 692600
rect 231624 692360 231864 692600
rect 231954 692360 232194 692600
rect 232284 692360 232524 692600
rect 227664 692030 227904 692270
rect 227994 692030 228234 692270
rect 228324 692030 228564 692270
rect 228654 692030 228894 692270
rect 228984 692030 229224 692270
rect 229314 692030 229554 692270
rect 229644 692030 229884 692270
rect 229974 692030 230214 692270
rect 230304 692030 230544 692270
rect 230634 692030 230874 692270
rect 230964 692030 231204 692270
rect 231294 692030 231534 692270
rect 231624 692030 231864 692270
rect 231954 692030 232194 692270
rect 232284 692030 232524 692270
rect 227664 691700 227904 691940
rect 227994 691700 228234 691940
rect 228324 691700 228564 691940
rect 228654 691700 228894 691940
rect 228984 691700 229224 691940
rect 229314 691700 229554 691940
rect 229644 691700 229884 691940
rect 229974 691700 230214 691940
rect 230304 691700 230544 691940
rect 230634 691700 230874 691940
rect 230964 691700 231204 691940
rect 231294 691700 231534 691940
rect 231624 691700 231864 691940
rect 231954 691700 232194 691940
rect 232284 691700 232524 691940
rect 227664 691370 227904 691610
rect 227994 691370 228234 691610
rect 228324 691370 228564 691610
rect 228654 691370 228894 691610
rect 228984 691370 229224 691610
rect 229314 691370 229554 691610
rect 229644 691370 229884 691610
rect 229974 691370 230214 691610
rect 230304 691370 230544 691610
rect 230634 691370 230874 691610
rect 230964 691370 231204 691610
rect 231294 691370 231534 691610
rect 231624 691370 231864 691610
rect 231954 691370 232194 691610
rect 232284 691370 232524 691610
rect 227664 691040 227904 691280
rect 227994 691040 228234 691280
rect 228324 691040 228564 691280
rect 228654 691040 228894 691280
rect 228984 691040 229224 691280
rect 229314 691040 229554 691280
rect 229644 691040 229884 691280
rect 229974 691040 230214 691280
rect 230304 691040 230544 691280
rect 230634 691040 230874 691280
rect 230964 691040 231204 691280
rect 231294 691040 231534 691280
rect 231624 691040 231864 691280
rect 231954 691040 232194 691280
rect 232284 691040 232524 691280
rect 227664 690710 227904 690950
rect 227994 690710 228234 690950
rect 228324 690710 228564 690950
rect 228654 690710 228894 690950
rect 228984 690710 229224 690950
rect 229314 690710 229554 690950
rect 229644 690710 229884 690950
rect 229974 690710 230214 690950
rect 230304 690710 230544 690950
rect 230634 690710 230874 690950
rect 230964 690710 231204 690950
rect 231294 690710 231534 690950
rect 231624 690710 231864 690950
rect 231954 690710 232194 690950
rect 232284 690710 232524 690950
rect 227664 690380 227904 690620
rect 227994 690380 228234 690620
rect 228324 690380 228564 690620
rect 228654 690380 228894 690620
rect 228984 690380 229224 690620
rect 229314 690380 229554 690620
rect 229644 690380 229884 690620
rect 229974 690380 230214 690620
rect 230304 690380 230544 690620
rect 230634 690380 230874 690620
rect 230964 690380 231204 690620
rect 231294 690380 231534 690620
rect 231624 690380 231864 690620
rect 231954 690380 232194 690620
rect 232284 690380 232524 690620
rect 227664 690050 227904 690290
rect 227994 690050 228234 690290
rect 228324 690050 228564 690290
rect 228654 690050 228894 690290
rect 228984 690050 229224 690290
rect 229314 690050 229554 690290
rect 229644 690050 229884 690290
rect 229974 690050 230214 690290
rect 230304 690050 230544 690290
rect 230634 690050 230874 690290
rect 230964 690050 231204 690290
rect 231294 690050 231534 690290
rect 231624 690050 231864 690290
rect 231954 690050 232194 690290
rect 232284 690050 232524 690290
rect 227664 689720 227904 689960
rect 227994 689720 228234 689960
rect 228324 689720 228564 689960
rect 228654 689720 228894 689960
rect 228984 689720 229224 689960
rect 229314 689720 229554 689960
rect 229644 689720 229884 689960
rect 229974 689720 230214 689960
rect 230304 689720 230544 689960
rect 230634 689720 230874 689960
rect 230964 689720 231204 689960
rect 231294 689720 231534 689960
rect 231624 689720 231864 689960
rect 231954 689720 232194 689960
rect 232284 689720 232524 689960
rect 227664 689390 227904 689630
rect 227994 689390 228234 689630
rect 228324 689390 228564 689630
rect 228654 689390 228894 689630
rect 228984 689390 229224 689630
rect 229314 689390 229554 689630
rect 229644 689390 229884 689630
rect 229974 689390 230214 689630
rect 230304 689390 230544 689630
rect 230634 689390 230874 689630
rect 230964 689390 231204 689630
rect 231294 689390 231534 689630
rect 231624 689390 231864 689630
rect 231954 689390 232194 689630
rect 232284 689390 232524 689630
rect 227664 689060 227904 689300
rect 227994 689060 228234 689300
rect 228324 689060 228564 689300
rect 228654 689060 228894 689300
rect 228984 689060 229224 689300
rect 229314 689060 229554 689300
rect 229644 689060 229884 689300
rect 229974 689060 230214 689300
rect 230304 689060 230544 689300
rect 230634 689060 230874 689300
rect 230964 689060 231204 689300
rect 231294 689060 231534 689300
rect 231624 689060 231864 689300
rect 231954 689060 232194 689300
rect 232284 689060 232524 689300
rect 227664 688730 227904 688970
rect 227994 688730 228234 688970
rect 228324 688730 228564 688970
rect 228654 688730 228894 688970
rect 228984 688730 229224 688970
rect 229314 688730 229554 688970
rect 229644 688730 229884 688970
rect 229974 688730 230214 688970
rect 230304 688730 230544 688970
rect 230634 688730 230874 688970
rect 230964 688730 231204 688970
rect 231294 688730 231534 688970
rect 231624 688730 231864 688970
rect 231954 688730 232194 688970
rect 232284 688730 232524 688970
rect 227664 688400 227904 688640
rect 227994 688400 228234 688640
rect 228324 688400 228564 688640
rect 228654 688400 228894 688640
rect 228984 688400 229224 688640
rect 229314 688400 229554 688640
rect 229644 688400 229884 688640
rect 229974 688400 230214 688640
rect 230304 688400 230544 688640
rect 230634 688400 230874 688640
rect 230964 688400 231204 688640
rect 231294 688400 231534 688640
rect 231624 688400 231864 688640
rect 231954 688400 232194 688640
rect 232284 688400 232524 688640
rect 227664 688070 227904 688310
rect 227994 688070 228234 688310
rect 228324 688070 228564 688310
rect 228654 688070 228894 688310
rect 228984 688070 229224 688310
rect 229314 688070 229554 688310
rect 229644 688070 229884 688310
rect 229974 688070 230214 688310
rect 230304 688070 230544 688310
rect 230634 688070 230874 688310
rect 230964 688070 231204 688310
rect 231294 688070 231534 688310
rect 231624 688070 231864 688310
rect 231954 688070 232194 688310
rect 232284 688070 232524 688310
rect 82750 668670 82990 668910
rect 83080 668670 83320 668910
rect 83410 668670 83650 668910
rect 83770 668670 84010 668910
rect 84100 668670 84340 668910
rect 84460 668670 84700 668910
rect 84790 668670 85030 668910
rect 82750 668340 82990 668580
rect 83080 668340 83320 668580
rect 83410 668340 83650 668580
rect 83770 668340 84010 668580
rect 84100 668340 84340 668580
rect 84460 668340 84700 668580
rect 84790 668340 85030 668580
rect 82750 668010 82990 668250
rect 83080 668010 83320 668250
rect 83410 668010 83650 668250
rect 83770 668010 84010 668250
rect 84100 668010 84340 668250
rect 84460 668010 84700 668250
rect 84790 668010 85030 668250
rect 82750 667650 82990 667890
rect 83080 667650 83320 667890
rect 83410 667650 83650 667890
rect 83770 667650 84010 667890
rect 84100 667650 84340 667890
rect 84460 667650 84700 667890
rect 84790 667650 85030 667890
rect 82750 667320 82990 667560
rect 83080 667320 83320 667560
rect 83410 667320 83650 667560
rect 83770 667320 84010 667560
rect 84100 667320 84340 667560
rect 84460 667320 84700 667560
rect 84790 667320 85030 667560
rect 82750 666960 82990 667200
rect 83080 666960 83320 667200
rect 83410 666960 83650 667200
rect 83770 666960 84010 667200
rect 84100 666960 84340 667200
rect 84460 666960 84700 667200
rect 84790 666960 85030 667200
rect 82750 666630 82990 666870
rect 83080 666630 83320 666870
rect 83410 666630 83650 666870
rect 83770 666630 84010 666870
rect 84100 666630 84340 666870
rect 84460 666630 84700 666870
rect 84790 666630 85030 666870
rect 82750 666270 82990 666510
rect 83080 666270 83320 666510
rect 83410 666270 83650 666510
rect 83770 666270 84010 666510
rect 84100 666270 84340 666510
rect 84460 666270 84700 666510
rect 84790 666270 85030 666510
rect 82750 665940 82990 666180
rect 83080 665940 83320 666180
rect 83410 665940 83650 666180
rect 83770 665940 84010 666180
rect 84100 665940 84340 666180
rect 84460 665940 84700 666180
rect 84790 665940 85030 666180
rect 82750 665580 82990 665820
rect 83080 665580 83320 665820
rect 83410 665580 83650 665820
rect 83770 665580 84010 665820
rect 84100 665580 84340 665820
rect 84460 665580 84700 665820
rect 84790 665580 85030 665820
rect 82750 665250 82990 665490
rect 83080 665250 83320 665490
rect 83410 665250 83650 665490
rect 83770 665250 84010 665490
rect 84100 665250 84340 665490
rect 84460 665250 84700 665490
rect 84790 665250 85030 665490
rect 82750 664890 82990 665130
rect 83080 664890 83320 665130
rect 83410 664890 83650 665130
rect 83770 664890 84010 665130
rect 84100 664890 84340 665130
rect 84460 664890 84700 665130
rect 84790 664890 85030 665130
rect 82750 664560 82990 664800
rect 83080 664560 83320 664800
rect 83410 664560 83650 664800
rect 83770 664560 84010 664800
rect 84100 664560 84340 664800
rect 84460 664560 84700 664800
rect 84790 664560 85030 664800
rect 82750 664230 82990 664470
rect 83080 664230 83320 664470
rect 83410 664230 83650 664470
rect 83770 664230 84010 664470
rect 84100 664230 84340 664470
rect 84460 664230 84700 664470
rect 84790 664230 85030 664470
rect 82750 656790 82990 657030
rect 83080 656790 83320 657030
rect 83410 656790 83650 657030
rect 83770 656790 84010 657030
rect 84100 656790 84340 657030
rect 84460 656790 84700 657030
rect 84790 656790 85030 657030
rect 82750 656460 82990 656700
rect 83080 656460 83320 656700
rect 83410 656460 83650 656700
rect 83770 656460 84010 656700
rect 84100 656460 84340 656700
rect 84460 656460 84700 656700
rect 84790 656460 85030 656700
rect 82750 656130 82990 656370
rect 83080 656130 83320 656370
rect 83410 656130 83650 656370
rect 83770 656130 84010 656370
rect 84100 656130 84340 656370
rect 84460 656130 84700 656370
rect 84790 656130 85030 656370
rect 3070 655690 3310 655930
rect 3400 655690 3640 655930
rect 3730 655690 3970 655930
rect 4060 655690 4300 655930
rect 4390 655690 4630 655930
rect 4720 655690 4960 655930
rect 5050 655690 5290 655930
rect 5380 655690 5620 655930
rect 5710 655690 5950 655930
rect 6040 655690 6280 655930
rect 6370 655690 6610 655930
rect 6700 655690 6940 655930
rect 7030 655690 7270 655930
rect 7360 655690 7600 655930
rect 7690 655690 7930 655930
rect 82750 655770 82990 656010
rect 83080 655770 83320 656010
rect 83410 655770 83650 656010
rect 83770 655770 84010 656010
rect 84100 655770 84340 656010
rect 84460 655770 84700 656010
rect 84790 655770 85030 656010
rect 3070 655360 3310 655600
rect 3400 655360 3640 655600
rect 3730 655360 3970 655600
rect 4060 655360 4300 655600
rect 4390 655360 4630 655600
rect 4720 655360 4960 655600
rect 5050 655360 5290 655600
rect 5380 655360 5620 655600
rect 5710 655360 5950 655600
rect 6040 655360 6280 655600
rect 6370 655360 6610 655600
rect 6700 655360 6940 655600
rect 7030 655360 7270 655600
rect 7360 655360 7600 655600
rect 7690 655360 7930 655600
rect 82750 655440 82990 655680
rect 83080 655440 83320 655680
rect 83410 655440 83650 655680
rect 83770 655440 84010 655680
rect 84100 655440 84340 655680
rect 84460 655440 84700 655680
rect 84790 655440 85030 655680
rect 3070 655030 3310 655270
rect 3400 655030 3640 655270
rect 3730 655030 3970 655270
rect 4060 655030 4300 655270
rect 4390 655030 4630 655270
rect 4720 655030 4960 655270
rect 5050 655030 5290 655270
rect 5380 655030 5620 655270
rect 5710 655030 5950 655270
rect 6040 655030 6280 655270
rect 6370 655030 6610 655270
rect 6700 655030 6940 655270
rect 7030 655030 7270 655270
rect 7360 655030 7600 655270
rect 7690 655030 7930 655270
rect 82750 655080 82990 655320
rect 83080 655080 83320 655320
rect 83410 655080 83650 655320
rect 83770 655080 84010 655320
rect 84100 655080 84340 655320
rect 84460 655080 84700 655320
rect 84790 655080 85030 655320
rect 3070 654700 3310 654940
rect 3400 654700 3640 654940
rect 3730 654700 3970 654940
rect 4060 654700 4300 654940
rect 4390 654700 4630 654940
rect 4720 654700 4960 654940
rect 5050 654700 5290 654940
rect 5380 654700 5620 654940
rect 5710 654700 5950 654940
rect 6040 654700 6280 654940
rect 6370 654700 6610 654940
rect 6700 654700 6940 654940
rect 7030 654700 7270 654940
rect 7360 654700 7600 654940
rect 7690 654700 7930 654940
rect 82750 654750 82990 654990
rect 83080 654750 83320 654990
rect 83410 654750 83650 654990
rect 83770 654750 84010 654990
rect 84100 654750 84340 654990
rect 84460 654750 84700 654990
rect 84790 654750 85030 654990
rect 3070 654370 3310 654610
rect 3400 654370 3640 654610
rect 3730 654370 3970 654610
rect 4060 654370 4300 654610
rect 4390 654370 4630 654610
rect 4720 654370 4960 654610
rect 5050 654370 5290 654610
rect 5380 654370 5620 654610
rect 5710 654370 5950 654610
rect 6040 654370 6280 654610
rect 6370 654370 6610 654610
rect 6700 654370 6940 654610
rect 7030 654370 7270 654610
rect 7360 654370 7600 654610
rect 7690 654370 7930 654610
rect 82750 654390 82990 654630
rect 83080 654390 83320 654630
rect 83410 654390 83650 654630
rect 83770 654390 84010 654630
rect 84100 654390 84340 654630
rect 84460 654390 84700 654630
rect 84790 654390 85030 654630
rect 3070 654040 3310 654280
rect 3400 654040 3640 654280
rect 3730 654040 3970 654280
rect 4060 654040 4300 654280
rect 4390 654040 4630 654280
rect 4720 654040 4960 654280
rect 5050 654040 5290 654280
rect 5380 654040 5620 654280
rect 5710 654040 5950 654280
rect 6040 654040 6280 654280
rect 6370 654040 6610 654280
rect 6700 654040 6940 654280
rect 7030 654040 7270 654280
rect 7360 654040 7600 654280
rect 7690 654040 7930 654280
rect 82750 654060 82990 654300
rect 83080 654060 83320 654300
rect 83410 654060 83650 654300
rect 83770 654060 84010 654300
rect 84100 654060 84340 654300
rect 84460 654060 84700 654300
rect 84790 654060 85030 654300
rect 3070 653710 3310 653950
rect 3400 653710 3640 653950
rect 3730 653710 3970 653950
rect 4060 653710 4300 653950
rect 4390 653710 4630 653950
rect 4720 653710 4960 653950
rect 5050 653710 5290 653950
rect 5380 653710 5620 653950
rect 5710 653710 5950 653950
rect 6040 653710 6280 653950
rect 6370 653710 6610 653950
rect 6700 653710 6940 653950
rect 7030 653710 7270 653950
rect 7360 653710 7600 653950
rect 7690 653710 7930 653950
rect 82750 653700 82990 653940
rect 83080 653700 83320 653940
rect 83410 653700 83650 653940
rect 83770 653700 84010 653940
rect 84100 653700 84340 653940
rect 84460 653700 84700 653940
rect 84790 653700 85030 653940
rect 3070 653380 3310 653620
rect 3400 653380 3640 653620
rect 3730 653380 3970 653620
rect 4060 653380 4300 653620
rect 4390 653380 4630 653620
rect 4720 653380 4960 653620
rect 5050 653380 5290 653620
rect 5380 653380 5620 653620
rect 5710 653380 5950 653620
rect 6040 653380 6280 653620
rect 6370 653380 6610 653620
rect 6700 653380 6940 653620
rect 7030 653380 7270 653620
rect 7360 653380 7600 653620
rect 7690 653380 7930 653620
rect 82750 653370 82990 653610
rect 83080 653370 83320 653610
rect 83410 653370 83650 653610
rect 83770 653370 84010 653610
rect 84100 653370 84340 653610
rect 84460 653370 84700 653610
rect 84790 653370 85030 653610
rect 3070 653050 3310 653290
rect 3400 653050 3640 653290
rect 3730 653050 3970 653290
rect 4060 653050 4300 653290
rect 4390 653050 4630 653290
rect 4720 653050 4960 653290
rect 5050 653050 5290 653290
rect 5380 653050 5620 653290
rect 5710 653050 5950 653290
rect 6040 653050 6280 653290
rect 6370 653050 6610 653290
rect 6700 653050 6940 653290
rect 7030 653050 7270 653290
rect 7360 653050 7600 653290
rect 7690 653050 7930 653290
rect 82750 653010 82990 653250
rect 83080 653010 83320 653250
rect 83410 653010 83650 653250
rect 83770 653010 84010 653250
rect 84100 653010 84340 653250
rect 84460 653010 84700 653250
rect 84790 653010 85030 653250
rect 3070 652720 3310 652960
rect 3400 652720 3640 652960
rect 3730 652720 3970 652960
rect 4060 652720 4300 652960
rect 4390 652720 4630 652960
rect 4720 652720 4960 652960
rect 5050 652720 5290 652960
rect 5380 652720 5620 652960
rect 5710 652720 5950 652960
rect 6040 652720 6280 652960
rect 6370 652720 6610 652960
rect 6700 652720 6940 652960
rect 7030 652720 7270 652960
rect 7360 652720 7600 652960
rect 7690 652720 7930 652960
rect 82750 652680 82990 652920
rect 83080 652680 83320 652920
rect 83410 652680 83650 652920
rect 83770 652680 84010 652920
rect 84100 652680 84340 652920
rect 84460 652680 84700 652920
rect 84790 652680 85030 652920
rect 3070 652390 3310 652630
rect 3400 652390 3640 652630
rect 3730 652390 3970 652630
rect 4060 652390 4300 652630
rect 4390 652390 4630 652630
rect 4720 652390 4960 652630
rect 5050 652390 5290 652630
rect 5380 652390 5620 652630
rect 5710 652390 5950 652630
rect 6040 652390 6280 652630
rect 6370 652390 6610 652630
rect 6700 652390 6940 652630
rect 7030 652390 7270 652630
rect 7360 652390 7600 652630
rect 7690 652390 7930 652630
rect 82750 652350 82990 652590
rect 83080 652350 83320 652590
rect 83410 652350 83650 652590
rect 83770 652350 84010 652590
rect 84100 652350 84340 652590
rect 84460 652350 84700 652590
rect 84790 652350 85030 652590
rect 3070 652060 3310 652300
rect 3400 652060 3640 652300
rect 3730 652060 3970 652300
rect 4060 652060 4300 652300
rect 4390 652060 4630 652300
rect 4720 652060 4960 652300
rect 5050 652060 5290 652300
rect 5380 652060 5620 652300
rect 5710 652060 5950 652300
rect 6040 652060 6280 652300
rect 6370 652060 6610 652300
rect 6700 652060 6940 652300
rect 7030 652060 7270 652300
rect 7360 652060 7600 652300
rect 7690 652060 7930 652300
rect 3070 651730 3310 651970
rect 3400 651730 3640 651970
rect 3730 651730 3970 651970
rect 4060 651730 4300 651970
rect 4390 651730 4630 651970
rect 4720 651730 4960 651970
rect 5050 651730 5290 651970
rect 5380 651730 5620 651970
rect 5710 651730 5950 651970
rect 6040 651730 6280 651970
rect 6370 651730 6610 651970
rect 6700 651730 6940 651970
rect 7030 651730 7270 651970
rect 7360 651730 7600 651970
rect 7690 651730 7930 651970
rect 3070 651400 3310 651640
rect 3400 651400 3640 651640
rect 3730 651400 3970 651640
rect 4060 651400 4300 651640
rect 4390 651400 4630 651640
rect 4720 651400 4960 651640
rect 5050 651400 5290 651640
rect 5380 651400 5620 651640
rect 5710 651400 5950 651640
rect 6040 651400 6280 651640
rect 6370 651400 6610 651640
rect 6700 651400 6940 651640
rect 7030 651400 7270 651640
rect 7360 651400 7600 651640
rect 7690 651400 7930 651640
rect 3070 651070 3310 651310
rect 3400 651070 3640 651310
rect 3730 651070 3970 651310
rect 4060 651070 4300 651310
rect 4390 651070 4630 651310
rect 4720 651070 4960 651310
rect 5050 651070 5290 651310
rect 5380 651070 5620 651310
rect 5710 651070 5950 651310
rect 6040 651070 6280 651310
rect 6370 651070 6610 651310
rect 6700 651070 6940 651310
rect 7030 651070 7270 651310
rect 7360 651070 7600 651310
rect 7690 651070 7930 651310
<< metal5 >>
rect 165594 701000 170594 704800
rect 175894 701000 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 3000 700930 581000 701000
rect 3000 700690 225164 700930
rect 225404 700690 225494 700930
rect 225734 700690 225824 700930
rect 226064 700690 226154 700930
rect 226394 700690 226484 700930
rect 226724 700690 226814 700930
rect 227054 700690 581000 700930
rect 3000 700600 581000 700690
rect 3000 700360 225164 700600
rect 225404 700360 225494 700600
rect 225734 700360 225824 700600
rect 226064 700360 226154 700600
rect 226394 700360 226484 700600
rect 226724 700360 226814 700600
rect 227054 700360 581000 700600
rect 3000 700270 581000 700360
rect 3000 700030 225164 700270
rect 225404 700030 225494 700270
rect 225734 700030 225824 700270
rect 226064 700030 226154 700270
rect 226394 700030 226484 700270
rect 226724 700030 226814 700270
rect 227054 700030 581000 700270
rect 3000 699940 581000 700030
rect 3000 699700 225164 699940
rect 225404 699700 225494 699940
rect 225734 699700 225824 699940
rect 226064 699700 226154 699940
rect 226394 699700 226484 699940
rect 226724 699700 226814 699940
rect 227054 699700 581000 699940
rect 3000 699610 581000 699700
rect 3000 699370 225164 699610
rect 225404 699370 225494 699610
rect 225734 699370 225824 699610
rect 226064 699370 226154 699610
rect 226394 699370 226484 699610
rect 226724 699370 226814 699610
rect 227054 699370 581000 699610
rect 3000 699280 581000 699370
rect 3000 699040 225164 699280
rect 225404 699040 225494 699280
rect 225734 699040 225824 699280
rect 226064 699040 226154 699280
rect 226394 699040 226484 699280
rect 226724 699040 226814 699280
rect 227054 699040 581000 699280
rect 3000 698950 581000 699040
rect 3000 698710 225164 698950
rect 225404 698710 225494 698950
rect 225734 698710 225824 698950
rect 226064 698710 226154 698950
rect 226394 698710 226484 698950
rect 226724 698710 226814 698950
rect 227054 698710 581000 698950
rect 3000 698620 581000 698710
rect 3000 698380 225164 698620
rect 225404 698380 225494 698620
rect 225734 698380 225824 698620
rect 226064 698380 226154 698620
rect 226394 698380 226484 698620
rect 226724 698380 226814 698620
rect 227054 698380 581000 698620
rect 3000 698290 581000 698380
rect 3000 698050 225164 698290
rect 225404 698050 225494 698290
rect 225734 698050 225824 698290
rect 226064 698050 226154 698290
rect 226394 698050 226484 698290
rect 226724 698050 226814 698290
rect 227054 698050 581000 698290
rect 3000 697960 581000 698050
rect 3000 697720 225164 697960
rect 225404 697720 225494 697960
rect 225734 697720 225824 697960
rect 226064 697720 226154 697960
rect 226394 697720 226484 697960
rect 226724 697720 226814 697960
rect 227054 697720 581000 697960
rect 3000 697630 581000 697720
rect 3000 697390 225164 697630
rect 225404 697390 225494 697630
rect 225734 697390 225824 697630
rect 226064 697390 226154 697630
rect 226394 697390 226484 697630
rect 226724 697390 226814 697630
rect 227054 697390 581000 697630
rect 3000 697300 581000 697390
rect 3000 697060 225164 697300
rect 225404 697060 225494 697300
rect 225734 697060 225824 697300
rect 226064 697060 226154 697300
rect 226394 697060 226484 697300
rect 226724 697060 226814 697300
rect 227054 697060 581000 697300
rect 3000 696970 581000 697060
rect 3000 696730 225164 696970
rect 225404 696730 225494 696970
rect 225734 696730 225824 696970
rect 226064 696730 226154 696970
rect 226394 696730 226484 696970
rect 226724 696730 226814 696970
rect 227054 696730 581000 696970
rect 3000 696640 581000 696730
rect 3000 696400 225164 696640
rect 225404 696400 225494 696640
rect 225734 696400 225824 696640
rect 226064 696400 226154 696640
rect 226394 696400 226484 696640
rect 226724 696400 226814 696640
rect 227054 696400 581000 696640
rect 3000 696310 581000 696400
rect 3000 696070 225164 696310
rect 225404 696070 225494 696310
rect 225734 696070 225824 696310
rect 226064 696070 226154 696310
rect 226394 696070 226484 696310
rect 226724 696070 226814 696310
rect 227054 696070 581000 696310
rect 3000 696000 581000 696070
rect 3000 655930 8000 696000
rect 3000 655690 3070 655930
rect 3310 655690 3400 655930
rect 3640 655690 3730 655930
rect 3970 655690 4060 655930
rect 4300 655690 4390 655930
rect 4630 655690 4720 655930
rect 4960 655690 5050 655930
rect 5290 655690 5380 655930
rect 5620 655690 5710 655930
rect 5950 655690 6040 655930
rect 6280 655690 6370 655930
rect 6610 655690 6700 655930
rect 6940 655690 7030 655930
rect 7270 655690 7360 655930
rect 7600 655690 7690 655930
rect 7930 655690 8000 655930
rect 3000 655600 8000 655690
rect 3000 655360 3070 655600
rect 3310 655360 3400 655600
rect 3640 655360 3730 655600
rect 3970 655360 4060 655600
rect 4300 655360 4390 655600
rect 4630 655360 4720 655600
rect 4960 655360 5050 655600
rect 5290 655360 5380 655600
rect 5620 655360 5710 655600
rect 5950 655360 6040 655600
rect 6280 655360 6370 655600
rect 6610 655360 6700 655600
rect 6940 655360 7030 655600
rect 7270 655360 7360 655600
rect 7600 655360 7690 655600
rect 7930 655360 8000 655600
rect 3000 655270 8000 655360
rect 3000 655030 3070 655270
rect 3310 655030 3400 655270
rect 3640 655030 3730 655270
rect 3970 655030 4060 655270
rect 4300 655030 4390 655270
rect 4630 655030 4720 655270
rect 4960 655030 5050 655270
rect 5290 655030 5380 655270
rect 5620 655030 5710 655270
rect 5950 655030 6040 655270
rect 6280 655030 6370 655270
rect 6610 655030 6700 655270
rect 6940 655030 7030 655270
rect 7270 655030 7360 655270
rect 7600 655030 7690 655270
rect 7930 655030 8000 655270
rect 3000 654940 8000 655030
rect 3000 654700 3070 654940
rect 3310 654700 3400 654940
rect 3640 654700 3730 654940
rect 3970 654700 4060 654940
rect 4300 654700 4390 654940
rect 4630 654700 4720 654940
rect 4960 654700 5050 654940
rect 5290 654700 5380 654940
rect 5620 654700 5710 654940
rect 5950 654700 6040 654940
rect 6280 654700 6370 654940
rect 6610 654700 6700 654940
rect 6940 654700 7030 654940
rect 7270 654700 7360 654940
rect 7600 654700 7690 654940
rect 7930 654700 8000 654940
rect 3000 654610 8000 654700
rect 3000 654370 3070 654610
rect 3310 654370 3400 654610
rect 3640 654370 3730 654610
rect 3970 654370 4060 654610
rect 4300 654370 4390 654610
rect 4630 654370 4720 654610
rect 4960 654370 5050 654610
rect 5290 654370 5380 654610
rect 5620 654370 5710 654610
rect 5950 654370 6040 654610
rect 6280 654370 6370 654610
rect 6610 654370 6700 654610
rect 6940 654370 7030 654610
rect 7270 654370 7360 654610
rect 7600 654370 7690 654610
rect 7930 654370 8000 654610
rect 3000 654280 8000 654370
rect 3000 654040 3070 654280
rect 3310 654040 3400 654280
rect 3640 654040 3730 654280
rect 3970 654040 4060 654280
rect 4300 654040 4390 654280
rect 4630 654040 4720 654280
rect 4960 654040 5050 654280
rect 5290 654040 5380 654280
rect 5620 654040 5710 654280
rect 5950 654040 6040 654280
rect 6280 654040 6370 654280
rect 6610 654040 6700 654280
rect 6940 654040 7030 654280
rect 7270 654040 7360 654280
rect 7600 654040 7690 654280
rect 7930 654040 8000 654280
rect 3000 653950 8000 654040
rect 3000 653710 3070 653950
rect 3310 653710 3400 653950
rect 3640 653710 3730 653950
rect 3970 653710 4060 653950
rect 4300 653710 4390 653950
rect 4630 653710 4720 653950
rect 4960 653710 5050 653950
rect 5290 653710 5380 653950
rect 5620 653710 5710 653950
rect 5950 653710 6040 653950
rect 6280 653710 6370 653950
rect 6610 653710 6700 653950
rect 6940 653710 7030 653950
rect 7270 653710 7360 653950
rect 7600 653710 7690 653950
rect 7930 653710 8000 653950
rect 3000 653620 8000 653710
rect 3000 653380 3070 653620
rect 3310 653380 3400 653620
rect 3640 653380 3730 653620
rect 3970 653380 4060 653620
rect 4300 653380 4390 653620
rect 4630 653380 4720 653620
rect 4960 653380 5050 653620
rect 5290 653380 5380 653620
rect 5620 653380 5710 653620
rect 5950 653380 6040 653620
rect 6280 653380 6370 653620
rect 6610 653380 6700 653620
rect 6940 653380 7030 653620
rect 7270 653380 7360 653620
rect 7600 653380 7690 653620
rect 7930 653380 8000 653620
rect 3000 653290 8000 653380
rect 3000 653050 3070 653290
rect 3310 653050 3400 653290
rect 3640 653050 3730 653290
rect 3970 653050 4060 653290
rect 4300 653050 4390 653290
rect 4630 653050 4720 653290
rect 4960 653050 5050 653290
rect 5290 653050 5380 653290
rect 5620 653050 5710 653290
rect 5950 653050 6040 653290
rect 6280 653050 6370 653290
rect 6610 653050 6700 653290
rect 6940 653050 7030 653290
rect 7270 653050 7360 653290
rect 7600 653050 7690 653290
rect 7930 653050 8000 653290
rect 3000 652960 8000 653050
rect 3000 652720 3070 652960
rect 3310 652720 3400 652960
rect 3640 652720 3730 652960
rect 3970 652720 4060 652960
rect 4300 652720 4390 652960
rect 4630 652720 4720 652960
rect 4960 652720 5050 652960
rect 5290 652720 5380 652960
rect 5620 652720 5710 652960
rect 5950 652720 6040 652960
rect 6280 652720 6370 652960
rect 6610 652720 6700 652960
rect 6940 652720 7030 652960
rect 7270 652720 7360 652960
rect 7600 652720 7690 652960
rect 7930 652720 8000 652960
rect 3000 652630 8000 652720
rect 3000 652390 3070 652630
rect 3310 652390 3400 652630
rect 3640 652390 3730 652630
rect 3970 652390 4060 652630
rect 4300 652390 4390 652630
rect 4630 652390 4720 652630
rect 4960 652390 5050 652630
rect 5290 652390 5380 652630
rect 5620 652390 5710 652630
rect 5950 652390 6040 652630
rect 6280 652390 6370 652630
rect 6610 652390 6700 652630
rect 6940 652390 7030 652630
rect 7270 652390 7360 652630
rect 7600 652390 7690 652630
rect 7930 652390 8000 652630
rect 3000 652300 8000 652390
rect 3000 652060 3070 652300
rect 3310 652060 3400 652300
rect 3640 652060 3730 652300
rect 3970 652060 4060 652300
rect 4300 652060 4390 652300
rect 4630 652060 4720 652300
rect 4960 652060 5050 652300
rect 5290 652060 5380 652300
rect 5620 652060 5710 652300
rect 5950 652060 6040 652300
rect 6280 652060 6370 652300
rect 6610 652060 6700 652300
rect 6940 652060 7030 652300
rect 7270 652060 7360 652300
rect 7600 652060 7690 652300
rect 7930 652060 8000 652300
rect 3000 651970 8000 652060
rect 3000 651730 3070 651970
rect 3310 651730 3400 651970
rect 3640 651730 3730 651970
rect 3970 651730 4060 651970
rect 4300 651730 4390 651970
rect 4630 651730 4720 651970
rect 4960 651730 5050 651970
rect 5290 651730 5380 651970
rect 5620 651730 5710 651970
rect 5950 651730 6040 651970
rect 6280 651730 6370 651970
rect 6610 651730 6700 651970
rect 6940 651730 7030 651970
rect 7270 651730 7360 651970
rect 7600 651730 7690 651970
rect 7930 651730 8000 651970
rect 3000 651640 8000 651730
rect 3000 651400 3070 651640
rect 3310 651400 3400 651640
rect 3640 651400 3730 651640
rect 3970 651400 4060 651640
rect 4300 651400 4390 651640
rect 4630 651400 4720 651640
rect 4960 651400 5050 651640
rect 5290 651400 5380 651640
rect 5620 651400 5710 651640
rect 5950 651400 6040 651640
rect 6280 651400 6370 651640
rect 6610 651400 6700 651640
rect 6940 651400 7030 651640
rect 7270 651400 7360 651640
rect 7600 651400 7690 651640
rect 7930 651400 8000 651640
rect 3000 651310 8000 651400
rect 3000 651070 3070 651310
rect 3310 651070 3400 651310
rect 3640 651070 3730 651310
rect 3970 651070 4060 651310
rect 4300 651070 4390 651310
rect 4630 651070 4720 651310
rect 4960 651070 5050 651310
rect 5290 651070 5380 651310
rect 5620 651070 5710 651310
rect 5950 651070 6040 651310
rect 6280 651070 6370 651310
rect 6610 651070 6700 651310
rect 6940 651070 7030 651310
rect 7270 651070 7360 651310
rect 7600 651070 7690 651310
rect 7930 651070 8000 651310
rect 3000 651000 8000 651070
rect 11000 692930 573000 693000
rect 11000 692690 170964 692930
rect 171204 692690 171294 692930
rect 171534 692690 171624 692930
rect 171864 692690 171954 692930
rect 172194 692690 172284 692930
rect 172524 692690 172614 692930
rect 172854 692690 217364 692930
rect 217604 692690 217694 692930
rect 217934 692690 218024 692930
rect 218264 692690 218354 692930
rect 218594 692690 218684 692930
rect 218924 692690 219014 692930
rect 219254 692690 219344 692930
rect 219584 692690 219674 692930
rect 219914 692690 220004 692930
rect 220244 692690 220334 692930
rect 220574 692690 220664 692930
rect 220904 692690 220994 692930
rect 221234 692690 221324 692930
rect 221564 692690 221654 692930
rect 221894 692690 221984 692930
rect 222224 692690 227664 692930
rect 227904 692690 227994 692930
rect 228234 692690 228324 692930
rect 228564 692690 228654 692930
rect 228894 692690 228984 692930
rect 229224 692690 229314 692930
rect 229554 692690 229644 692930
rect 229884 692690 229974 692930
rect 230214 692690 230304 692930
rect 230544 692690 230634 692930
rect 230874 692690 230964 692930
rect 231204 692690 231294 692930
rect 231534 692690 231624 692930
rect 231864 692690 231954 692930
rect 232194 692690 232284 692930
rect 232524 692690 573000 692930
rect 11000 692600 573000 692690
rect 11000 692360 170964 692600
rect 171204 692360 171294 692600
rect 171534 692360 171624 692600
rect 171864 692360 171954 692600
rect 172194 692360 172284 692600
rect 172524 692360 172614 692600
rect 172854 692360 217364 692600
rect 217604 692360 217694 692600
rect 217934 692360 218024 692600
rect 218264 692360 218354 692600
rect 218594 692360 218684 692600
rect 218924 692360 219014 692600
rect 219254 692360 219344 692600
rect 219584 692360 219674 692600
rect 219914 692360 220004 692600
rect 220244 692360 220334 692600
rect 220574 692360 220664 692600
rect 220904 692360 220994 692600
rect 221234 692360 221324 692600
rect 221564 692360 221654 692600
rect 221894 692360 221984 692600
rect 222224 692360 227664 692600
rect 227904 692360 227994 692600
rect 228234 692360 228324 692600
rect 228564 692360 228654 692600
rect 228894 692360 228984 692600
rect 229224 692360 229314 692600
rect 229554 692360 229644 692600
rect 229884 692360 229974 692600
rect 230214 692360 230304 692600
rect 230544 692360 230634 692600
rect 230874 692360 230964 692600
rect 231204 692360 231294 692600
rect 231534 692360 231624 692600
rect 231864 692360 231954 692600
rect 232194 692360 232284 692600
rect 232524 692360 573000 692600
rect 11000 692270 573000 692360
rect 11000 692030 170964 692270
rect 171204 692030 171294 692270
rect 171534 692030 171624 692270
rect 171864 692030 171954 692270
rect 172194 692030 172284 692270
rect 172524 692030 172614 692270
rect 172854 692030 217364 692270
rect 217604 692030 217694 692270
rect 217934 692030 218024 692270
rect 218264 692030 218354 692270
rect 218594 692030 218684 692270
rect 218924 692030 219014 692270
rect 219254 692030 219344 692270
rect 219584 692030 219674 692270
rect 219914 692030 220004 692270
rect 220244 692030 220334 692270
rect 220574 692030 220664 692270
rect 220904 692030 220994 692270
rect 221234 692030 221324 692270
rect 221564 692030 221654 692270
rect 221894 692030 221984 692270
rect 222224 692030 227664 692270
rect 227904 692030 227994 692270
rect 228234 692030 228324 692270
rect 228564 692030 228654 692270
rect 228894 692030 228984 692270
rect 229224 692030 229314 692270
rect 229554 692030 229644 692270
rect 229884 692030 229974 692270
rect 230214 692030 230304 692270
rect 230544 692030 230634 692270
rect 230874 692030 230964 692270
rect 231204 692030 231294 692270
rect 231534 692030 231624 692270
rect 231864 692030 231954 692270
rect 232194 692030 232284 692270
rect 232524 692030 573000 692270
rect 11000 691940 573000 692030
rect 11000 691700 170964 691940
rect 171204 691700 171294 691940
rect 171534 691700 171624 691940
rect 171864 691700 171954 691940
rect 172194 691700 172284 691940
rect 172524 691700 172614 691940
rect 172854 691700 217364 691940
rect 217604 691700 217694 691940
rect 217934 691700 218024 691940
rect 218264 691700 218354 691940
rect 218594 691700 218684 691940
rect 218924 691700 219014 691940
rect 219254 691700 219344 691940
rect 219584 691700 219674 691940
rect 219914 691700 220004 691940
rect 220244 691700 220334 691940
rect 220574 691700 220664 691940
rect 220904 691700 220994 691940
rect 221234 691700 221324 691940
rect 221564 691700 221654 691940
rect 221894 691700 221984 691940
rect 222224 691700 227664 691940
rect 227904 691700 227994 691940
rect 228234 691700 228324 691940
rect 228564 691700 228654 691940
rect 228894 691700 228984 691940
rect 229224 691700 229314 691940
rect 229554 691700 229644 691940
rect 229884 691700 229974 691940
rect 230214 691700 230304 691940
rect 230544 691700 230634 691940
rect 230874 691700 230964 691940
rect 231204 691700 231294 691940
rect 231534 691700 231624 691940
rect 231864 691700 231954 691940
rect 232194 691700 232284 691940
rect 232524 691700 573000 691940
rect 11000 691610 573000 691700
rect 11000 691370 170964 691610
rect 171204 691370 171294 691610
rect 171534 691370 171624 691610
rect 171864 691370 171954 691610
rect 172194 691370 172284 691610
rect 172524 691370 172614 691610
rect 172854 691370 217364 691610
rect 217604 691370 217694 691610
rect 217934 691370 218024 691610
rect 218264 691370 218354 691610
rect 218594 691370 218684 691610
rect 218924 691370 219014 691610
rect 219254 691370 219344 691610
rect 219584 691370 219674 691610
rect 219914 691370 220004 691610
rect 220244 691370 220334 691610
rect 220574 691370 220664 691610
rect 220904 691370 220994 691610
rect 221234 691370 221324 691610
rect 221564 691370 221654 691610
rect 221894 691370 221984 691610
rect 222224 691370 227664 691610
rect 227904 691370 227994 691610
rect 228234 691370 228324 691610
rect 228564 691370 228654 691610
rect 228894 691370 228984 691610
rect 229224 691370 229314 691610
rect 229554 691370 229644 691610
rect 229884 691370 229974 691610
rect 230214 691370 230304 691610
rect 230544 691370 230634 691610
rect 230874 691370 230964 691610
rect 231204 691370 231294 691610
rect 231534 691370 231624 691610
rect 231864 691370 231954 691610
rect 232194 691370 232284 691610
rect 232524 691370 573000 691610
rect 11000 691280 573000 691370
rect 11000 691040 170964 691280
rect 171204 691040 171294 691280
rect 171534 691040 171624 691280
rect 171864 691040 171954 691280
rect 172194 691040 172284 691280
rect 172524 691040 172614 691280
rect 172854 691040 217364 691280
rect 217604 691040 217694 691280
rect 217934 691040 218024 691280
rect 218264 691040 218354 691280
rect 218594 691040 218684 691280
rect 218924 691040 219014 691280
rect 219254 691040 219344 691280
rect 219584 691040 219674 691280
rect 219914 691040 220004 691280
rect 220244 691040 220334 691280
rect 220574 691040 220664 691280
rect 220904 691040 220994 691280
rect 221234 691040 221324 691280
rect 221564 691040 221654 691280
rect 221894 691040 221984 691280
rect 222224 691040 227664 691280
rect 227904 691040 227994 691280
rect 228234 691040 228324 691280
rect 228564 691040 228654 691280
rect 228894 691040 228984 691280
rect 229224 691040 229314 691280
rect 229554 691040 229644 691280
rect 229884 691040 229974 691280
rect 230214 691040 230304 691280
rect 230544 691040 230634 691280
rect 230874 691040 230964 691280
rect 231204 691040 231294 691280
rect 231534 691040 231624 691280
rect 231864 691040 231954 691280
rect 232194 691040 232284 691280
rect 232524 691040 573000 691280
rect 11000 690950 573000 691040
rect 11000 690710 170964 690950
rect 171204 690710 171294 690950
rect 171534 690710 171624 690950
rect 171864 690710 171954 690950
rect 172194 690710 172284 690950
rect 172524 690710 172614 690950
rect 172854 690710 217364 690950
rect 217604 690710 217694 690950
rect 217934 690710 218024 690950
rect 218264 690710 218354 690950
rect 218594 690710 218684 690950
rect 218924 690710 219014 690950
rect 219254 690710 219344 690950
rect 219584 690710 219674 690950
rect 219914 690710 220004 690950
rect 220244 690710 220334 690950
rect 220574 690710 220664 690950
rect 220904 690710 220994 690950
rect 221234 690710 221324 690950
rect 221564 690710 221654 690950
rect 221894 690710 221984 690950
rect 222224 690710 227664 690950
rect 227904 690710 227994 690950
rect 228234 690710 228324 690950
rect 228564 690710 228654 690950
rect 228894 690710 228984 690950
rect 229224 690710 229314 690950
rect 229554 690710 229644 690950
rect 229884 690710 229974 690950
rect 230214 690710 230304 690950
rect 230544 690710 230634 690950
rect 230874 690710 230964 690950
rect 231204 690710 231294 690950
rect 231534 690710 231624 690950
rect 231864 690710 231954 690950
rect 232194 690710 232284 690950
rect 232524 690710 573000 690950
rect 11000 690620 573000 690710
rect 11000 690380 170964 690620
rect 171204 690380 171294 690620
rect 171534 690380 171624 690620
rect 171864 690380 171954 690620
rect 172194 690380 172284 690620
rect 172524 690380 172614 690620
rect 172854 690380 217364 690620
rect 217604 690380 217694 690620
rect 217934 690380 218024 690620
rect 218264 690380 218354 690620
rect 218594 690380 218684 690620
rect 218924 690380 219014 690620
rect 219254 690380 219344 690620
rect 219584 690380 219674 690620
rect 219914 690380 220004 690620
rect 220244 690380 220334 690620
rect 220574 690380 220664 690620
rect 220904 690380 220994 690620
rect 221234 690380 221324 690620
rect 221564 690380 221654 690620
rect 221894 690380 221984 690620
rect 222224 690380 227664 690620
rect 227904 690380 227994 690620
rect 228234 690380 228324 690620
rect 228564 690380 228654 690620
rect 228894 690380 228984 690620
rect 229224 690380 229314 690620
rect 229554 690380 229644 690620
rect 229884 690380 229974 690620
rect 230214 690380 230304 690620
rect 230544 690380 230634 690620
rect 230874 690380 230964 690620
rect 231204 690380 231294 690620
rect 231534 690380 231624 690620
rect 231864 690380 231954 690620
rect 232194 690380 232284 690620
rect 232524 690380 573000 690620
rect 11000 690290 573000 690380
rect 11000 690050 170964 690290
rect 171204 690050 171294 690290
rect 171534 690050 171624 690290
rect 171864 690050 171954 690290
rect 172194 690050 172284 690290
rect 172524 690050 172614 690290
rect 172854 690050 217364 690290
rect 217604 690050 217694 690290
rect 217934 690050 218024 690290
rect 218264 690050 218354 690290
rect 218594 690050 218684 690290
rect 218924 690050 219014 690290
rect 219254 690050 219344 690290
rect 219584 690050 219674 690290
rect 219914 690050 220004 690290
rect 220244 690050 220334 690290
rect 220574 690050 220664 690290
rect 220904 690050 220994 690290
rect 221234 690050 221324 690290
rect 221564 690050 221654 690290
rect 221894 690050 221984 690290
rect 222224 690050 227664 690290
rect 227904 690050 227994 690290
rect 228234 690050 228324 690290
rect 228564 690050 228654 690290
rect 228894 690050 228984 690290
rect 229224 690050 229314 690290
rect 229554 690050 229644 690290
rect 229884 690050 229974 690290
rect 230214 690050 230304 690290
rect 230544 690050 230634 690290
rect 230874 690050 230964 690290
rect 231204 690050 231294 690290
rect 231534 690050 231624 690290
rect 231864 690050 231954 690290
rect 232194 690050 232284 690290
rect 232524 690050 573000 690290
rect 11000 689960 573000 690050
rect 11000 689720 170964 689960
rect 171204 689720 171294 689960
rect 171534 689720 171624 689960
rect 171864 689720 171954 689960
rect 172194 689720 172284 689960
rect 172524 689720 172614 689960
rect 172854 689720 217364 689960
rect 217604 689720 217694 689960
rect 217934 689720 218024 689960
rect 218264 689720 218354 689960
rect 218594 689720 218684 689960
rect 218924 689720 219014 689960
rect 219254 689720 219344 689960
rect 219584 689720 219674 689960
rect 219914 689720 220004 689960
rect 220244 689720 220334 689960
rect 220574 689720 220664 689960
rect 220904 689720 220994 689960
rect 221234 689720 221324 689960
rect 221564 689720 221654 689960
rect 221894 689720 221984 689960
rect 222224 689720 227664 689960
rect 227904 689720 227994 689960
rect 228234 689720 228324 689960
rect 228564 689720 228654 689960
rect 228894 689720 228984 689960
rect 229224 689720 229314 689960
rect 229554 689720 229644 689960
rect 229884 689720 229974 689960
rect 230214 689720 230304 689960
rect 230544 689720 230634 689960
rect 230874 689720 230964 689960
rect 231204 689720 231294 689960
rect 231534 689720 231624 689960
rect 231864 689720 231954 689960
rect 232194 689720 232284 689960
rect 232524 689720 573000 689960
rect 11000 689630 573000 689720
rect 11000 689390 170964 689630
rect 171204 689390 171294 689630
rect 171534 689390 171624 689630
rect 171864 689390 171954 689630
rect 172194 689390 172284 689630
rect 172524 689390 172614 689630
rect 172854 689390 217364 689630
rect 217604 689390 217694 689630
rect 217934 689390 218024 689630
rect 218264 689390 218354 689630
rect 218594 689390 218684 689630
rect 218924 689390 219014 689630
rect 219254 689390 219344 689630
rect 219584 689390 219674 689630
rect 219914 689390 220004 689630
rect 220244 689390 220334 689630
rect 220574 689390 220664 689630
rect 220904 689390 220994 689630
rect 221234 689390 221324 689630
rect 221564 689390 221654 689630
rect 221894 689390 221984 689630
rect 222224 689390 227664 689630
rect 227904 689390 227994 689630
rect 228234 689390 228324 689630
rect 228564 689390 228654 689630
rect 228894 689390 228984 689630
rect 229224 689390 229314 689630
rect 229554 689390 229644 689630
rect 229884 689390 229974 689630
rect 230214 689390 230304 689630
rect 230544 689390 230634 689630
rect 230874 689390 230964 689630
rect 231204 689390 231294 689630
rect 231534 689390 231624 689630
rect 231864 689390 231954 689630
rect 232194 689390 232284 689630
rect 232524 689390 573000 689630
rect 11000 689300 573000 689390
rect 11000 689060 170964 689300
rect 171204 689060 171294 689300
rect 171534 689060 171624 689300
rect 171864 689060 171954 689300
rect 172194 689060 172284 689300
rect 172524 689060 172614 689300
rect 172854 689060 217364 689300
rect 217604 689060 217694 689300
rect 217934 689060 218024 689300
rect 218264 689060 218354 689300
rect 218594 689060 218684 689300
rect 218924 689060 219014 689300
rect 219254 689060 219344 689300
rect 219584 689060 219674 689300
rect 219914 689060 220004 689300
rect 220244 689060 220334 689300
rect 220574 689060 220664 689300
rect 220904 689060 220994 689300
rect 221234 689060 221324 689300
rect 221564 689060 221654 689300
rect 221894 689060 221984 689300
rect 222224 689060 227664 689300
rect 227904 689060 227994 689300
rect 228234 689060 228324 689300
rect 228564 689060 228654 689300
rect 228894 689060 228984 689300
rect 229224 689060 229314 689300
rect 229554 689060 229644 689300
rect 229884 689060 229974 689300
rect 230214 689060 230304 689300
rect 230544 689060 230634 689300
rect 230874 689060 230964 689300
rect 231204 689060 231294 689300
rect 231534 689060 231624 689300
rect 231864 689060 231954 689300
rect 232194 689060 232284 689300
rect 232524 689060 573000 689300
rect 11000 688970 573000 689060
rect 11000 688730 170964 688970
rect 171204 688730 171294 688970
rect 171534 688730 171624 688970
rect 171864 688730 171954 688970
rect 172194 688730 172284 688970
rect 172524 688730 172614 688970
rect 172854 688730 217364 688970
rect 217604 688730 217694 688970
rect 217934 688730 218024 688970
rect 218264 688730 218354 688970
rect 218594 688730 218684 688970
rect 218924 688730 219014 688970
rect 219254 688730 219344 688970
rect 219584 688730 219674 688970
rect 219914 688730 220004 688970
rect 220244 688730 220334 688970
rect 220574 688730 220664 688970
rect 220904 688730 220994 688970
rect 221234 688730 221324 688970
rect 221564 688730 221654 688970
rect 221894 688730 221984 688970
rect 222224 688730 227664 688970
rect 227904 688730 227994 688970
rect 228234 688730 228324 688970
rect 228564 688730 228654 688970
rect 228894 688730 228984 688970
rect 229224 688730 229314 688970
rect 229554 688730 229644 688970
rect 229884 688730 229974 688970
rect 230214 688730 230304 688970
rect 230544 688730 230634 688970
rect 230874 688730 230964 688970
rect 231204 688730 231294 688970
rect 231534 688730 231624 688970
rect 231864 688730 231954 688970
rect 232194 688730 232284 688970
rect 232524 688730 573000 688970
rect 11000 688640 573000 688730
rect 11000 688400 170964 688640
rect 171204 688400 171294 688640
rect 171534 688400 171624 688640
rect 171864 688400 171954 688640
rect 172194 688400 172284 688640
rect 172524 688400 172614 688640
rect 172854 688400 217364 688640
rect 217604 688400 217694 688640
rect 217934 688400 218024 688640
rect 218264 688400 218354 688640
rect 218594 688400 218684 688640
rect 218924 688400 219014 688640
rect 219254 688400 219344 688640
rect 219584 688400 219674 688640
rect 219914 688400 220004 688640
rect 220244 688400 220334 688640
rect 220574 688400 220664 688640
rect 220904 688400 220994 688640
rect 221234 688400 221324 688640
rect 221564 688400 221654 688640
rect 221894 688400 221984 688640
rect 222224 688400 227664 688640
rect 227904 688400 227994 688640
rect 228234 688400 228324 688640
rect 228564 688400 228654 688640
rect 228894 688400 228984 688640
rect 229224 688400 229314 688640
rect 229554 688400 229644 688640
rect 229884 688400 229974 688640
rect 230214 688400 230304 688640
rect 230544 688400 230634 688640
rect 230874 688400 230964 688640
rect 231204 688400 231294 688640
rect 231534 688400 231624 688640
rect 231864 688400 231954 688640
rect 232194 688400 232284 688640
rect 232524 688400 573000 688640
rect 11000 688310 573000 688400
rect 11000 688070 170964 688310
rect 171204 688070 171294 688310
rect 171534 688070 171624 688310
rect 171864 688070 171954 688310
rect 172194 688070 172284 688310
rect 172524 688070 172614 688310
rect 172854 688070 217364 688310
rect 217604 688070 217694 688310
rect 217934 688070 218024 688310
rect 218264 688070 218354 688310
rect 218594 688070 218684 688310
rect 218924 688070 219014 688310
rect 219254 688070 219344 688310
rect 219584 688070 219674 688310
rect 219914 688070 220004 688310
rect 220244 688070 220334 688310
rect 220574 688070 220664 688310
rect 220904 688070 220994 688310
rect 221234 688070 221324 688310
rect 221564 688070 221654 688310
rect 221894 688070 221984 688310
rect 222224 688070 227664 688310
rect 227904 688070 227994 688310
rect 228234 688070 228324 688310
rect 228564 688070 228654 688310
rect 228894 688070 228984 688310
rect 229224 688070 229314 688310
rect 229554 688070 229644 688310
rect 229884 688070 229974 688310
rect 230214 688070 230304 688310
rect 230544 688070 230634 688310
rect 230874 688070 230964 688310
rect 231204 688070 231294 688310
rect 231534 688070 231624 688310
rect 231864 688070 231954 688310
rect 232194 688070 232284 688310
rect 232524 688070 573000 688310
rect 11000 688000 573000 688070
rect 11000 664122 16000 688000
rect 568000 670556 573000 688000
rect 576000 670556 581000 696000
rect 82720 668910 85310 669190
rect 82720 668670 82750 668910
rect 82990 668670 83080 668910
rect 83320 668670 83410 668910
rect 83650 668670 83770 668910
rect 84010 668670 84100 668910
rect 84340 668670 84460 668910
rect 84700 668670 84790 668910
rect 85030 668670 85310 668910
rect 82720 668580 85310 668670
rect 82720 668340 82750 668580
rect 82990 668340 83080 668580
rect 83320 668340 83410 668580
rect 83650 668340 83770 668580
rect 84010 668340 84100 668580
rect 84340 668340 84460 668580
rect 84700 668340 84790 668580
rect 85030 668340 85310 668580
rect 82720 668250 85310 668340
rect 82720 668010 82750 668250
rect 82990 668010 83080 668250
rect 83320 668010 83410 668250
rect 83650 668010 83770 668250
rect 84010 668010 84100 668250
rect 84340 668010 84460 668250
rect 84700 668010 84790 668250
rect 85030 668010 85310 668250
rect 82720 667890 85310 668010
rect 82720 667650 82750 667890
rect 82990 667650 83080 667890
rect 83320 667650 83410 667890
rect 83650 667650 83770 667890
rect 84010 667650 84100 667890
rect 84340 667650 84460 667890
rect 84700 667650 84790 667890
rect 85030 667650 85310 667890
rect 82720 667560 85310 667650
rect 82720 667320 82750 667560
rect 82990 667320 83080 667560
rect 83320 667320 83410 667560
rect 83650 667320 83770 667560
rect 84010 667320 84100 667560
rect 84340 667320 84460 667560
rect 84700 667320 84790 667560
rect 85030 667320 85310 667560
rect 82720 667200 85310 667320
rect 82720 666960 82750 667200
rect 82990 666960 83080 667200
rect 83320 666960 83410 667200
rect 83650 666960 83770 667200
rect 84010 666960 84100 667200
rect 84340 666960 84460 667200
rect 84700 666960 84790 667200
rect 85030 666960 85310 667200
rect 82720 666870 85310 666960
rect 82720 666630 82750 666870
rect 82990 666630 83080 666870
rect 83320 666630 83410 666870
rect 83650 666630 83770 666870
rect 84010 666630 84100 666870
rect 84340 666630 84460 666870
rect 84700 666630 84790 666870
rect 85030 666630 85310 666870
rect 82720 666510 85310 666630
rect 82720 666270 82750 666510
rect 82990 666270 83080 666510
rect 83320 666270 83410 666510
rect 83650 666270 83770 666510
rect 84010 666270 84100 666510
rect 84340 666270 84460 666510
rect 84700 666270 84790 666510
rect 85030 666270 85310 666510
rect 82720 666180 85310 666270
rect 82720 665940 82750 666180
rect 82990 665940 83080 666180
rect 83320 665940 83410 666180
rect 83650 665940 83770 666180
rect 84010 665940 84100 666180
rect 84340 665940 84460 666180
rect 84700 665940 84790 666180
rect 85030 665940 85310 666180
rect 82720 665820 85310 665940
rect 82720 665580 82750 665820
rect 82990 665580 83080 665820
rect 83320 665580 83410 665820
rect 83650 665580 83770 665820
rect 84010 665580 84100 665820
rect 84340 665580 84460 665820
rect 84700 665580 84790 665820
rect 85030 665580 85310 665820
rect 82720 665490 85310 665580
rect 82720 665250 82750 665490
rect 82990 665250 83080 665490
rect 83320 665250 83410 665490
rect 83650 665250 83770 665490
rect 84010 665250 84100 665490
rect 84340 665250 84460 665490
rect 84700 665250 84790 665490
rect 85030 665250 85310 665490
rect 82720 665130 85310 665250
rect 82720 664890 82750 665130
rect 82990 664890 83080 665130
rect 83320 664890 83410 665130
rect 83650 664890 83770 665130
rect 84010 664890 84100 665130
rect 84340 664890 84460 665130
rect 84700 664890 84790 665130
rect 85030 664890 85310 665130
rect 82720 664800 85310 664890
rect 82720 664560 82750 664800
rect 82990 664560 83080 664800
rect 83320 664560 83410 664800
rect 83650 664560 83770 664800
rect 84010 664560 84100 664800
rect 84340 664560 84460 664800
rect 84700 664560 84790 664800
rect 85030 664560 85310 664800
rect 82720 664470 85310 664560
rect 82720 664230 82750 664470
rect 82990 664230 83080 664470
rect 83320 664230 83410 664470
rect 83650 664230 83770 664470
rect 84010 664230 84100 664470
rect 84340 664230 84460 664470
rect 84700 664230 84790 664470
rect 85030 664230 85310 664470
rect 82720 664190 85310 664230
rect 11000 659122 78838 664122
rect 11000 639480 16000 659122
rect 82720 657030 85320 657320
rect 82720 656790 82750 657030
rect 82990 656790 83080 657030
rect 83320 656790 83410 657030
rect 83650 656790 83770 657030
rect 84010 656790 84100 657030
rect 84340 656790 84460 657030
rect 84700 656790 84790 657030
rect 85030 656790 85320 657030
rect 82720 656700 85320 656790
rect 82720 656460 82750 656700
rect 82990 656460 83080 656700
rect 83320 656460 83410 656700
rect 83650 656460 83770 656700
rect 84010 656460 84100 656700
rect 84340 656460 84460 656700
rect 84700 656460 84790 656700
rect 85030 656460 85320 656700
rect 82720 656370 85320 656460
rect 82720 656130 82750 656370
rect 82990 656130 83080 656370
rect 83320 656130 83410 656370
rect 83650 656130 83770 656370
rect 84010 656130 84100 656370
rect 84340 656130 84460 656370
rect 84700 656130 84790 656370
rect 85030 656130 85320 656370
rect 82720 656010 85320 656130
rect 82720 655770 82750 656010
rect 82990 655770 83080 656010
rect 83320 655770 83410 656010
rect 83650 655770 83770 656010
rect 84010 655770 84100 656010
rect 84340 655770 84460 656010
rect 84700 655770 84790 656010
rect 85030 655770 85320 656010
rect 82720 655680 85320 655770
rect 82720 655440 82750 655680
rect 82990 655440 83080 655680
rect 83320 655440 83410 655680
rect 83650 655440 83770 655680
rect 84010 655440 84100 655680
rect 84340 655440 84460 655680
rect 84700 655440 84790 655680
rect 85030 655440 85320 655680
rect 82720 655320 85320 655440
rect 82720 655080 82750 655320
rect 82990 655080 83080 655320
rect 83320 655080 83410 655320
rect 83650 655080 83770 655320
rect 84010 655080 84100 655320
rect 84340 655080 84460 655320
rect 84700 655080 84790 655320
rect 85030 655080 85320 655320
rect 82720 654990 85320 655080
rect 82720 654750 82750 654990
rect 82990 654750 83080 654990
rect 83320 654750 83410 654990
rect 83650 654750 83770 654990
rect 84010 654750 84100 654990
rect 84340 654750 84460 654990
rect 84700 654750 84790 654990
rect 85030 654750 85320 654990
rect 82720 654630 85320 654750
rect 82720 654390 82750 654630
rect 82990 654390 83080 654630
rect 83320 654390 83410 654630
rect 83650 654390 83770 654630
rect 84010 654390 84100 654630
rect 84340 654390 84460 654630
rect 84700 654390 84790 654630
rect 85030 654390 85320 654630
rect 82720 654300 85320 654390
rect 82720 654060 82750 654300
rect 82990 654060 83080 654300
rect 83320 654060 83410 654300
rect 83650 654060 83770 654300
rect 84010 654060 84100 654300
rect 84340 654060 84460 654300
rect 84700 654060 84790 654300
rect 85030 654060 85320 654300
rect 82720 653940 85320 654060
rect 82720 653700 82750 653940
rect 82990 653700 83080 653940
rect 83320 653700 83410 653940
rect 83650 653700 83770 653940
rect 84010 653700 84100 653940
rect 84340 653700 84460 653940
rect 84700 653700 84790 653940
rect 85030 653700 85320 653940
rect 82720 653610 85320 653700
rect 82720 653370 82750 653610
rect 82990 653370 83080 653610
rect 83320 653370 83410 653610
rect 83650 653370 83770 653610
rect 84010 653370 84100 653610
rect 84340 653370 84460 653610
rect 84700 653370 84790 653610
rect 85030 653370 85320 653610
rect 82720 653250 85320 653370
rect 82720 653010 82750 653250
rect 82990 653010 83080 653250
rect 83320 653010 83410 653250
rect 83650 653010 83770 653250
rect 84010 653010 84100 653250
rect 84340 653010 84460 653250
rect 84700 653010 84790 653250
rect 85030 653010 85320 653250
rect 82720 652920 85320 653010
rect 82720 652680 82750 652920
rect 82990 652680 83080 652920
rect 83320 652680 83410 652920
rect 83650 652680 83770 652920
rect 84010 652680 84100 652920
rect 84340 652680 84460 652920
rect 84700 652680 84790 652920
rect 85030 652680 85320 652920
rect 82720 652590 85320 652680
rect 82720 652350 82750 652590
rect 82990 652350 83080 652590
rect 83320 652350 83410 652590
rect 83650 652350 83770 652590
rect 84010 652350 84100 652590
rect 84340 652350 84460 652590
rect 84700 652350 84790 652590
rect 85030 652350 85320 652590
rect 82720 652300 85320 652350
rect 11000 634480 110854 639480
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use esd_wide  esd_wide_3
timestamp 1637690973
transform 0 -1 24350 1 0 664950
box 11570 11470 24390 18230
use esd_wide  esd_wide_2
timestamp 1637690973
transform 1 0 870 0 1 679650
box 11570 11470 24390 18230
use big_cap  big_cap_0
timestamp 1636526374
transform 1 0 -27430 0 1 658600
box 60730 -31110 106740 14450
use top  top_0
timestamp 1637733805
transform 1 0 89244 0 1 662150
box -6530 -24030 39650 21850
use esd_half  esd_half_0
timestamp 1637734524
transform 1 0 52890 0 1 679650
box 11570 11470 18780 18230
use esd_half  esd_half_1
timestamp 1637734524
transform -1 0 140498 0 1 679650
box 11570 11470 18780 18230
use esd  esd_0
timestamp 1637690859
transform 1 0 304030 0 1 679650
box 11570 11470 23360 18230
use esd  esd_1
timestamp 1637690859
transform 1 0 398430 0 1 679650
box 11570 11470 23360 18230
use esd  esd_2
timestamp 1637690859
transform 1 0 450430 0 1 679650
box 11570 11470 23360 18230
use esd  esd_3
timestamp 1637690859
transform 1 0 549540 0 1 679650
box 11570 11470 23360 18230
use esd  esd_4
timestamp 1637690859
transform 0 1 559650 -1 0 696716
box 11570 11470 23360 18230
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
