magic
tech sky130A
magscale 1 2
timestamp 1637690973
<< nwell >>
rect 11630 16000 17124 17368
rect 18836 16000 24330 17368
<< pwell >>
rect 11630 12313 17124 13671
rect 18836 12313 24330 13671
<< pmoslvt >>
rect 11826 16220 12026 17220
rect 12084 16220 12284 17220
rect 12342 16220 12542 17220
rect 12600 16220 12800 17220
rect 12858 16220 13058 17220
rect 13116 16220 13316 17220
rect 13374 16220 13574 17220
rect 13632 16220 13832 17220
rect 13890 16220 14090 17220
rect 14148 16220 14348 17220
rect 14406 16220 14606 17220
rect 14664 16220 14864 17220
rect 14922 16220 15122 17220
rect 15180 16220 15380 17220
rect 15438 16220 15638 17220
rect 15696 16220 15896 17220
rect 15954 16220 16154 17220
rect 16212 16220 16412 17220
rect 16470 16220 16670 17220
rect 16728 16220 16928 17220
rect 19032 16220 19232 17220
rect 19290 16220 19490 17220
rect 19548 16220 19748 17220
rect 19806 16220 20006 17220
rect 20064 16220 20264 17220
rect 20322 16220 20522 17220
rect 20580 16220 20780 17220
rect 20838 16220 21038 17220
rect 21096 16220 21296 17220
rect 21354 16220 21554 17220
rect 21612 16220 21812 17220
rect 21870 16220 22070 17220
rect 22128 16220 22328 17220
rect 22386 16220 22586 17220
rect 22644 16220 22844 17220
rect 22902 16220 23102 17220
rect 23160 16220 23360 17220
rect 23418 16220 23618 17220
rect 23676 16220 23876 17220
rect 23934 16220 24134 17220
<< nmoslvt >>
rect 11826 12461 12026 13461
rect 12084 12461 12284 13461
rect 12342 12461 12542 13461
rect 12600 12461 12800 13461
rect 12858 12461 13058 13461
rect 13116 12461 13316 13461
rect 13374 12461 13574 13461
rect 13632 12461 13832 13461
rect 13890 12461 14090 13461
rect 14148 12461 14348 13461
rect 14406 12461 14606 13461
rect 14664 12461 14864 13461
rect 14922 12461 15122 13461
rect 15180 12461 15380 13461
rect 15438 12461 15638 13461
rect 15696 12461 15896 13461
rect 15954 12461 16154 13461
rect 16212 12461 16412 13461
rect 16470 12461 16670 13461
rect 16728 12461 16928 13461
rect 19032 12461 19232 13461
rect 19290 12461 19490 13461
rect 19548 12461 19748 13461
rect 19806 12461 20006 13461
rect 20064 12461 20264 13461
rect 20322 12461 20522 13461
rect 20580 12461 20780 13461
rect 20838 12461 21038 13461
rect 21096 12461 21296 13461
rect 21354 12461 21554 13461
rect 21612 12461 21812 13461
rect 21870 12461 22070 13461
rect 22128 12461 22328 13461
rect 22386 12461 22586 13461
rect 22644 12461 22844 13461
rect 22902 12461 23102 13461
rect 23160 12461 23360 13461
rect 23418 12461 23618 13461
rect 23676 12461 23876 13461
rect 23934 12461 24134 13461
<< ndiff >>
rect 11768 13449 11826 13461
rect 11768 12473 11780 13449
rect 11814 12473 11826 13449
rect 11768 12461 11826 12473
rect 12026 13449 12084 13461
rect 12026 12473 12038 13449
rect 12072 12473 12084 13449
rect 12026 12461 12084 12473
rect 12284 13449 12342 13461
rect 12284 12473 12296 13449
rect 12330 12473 12342 13449
rect 12284 12461 12342 12473
rect 12542 13449 12600 13461
rect 12542 12473 12554 13449
rect 12588 12473 12600 13449
rect 12542 12461 12600 12473
rect 12800 13449 12858 13461
rect 12800 12473 12812 13449
rect 12846 12473 12858 13449
rect 12800 12461 12858 12473
rect 13058 13449 13116 13461
rect 13058 12473 13070 13449
rect 13104 12473 13116 13449
rect 13058 12461 13116 12473
rect 13316 13449 13374 13461
rect 13316 12473 13328 13449
rect 13362 12473 13374 13449
rect 13316 12461 13374 12473
rect 13574 13449 13632 13461
rect 13574 12473 13586 13449
rect 13620 12473 13632 13449
rect 13574 12461 13632 12473
rect 13832 13449 13890 13461
rect 13832 12473 13844 13449
rect 13878 12473 13890 13449
rect 13832 12461 13890 12473
rect 14090 13449 14148 13461
rect 14090 12473 14102 13449
rect 14136 12473 14148 13449
rect 14090 12461 14148 12473
rect 14348 13449 14406 13461
rect 14348 12473 14360 13449
rect 14394 12473 14406 13449
rect 14348 12461 14406 12473
rect 14606 13449 14664 13461
rect 14606 12473 14618 13449
rect 14652 12473 14664 13449
rect 14606 12461 14664 12473
rect 14864 13449 14922 13461
rect 14864 12473 14876 13449
rect 14910 12473 14922 13449
rect 14864 12461 14922 12473
rect 15122 13449 15180 13461
rect 15122 12473 15134 13449
rect 15168 12473 15180 13449
rect 15122 12461 15180 12473
rect 15380 13449 15438 13461
rect 15380 12473 15392 13449
rect 15426 12473 15438 13449
rect 15380 12461 15438 12473
rect 15638 13449 15696 13461
rect 15638 12473 15650 13449
rect 15684 12473 15696 13449
rect 15638 12461 15696 12473
rect 15896 13449 15954 13461
rect 15896 12473 15908 13449
rect 15942 12473 15954 13449
rect 15896 12461 15954 12473
rect 16154 13449 16212 13461
rect 16154 12473 16166 13449
rect 16200 12473 16212 13449
rect 16154 12461 16212 12473
rect 16412 13449 16470 13461
rect 16412 12473 16424 13449
rect 16458 12473 16470 13449
rect 16412 12461 16470 12473
rect 16670 13449 16728 13461
rect 16670 12473 16682 13449
rect 16716 12473 16728 13449
rect 16670 12461 16728 12473
rect 16928 13449 16986 13461
rect 16928 12473 16940 13449
rect 16974 12473 16986 13449
rect 16928 12461 16986 12473
rect 18974 13449 19032 13461
rect 18974 12473 18986 13449
rect 19020 12473 19032 13449
rect 18974 12461 19032 12473
rect 19232 13449 19290 13461
rect 19232 12473 19244 13449
rect 19278 12473 19290 13449
rect 19232 12461 19290 12473
rect 19490 13449 19548 13461
rect 19490 12473 19502 13449
rect 19536 12473 19548 13449
rect 19490 12461 19548 12473
rect 19748 13449 19806 13461
rect 19748 12473 19760 13449
rect 19794 12473 19806 13449
rect 19748 12461 19806 12473
rect 20006 13449 20064 13461
rect 20006 12473 20018 13449
rect 20052 12473 20064 13449
rect 20006 12461 20064 12473
rect 20264 13449 20322 13461
rect 20264 12473 20276 13449
rect 20310 12473 20322 13449
rect 20264 12461 20322 12473
rect 20522 13449 20580 13461
rect 20522 12473 20534 13449
rect 20568 12473 20580 13449
rect 20522 12461 20580 12473
rect 20780 13449 20838 13461
rect 20780 12473 20792 13449
rect 20826 12473 20838 13449
rect 20780 12461 20838 12473
rect 21038 13449 21096 13461
rect 21038 12473 21050 13449
rect 21084 12473 21096 13449
rect 21038 12461 21096 12473
rect 21296 13449 21354 13461
rect 21296 12473 21308 13449
rect 21342 12473 21354 13449
rect 21296 12461 21354 12473
rect 21554 13449 21612 13461
rect 21554 12473 21566 13449
rect 21600 12473 21612 13449
rect 21554 12461 21612 12473
rect 21812 13449 21870 13461
rect 21812 12473 21824 13449
rect 21858 12473 21870 13449
rect 21812 12461 21870 12473
rect 22070 13449 22128 13461
rect 22070 12473 22082 13449
rect 22116 12473 22128 13449
rect 22070 12461 22128 12473
rect 22328 13449 22386 13461
rect 22328 12473 22340 13449
rect 22374 12473 22386 13449
rect 22328 12461 22386 12473
rect 22586 13449 22644 13461
rect 22586 12473 22598 13449
rect 22632 12473 22644 13449
rect 22586 12461 22644 12473
rect 22844 13449 22902 13461
rect 22844 12473 22856 13449
rect 22890 12473 22902 13449
rect 22844 12461 22902 12473
rect 23102 13449 23160 13461
rect 23102 12473 23114 13449
rect 23148 12473 23160 13449
rect 23102 12461 23160 12473
rect 23360 13449 23418 13461
rect 23360 12473 23372 13449
rect 23406 12473 23418 13449
rect 23360 12461 23418 12473
rect 23618 13449 23676 13461
rect 23618 12473 23630 13449
rect 23664 12473 23676 13449
rect 23618 12461 23676 12473
rect 23876 13449 23934 13461
rect 23876 12473 23888 13449
rect 23922 12473 23934 13449
rect 23876 12461 23934 12473
rect 24134 13449 24192 13461
rect 24134 12473 24146 13449
rect 24180 12473 24192 13449
rect 24134 12461 24192 12473
<< pdiff >>
rect 11768 17208 11826 17220
rect 11768 16232 11780 17208
rect 11814 16232 11826 17208
rect 11768 16220 11826 16232
rect 12026 17208 12084 17220
rect 12026 16232 12038 17208
rect 12072 16232 12084 17208
rect 12026 16220 12084 16232
rect 12284 17208 12342 17220
rect 12284 16232 12296 17208
rect 12330 16232 12342 17208
rect 12284 16220 12342 16232
rect 12542 17208 12600 17220
rect 12542 16232 12554 17208
rect 12588 16232 12600 17208
rect 12542 16220 12600 16232
rect 12800 17208 12858 17220
rect 12800 16232 12812 17208
rect 12846 16232 12858 17208
rect 12800 16220 12858 16232
rect 13058 17208 13116 17220
rect 13058 16232 13070 17208
rect 13104 16232 13116 17208
rect 13058 16220 13116 16232
rect 13316 17208 13374 17220
rect 13316 16232 13328 17208
rect 13362 16232 13374 17208
rect 13316 16220 13374 16232
rect 13574 17208 13632 17220
rect 13574 16232 13586 17208
rect 13620 16232 13632 17208
rect 13574 16220 13632 16232
rect 13832 17208 13890 17220
rect 13832 16232 13844 17208
rect 13878 16232 13890 17208
rect 13832 16220 13890 16232
rect 14090 17208 14148 17220
rect 14090 16232 14102 17208
rect 14136 16232 14148 17208
rect 14090 16220 14148 16232
rect 14348 17208 14406 17220
rect 14348 16232 14360 17208
rect 14394 16232 14406 17208
rect 14348 16220 14406 16232
rect 14606 17208 14664 17220
rect 14606 16232 14618 17208
rect 14652 16232 14664 17208
rect 14606 16220 14664 16232
rect 14864 17208 14922 17220
rect 14864 16232 14876 17208
rect 14910 16232 14922 17208
rect 14864 16220 14922 16232
rect 15122 17208 15180 17220
rect 15122 16232 15134 17208
rect 15168 16232 15180 17208
rect 15122 16220 15180 16232
rect 15380 17208 15438 17220
rect 15380 16232 15392 17208
rect 15426 16232 15438 17208
rect 15380 16220 15438 16232
rect 15638 17208 15696 17220
rect 15638 16232 15650 17208
rect 15684 16232 15696 17208
rect 15638 16220 15696 16232
rect 15896 17208 15954 17220
rect 15896 16232 15908 17208
rect 15942 16232 15954 17208
rect 15896 16220 15954 16232
rect 16154 17208 16212 17220
rect 16154 16232 16166 17208
rect 16200 16232 16212 17208
rect 16154 16220 16212 16232
rect 16412 17208 16470 17220
rect 16412 16232 16424 17208
rect 16458 16232 16470 17208
rect 16412 16220 16470 16232
rect 16670 17208 16728 17220
rect 16670 16232 16682 17208
rect 16716 16232 16728 17208
rect 16670 16220 16728 16232
rect 16928 17208 16986 17220
rect 16928 16232 16940 17208
rect 16974 16232 16986 17208
rect 16928 16220 16986 16232
rect 18974 17208 19032 17220
rect 18974 16232 18986 17208
rect 19020 16232 19032 17208
rect 18974 16220 19032 16232
rect 19232 17208 19290 17220
rect 19232 16232 19244 17208
rect 19278 16232 19290 17208
rect 19232 16220 19290 16232
rect 19490 17208 19548 17220
rect 19490 16232 19502 17208
rect 19536 16232 19548 17208
rect 19490 16220 19548 16232
rect 19748 17208 19806 17220
rect 19748 16232 19760 17208
rect 19794 16232 19806 17208
rect 19748 16220 19806 16232
rect 20006 17208 20064 17220
rect 20006 16232 20018 17208
rect 20052 16232 20064 17208
rect 20006 16220 20064 16232
rect 20264 17208 20322 17220
rect 20264 16232 20276 17208
rect 20310 16232 20322 17208
rect 20264 16220 20322 16232
rect 20522 17208 20580 17220
rect 20522 16232 20534 17208
rect 20568 16232 20580 17208
rect 20522 16220 20580 16232
rect 20780 17208 20838 17220
rect 20780 16232 20792 17208
rect 20826 16232 20838 17208
rect 20780 16220 20838 16232
rect 21038 17208 21096 17220
rect 21038 16232 21050 17208
rect 21084 16232 21096 17208
rect 21038 16220 21096 16232
rect 21296 17208 21354 17220
rect 21296 16232 21308 17208
rect 21342 16232 21354 17208
rect 21296 16220 21354 16232
rect 21554 17208 21612 17220
rect 21554 16232 21566 17208
rect 21600 16232 21612 17208
rect 21554 16220 21612 16232
rect 21812 17208 21870 17220
rect 21812 16232 21824 17208
rect 21858 16232 21870 17208
rect 21812 16220 21870 16232
rect 22070 17208 22128 17220
rect 22070 16232 22082 17208
rect 22116 16232 22128 17208
rect 22070 16220 22128 16232
rect 22328 17208 22386 17220
rect 22328 16232 22340 17208
rect 22374 16232 22386 17208
rect 22328 16220 22386 16232
rect 22586 17208 22644 17220
rect 22586 16232 22598 17208
rect 22632 16232 22644 17208
rect 22586 16220 22644 16232
rect 22844 17208 22902 17220
rect 22844 16232 22856 17208
rect 22890 16232 22902 17208
rect 22844 16220 22902 16232
rect 23102 17208 23160 17220
rect 23102 16232 23114 17208
rect 23148 16232 23160 17208
rect 23102 16220 23160 16232
rect 23360 17208 23418 17220
rect 23360 16232 23372 17208
rect 23406 16232 23418 17208
rect 23360 16220 23418 16232
rect 23618 17208 23676 17220
rect 23618 16232 23630 17208
rect 23664 16232 23676 17208
rect 23618 16220 23676 16232
rect 23876 17208 23934 17220
rect 23876 16232 23888 17208
rect 23922 16232 23934 17208
rect 23876 16220 23934 16232
rect 24134 17208 24192 17220
rect 24134 16232 24146 17208
rect 24180 16232 24192 17208
rect 24134 16220 24192 16232
<< ndiffc >>
rect 11780 12473 11814 13449
rect 12038 12473 12072 13449
rect 12296 12473 12330 13449
rect 12554 12473 12588 13449
rect 12812 12473 12846 13449
rect 13070 12473 13104 13449
rect 13328 12473 13362 13449
rect 13586 12473 13620 13449
rect 13844 12473 13878 13449
rect 14102 12473 14136 13449
rect 14360 12473 14394 13449
rect 14618 12473 14652 13449
rect 14876 12473 14910 13449
rect 15134 12473 15168 13449
rect 15392 12473 15426 13449
rect 15650 12473 15684 13449
rect 15908 12473 15942 13449
rect 16166 12473 16200 13449
rect 16424 12473 16458 13449
rect 16682 12473 16716 13449
rect 16940 12473 16974 13449
rect 18986 12473 19020 13449
rect 19244 12473 19278 13449
rect 19502 12473 19536 13449
rect 19760 12473 19794 13449
rect 20018 12473 20052 13449
rect 20276 12473 20310 13449
rect 20534 12473 20568 13449
rect 20792 12473 20826 13449
rect 21050 12473 21084 13449
rect 21308 12473 21342 13449
rect 21566 12473 21600 13449
rect 21824 12473 21858 13449
rect 22082 12473 22116 13449
rect 22340 12473 22374 13449
rect 22598 12473 22632 13449
rect 22856 12473 22890 13449
rect 23114 12473 23148 13449
rect 23372 12473 23406 13449
rect 23630 12473 23664 13449
rect 23888 12473 23922 13449
rect 24146 12473 24180 13449
<< pdiffc >>
rect 11780 16232 11814 17208
rect 12038 16232 12072 17208
rect 12296 16232 12330 17208
rect 12554 16232 12588 17208
rect 12812 16232 12846 17208
rect 13070 16232 13104 17208
rect 13328 16232 13362 17208
rect 13586 16232 13620 17208
rect 13844 16232 13878 17208
rect 14102 16232 14136 17208
rect 14360 16232 14394 17208
rect 14618 16232 14652 17208
rect 14876 16232 14910 17208
rect 15134 16232 15168 17208
rect 15392 16232 15426 17208
rect 15650 16232 15684 17208
rect 15908 16232 15942 17208
rect 16166 16232 16200 17208
rect 16424 16232 16458 17208
rect 16682 16232 16716 17208
rect 16940 16232 16974 17208
rect 18986 16232 19020 17208
rect 19244 16232 19278 17208
rect 19502 16232 19536 17208
rect 19760 16232 19794 17208
rect 20018 16232 20052 17208
rect 20276 16232 20310 17208
rect 20534 16232 20568 17208
rect 20792 16232 20826 17208
rect 21050 16232 21084 17208
rect 21308 16232 21342 17208
rect 21566 16232 21600 17208
rect 21824 16232 21858 17208
rect 22082 16232 22116 17208
rect 22340 16232 22374 17208
rect 22598 16232 22632 17208
rect 22856 16232 22890 17208
rect 23114 16232 23148 17208
rect 23372 16232 23406 17208
rect 23630 16232 23664 17208
rect 23888 16232 23922 17208
rect 24146 16232 24180 17208
<< psubdiff >>
rect 11666 13601 11762 13635
rect 16992 13601 17088 13635
rect 11666 13539 11700 13601
rect 17054 13539 17088 13601
rect 11666 12383 11700 12445
rect 17054 12383 17088 12445
rect 11666 12349 11762 12383
rect 16992 12349 17088 12383
rect 18872 13601 18968 13635
rect 24198 13601 24294 13635
rect 18872 13539 18906 13601
rect 24260 13539 24294 13601
rect 18872 12383 18906 12445
rect 24260 12383 24294 12445
rect 18872 12349 18968 12383
rect 24198 12349 24294 12383
<< nsubdiff >>
rect 11666 17298 11762 17332
rect 16992 17298 17088 17332
rect 11666 17235 11700 17298
rect 17054 17235 17088 17298
rect 11666 16070 11700 16133
rect 17054 16070 17088 16133
rect 11666 16036 11762 16070
rect 16992 16036 17088 16070
rect 18872 17298 18968 17332
rect 24198 17298 24294 17332
rect 18872 17235 18906 17298
rect 24260 17235 24294 17298
rect 18872 16070 18906 16133
rect 24260 16070 24294 16133
rect 18872 16036 18968 16070
rect 24198 16036 24294 16070
<< psubdiffcont >>
rect 11762 13601 16992 13635
rect 11666 12445 11700 13539
rect 17054 12445 17088 13539
rect 11762 12349 16992 12383
rect 18968 13601 24198 13635
rect 18872 12445 18906 13539
rect 24260 12445 24294 13539
rect 18968 12349 24198 12383
<< nsubdiffcont >>
rect 11762 17298 16992 17332
rect 11666 16133 11700 17235
rect 17054 16133 17088 17235
rect 11762 16036 16992 16070
rect 18968 17298 24198 17332
rect 18872 16133 18906 17235
rect 24260 16133 24294 17235
rect 18968 16036 24198 16070
<< poly >>
rect 11826 17220 12026 17246
rect 12084 17220 12284 17246
rect 12342 17220 12542 17246
rect 12600 17220 12800 17246
rect 12858 17220 13058 17246
rect 13116 17220 13316 17246
rect 13374 17220 13574 17246
rect 13632 17220 13832 17246
rect 13890 17220 14090 17246
rect 14148 17220 14348 17246
rect 14406 17220 14606 17246
rect 14664 17220 14864 17246
rect 14922 17220 15122 17246
rect 15180 17220 15380 17246
rect 15438 17220 15638 17246
rect 15696 17220 15896 17246
rect 15954 17220 16154 17246
rect 16212 17220 16412 17246
rect 16470 17220 16670 17246
rect 16728 17220 16928 17246
rect 11826 16173 12026 16220
rect 11826 16139 11842 16173
rect 12010 16139 12026 16173
rect 11826 16123 12026 16139
rect 12084 16173 12284 16220
rect 12084 16139 12100 16173
rect 12268 16139 12284 16173
rect 12084 16123 12284 16139
rect 12342 16173 12542 16220
rect 12342 16139 12358 16173
rect 12526 16139 12542 16173
rect 12342 16123 12542 16139
rect 12600 16173 12800 16220
rect 12600 16139 12616 16173
rect 12784 16139 12800 16173
rect 12600 16123 12800 16139
rect 12858 16173 13058 16220
rect 12858 16139 12874 16173
rect 13042 16139 13058 16173
rect 12858 16123 13058 16139
rect 13116 16173 13316 16220
rect 13116 16139 13132 16173
rect 13300 16139 13316 16173
rect 13116 16123 13316 16139
rect 13374 16173 13574 16220
rect 13374 16139 13390 16173
rect 13558 16139 13574 16173
rect 13374 16123 13574 16139
rect 13632 16173 13832 16220
rect 13632 16139 13648 16173
rect 13816 16139 13832 16173
rect 13632 16123 13832 16139
rect 13890 16173 14090 16220
rect 13890 16139 13906 16173
rect 14074 16139 14090 16173
rect 13890 16123 14090 16139
rect 14148 16173 14348 16220
rect 14148 16139 14164 16173
rect 14332 16139 14348 16173
rect 14148 16123 14348 16139
rect 14406 16173 14606 16220
rect 14406 16139 14422 16173
rect 14590 16139 14606 16173
rect 14406 16123 14606 16139
rect 14664 16173 14864 16220
rect 14664 16139 14680 16173
rect 14848 16139 14864 16173
rect 14664 16123 14864 16139
rect 14922 16173 15122 16220
rect 14922 16139 14938 16173
rect 15106 16139 15122 16173
rect 14922 16123 15122 16139
rect 15180 16173 15380 16220
rect 15180 16139 15196 16173
rect 15364 16139 15380 16173
rect 15180 16123 15380 16139
rect 15438 16173 15638 16220
rect 15438 16139 15454 16173
rect 15622 16139 15638 16173
rect 15438 16123 15638 16139
rect 15696 16173 15896 16220
rect 15696 16139 15712 16173
rect 15880 16139 15896 16173
rect 15696 16123 15896 16139
rect 15954 16173 16154 16220
rect 15954 16139 15970 16173
rect 16138 16139 16154 16173
rect 15954 16123 16154 16139
rect 16212 16173 16412 16220
rect 16212 16139 16228 16173
rect 16396 16139 16412 16173
rect 16212 16123 16412 16139
rect 16470 16173 16670 16220
rect 16470 16139 16486 16173
rect 16654 16139 16670 16173
rect 16470 16123 16670 16139
rect 16728 16173 16928 16220
rect 16728 16139 16744 16173
rect 16912 16139 16928 16173
rect 16728 16123 16928 16139
rect 19032 17220 19232 17246
rect 19290 17220 19490 17246
rect 19548 17220 19748 17246
rect 19806 17220 20006 17246
rect 20064 17220 20264 17246
rect 20322 17220 20522 17246
rect 20580 17220 20780 17246
rect 20838 17220 21038 17246
rect 21096 17220 21296 17246
rect 21354 17220 21554 17246
rect 21612 17220 21812 17246
rect 21870 17220 22070 17246
rect 22128 17220 22328 17246
rect 22386 17220 22586 17246
rect 22644 17220 22844 17246
rect 22902 17220 23102 17246
rect 23160 17220 23360 17246
rect 23418 17220 23618 17246
rect 23676 17220 23876 17246
rect 23934 17220 24134 17246
rect 19032 16173 19232 16220
rect 19032 16139 19048 16173
rect 19216 16139 19232 16173
rect 19032 16123 19232 16139
rect 19290 16173 19490 16220
rect 19290 16139 19306 16173
rect 19474 16139 19490 16173
rect 19290 16123 19490 16139
rect 19548 16173 19748 16220
rect 19548 16139 19564 16173
rect 19732 16139 19748 16173
rect 19548 16123 19748 16139
rect 19806 16173 20006 16220
rect 19806 16139 19822 16173
rect 19990 16139 20006 16173
rect 19806 16123 20006 16139
rect 20064 16173 20264 16220
rect 20064 16139 20080 16173
rect 20248 16139 20264 16173
rect 20064 16123 20264 16139
rect 20322 16173 20522 16220
rect 20322 16139 20338 16173
rect 20506 16139 20522 16173
rect 20322 16123 20522 16139
rect 20580 16173 20780 16220
rect 20580 16139 20596 16173
rect 20764 16139 20780 16173
rect 20580 16123 20780 16139
rect 20838 16173 21038 16220
rect 20838 16139 20854 16173
rect 21022 16139 21038 16173
rect 20838 16123 21038 16139
rect 21096 16173 21296 16220
rect 21096 16139 21112 16173
rect 21280 16139 21296 16173
rect 21096 16123 21296 16139
rect 21354 16173 21554 16220
rect 21354 16139 21370 16173
rect 21538 16139 21554 16173
rect 21354 16123 21554 16139
rect 21612 16173 21812 16220
rect 21612 16139 21628 16173
rect 21796 16139 21812 16173
rect 21612 16123 21812 16139
rect 21870 16173 22070 16220
rect 21870 16139 21886 16173
rect 22054 16139 22070 16173
rect 21870 16123 22070 16139
rect 22128 16173 22328 16220
rect 22128 16139 22144 16173
rect 22312 16139 22328 16173
rect 22128 16123 22328 16139
rect 22386 16173 22586 16220
rect 22386 16139 22402 16173
rect 22570 16139 22586 16173
rect 22386 16123 22586 16139
rect 22644 16173 22844 16220
rect 22644 16139 22660 16173
rect 22828 16139 22844 16173
rect 22644 16123 22844 16139
rect 22902 16173 23102 16220
rect 22902 16139 22918 16173
rect 23086 16139 23102 16173
rect 22902 16123 23102 16139
rect 23160 16173 23360 16220
rect 23160 16139 23176 16173
rect 23344 16139 23360 16173
rect 23160 16123 23360 16139
rect 23418 16173 23618 16220
rect 23418 16139 23434 16173
rect 23602 16139 23618 16173
rect 23418 16123 23618 16139
rect 23676 16173 23876 16220
rect 23676 16139 23692 16173
rect 23860 16139 23876 16173
rect 23676 16123 23876 16139
rect 23934 16173 24134 16220
rect 23934 16139 23950 16173
rect 24118 16139 24134 16173
rect 23934 16123 24134 16139
rect 11826 13533 12026 13549
rect 11826 13499 11842 13533
rect 12010 13499 12026 13533
rect 11826 13461 12026 13499
rect 12084 13533 12284 13549
rect 12084 13499 12100 13533
rect 12268 13499 12284 13533
rect 12084 13461 12284 13499
rect 12342 13533 12542 13549
rect 12342 13499 12358 13533
rect 12526 13499 12542 13533
rect 12342 13461 12542 13499
rect 12600 13533 12800 13549
rect 12600 13499 12616 13533
rect 12784 13499 12800 13533
rect 12600 13461 12800 13499
rect 12858 13533 13058 13549
rect 12858 13499 12874 13533
rect 13042 13499 13058 13533
rect 12858 13461 13058 13499
rect 13116 13533 13316 13549
rect 13116 13499 13132 13533
rect 13300 13499 13316 13533
rect 13116 13461 13316 13499
rect 13374 13533 13574 13549
rect 13374 13499 13390 13533
rect 13558 13499 13574 13533
rect 13374 13461 13574 13499
rect 13632 13533 13832 13549
rect 13632 13499 13648 13533
rect 13816 13499 13832 13533
rect 13632 13461 13832 13499
rect 13890 13533 14090 13549
rect 13890 13499 13906 13533
rect 14074 13499 14090 13533
rect 13890 13461 14090 13499
rect 14148 13533 14348 13549
rect 14148 13499 14164 13533
rect 14332 13499 14348 13533
rect 14148 13461 14348 13499
rect 14406 13533 14606 13549
rect 14406 13499 14422 13533
rect 14590 13499 14606 13533
rect 14406 13461 14606 13499
rect 14664 13533 14864 13549
rect 14664 13499 14680 13533
rect 14848 13499 14864 13533
rect 14664 13461 14864 13499
rect 14922 13533 15122 13549
rect 14922 13499 14938 13533
rect 15106 13499 15122 13533
rect 14922 13461 15122 13499
rect 15180 13533 15380 13549
rect 15180 13499 15196 13533
rect 15364 13499 15380 13533
rect 15180 13461 15380 13499
rect 15438 13533 15638 13549
rect 15438 13499 15454 13533
rect 15622 13499 15638 13533
rect 15438 13461 15638 13499
rect 15696 13533 15896 13549
rect 15696 13499 15712 13533
rect 15880 13499 15896 13533
rect 15696 13461 15896 13499
rect 15954 13533 16154 13549
rect 15954 13499 15970 13533
rect 16138 13499 16154 13533
rect 15954 13461 16154 13499
rect 16212 13533 16412 13549
rect 16212 13499 16228 13533
rect 16396 13499 16412 13533
rect 16212 13461 16412 13499
rect 16470 13533 16670 13549
rect 16470 13499 16486 13533
rect 16654 13499 16670 13533
rect 16470 13461 16670 13499
rect 16728 13533 16928 13549
rect 16728 13499 16744 13533
rect 16912 13499 16928 13533
rect 16728 13461 16928 13499
rect 11826 12435 12026 12461
rect 12084 12435 12284 12461
rect 12342 12435 12542 12461
rect 12600 12435 12800 12461
rect 12858 12435 13058 12461
rect 13116 12435 13316 12461
rect 13374 12435 13574 12461
rect 13632 12435 13832 12461
rect 13890 12435 14090 12461
rect 14148 12435 14348 12461
rect 14406 12435 14606 12461
rect 14664 12435 14864 12461
rect 14922 12435 15122 12461
rect 15180 12435 15380 12461
rect 15438 12435 15638 12461
rect 15696 12435 15896 12461
rect 15954 12435 16154 12461
rect 16212 12435 16412 12461
rect 16470 12435 16670 12461
rect 16728 12435 16928 12461
rect 19032 13533 19232 13549
rect 19032 13499 19048 13533
rect 19216 13499 19232 13533
rect 19032 13461 19232 13499
rect 19290 13533 19490 13549
rect 19290 13499 19306 13533
rect 19474 13499 19490 13533
rect 19290 13461 19490 13499
rect 19548 13533 19748 13549
rect 19548 13499 19564 13533
rect 19732 13499 19748 13533
rect 19548 13461 19748 13499
rect 19806 13533 20006 13549
rect 19806 13499 19822 13533
rect 19990 13499 20006 13533
rect 19806 13461 20006 13499
rect 20064 13533 20264 13549
rect 20064 13499 20080 13533
rect 20248 13499 20264 13533
rect 20064 13461 20264 13499
rect 20322 13533 20522 13549
rect 20322 13499 20338 13533
rect 20506 13499 20522 13533
rect 20322 13461 20522 13499
rect 20580 13533 20780 13549
rect 20580 13499 20596 13533
rect 20764 13499 20780 13533
rect 20580 13461 20780 13499
rect 20838 13533 21038 13549
rect 20838 13499 20854 13533
rect 21022 13499 21038 13533
rect 20838 13461 21038 13499
rect 21096 13533 21296 13549
rect 21096 13499 21112 13533
rect 21280 13499 21296 13533
rect 21096 13461 21296 13499
rect 21354 13533 21554 13549
rect 21354 13499 21370 13533
rect 21538 13499 21554 13533
rect 21354 13461 21554 13499
rect 21612 13533 21812 13549
rect 21612 13499 21628 13533
rect 21796 13499 21812 13533
rect 21612 13461 21812 13499
rect 21870 13533 22070 13549
rect 21870 13499 21886 13533
rect 22054 13499 22070 13533
rect 21870 13461 22070 13499
rect 22128 13533 22328 13549
rect 22128 13499 22144 13533
rect 22312 13499 22328 13533
rect 22128 13461 22328 13499
rect 22386 13533 22586 13549
rect 22386 13499 22402 13533
rect 22570 13499 22586 13533
rect 22386 13461 22586 13499
rect 22644 13533 22844 13549
rect 22644 13499 22660 13533
rect 22828 13499 22844 13533
rect 22644 13461 22844 13499
rect 22902 13533 23102 13549
rect 22902 13499 22918 13533
rect 23086 13499 23102 13533
rect 22902 13461 23102 13499
rect 23160 13533 23360 13549
rect 23160 13499 23176 13533
rect 23344 13499 23360 13533
rect 23160 13461 23360 13499
rect 23418 13533 23618 13549
rect 23418 13499 23434 13533
rect 23602 13499 23618 13533
rect 23418 13461 23618 13499
rect 23676 13533 23876 13549
rect 23676 13499 23692 13533
rect 23860 13499 23876 13533
rect 23676 13461 23876 13499
rect 23934 13533 24134 13549
rect 23934 13499 23950 13533
rect 24118 13499 24134 13533
rect 23934 13461 24134 13499
rect 19032 12435 19232 12461
rect 19290 12435 19490 12461
rect 19548 12435 19748 12461
rect 19806 12435 20006 12461
rect 20064 12435 20264 12461
rect 20322 12435 20522 12461
rect 20580 12435 20780 12461
rect 20838 12435 21038 12461
rect 21096 12435 21296 12461
rect 21354 12435 21554 12461
rect 21612 12435 21812 12461
rect 21870 12435 22070 12461
rect 22128 12435 22328 12461
rect 22386 12435 22586 12461
rect 22644 12435 22844 12461
rect 22902 12435 23102 12461
rect 23160 12435 23360 12461
rect 23418 12435 23618 12461
rect 23676 12435 23876 12461
rect 23934 12435 24134 12461
<< polycont >>
rect 11842 16139 12010 16173
rect 12100 16139 12268 16173
rect 12358 16139 12526 16173
rect 12616 16139 12784 16173
rect 12874 16139 13042 16173
rect 13132 16139 13300 16173
rect 13390 16139 13558 16173
rect 13648 16139 13816 16173
rect 13906 16139 14074 16173
rect 14164 16139 14332 16173
rect 14422 16139 14590 16173
rect 14680 16139 14848 16173
rect 14938 16139 15106 16173
rect 15196 16139 15364 16173
rect 15454 16139 15622 16173
rect 15712 16139 15880 16173
rect 15970 16139 16138 16173
rect 16228 16139 16396 16173
rect 16486 16139 16654 16173
rect 16744 16139 16912 16173
rect 19048 16139 19216 16173
rect 19306 16139 19474 16173
rect 19564 16139 19732 16173
rect 19822 16139 19990 16173
rect 20080 16139 20248 16173
rect 20338 16139 20506 16173
rect 20596 16139 20764 16173
rect 20854 16139 21022 16173
rect 21112 16139 21280 16173
rect 21370 16139 21538 16173
rect 21628 16139 21796 16173
rect 21886 16139 22054 16173
rect 22144 16139 22312 16173
rect 22402 16139 22570 16173
rect 22660 16139 22828 16173
rect 22918 16139 23086 16173
rect 23176 16139 23344 16173
rect 23434 16139 23602 16173
rect 23692 16139 23860 16173
rect 23950 16139 24118 16173
rect 11842 13499 12010 13533
rect 12100 13499 12268 13533
rect 12358 13499 12526 13533
rect 12616 13499 12784 13533
rect 12874 13499 13042 13533
rect 13132 13499 13300 13533
rect 13390 13499 13558 13533
rect 13648 13499 13816 13533
rect 13906 13499 14074 13533
rect 14164 13499 14332 13533
rect 14422 13499 14590 13533
rect 14680 13499 14848 13533
rect 14938 13499 15106 13533
rect 15196 13499 15364 13533
rect 15454 13499 15622 13533
rect 15712 13499 15880 13533
rect 15970 13499 16138 13533
rect 16228 13499 16396 13533
rect 16486 13499 16654 13533
rect 16744 13499 16912 13533
rect 19048 13499 19216 13533
rect 19306 13499 19474 13533
rect 19564 13499 19732 13533
rect 19822 13499 19990 13533
rect 20080 13499 20248 13533
rect 20338 13499 20506 13533
rect 20596 13499 20764 13533
rect 20854 13499 21022 13533
rect 21112 13499 21280 13533
rect 21370 13499 21538 13533
rect 21628 13499 21796 13533
rect 21886 13499 22054 13533
rect 22144 13499 22312 13533
rect 22402 13499 22570 13533
rect 22660 13499 22828 13533
rect 22918 13499 23086 13533
rect 23176 13499 23344 13533
rect 23434 13499 23602 13533
rect 23692 13499 23860 13533
rect 23950 13499 24118 13533
<< xpolycontact >>
rect 17690 14980 18260 15460
rect 17690 14240 18260 14720
<< ppolyres >>
rect 17690 14720 18260 14980
<< locali >>
rect 11666 17235 11700 17332
rect 17054 17235 17088 17332
rect 11780 17208 11814 17224
rect 11780 16216 11814 16232
rect 12038 17208 12072 17224
rect 12038 16173 12072 16232
rect 12296 17208 12330 17224
rect 12296 16216 12330 16232
rect 12554 17208 12588 17224
rect 12554 16173 12588 16232
rect 12812 17208 12846 17224
rect 12812 16216 12846 16232
rect 13070 17208 13104 17224
rect 13070 16173 13104 16232
rect 13328 17208 13362 17224
rect 13328 16216 13362 16232
rect 13586 17208 13620 17224
rect 13586 16173 13620 16232
rect 13844 17208 13878 17224
rect 13844 16216 13878 16232
rect 14102 17208 14136 17224
rect 14102 16173 14136 16232
rect 14360 17208 14394 17224
rect 14360 16216 14394 16232
rect 14618 17208 14652 17224
rect 14618 16173 14652 16232
rect 14876 17208 14910 17224
rect 14876 16216 14910 16232
rect 15134 17208 15168 17224
rect 15134 16173 15168 16232
rect 15392 17208 15426 17224
rect 15392 16216 15426 16232
rect 15650 17208 15684 17224
rect 15650 16173 15684 16232
rect 15908 17208 15942 17224
rect 15908 16216 15942 16232
rect 16166 17208 16200 17224
rect 16166 16173 16200 16232
rect 16424 17208 16458 17224
rect 16424 16216 16458 16232
rect 16682 17208 16716 17224
rect 16682 16173 16716 16232
rect 16940 17208 16974 17224
rect 16940 16216 16974 16232
rect 11780 16139 11842 16173
rect 12010 16139 12100 16173
rect 12268 16139 12358 16173
rect 12526 16139 12616 16173
rect 12784 16139 12874 16173
rect 13042 16139 13132 16173
rect 13300 16139 13390 16173
rect 13558 16139 13648 16173
rect 13816 16139 13906 16173
rect 14074 16139 14164 16173
rect 14332 16139 14422 16173
rect 14590 16139 14680 16173
rect 14848 16139 14938 16173
rect 15106 16139 15196 16173
rect 15364 16139 15454 16173
rect 15622 16139 15712 16173
rect 15880 16139 15970 16173
rect 16138 16139 16228 16173
rect 16396 16139 16486 16173
rect 16654 16139 16744 16173
rect 16912 16139 16974 16173
rect 11666 16070 11700 16133
rect 17054 16070 17088 16133
rect 11666 16036 11762 16070
rect 16992 16036 17088 16070
rect 18872 17235 18906 17332
rect 24260 17235 24294 17332
rect 18986 17208 19020 17224
rect 18986 16216 19020 16232
rect 19244 17208 19278 17224
rect 19244 16173 19278 16232
rect 19502 17208 19536 17224
rect 19502 16216 19536 16232
rect 19760 17208 19794 17224
rect 19760 16173 19794 16232
rect 20018 17208 20052 17224
rect 20018 16216 20052 16232
rect 20276 17208 20310 17224
rect 20276 16173 20310 16232
rect 20534 17208 20568 17224
rect 20534 16216 20568 16232
rect 20792 17208 20826 17224
rect 20792 16173 20826 16232
rect 21050 17208 21084 17224
rect 21050 16216 21084 16232
rect 21308 17208 21342 17224
rect 21308 16173 21342 16232
rect 21566 17208 21600 17224
rect 21566 16216 21600 16232
rect 21824 17208 21858 17224
rect 21824 16173 21858 16232
rect 22082 17208 22116 17224
rect 22082 16216 22116 16232
rect 22340 17208 22374 17224
rect 22340 16173 22374 16232
rect 22598 17208 22632 17224
rect 22598 16216 22632 16232
rect 22856 17208 22890 17224
rect 22856 16173 22890 16232
rect 23114 17208 23148 17224
rect 23114 16216 23148 16232
rect 23372 17208 23406 17224
rect 23372 16173 23406 16232
rect 23630 17208 23664 17224
rect 23630 16216 23664 16232
rect 23888 17208 23922 17224
rect 23888 16173 23922 16232
rect 24146 17208 24180 17224
rect 24146 16216 24180 16232
rect 18986 16139 19048 16173
rect 19216 16139 19306 16173
rect 19474 16139 19564 16173
rect 19732 16139 19822 16173
rect 19990 16139 20080 16173
rect 20248 16139 20338 16173
rect 20506 16139 20596 16173
rect 20764 16139 20854 16173
rect 21022 16139 21112 16173
rect 21280 16139 21370 16173
rect 21538 16139 21628 16173
rect 21796 16139 21886 16173
rect 22054 16139 22144 16173
rect 22312 16139 22402 16173
rect 22570 16139 22660 16173
rect 22828 16139 22918 16173
rect 23086 16139 23176 16173
rect 23344 16139 23434 16173
rect 23602 16139 23692 16173
rect 23860 16139 23950 16173
rect 24118 16139 24180 16173
rect 18872 16070 18906 16133
rect 24260 16070 24294 16133
rect 18872 16036 18968 16070
rect 24198 16036 24294 16070
rect 11666 13601 11762 13635
rect 16992 13601 17088 13635
rect 11666 13539 11700 13601
rect 17054 13539 17088 13601
rect 11778 13499 11842 13533
rect 12010 13499 12100 13533
rect 12268 13499 12358 13533
rect 12526 13499 12616 13533
rect 12784 13499 12874 13533
rect 13042 13499 13132 13533
rect 13300 13499 13390 13533
rect 13558 13499 13648 13533
rect 13816 13499 13906 13533
rect 14074 13499 14164 13533
rect 14332 13499 14422 13533
rect 14590 13499 14680 13533
rect 14848 13499 14938 13533
rect 15106 13499 15196 13533
rect 15364 13499 15454 13533
rect 15622 13499 15712 13533
rect 15880 13499 15970 13533
rect 16138 13499 16228 13533
rect 16396 13499 16486 13533
rect 16654 13499 16744 13533
rect 16912 13499 16975 13533
rect 11780 13449 11814 13465
rect 11780 12457 11814 12473
rect 12038 13449 12072 13499
rect 12038 12457 12072 12473
rect 12296 13449 12330 13465
rect 12296 12457 12330 12473
rect 12554 13449 12588 13499
rect 12554 12457 12588 12473
rect 12812 13449 12846 13465
rect 12812 12457 12846 12473
rect 13070 13449 13104 13499
rect 13070 12457 13104 12473
rect 13328 13449 13362 13465
rect 13328 12457 13362 12473
rect 13586 13449 13620 13499
rect 13586 12457 13620 12473
rect 13844 13449 13878 13465
rect 13844 12457 13878 12473
rect 14102 13449 14136 13499
rect 14102 12457 14136 12473
rect 14360 13449 14394 13465
rect 14360 12457 14394 12473
rect 14618 13449 14652 13499
rect 14618 12457 14652 12473
rect 14876 13449 14910 13465
rect 14876 12457 14910 12473
rect 15134 13449 15168 13499
rect 15134 12457 15168 12473
rect 15392 13449 15426 13465
rect 15392 12457 15426 12473
rect 15650 13449 15684 13499
rect 15650 12457 15684 12473
rect 15908 13449 15942 13465
rect 15908 12457 15942 12473
rect 16166 13449 16200 13499
rect 16166 12457 16200 12473
rect 16424 13449 16458 13465
rect 16424 12457 16458 12473
rect 16682 13449 16716 13499
rect 16682 12457 16716 12473
rect 16940 13449 16974 13465
rect 16940 12457 16974 12473
rect 11666 12349 11700 12445
rect 17054 12349 17088 12445
rect 18872 13601 18968 13635
rect 24198 13601 24294 13635
rect 18872 13539 18906 13601
rect 24260 13539 24294 13601
rect 18985 13499 19048 13533
rect 19216 13499 19306 13533
rect 19474 13499 19564 13533
rect 19732 13499 19822 13533
rect 19990 13499 20080 13533
rect 20248 13499 20338 13533
rect 20506 13499 20596 13533
rect 20764 13499 20854 13533
rect 21022 13499 21112 13533
rect 21280 13499 21370 13533
rect 21538 13499 21628 13533
rect 21796 13499 21886 13533
rect 22054 13499 22144 13533
rect 22312 13499 22402 13533
rect 22570 13499 22660 13533
rect 22828 13499 22918 13533
rect 23086 13499 23176 13533
rect 23344 13499 23434 13533
rect 23602 13499 23692 13533
rect 23860 13499 23950 13533
rect 24118 13499 24182 13533
rect 18986 13449 19020 13465
rect 18986 12457 19020 12473
rect 19244 13449 19278 13499
rect 19244 12457 19278 12473
rect 19502 13449 19536 13465
rect 19502 12457 19536 12473
rect 19760 13449 19794 13499
rect 19760 12457 19794 12473
rect 20018 13449 20052 13465
rect 20018 12457 20052 12473
rect 20276 13449 20310 13499
rect 20276 12457 20310 12473
rect 20534 13449 20568 13465
rect 20534 12457 20568 12473
rect 20792 13449 20826 13499
rect 20792 12457 20826 12473
rect 21050 13449 21084 13465
rect 21050 12457 21084 12473
rect 21308 13449 21342 13499
rect 21308 12457 21342 12473
rect 21566 13449 21600 13465
rect 21566 12457 21600 12473
rect 21824 13449 21858 13499
rect 21824 12457 21858 12473
rect 22082 13449 22116 13465
rect 22082 12457 22116 12473
rect 22340 13449 22374 13499
rect 22340 12457 22374 12473
rect 22598 13449 22632 13465
rect 22598 12457 22632 12473
rect 22856 13449 22890 13499
rect 22856 12457 22890 12473
rect 23114 13449 23148 13465
rect 23114 12457 23148 12473
rect 23372 13449 23406 13499
rect 23372 12457 23406 12473
rect 23630 13449 23664 13465
rect 23630 12457 23664 12473
rect 23888 13449 23922 13499
rect 23888 12457 23922 12473
rect 24146 13449 24180 13465
rect 24146 12457 24180 12473
rect 18872 12349 18906 12445
rect 24260 12349 24294 12445
<< viali >>
rect 11700 17298 11762 17332
rect 11762 17298 16992 17332
rect 16992 17298 17054 17332
rect 11666 16193 11700 17175
rect 11780 16232 11814 17208
rect 12038 16232 12072 17208
rect 12296 16232 12330 17208
rect 12554 16232 12588 17208
rect 12812 16232 12846 17208
rect 13070 16232 13104 17208
rect 13328 16232 13362 17208
rect 13586 16232 13620 17208
rect 13844 16232 13878 17208
rect 14102 16232 14136 17208
rect 14360 16232 14394 17208
rect 14618 16232 14652 17208
rect 14876 16232 14910 17208
rect 15134 16232 15168 17208
rect 15392 16232 15426 17208
rect 15650 16232 15684 17208
rect 15908 16232 15942 17208
rect 16166 16232 16200 17208
rect 16424 16232 16458 17208
rect 16682 16232 16716 17208
rect 16940 16232 16974 17208
rect 17054 16193 17088 17175
rect 11884 16139 11968 16173
rect 12142 16139 12226 16173
rect 12400 16139 12484 16173
rect 12658 16139 12742 16173
rect 12916 16139 13000 16173
rect 13174 16139 13258 16173
rect 13432 16139 13516 16173
rect 13690 16139 13774 16173
rect 13948 16139 14032 16173
rect 14206 16139 14290 16173
rect 14464 16139 14548 16173
rect 14722 16139 14806 16173
rect 14980 16139 15064 16173
rect 15238 16139 15322 16173
rect 15496 16139 15580 16173
rect 15754 16139 15838 16173
rect 16012 16139 16096 16173
rect 16270 16139 16354 16173
rect 16528 16139 16612 16173
rect 16786 16139 16870 16173
rect 18906 17298 18968 17332
rect 18968 17298 24198 17332
rect 24198 17298 24260 17332
rect 18872 16193 18906 17175
rect 18986 16232 19020 17208
rect 19244 16232 19278 17208
rect 19502 16232 19536 17208
rect 19760 16232 19794 17208
rect 20018 16232 20052 17208
rect 20276 16232 20310 17208
rect 20534 16232 20568 17208
rect 20792 16232 20826 17208
rect 21050 16232 21084 17208
rect 21308 16232 21342 17208
rect 21566 16232 21600 17208
rect 21824 16232 21858 17208
rect 22082 16232 22116 17208
rect 22340 16232 22374 17208
rect 22598 16232 22632 17208
rect 22856 16232 22890 17208
rect 23114 16232 23148 17208
rect 23372 16232 23406 17208
rect 23630 16232 23664 17208
rect 23888 16232 23922 17208
rect 24146 16232 24180 17208
rect 24260 16193 24294 17175
rect 19090 16139 19174 16173
rect 19348 16139 19432 16173
rect 19606 16139 19690 16173
rect 19864 16139 19948 16173
rect 20122 16139 20206 16173
rect 20380 16139 20464 16173
rect 20638 16139 20722 16173
rect 20896 16139 20980 16173
rect 21154 16139 21238 16173
rect 21412 16139 21496 16173
rect 21670 16139 21754 16173
rect 21928 16139 22012 16173
rect 22186 16139 22270 16173
rect 22444 16139 22528 16173
rect 22702 16139 22786 16173
rect 22960 16139 23044 16173
rect 23218 16139 23302 16173
rect 23476 16139 23560 16173
rect 23734 16139 23818 16173
rect 23992 16139 24076 16173
rect 17710 15400 17750 15440
rect 17790 15400 17830 15440
rect 17870 15400 17910 15440
rect 17950 15400 18000 15440
rect 18040 15400 18080 15440
rect 18120 15400 18160 15440
rect 18200 15400 18240 15440
rect 17710 15320 17750 15360
rect 17790 15320 17830 15360
rect 17870 15320 17910 15360
rect 17950 15320 18000 15360
rect 18040 15320 18080 15360
rect 18120 15320 18160 15360
rect 18200 15320 18240 15360
rect 17710 15240 17750 15280
rect 17790 15240 17830 15280
rect 17870 15240 17910 15280
rect 17950 15240 18000 15280
rect 18040 15240 18080 15280
rect 18120 15240 18160 15280
rect 18200 15240 18240 15280
rect 17710 15160 17750 15200
rect 17790 15160 17830 15200
rect 17870 15160 17910 15200
rect 17950 15160 18000 15200
rect 18040 15160 18080 15200
rect 18120 15160 18160 15200
rect 18200 15160 18240 15200
rect 17710 15080 17750 15120
rect 17790 15080 17830 15120
rect 17870 15080 17910 15120
rect 17950 15080 18000 15120
rect 18040 15080 18080 15120
rect 18120 15080 18160 15120
rect 18200 15080 18240 15120
rect 17710 15000 17750 15040
rect 17790 15000 17830 15040
rect 17870 15000 17910 15040
rect 17950 15000 18000 15040
rect 18040 15000 18080 15040
rect 18120 15000 18160 15040
rect 18200 15000 18240 15040
rect 17710 14660 17750 14700
rect 17790 14660 17830 14700
rect 17870 14660 17910 14700
rect 17950 14660 18000 14700
rect 18040 14660 18080 14700
rect 18120 14660 18160 14700
rect 18200 14660 18240 14700
rect 17710 14580 17750 14620
rect 17790 14580 17830 14620
rect 17870 14580 17910 14620
rect 17950 14580 18000 14620
rect 18040 14580 18080 14620
rect 18120 14580 18160 14620
rect 18200 14580 18240 14620
rect 17710 14500 17750 14540
rect 17790 14500 17830 14540
rect 17870 14500 17910 14540
rect 17950 14500 18000 14540
rect 18040 14500 18080 14540
rect 18120 14500 18160 14540
rect 18200 14500 18240 14540
rect 17710 14420 17750 14460
rect 17790 14420 17830 14460
rect 17870 14420 17910 14460
rect 17950 14420 18000 14460
rect 18040 14420 18080 14460
rect 18120 14420 18160 14460
rect 18200 14420 18240 14460
rect 17710 14340 17750 14380
rect 17790 14340 17830 14380
rect 17870 14340 17910 14380
rect 17950 14340 18000 14380
rect 18040 14340 18080 14380
rect 18120 14340 18160 14380
rect 18200 14340 18240 14380
rect 17710 14260 17750 14300
rect 17790 14260 17830 14300
rect 17870 14260 17910 14300
rect 17950 14260 18000 14300
rect 18040 14260 18080 14300
rect 18120 14260 18160 14300
rect 18200 14260 18240 14300
rect 11884 13499 11968 13533
rect 12142 13499 12226 13533
rect 12400 13499 12484 13533
rect 12658 13499 12742 13533
rect 12916 13499 13000 13533
rect 13174 13499 13258 13533
rect 13432 13499 13516 13533
rect 13690 13499 13774 13533
rect 13948 13499 14032 13533
rect 14206 13499 14290 13533
rect 14464 13499 14548 13533
rect 14722 13499 14806 13533
rect 14980 13499 15064 13533
rect 15238 13499 15322 13533
rect 15496 13499 15580 13533
rect 15754 13499 15838 13533
rect 16012 13499 16096 13533
rect 16270 13499 16354 13533
rect 16528 13499 16612 13533
rect 16786 13499 16870 13533
rect 11666 12505 11700 13479
rect 11780 12473 11814 13449
rect 12038 12473 12072 13449
rect 12296 12473 12330 13449
rect 12554 12473 12588 13449
rect 12812 12473 12846 13449
rect 13070 12473 13104 13449
rect 13328 12473 13362 13449
rect 13586 12473 13620 13449
rect 13844 12473 13878 13449
rect 14102 12473 14136 13449
rect 14360 12473 14394 13449
rect 14618 12473 14652 13449
rect 14876 12473 14910 13449
rect 15134 12473 15168 13449
rect 15392 12473 15426 13449
rect 15650 12473 15684 13449
rect 15908 12473 15942 13449
rect 16166 12473 16200 13449
rect 16424 12473 16458 13449
rect 16682 12473 16716 13449
rect 16940 12473 16974 13449
rect 17054 12505 17088 13479
rect 11700 12349 11762 12383
rect 11762 12349 16992 12383
rect 16992 12349 17054 12383
rect 19090 13499 19174 13533
rect 19348 13499 19432 13533
rect 19606 13499 19690 13533
rect 19864 13499 19948 13533
rect 20122 13499 20206 13533
rect 20380 13499 20464 13533
rect 20638 13499 20722 13533
rect 20896 13499 20980 13533
rect 21154 13499 21238 13533
rect 21412 13499 21496 13533
rect 21670 13499 21754 13533
rect 21928 13499 22012 13533
rect 22186 13499 22270 13533
rect 22444 13499 22528 13533
rect 22702 13499 22786 13533
rect 22960 13499 23044 13533
rect 23218 13499 23302 13533
rect 23476 13499 23560 13533
rect 23734 13499 23818 13533
rect 23992 13499 24076 13533
rect 18872 12505 18906 13479
rect 18986 12473 19020 13449
rect 19244 12473 19278 13449
rect 19502 12473 19536 13449
rect 19760 12473 19794 13449
rect 20018 12473 20052 13449
rect 20276 12473 20310 13449
rect 20534 12473 20568 13449
rect 20792 12473 20826 13449
rect 21050 12473 21084 13449
rect 21308 12473 21342 13449
rect 21566 12473 21600 13449
rect 21824 12473 21858 13449
rect 22082 12473 22116 13449
rect 22340 12473 22374 13449
rect 22598 12473 22632 13449
rect 22856 12473 22890 13449
rect 23114 12473 23148 13449
rect 23372 12473 23406 13449
rect 23630 12473 23664 13449
rect 23888 12473 23922 13449
rect 24146 12473 24180 13449
rect 24260 12505 24294 13479
rect 18906 12349 18968 12383
rect 18968 12349 24198 12383
rect 24198 12349 24260 12383
<< metal1 >>
rect 11690 17590 11930 17610
rect 12020 17590 12260 17610
rect 12350 17590 12590 17610
rect 12680 17590 12920 17610
rect 13010 17590 13250 17610
rect 13340 17590 13580 17610
rect 13670 17590 13910 17610
rect 14000 17590 14240 17610
rect 14330 17590 14570 17610
rect 14660 17590 14900 17610
rect 14990 17590 15230 17610
rect 15320 17590 15560 17610
rect 15650 17590 15890 17610
rect 15980 17590 16220 17610
rect 16310 17590 16550 17610
rect 16640 17590 16880 17610
rect 19080 17590 19320 17610
rect 19410 17590 19650 17610
rect 19740 17590 19980 17610
rect 20070 17590 20310 17610
rect 20400 17590 20640 17610
rect 20730 17590 20970 17610
rect 21060 17590 21300 17610
rect 21390 17590 21630 17610
rect 21720 17590 21960 17610
rect 22050 17590 22290 17610
rect 22380 17590 22620 17610
rect 22710 17590 22950 17610
rect 23040 17590 23280 17610
rect 23370 17590 23610 17610
rect 23700 17590 23940 17610
rect 24030 17590 24270 17610
rect 11660 17570 17094 17590
rect 11660 17560 14660 17570
rect 11660 17490 11690 17560
rect 11760 17490 11810 17560
rect 11880 17490 12020 17560
rect 12090 17490 12140 17560
rect 12210 17490 12350 17560
rect 12420 17490 12470 17560
rect 12540 17490 12680 17560
rect 12750 17490 12800 17560
rect 12870 17490 13010 17560
rect 13080 17490 13130 17560
rect 13200 17490 13340 17560
rect 13410 17490 13460 17560
rect 13530 17490 13670 17560
rect 13740 17490 13790 17560
rect 13860 17490 14000 17560
rect 14070 17490 14120 17560
rect 14190 17490 14330 17560
rect 14400 17490 14450 17560
rect 14520 17500 14660 17560
rect 14730 17500 14780 17570
rect 14850 17500 14990 17570
rect 15060 17500 15110 17570
rect 15180 17500 15320 17570
rect 15390 17500 15440 17570
rect 15510 17560 17094 17570
rect 15510 17500 15650 17560
rect 14520 17490 15650 17500
rect 15720 17490 15770 17560
rect 15840 17490 15980 17560
rect 16050 17490 16100 17560
rect 16170 17490 16310 17560
rect 16380 17490 16430 17560
rect 16500 17490 16640 17560
rect 16710 17490 16760 17560
rect 16830 17490 17094 17560
rect 11660 17450 17094 17490
rect 11660 17440 14660 17450
rect 11660 17370 11690 17440
rect 11760 17370 11810 17440
rect 11880 17370 12020 17440
rect 12090 17370 12140 17440
rect 12210 17370 12350 17440
rect 12420 17370 12470 17440
rect 12540 17370 12680 17440
rect 12750 17370 12800 17440
rect 12870 17370 13010 17440
rect 13080 17370 13130 17440
rect 13200 17370 13340 17440
rect 13410 17370 13460 17440
rect 13530 17370 13670 17440
rect 13740 17370 13790 17440
rect 13860 17370 14000 17440
rect 14070 17370 14120 17440
rect 14190 17370 14330 17440
rect 14400 17370 14450 17440
rect 14520 17380 14660 17440
rect 14730 17380 14780 17450
rect 14850 17380 14990 17450
rect 15060 17380 15110 17450
rect 15180 17380 15320 17450
rect 15390 17380 15440 17450
rect 15510 17440 17094 17450
rect 15510 17380 15650 17440
rect 14520 17370 15650 17380
rect 15720 17370 15770 17440
rect 15840 17370 15980 17440
rect 16050 17370 16100 17440
rect 16170 17370 16310 17440
rect 16380 17370 16430 17440
rect 16500 17370 16640 17440
rect 16710 17370 16760 17440
rect 16830 17370 17094 17440
rect 11660 17332 17094 17370
rect 11660 17298 11700 17332
rect 17054 17298 17094 17332
rect 11660 17292 17094 17298
rect 11660 17175 11706 17292
rect 11660 16193 11666 17175
rect 11700 16193 11706 17175
rect 11660 16181 11706 16193
rect 11774 17208 11820 17220
rect 11774 16232 11780 17208
rect 11814 16232 11820 17208
rect 11774 16100 11820 16232
rect 12032 17208 12078 17292
rect 12032 16232 12038 17208
rect 12072 16232 12078 17208
rect 12032 16220 12078 16232
rect 12290 17208 12336 17220
rect 12290 16232 12296 17208
rect 12330 16232 12336 17208
rect 11872 16173 11980 16179
rect 11872 16139 11884 16173
rect 11968 16139 11980 16173
rect 11872 16133 11980 16139
rect 12130 16173 12238 16179
rect 12130 16139 12142 16173
rect 12226 16139 12238 16173
rect 12130 16133 12238 16139
rect 12290 16100 12336 16232
rect 12548 17208 12594 17292
rect 12548 16232 12554 17208
rect 12588 16232 12594 17208
rect 12548 16220 12594 16232
rect 12806 17208 12852 17220
rect 12806 16232 12812 17208
rect 12846 16232 12852 17208
rect 12388 16173 12496 16179
rect 12388 16139 12400 16173
rect 12484 16139 12496 16173
rect 12388 16133 12496 16139
rect 12646 16173 12754 16179
rect 12646 16139 12658 16173
rect 12742 16139 12754 16173
rect 12646 16133 12754 16139
rect 12806 16100 12852 16232
rect 13064 17208 13110 17292
rect 13064 16232 13070 17208
rect 13104 16232 13110 17208
rect 13064 16220 13110 16232
rect 13322 17208 13368 17220
rect 13322 16232 13328 17208
rect 13362 16232 13368 17208
rect 12904 16173 13012 16179
rect 12904 16139 12916 16173
rect 13000 16139 13012 16173
rect 12904 16133 13012 16139
rect 13162 16173 13270 16179
rect 13162 16139 13174 16173
rect 13258 16139 13270 16173
rect 13162 16133 13270 16139
rect 13322 16100 13368 16232
rect 13580 17208 13626 17292
rect 13580 16232 13586 17208
rect 13620 16232 13626 17208
rect 13580 16220 13626 16232
rect 13838 17208 13884 17220
rect 13838 16232 13844 17208
rect 13878 16232 13884 17208
rect 13420 16173 13528 16179
rect 13420 16139 13432 16173
rect 13516 16139 13528 16173
rect 13420 16133 13528 16139
rect 13678 16173 13786 16179
rect 13678 16139 13690 16173
rect 13774 16139 13786 16173
rect 13678 16133 13786 16139
rect 13838 16100 13884 16232
rect 14096 17208 14142 17292
rect 14096 16232 14102 17208
rect 14136 16232 14142 17208
rect 14096 16220 14142 16232
rect 14354 17208 14400 17220
rect 14354 16232 14360 17208
rect 14394 16232 14400 17208
rect 13936 16173 14044 16179
rect 13936 16139 13948 16173
rect 14032 16139 14044 16173
rect 13936 16133 14044 16139
rect 14194 16173 14302 16179
rect 14194 16139 14206 16173
rect 14290 16139 14302 16173
rect 14194 16133 14302 16139
rect 14354 16100 14400 16232
rect 14612 17208 14658 17292
rect 14612 16232 14618 17208
rect 14652 16232 14658 17208
rect 14612 16220 14658 16232
rect 14870 17208 14916 17220
rect 14870 16232 14876 17208
rect 14910 16232 14916 17208
rect 14452 16173 14560 16179
rect 14452 16139 14464 16173
rect 14548 16139 14560 16173
rect 14452 16133 14560 16139
rect 14710 16173 14818 16179
rect 14710 16139 14722 16173
rect 14806 16139 14818 16173
rect 14710 16133 14818 16139
rect 14870 16100 14916 16232
rect 15128 17208 15174 17292
rect 15128 16232 15134 17208
rect 15168 16232 15174 17208
rect 15128 16220 15174 16232
rect 15386 17208 15432 17220
rect 15386 16232 15392 17208
rect 15426 16232 15432 17208
rect 14968 16173 15076 16179
rect 14968 16139 14980 16173
rect 15064 16139 15076 16173
rect 14968 16133 15076 16139
rect 15226 16173 15334 16179
rect 15226 16139 15238 16173
rect 15322 16139 15334 16173
rect 15226 16133 15334 16139
rect 15386 16100 15432 16232
rect 15644 17208 15690 17292
rect 15644 16232 15650 17208
rect 15684 16232 15690 17208
rect 15644 16220 15690 16232
rect 15902 17208 15948 17220
rect 15902 16232 15908 17208
rect 15942 16232 15948 17208
rect 15484 16173 15592 16179
rect 15484 16139 15496 16173
rect 15580 16139 15592 16173
rect 15484 16133 15592 16139
rect 15742 16173 15850 16179
rect 15742 16139 15754 16173
rect 15838 16139 15850 16173
rect 15742 16133 15850 16139
rect 15902 16100 15948 16232
rect 16160 17208 16206 17292
rect 16160 16232 16166 17208
rect 16200 16232 16206 17208
rect 16160 16220 16206 16232
rect 16418 17208 16464 17220
rect 16418 16232 16424 17208
rect 16458 16232 16464 17208
rect 16000 16173 16108 16179
rect 16000 16139 16012 16173
rect 16096 16139 16108 16173
rect 16000 16133 16108 16139
rect 16258 16173 16366 16179
rect 16258 16139 16270 16173
rect 16354 16139 16366 16173
rect 16258 16133 16366 16139
rect 16418 16100 16464 16232
rect 16676 17208 16722 17292
rect 16676 16232 16682 17208
rect 16716 16232 16722 17208
rect 16676 16220 16722 16232
rect 16934 17208 16980 17220
rect 16934 16232 16940 17208
rect 16974 16232 16980 17208
rect 16516 16173 16624 16179
rect 16516 16139 16528 16173
rect 16612 16139 16624 16173
rect 16516 16133 16624 16139
rect 16774 16173 16882 16179
rect 16774 16139 16786 16173
rect 16870 16139 16882 16173
rect 16774 16133 16882 16139
rect 16934 16100 16980 16232
rect 17048 17175 17094 17292
rect 17048 16193 17054 17175
rect 17088 16193 17094 17175
rect 17048 16181 17094 16193
rect 18866 17570 24300 17590
rect 18866 17560 20450 17570
rect 18866 17490 19130 17560
rect 19200 17490 19250 17560
rect 19320 17490 19460 17560
rect 19530 17490 19580 17560
rect 19650 17490 19790 17560
rect 19860 17490 19910 17560
rect 19980 17490 20120 17560
rect 20190 17490 20240 17560
rect 20310 17500 20450 17560
rect 20520 17500 20570 17570
rect 20640 17500 20780 17570
rect 20850 17500 20900 17570
rect 20970 17500 21110 17570
rect 21180 17500 21230 17570
rect 21300 17560 24300 17570
rect 21300 17500 21440 17560
rect 20310 17490 21440 17500
rect 21510 17490 21560 17560
rect 21630 17490 21770 17560
rect 21840 17490 21890 17560
rect 21960 17490 22100 17560
rect 22170 17490 22220 17560
rect 22290 17490 22430 17560
rect 22500 17490 22550 17560
rect 22620 17490 22760 17560
rect 22830 17490 22880 17560
rect 22950 17490 23090 17560
rect 23160 17490 23210 17560
rect 23280 17490 23420 17560
rect 23490 17490 23540 17560
rect 23610 17490 23750 17560
rect 23820 17490 23870 17560
rect 23940 17490 24080 17560
rect 24150 17490 24200 17560
rect 24270 17490 24300 17560
rect 18866 17450 24300 17490
rect 18866 17440 20450 17450
rect 18866 17370 19130 17440
rect 19200 17370 19250 17440
rect 19320 17370 19460 17440
rect 19530 17370 19580 17440
rect 19650 17370 19790 17440
rect 19860 17370 19910 17440
rect 19980 17370 20120 17440
rect 20190 17370 20240 17440
rect 20310 17380 20450 17440
rect 20520 17380 20570 17450
rect 20640 17380 20780 17450
rect 20850 17380 20900 17450
rect 20970 17380 21110 17450
rect 21180 17380 21230 17450
rect 21300 17440 24300 17450
rect 21300 17380 21440 17440
rect 20310 17370 21440 17380
rect 21510 17370 21560 17440
rect 21630 17370 21770 17440
rect 21840 17370 21890 17440
rect 21960 17370 22100 17440
rect 22170 17370 22220 17440
rect 22290 17370 22430 17440
rect 22500 17370 22550 17440
rect 22620 17370 22760 17440
rect 22830 17370 22880 17440
rect 22950 17370 23090 17440
rect 23160 17370 23210 17440
rect 23280 17370 23420 17440
rect 23490 17370 23540 17440
rect 23610 17370 23750 17440
rect 23820 17370 23870 17440
rect 23940 17370 24080 17440
rect 24150 17370 24200 17440
rect 24270 17370 24300 17440
rect 18866 17332 24300 17370
rect 18866 17298 18906 17332
rect 24260 17298 24300 17332
rect 18866 17292 24300 17298
rect 18866 17175 18912 17292
rect 18866 16193 18872 17175
rect 18906 16193 18912 17175
rect 18866 16181 18912 16193
rect 18980 17208 19026 17220
rect 18980 16232 18986 17208
rect 19020 16232 19026 17208
rect 18980 16100 19026 16232
rect 19238 17208 19284 17292
rect 19238 16232 19244 17208
rect 19278 16232 19284 17208
rect 19238 16220 19284 16232
rect 19496 17208 19542 17220
rect 19496 16232 19502 17208
rect 19536 16232 19542 17208
rect 19078 16173 19186 16179
rect 19078 16139 19090 16173
rect 19174 16139 19186 16173
rect 19078 16133 19186 16139
rect 19336 16173 19444 16179
rect 19336 16139 19348 16173
rect 19432 16139 19444 16173
rect 19336 16133 19444 16139
rect 19496 16100 19542 16232
rect 19754 17208 19800 17292
rect 19754 16232 19760 17208
rect 19794 16232 19800 17208
rect 19754 16220 19800 16232
rect 20012 17208 20058 17220
rect 20012 16232 20018 17208
rect 20052 16232 20058 17208
rect 19594 16173 19702 16179
rect 19594 16139 19606 16173
rect 19690 16139 19702 16173
rect 19594 16133 19702 16139
rect 19852 16173 19960 16179
rect 19852 16139 19864 16173
rect 19948 16139 19960 16173
rect 19852 16133 19960 16139
rect 20012 16100 20058 16232
rect 20270 17208 20316 17292
rect 20270 16232 20276 17208
rect 20310 16232 20316 17208
rect 20270 16220 20316 16232
rect 20528 17208 20574 17220
rect 20528 16232 20534 17208
rect 20568 16232 20574 17208
rect 20110 16173 20218 16179
rect 20110 16139 20122 16173
rect 20206 16139 20218 16173
rect 20110 16133 20218 16139
rect 20368 16173 20476 16179
rect 20368 16139 20380 16173
rect 20464 16139 20476 16173
rect 20368 16133 20476 16139
rect 20528 16100 20574 16232
rect 20786 17208 20832 17292
rect 20786 16232 20792 17208
rect 20826 16232 20832 17208
rect 20786 16220 20832 16232
rect 21044 17208 21090 17220
rect 21044 16232 21050 17208
rect 21084 16232 21090 17208
rect 20626 16173 20734 16179
rect 20626 16139 20638 16173
rect 20722 16139 20734 16173
rect 20626 16133 20734 16139
rect 20884 16173 20992 16179
rect 20884 16139 20896 16173
rect 20980 16139 20992 16173
rect 20884 16133 20992 16139
rect 21044 16100 21090 16232
rect 21302 17208 21348 17292
rect 21302 16232 21308 17208
rect 21342 16232 21348 17208
rect 21302 16220 21348 16232
rect 21560 17208 21606 17220
rect 21560 16232 21566 17208
rect 21600 16232 21606 17208
rect 21142 16173 21250 16179
rect 21142 16139 21154 16173
rect 21238 16139 21250 16173
rect 21142 16133 21250 16139
rect 21400 16173 21508 16179
rect 21400 16139 21412 16173
rect 21496 16139 21508 16173
rect 21400 16133 21508 16139
rect 21560 16100 21606 16232
rect 21818 17208 21864 17292
rect 21818 16232 21824 17208
rect 21858 16232 21864 17208
rect 21818 16220 21864 16232
rect 22076 17208 22122 17220
rect 22076 16232 22082 17208
rect 22116 16232 22122 17208
rect 21658 16173 21766 16179
rect 21658 16139 21670 16173
rect 21754 16139 21766 16173
rect 21658 16133 21766 16139
rect 21916 16173 22024 16179
rect 21916 16139 21928 16173
rect 22012 16139 22024 16173
rect 21916 16133 22024 16139
rect 22076 16100 22122 16232
rect 22334 17208 22380 17292
rect 22334 16232 22340 17208
rect 22374 16232 22380 17208
rect 22334 16220 22380 16232
rect 22592 17208 22638 17220
rect 22592 16232 22598 17208
rect 22632 16232 22638 17208
rect 22174 16173 22282 16179
rect 22174 16139 22186 16173
rect 22270 16139 22282 16173
rect 22174 16133 22282 16139
rect 22432 16173 22540 16179
rect 22432 16139 22444 16173
rect 22528 16139 22540 16173
rect 22432 16133 22540 16139
rect 22592 16100 22638 16232
rect 22850 17208 22896 17292
rect 22850 16232 22856 17208
rect 22890 16232 22896 17208
rect 22850 16220 22896 16232
rect 23108 17208 23154 17220
rect 23108 16232 23114 17208
rect 23148 16232 23154 17208
rect 22690 16173 22798 16179
rect 22690 16139 22702 16173
rect 22786 16139 22798 16173
rect 22690 16133 22798 16139
rect 22948 16173 23056 16179
rect 22948 16139 22960 16173
rect 23044 16139 23056 16173
rect 22948 16133 23056 16139
rect 23108 16100 23154 16232
rect 23366 17208 23412 17292
rect 23366 16232 23372 17208
rect 23406 16232 23412 17208
rect 23366 16220 23412 16232
rect 23624 17208 23670 17220
rect 23624 16232 23630 17208
rect 23664 16232 23670 17208
rect 23206 16173 23314 16179
rect 23206 16139 23218 16173
rect 23302 16139 23314 16173
rect 23206 16133 23314 16139
rect 23464 16173 23572 16179
rect 23464 16139 23476 16173
rect 23560 16139 23572 16173
rect 23464 16133 23572 16139
rect 23624 16100 23670 16232
rect 23882 17208 23928 17292
rect 23882 16232 23888 17208
rect 23922 16232 23928 17208
rect 23882 16220 23928 16232
rect 24140 17208 24186 17220
rect 24140 16232 24146 17208
rect 24180 16232 24186 17208
rect 23722 16173 23830 16179
rect 23722 16139 23734 16173
rect 23818 16139 23830 16173
rect 23722 16133 23830 16139
rect 23980 16173 24088 16179
rect 23980 16139 23992 16173
rect 24076 16139 24088 16173
rect 23980 16133 24088 16139
rect 24140 16100 24186 16232
rect 24254 17175 24300 17292
rect 24254 16193 24260 17175
rect 24294 16193 24300 17175
rect 24254 16181 24300 16193
rect 11630 16070 18260 16100
rect 11630 15990 17740 16070
rect 11630 15930 11650 15990
rect 11710 15930 11740 15990
rect 11800 15930 11830 15990
rect 11890 15930 11920 15990
rect 11980 15930 12010 15990
rect 12070 15930 12100 15990
rect 12160 15930 12190 15990
rect 12250 15930 12280 15990
rect 12340 15930 12370 15990
rect 12430 15930 12460 15990
rect 12520 15930 12550 15990
rect 12610 15930 12640 15990
rect 12700 15930 12730 15990
rect 12790 15930 12820 15990
rect 12880 15930 12910 15990
rect 12970 15930 13000 15990
rect 13060 15930 13090 15990
rect 13150 15930 13180 15990
rect 13240 15930 13270 15990
rect 13330 15930 13360 15990
rect 13420 15930 13450 15990
rect 13510 15930 13540 15990
rect 13600 15930 13630 15990
rect 13690 15930 13720 15990
rect 13780 15930 13810 15990
rect 13870 15930 13900 15990
rect 13960 15930 13990 15990
rect 14050 15930 14080 15990
rect 14140 15930 14170 15990
rect 14230 15930 14260 15990
rect 14320 15930 14350 15990
rect 14410 15930 14440 15990
rect 14500 15930 14530 15990
rect 14590 15930 14620 15990
rect 14680 15930 14710 15990
rect 14770 15930 14800 15990
rect 14860 15930 14890 15990
rect 14950 15930 14980 15990
rect 15040 15930 15070 15990
rect 15130 15930 15160 15990
rect 15220 15930 15250 15990
rect 15310 15930 15340 15990
rect 15400 15930 15430 15990
rect 15490 15930 15520 15990
rect 15580 15930 15610 15990
rect 15670 15930 15700 15990
rect 15760 15930 15790 15990
rect 15850 15930 15880 15990
rect 15940 15930 15970 15990
rect 16030 15930 16060 15990
rect 16120 15930 16150 15990
rect 16210 15930 16240 15990
rect 16300 15930 16330 15990
rect 16390 15930 16420 15990
rect 16480 15930 16510 15990
rect 16570 15930 16600 15990
rect 16660 15930 16690 15990
rect 16750 15930 16780 15990
rect 16840 15930 16870 15990
rect 16930 15930 16960 15990
rect 17020 15930 17050 15990
rect 17110 15980 17740 15990
rect 17810 15980 17840 16070
rect 17910 15980 17940 16070
rect 18010 15980 18040 16070
rect 18110 15980 18140 16070
rect 18210 15980 18260 16070
rect 17110 15940 18260 15980
rect 17110 15930 17740 15940
rect 11630 15900 17740 15930
rect 11630 15840 11650 15900
rect 11710 15840 11740 15900
rect 11800 15840 11830 15900
rect 11890 15840 11920 15900
rect 11980 15840 12010 15900
rect 12070 15840 12100 15900
rect 12160 15840 12190 15900
rect 12250 15840 12280 15900
rect 12340 15840 12370 15900
rect 12430 15840 12460 15900
rect 12520 15840 12550 15900
rect 12610 15840 12640 15900
rect 12700 15840 12730 15900
rect 12790 15840 12820 15900
rect 12880 15840 12910 15900
rect 12970 15840 13000 15900
rect 13060 15840 13090 15900
rect 13150 15840 13180 15900
rect 13240 15840 13270 15900
rect 13330 15840 13360 15900
rect 13420 15840 13450 15900
rect 13510 15840 13540 15900
rect 13600 15840 13630 15900
rect 13690 15840 13720 15900
rect 13780 15840 13810 15900
rect 13870 15840 13900 15900
rect 13960 15840 13990 15900
rect 14050 15840 14080 15900
rect 14140 15840 14170 15900
rect 14230 15840 14260 15900
rect 14320 15840 14350 15900
rect 14410 15840 14440 15900
rect 14500 15840 14530 15900
rect 14590 15840 14620 15900
rect 14680 15840 14710 15900
rect 14770 15840 14800 15900
rect 14860 15840 14890 15900
rect 14950 15840 14980 15900
rect 15040 15840 15070 15900
rect 15130 15840 15160 15900
rect 15220 15840 15250 15900
rect 15310 15840 15340 15900
rect 15400 15840 15430 15900
rect 15490 15840 15520 15900
rect 15580 15840 15610 15900
rect 15670 15840 15700 15900
rect 15760 15840 15790 15900
rect 15850 15840 15880 15900
rect 15940 15840 15970 15900
rect 16030 15840 16060 15900
rect 16120 15840 16150 15900
rect 16210 15840 16240 15900
rect 16300 15840 16330 15900
rect 16390 15840 16420 15900
rect 16480 15840 16510 15900
rect 16570 15840 16600 15900
rect 16660 15840 16690 15900
rect 16750 15840 16780 15900
rect 16840 15840 16870 15900
rect 16930 15840 16960 15900
rect 17020 15840 17050 15900
rect 17110 15850 17740 15900
rect 17810 15850 17840 15940
rect 17910 15850 17940 15940
rect 18010 15850 18040 15940
rect 18110 15850 18140 15940
rect 18210 15850 18260 15940
rect 17110 15840 18260 15850
rect 11630 15820 18260 15840
rect 18980 15990 24330 16100
rect 18980 15930 19030 15990
rect 19090 15930 19120 15990
rect 19180 15930 19210 15990
rect 19270 15930 19300 15990
rect 19360 15930 19390 15990
rect 19450 15930 19480 15990
rect 19540 15930 19570 15990
rect 19630 15930 19660 15990
rect 19720 15930 19750 15990
rect 19810 15930 19840 15990
rect 19900 15930 19930 15990
rect 19990 15930 20020 15990
rect 20080 15930 20110 15990
rect 20170 15930 20200 15990
rect 20260 15930 20290 15990
rect 20350 15930 20380 15990
rect 20440 15930 20470 15990
rect 20530 15930 20560 15990
rect 20620 15930 20650 15990
rect 20710 15930 20740 15990
rect 20800 15930 20830 15990
rect 20890 15930 20920 15990
rect 20980 15930 21010 15990
rect 21070 15930 21100 15990
rect 21160 15930 21190 15990
rect 21250 15930 21280 15990
rect 21340 15930 21370 15990
rect 21430 15930 21460 15990
rect 21520 15930 21550 15990
rect 21610 15930 21640 15990
rect 21700 15930 21730 15990
rect 21790 15930 21820 15990
rect 21880 15930 21910 15990
rect 21970 15930 22000 15990
rect 22060 15930 22090 15990
rect 22150 15930 22180 15990
rect 22240 15930 22270 15990
rect 22330 15930 22360 15990
rect 22420 15930 22450 15990
rect 22510 15930 22540 15990
rect 22600 15930 22630 15990
rect 22690 15930 22720 15990
rect 22780 15930 22810 15990
rect 22870 15930 22900 15990
rect 22960 15930 22990 15990
rect 23050 15930 23080 15990
rect 23140 15930 23170 15990
rect 23230 15930 23260 15990
rect 23320 15930 23350 15990
rect 23410 15930 23440 15990
rect 23500 15930 23530 15990
rect 23590 15930 23620 15990
rect 23680 15930 23710 15990
rect 23770 15930 23800 15990
rect 23860 15930 23890 15990
rect 23950 15930 23980 15990
rect 24040 15930 24070 15990
rect 24130 15930 24160 15990
rect 24220 15930 24250 15990
rect 24310 15930 24330 15990
rect 18980 15900 24330 15930
rect 18980 15840 19030 15900
rect 19090 15840 19120 15900
rect 19180 15840 19210 15900
rect 19270 15840 19300 15900
rect 19360 15840 19390 15900
rect 19450 15840 19480 15900
rect 19540 15840 19570 15900
rect 19630 15840 19660 15900
rect 19720 15840 19750 15900
rect 19810 15840 19840 15900
rect 19900 15840 19930 15900
rect 19990 15840 20020 15900
rect 20080 15840 20110 15900
rect 20170 15840 20200 15900
rect 20260 15840 20290 15900
rect 20350 15840 20380 15900
rect 20440 15840 20470 15900
rect 20530 15840 20560 15900
rect 20620 15840 20650 15900
rect 20710 15840 20740 15900
rect 20800 15840 20830 15900
rect 20890 15840 20920 15900
rect 20980 15840 21010 15900
rect 21070 15840 21100 15900
rect 21160 15840 21190 15900
rect 21250 15840 21280 15900
rect 21340 15840 21370 15900
rect 21430 15840 21460 15900
rect 21520 15840 21550 15900
rect 21610 15840 21640 15900
rect 21700 15840 21730 15900
rect 21790 15840 21820 15900
rect 21880 15840 21910 15900
rect 21970 15840 22000 15900
rect 22060 15840 22090 15900
rect 22150 15840 22180 15900
rect 22240 15840 22270 15900
rect 22330 15840 22360 15900
rect 22420 15840 22450 15900
rect 22510 15840 22540 15900
rect 22600 15840 22630 15900
rect 22690 15840 22720 15900
rect 22780 15840 22810 15900
rect 22870 15840 22900 15900
rect 22960 15840 22990 15900
rect 23050 15840 23080 15900
rect 23140 15840 23170 15900
rect 23230 15840 23260 15900
rect 23320 15840 23350 15900
rect 23410 15840 23440 15900
rect 23500 15840 23530 15900
rect 23590 15840 23620 15900
rect 23680 15840 23710 15900
rect 23770 15840 23800 15900
rect 23860 15840 23890 15900
rect 23950 15840 23980 15900
rect 24040 15840 24070 15900
rect 24130 15840 24160 15900
rect 24220 15840 24250 15900
rect 24310 15840 24330 15900
rect 18980 15820 24330 15840
rect 17690 15440 18260 15820
rect 17690 15400 17710 15440
rect 17750 15400 17790 15440
rect 17830 15400 17870 15440
rect 17910 15400 17950 15440
rect 18000 15400 18040 15440
rect 18080 15400 18120 15440
rect 18160 15400 18200 15440
rect 18240 15400 18260 15440
rect 17690 15360 18260 15400
rect 17690 15320 17710 15360
rect 17750 15320 17790 15360
rect 17830 15320 17870 15360
rect 17910 15320 17950 15360
rect 18000 15320 18040 15360
rect 18080 15320 18120 15360
rect 18160 15320 18200 15360
rect 18240 15320 18260 15360
rect 17690 15280 18260 15320
rect 17690 15240 17710 15280
rect 17750 15240 17790 15280
rect 17830 15240 17870 15280
rect 17910 15240 17950 15280
rect 18000 15240 18040 15280
rect 18080 15240 18120 15280
rect 18160 15240 18200 15280
rect 18240 15240 18260 15280
rect 17690 15200 18260 15240
rect 17690 15160 17710 15200
rect 17750 15160 17790 15200
rect 17830 15160 17870 15200
rect 17910 15160 17950 15200
rect 18000 15160 18040 15200
rect 18080 15160 18120 15200
rect 18160 15160 18200 15200
rect 18240 15160 18260 15200
rect 17690 15120 18260 15160
rect 17690 15080 17710 15120
rect 17750 15080 17790 15120
rect 17830 15080 17870 15120
rect 17910 15080 17950 15120
rect 18000 15080 18040 15120
rect 18080 15080 18120 15120
rect 18160 15080 18200 15120
rect 18240 15080 18260 15120
rect 17690 15040 18260 15080
rect 17690 15000 17710 15040
rect 17750 15000 17790 15040
rect 17830 15000 17870 15040
rect 17910 15000 17950 15040
rect 18000 15000 18040 15040
rect 18080 15000 18120 15040
rect 18160 15000 18200 15040
rect 18240 15000 18260 15040
rect 17690 14980 18260 15000
rect 17690 14700 18260 14720
rect 17690 14660 17710 14700
rect 17750 14660 17790 14700
rect 17830 14660 17870 14700
rect 17910 14660 17950 14700
rect 18000 14660 18040 14700
rect 18080 14660 18120 14700
rect 18160 14660 18200 14700
rect 18240 14660 18260 14700
rect 17690 14620 18260 14660
rect 17690 14580 17710 14620
rect 17750 14580 17790 14620
rect 17830 14580 17870 14620
rect 17910 14580 17950 14620
rect 18000 14580 18040 14620
rect 18080 14580 18120 14620
rect 18160 14580 18200 14620
rect 18240 14580 18260 14620
rect 17690 14540 18260 14580
rect 17690 14500 17710 14540
rect 17750 14500 17790 14540
rect 17830 14500 17870 14540
rect 17910 14500 17950 14540
rect 18000 14500 18040 14540
rect 18080 14500 18120 14540
rect 18160 14500 18200 14540
rect 18240 14500 18260 14540
rect 17690 14460 18260 14500
rect 17690 14420 17710 14460
rect 17750 14420 17790 14460
rect 17830 14420 17870 14460
rect 17910 14420 17950 14460
rect 18000 14420 18040 14460
rect 18080 14420 18120 14460
rect 18160 14420 18200 14460
rect 18240 14420 18260 14460
rect 17690 14380 18260 14420
rect 17690 14340 17710 14380
rect 17750 14340 17790 14380
rect 17830 14340 17870 14380
rect 17910 14340 17950 14380
rect 18000 14340 18040 14380
rect 18080 14340 18120 14380
rect 18160 14340 18200 14380
rect 18240 14340 18260 14380
rect 17690 14300 18260 14340
rect 17690 14260 17710 14300
rect 17750 14260 17790 14300
rect 17830 14260 17870 14300
rect 17910 14260 17950 14300
rect 18000 14260 18040 14300
rect 18080 14260 18120 14300
rect 18160 14260 18200 14300
rect 18240 14260 18260 14300
rect 17690 13880 18260 14260
rect 11630 13860 16980 13880
rect 11630 13800 11650 13860
rect 11710 13800 11740 13860
rect 11800 13800 11830 13860
rect 11890 13800 11920 13860
rect 11980 13800 12010 13860
rect 12070 13800 12100 13860
rect 12160 13800 12190 13860
rect 12250 13800 12280 13860
rect 12340 13800 12370 13860
rect 12430 13800 12460 13860
rect 12520 13800 12550 13860
rect 12610 13800 12640 13860
rect 12700 13800 12730 13860
rect 12790 13800 12820 13860
rect 12880 13800 12910 13860
rect 12970 13800 13000 13860
rect 13060 13800 13090 13860
rect 13150 13800 13180 13860
rect 13240 13800 13270 13860
rect 13330 13800 13360 13860
rect 13420 13800 13450 13860
rect 13510 13800 13540 13860
rect 13600 13800 13630 13860
rect 13690 13800 13720 13860
rect 13780 13800 13810 13860
rect 13870 13800 13900 13860
rect 13960 13800 13990 13860
rect 14050 13800 14080 13860
rect 14140 13800 14170 13860
rect 14230 13800 14260 13860
rect 14320 13800 14350 13860
rect 14410 13800 14440 13860
rect 14500 13800 14530 13860
rect 14590 13800 14620 13860
rect 14680 13800 14710 13860
rect 14770 13800 14800 13860
rect 14860 13800 14890 13860
rect 14950 13800 14980 13860
rect 15040 13800 15070 13860
rect 15130 13800 15160 13860
rect 15220 13800 15250 13860
rect 15310 13800 15340 13860
rect 15400 13800 15430 13860
rect 15490 13800 15520 13860
rect 15580 13800 15610 13860
rect 15670 13800 15700 13860
rect 15760 13800 15790 13860
rect 15850 13800 15880 13860
rect 15940 13800 15970 13860
rect 16030 13800 16060 13860
rect 16120 13800 16150 13860
rect 16210 13800 16240 13860
rect 16300 13800 16330 13860
rect 16390 13800 16420 13860
rect 16480 13800 16510 13860
rect 16570 13800 16600 13860
rect 16660 13800 16690 13860
rect 16750 13800 16780 13860
rect 16840 13800 16870 13860
rect 16930 13800 16980 13860
rect 11630 13770 16980 13800
rect 11630 13710 11650 13770
rect 11710 13710 11740 13770
rect 11800 13710 11830 13770
rect 11890 13710 11920 13770
rect 11980 13710 12010 13770
rect 12070 13710 12100 13770
rect 12160 13710 12190 13770
rect 12250 13710 12280 13770
rect 12340 13710 12370 13770
rect 12430 13710 12460 13770
rect 12520 13710 12550 13770
rect 12610 13710 12640 13770
rect 12700 13710 12730 13770
rect 12790 13710 12820 13770
rect 12880 13710 12910 13770
rect 12970 13710 13000 13770
rect 13060 13710 13090 13770
rect 13150 13710 13180 13770
rect 13240 13710 13270 13770
rect 13330 13710 13360 13770
rect 13420 13710 13450 13770
rect 13510 13710 13540 13770
rect 13600 13710 13630 13770
rect 13690 13710 13720 13770
rect 13780 13710 13810 13770
rect 13870 13710 13900 13770
rect 13960 13710 13990 13770
rect 14050 13710 14080 13770
rect 14140 13710 14170 13770
rect 14230 13710 14260 13770
rect 14320 13710 14350 13770
rect 14410 13710 14440 13770
rect 14500 13710 14530 13770
rect 14590 13710 14620 13770
rect 14680 13710 14710 13770
rect 14770 13710 14800 13770
rect 14860 13710 14890 13770
rect 14950 13710 14980 13770
rect 15040 13710 15070 13770
rect 15130 13710 15160 13770
rect 15220 13710 15250 13770
rect 15310 13710 15340 13770
rect 15400 13710 15430 13770
rect 15490 13710 15520 13770
rect 15580 13710 15610 13770
rect 15670 13710 15700 13770
rect 15760 13710 15790 13770
rect 15850 13710 15880 13770
rect 15940 13710 15970 13770
rect 16030 13710 16060 13770
rect 16120 13710 16150 13770
rect 16210 13710 16240 13770
rect 16300 13710 16330 13770
rect 16390 13710 16420 13770
rect 16480 13710 16510 13770
rect 16570 13710 16600 13770
rect 16660 13710 16690 13770
rect 16750 13710 16780 13770
rect 16840 13710 16870 13770
rect 16930 13710 16980 13770
rect 11630 13600 16980 13710
rect 17690 13860 24330 13880
rect 17690 13850 18850 13860
rect 17690 13760 17740 13850
rect 17810 13760 17840 13850
rect 17910 13760 17940 13850
rect 18010 13760 18040 13850
rect 18110 13760 18140 13850
rect 18210 13800 18850 13850
rect 18910 13800 18940 13860
rect 19000 13800 19030 13860
rect 19090 13800 19120 13860
rect 19180 13800 19210 13860
rect 19270 13800 19300 13860
rect 19360 13800 19390 13860
rect 19450 13800 19480 13860
rect 19540 13800 19570 13860
rect 19630 13800 19660 13860
rect 19720 13800 19750 13860
rect 19810 13800 19840 13860
rect 19900 13800 19930 13860
rect 19990 13800 20020 13860
rect 20080 13800 20110 13860
rect 20170 13800 20200 13860
rect 20260 13800 20290 13860
rect 20350 13800 20380 13860
rect 20440 13800 20470 13860
rect 20530 13800 20560 13860
rect 20620 13800 20650 13860
rect 20710 13800 20740 13860
rect 20800 13800 20830 13860
rect 20890 13800 20920 13860
rect 20980 13800 21010 13860
rect 21070 13800 21100 13860
rect 21160 13800 21190 13860
rect 21250 13800 21280 13860
rect 21340 13800 21370 13860
rect 21430 13800 21460 13860
rect 21520 13800 21550 13860
rect 21610 13800 21640 13860
rect 21700 13800 21730 13860
rect 21790 13800 21820 13860
rect 21880 13800 21910 13860
rect 21970 13800 22000 13860
rect 22060 13800 22090 13860
rect 22150 13800 22180 13860
rect 22240 13800 22270 13860
rect 22330 13800 22360 13860
rect 22420 13800 22450 13860
rect 22510 13800 22540 13860
rect 22600 13800 22630 13860
rect 22690 13800 22720 13860
rect 22780 13800 22810 13860
rect 22870 13800 22900 13860
rect 22960 13800 22990 13860
rect 23050 13800 23080 13860
rect 23140 13800 23170 13860
rect 23230 13800 23260 13860
rect 23320 13800 23350 13860
rect 23410 13800 23440 13860
rect 23500 13800 23530 13860
rect 23590 13800 23620 13860
rect 23680 13800 23710 13860
rect 23770 13800 23800 13860
rect 23860 13800 23890 13860
rect 23950 13800 23980 13860
rect 24040 13800 24070 13860
rect 24130 13800 24160 13860
rect 24220 13800 24250 13860
rect 24310 13800 24330 13860
rect 18210 13770 24330 13800
rect 18210 13760 18850 13770
rect 17690 13720 18850 13760
rect 17690 13630 17740 13720
rect 17810 13630 17840 13720
rect 17910 13630 17940 13720
rect 18010 13630 18040 13720
rect 18110 13630 18140 13720
rect 18210 13710 18850 13720
rect 18910 13710 18940 13770
rect 19000 13710 19030 13770
rect 19090 13710 19120 13770
rect 19180 13710 19210 13770
rect 19270 13710 19300 13770
rect 19360 13710 19390 13770
rect 19450 13710 19480 13770
rect 19540 13710 19570 13770
rect 19630 13710 19660 13770
rect 19720 13710 19750 13770
rect 19810 13710 19840 13770
rect 19900 13710 19930 13770
rect 19990 13710 20020 13770
rect 20080 13710 20110 13770
rect 20170 13710 20200 13770
rect 20260 13710 20290 13770
rect 20350 13710 20380 13770
rect 20440 13710 20470 13770
rect 20530 13710 20560 13770
rect 20620 13710 20650 13770
rect 20710 13710 20740 13770
rect 20800 13710 20830 13770
rect 20890 13710 20920 13770
rect 20980 13710 21010 13770
rect 21070 13710 21100 13770
rect 21160 13710 21190 13770
rect 21250 13710 21280 13770
rect 21340 13710 21370 13770
rect 21430 13710 21460 13770
rect 21520 13710 21550 13770
rect 21610 13710 21640 13770
rect 21700 13710 21730 13770
rect 21790 13710 21820 13770
rect 21880 13710 21910 13770
rect 21970 13710 22000 13770
rect 22060 13710 22090 13770
rect 22150 13710 22180 13770
rect 22240 13710 22270 13770
rect 22330 13710 22360 13770
rect 22420 13710 22450 13770
rect 22510 13710 22540 13770
rect 22600 13710 22630 13770
rect 22690 13710 22720 13770
rect 22780 13710 22810 13770
rect 22870 13710 22900 13770
rect 22960 13710 22990 13770
rect 23050 13710 23080 13770
rect 23140 13710 23170 13770
rect 23230 13710 23260 13770
rect 23320 13710 23350 13770
rect 23410 13710 23440 13770
rect 23500 13710 23530 13770
rect 23590 13710 23620 13770
rect 23680 13710 23710 13770
rect 23770 13710 23800 13770
rect 23860 13710 23890 13770
rect 23950 13710 23980 13770
rect 24040 13710 24070 13770
rect 24130 13710 24160 13770
rect 24220 13710 24250 13770
rect 24310 13710 24330 13770
rect 18210 13630 24330 13710
rect 17690 13600 24330 13630
rect 11660 13479 11706 13491
rect 11660 12505 11666 13479
rect 11700 12505 11706 13479
rect 11660 12423 11706 12505
rect 11774 13449 11820 13600
rect 11872 13533 11980 13539
rect 11872 13499 11884 13533
rect 11968 13499 11980 13533
rect 11872 13493 11980 13499
rect 12130 13533 12238 13539
rect 12130 13499 12142 13533
rect 12226 13499 12238 13533
rect 12130 13493 12238 13499
rect 11774 12473 11780 13449
rect 11814 12473 11820 13449
rect 11774 12461 11820 12473
rect 12032 13449 12078 13461
rect 12032 12473 12038 13449
rect 12072 12473 12078 13449
rect 12032 12461 12078 12473
rect 12290 13449 12336 13600
rect 12388 13533 12496 13539
rect 12388 13499 12400 13533
rect 12484 13499 12496 13533
rect 12388 13493 12496 13499
rect 12646 13533 12754 13539
rect 12646 13499 12658 13533
rect 12742 13499 12754 13533
rect 12646 13493 12754 13499
rect 12290 12473 12296 13449
rect 12330 12473 12336 13449
rect 12290 12461 12336 12473
rect 12548 13449 12594 13461
rect 12548 12473 12554 13449
rect 12588 12473 12594 13449
rect 12548 12461 12594 12473
rect 12806 13449 12852 13600
rect 12904 13533 13012 13539
rect 12904 13499 12916 13533
rect 13000 13499 13012 13533
rect 12904 13493 13012 13499
rect 13162 13533 13270 13539
rect 13162 13499 13174 13533
rect 13258 13499 13270 13533
rect 13162 13493 13270 13499
rect 12806 12473 12812 13449
rect 12846 12473 12852 13449
rect 12806 12461 12852 12473
rect 13064 13449 13110 13461
rect 13064 12473 13070 13449
rect 13104 12473 13110 13449
rect 13064 12461 13110 12473
rect 13322 13449 13368 13600
rect 13420 13533 13528 13539
rect 13420 13499 13432 13533
rect 13516 13499 13528 13533
rect 13420 13493 13528 13499
rect 13678 13533 13786 13539
rect 13678 13499 13690 13533
rect 13774 13499 13786 13533
rect 13678 13493 13786 13499
rect 13322 12473 13328 13449
rect 13362 12473 13368 13449
rect 13322 12461 13368 12473
rect 13580 13449 13626 13461
rect 13580 12473 13586 13449
rect 13620 12473 13626 13449
rect 13580 12461 13626 12473
rect 13838 13449 13884 13600
rect 13936 13533 14044 13539
rect 13936 13499 13948 13533
rect 14032 13499 14044 13533
rect 13936 13493 14044 13499
rect 14194 13533 14302 13539
rect 14194 13499 14206 13533
rect 14290 13499 14302 13533
rect 14194 13493 14302 13499
rect 13838 12473 13844 13449
rect 13878 12473 13884 13449
rect 13838 12461 13884 12473
rect 14096 13449 14142 13461
rect 14096 12473 14102 13449
rect 14136 12473 14142 13449
rect 14096 12461 14142 12473
rect 14354 13449 14400 13600
rect 14452 13533 14560 13539
rect 14452 13499 14464 13533
rect 14548 13499 14560 13533
rect 14452 13493 14560 13499
rect 14710 13533 14818 13539
rect 14710 13499 14722 13533
rect 14806 13499 14818 13533
rect 14710 13493 14818 13499
rect 14354 12473 14360 13449
rect 14394 12473 14400 13449
rect 14354 12461 14400 12473
rect 14612 13449 14658 13461
rect 14612 12473 14618 13449
rect 14652 12473 14658 13449
rect 14612 12461 14658 12473
rect 14870 13449 14916 13600
rect 14968 13533 15076 13539
rect 14968 13499 14980 13533
rect 15064 13499 15076 13533
rect 14968 13493 15076 13499
rect 15226 13533 15334 13539
rect 15226 13499 15238 13533
rect 15322 13499 15334 13533
rect 15226 13493 15334 13499
rect 14870 12473 14876 13449
rect 14910 12473 14916 13449
rect 14870 12461 14916 12473
rect 15128 13449 15174 13461
rect 15128 12473 15134 13449
rect 15168 12473 15174 13449
rect 15128 12461 15174 12473
rect 15386 13449 15432 13600
rect 15484 13533 15592 13539
rect 15484 13499 15496 13533
rect 15580 13499 15592 13533
rect 15484 13493 15592 13499
rect 15742 13533 15850 13539
rect 15742 13499 15754 13533
rect 15838 13499 15850 13533
rect 15742 13493 15850 13499
rect 15386 12473 15392 13449
rect 15426 12473 15432 13449
rect 15386 12461 15432 12473
rect 15644 13449 15690 13461
rect 15644 12473 15650 13449
rect 15684 12473 15690 13449
rect 15644 12461 15690 12473
rect 15902 13449 15948 13600
rect 16000 13533 16108 13539
rect 16000 13499 16012 13533
rect 16096 13499 16108 13533
rect 16000 13493 16108 13499
rect 16258 13533 16366 13539
rect 16258 13499 16270 13533
rect 16354 13499 16366 13533
rect 16258 13493 16366 13499
rect 15902 12473 15908 13449
rect 15942 12473 15948 13449
rect 15902 12461 15948 12473
rect 16160 13449 16206 13461
rect 16160 12473 16166 13449
rect 16200 12473 16206 13449
rect 16160 12461 16206 12473
rect 16418 13449 16464 13600
rect 16516 13533 16624 13539
rect 16516 13499 16528 13533
rect 16612 13499 16624 13533
rect 16516 13493 16624 13499
rect 16774 13533 16882 13539
rect 16774 13499 16786 13533
rect 16870 13499 16882 13533
rect 16774 13493 16882 13499
rect 16418 12473 16424 13449
rect 16458 12473 16464 13449
rect 16418 12461 16464 12473
rect 16676 13449 16722 13461
rect 16676 12473 16682 13449
rect 16716 12473 16722 13449
rect 16676 12461 16722 12473
rect 16934 13449 16980 13600
rect 16934 12473 16940 13449
rect 16974 12473 16980 13449
rect 16934 12461 16980 12473
rect 17048 13479 17094 13491
rect 17048 12505 17054 13479
rect 17088 12505 17094 13479
rect 12038 12423 12072 12461
rect 12554 12423 12588 12461
rect 13070 12423 13104 12461
rect 13586 12423 13620 12461
rect 14102 12423 14136 12461
rect 14618 12423 14652 12461
rect 15134 12423 15168 12461
rect 15650 12423 15684 12461
rect 16166 12423 16200 12461
rect 16682 12423 16716 12461
rect 17048 12423 17094 12505
rect 11660 12383 17094 12423
rect 11660 12349 11700 12383
rect 17054 12349 17094 12383
rect 11660 12310 17094 12349
rect 11660 12240 11690 12310
rect 11760 12240 11810 12310
rect 11880 12240 12020 12310
rect 12090 12240 12140 12310
rect 12210 12240 12350 12310
rect 12420 12240 12470 12310
rect 12540 12240 12680 12310
rect 12750 12240 12800 12310
rect 12870 12240 13010 12310
rect 13080 12240 13130 12310
rect 13200 12240 13340 12310
rect 13410 12240 13460 12310
rect 13530 12240 13670 12310
rect 13740 12240 13790 12310
rect 13860 12240 14000 12310
rect 14070 12240 14120 12310
rect 14190 12240 14330 12310
rect 14400 12240 14450 12310
rect 14520 12300 15650 12310
rect 14520 12240 14660 12300
rect 11660 12230 14660 12240
rect 14730 12230 14780 12300
rect 14850 12230 14990 12300
rect 15060 12230 15110 12300
rect 15180 12230 15320 12300
rect 15390 12230 15440 12300
rect 15510 12240 15650 12300
rect 15720 12240 15770 12310
rect 15840 12240 15980 12310
rect 16050 12240 16100 12310
rect 16170 12240 16310 12310
rect 16380 12240 16430 12310
rect 16500 12240 16640 12310
rect 16710 12240 16760 12310
rect 16830 12240 17094 12310
rect 15510 12230 17094 12240
rect 11660 12190 17094 12230
rect 11660 12120 11690 12190
rect 11760 12120 11810 12190
rect 11880 12120 12020 12190
rect 12090 12120 12140 12190
rect 12210 12120 12350 12190
rect 12420 12120 12470 12190
rect 12540 12120 12680 12190
rect 12750 12120 12800 12190
rect 12870 12120 13010 12190
rect 13080 12120 13130 12190
rect 13200 12120 13340 12190
rect 13410 12120 13460 12190
rect 13530 12120 13670 12190
rect 13740 12120 13790 12190
rect 13860 12120 14000 12190
rect 14070 12120 14120 12190
rect 14190 12120 14330 12190
rect 14400 12120 14450 12190
rect 14520 12180 15650 12190
rect 14520 12120 14660 12180
rect 11660 12110 14660 12120
rect 14730 12110 14780 12180
rect 14850 12110 14990 12180
rect 15060 12110 15110 12180
rect 15180 12110 15320 12180
rect 15390 12110 15440 12180
rect 15510 12120 15650 12180
rect 15720 12120 15770 12190
rect 15840 12120 15980 12190
rect 16050 12120 16100 12190
rect 16170 12120 16310 12190
rect 16380 12120 16430 12190
rect 16500 12120 16640 12190
rect 16710 12120 16760 12190
rect 16830 12130 17094 12190
rect 18866 13479 18912 13491
rect 18866 12505 18872 13479
rect 18906 12505 18912 13479
rect 18866 12423 18912 12505
rect 18980 13449 19026 13600
rect 19078 13533 19186 13539
rect 19078 13499 19090 13533
rect 19174 13499 19186 13533
rect 19078 13493 19186 13499
rect 19336 13533 19444 13539
rect 19336 13499 19348 13533
rect 19432 13499 19444 13533
rect 19336 13493 19444 13499
rect 18980 12473 18986 13449
rect 19020 12473 19026 13449
rect 18980 12461 19026 12473
rect 19238 13449 19284 13461
rect 19238 12473 19244 13449
rect 19278 12473 19284 13449
rect 19238 12461 19284 12473
rect 19496 13449 19542 13600
rect 19594 13533 19702 13539
rect 19594 13499 19606 13533
rect 19690 13499 19702 13533
rect 19594 13493 19702 13499
rect 19852 13533 19960 13539
rect 19852 13499 19864 13533
rect 19948 13499 19960 13533
rect 19852 13493 19960 13499
rect 19496 12473 19502 13449
rect 19536 12473 19542 13449
rect 19496 12461 19542 12473
rect 19754 13449 19800 13461
rect 19754 12473 19760 13449
rect 19794 12473 19800 13449
rect 19754 12461 19800 12473
rect 20012 13449 20058 13600
rect 20110 13533 20218 13539
rect 20110 13499 20122 13533
rect 20206 13499 20218 13533
rect 20110 13493 20218 13499
rect 20368 13533 20476 13539
rect 20368 13499 20380 13533
rect 20464 13499 20476 13533
rect 20368 13493 20476 13499
rect 20012 12473 20018 13449
rect 20052 12473 20058 13449
rect 20012 12461 20058 12473
rect 20270 13449 20316 13461
rect 20270 12473 20276 13449
rect 20310 12473 20316 13449
rect 20270 12461 20316 12473
rect 20528 13449 20574 13600
rect 20626 13533 20734 13539
rect 20626 13499 20638 13533
rect 20722 13499 20734 13533
rect 20626 13493 20734 13499
rect 20884 13533 20992 13539
rect 20884 13499 20896 13533
rect 20980 13499 20992 13533
rect 20884 13493 20992 13499
rect 20528 12473 20534 13449
rect 20568 12473 20574 13449
rect 20528 12461 20574 12473
rect 20786 13449 20832 13461
rect 20786 12473 20792 13449
rect 20826 12473 20832 13449
rect 20786 12461 20832 12473
rect 21044 13449 21090 13600
rect 21142 13533 21250 13539
rect 21142 13499 21154 13533
rect 21238 13499 21250 13533
rect 21142 13493 21250 13499
rect 21400 13533 21508 13539
rect 21400 13499 21412 13533
rect 21496 13499 21508 13533
rect 21400 13493 21508 13499
rect 21044 12473 21050 13449
rect 21084 12473 21090 13449
rect 21044 12461 21090 12473
rect 21302 13449 21348 13461
rect 21302 12473 21308 13449
rect 21342 12473 21348 13449
rect 21302 12461 21348 12473
rect 21560 13449 21606 13600
rect 21658 13533 21766 13539
rect 21658 13499 21670 13533
rect 21754 13499 21766 13533
rect 21658 13493 21766 13499
rect 21916 13533 22024 13539
rect 21916 13499 21928 13533
rect 22012 13499 22024 13533
rect 21916 13493 22024 13499
rect 21560 12473 21566 13449
rect 21600 12473 21606 13449
rect 21560 12461 21606 12473
rect 21818 13449 21864 13461
rect 21818 12473 21824 13449
rect 21858 12473 21864 13449
rect 21818 12461 21864 12473
rect 22076 13449 22122 13600
rect 22174 13533 22282 13539
rect 22174 13499 22186 13533
rect 22270 13499 22282 13533
rect 22174 13493 22282 13499
rect 22432 13533 22540 13539
rect 22432 13499 22444 13533
rect 22528 13499 22540 13533
rect 22432 13493 22540 13499
rect 22076 12473 22082 13449
rect 22116 12473 22122 13449
rect 22076 12461 22122 12473
rect 22334 13449 22380 13461
rect 22334 12473 22340 13449
rect 22374 12473 22380 13449
rect 22334 12461 22380 12473
rect 22592 13449 22638 13600
rect 22690 13533 22798 13539
rect 22690 13499 22702 13533
rect 22786 13499 22798 13533
rect 22690 13493 22798 13499
rect 22948 13533 23056 13539
rect 22948 13499 22960 13533
rect 23044 13499 23056 13533
rect 22948 13493 23056 13499
rect 22592 12473 22598 13449
rect 22632 12473 22638 13449
rect 22592 12461 22638 12473
rect 22850 13449 22896 13461
rect 22850 12473 22856 13449
rect 22890 12473 22896 13449
rect 22850 12461 22896 12473
rect 23108 13449 23154 13600
rect 23206 13533 23314 13539
rect 23206 13499 23218 13533
rect 23302 13499 23314 13533
rect 23206 13493 23314 13499
rect 23464 13533 23572 13539
rect 23464 13499 23476 13533
rect 23560 13499 23572 13533
rect 23464 13493 23572 13499
rect 23108 12473 23114 13449
rect 23148 12473 23154 13449
rect 23108 12461 23154 12473
rect 23366 13449 23412 13461
rect 23366 12473 23372 13449
rect 23406 12473 23412 13449
rect 23366 12461 23412 12473
rect 23624 13449 23670 13600
rect 23722 13533 23830 13539
rect 23722 13499 23734 13533
rect 23818 13499 23830 13533
rect 23722 13493 23830 13499
rect 23980 13533 24088 13539
rect 23980 13499 23992 13533
rect 24076 13499 24088 13533
rect 23980 13493 24088 13499
rect 23624 12473 23630 13449
rect 23664 12473 23670 13449
rect 23624 12461 23670 12473
rect 23882 13449 23928 13461
rect 23882 12473 23888 13449
rect 23922 12473 23928 13449
rect 23882 12461 23928 12473
rect 24140 13449 24186 13600
rect 24140 12473 24146 13449
rect 24180 12473 24186 13449
rect 24140 12461 24186 12473
rect 24254 13479 24300 13491
rect 24254 12505 24260 13479
rect 24294 12505 24300 13479
rect 19244 12423 19278 12461
rect 19760 12423 19794 12461
rect 20276 12423 20310 12461
rect 20792 12423 20826 12461
rect 21308 12423 21342 12461
rect 21824 12423 21858 12461
rect 22340 12423 22374 12461
rect 22856 12423 22890 12461
rect 23372 12423 23406 12461
rect 23888 12423 23922 12461
rect 24254 12423 24300 12505
rect 18866 12383 24300 12423
rect 18866 12349 18906 12383
rect 24260 12349 24300 12383
rect 18866 12310 24300 12349
rect 18866 12240 19130 12310
rect 19200 12240 19250 12310
rect 19320 12240 19460 12310
rect 19530 12240 19580 12310
rect 19650 12240 19790 12310
rect 19860 12240 19910 12310
rect 19980 12240 20120 12310
rect 20190 12240 20240 12310
rect 20310 12300 21440 12310
rect 20310 12240 20450 12300
rect 18866 12230 20450 12240
rect 20520 12230 20570 12300
rect 20640 12230 20780 12300
rect 20850 12230 20900 12300
rect 20970 12230 21110 12300
rect 21180 12230 21230 12300
rect 21300 12240 21440 12300
rect 21510 12240 21560 12310
rect 21630 12240 21770 12310
rect 21840 12240 21890 12310
rect 21960 12240 22100 12310
rect 22170 12240 22220 12310
rect 22290 12240 22430 12310
rect 22500 12240 22550 12310
rect 22620 12240 22760 12310
rect 22830 12240 22880 12310
rect 22950 12240 23090 12310
rect 23160 12240 23210 12310
rect 23280 12240 23420 12310
rect 23490 12240 23540 12310
rect 23610 12240 23750 12310
rect 23820 12240 23870 12310
rect 23940 12240 24080 12310
rect 24150 12240 24200 12310
rect 24270 12240 24300 12310
rect 21300 12230 24300 12240
rect 18866 12190 24300 12230
rect 18866 12130 19130 12190
rect 16830 12120 17090 12130
rect 15510 12110 17090 12120
rect 11660 12090 17090 12110
rect 18870 12120 19130 12130
rect 19200 12120 19250 12190
rect 19320 12120 19460 12190
rect 19530 12120 19580 12190
rect 19650 12120 19790 12190
rect 19860 12120 19910 12190
rect 19980 12120 20120 12190
rect 20190 12120 20240 12190
rect 20310 12180 21440 12190
rect 20310 12120 20450 12180
rect 18870 12110 20450 12120
rect 20520 12110 20570 12180
rect 20640 12110 20780 12180
rect 20850 12110 20900 12180
rect 20970 12110 21110 12180
rect 21180 12110 21230 12180
rect 21300 12120 21440 12180
rect 21510 12120 21560 12190
rect 21630 12120 21770 12190
rect 21840 12120 21890 12190
rect 21960 12120 22100 12190
rect 22170 12120 22220 12190
rect 22290 12120 22430 12190
rect 22500 12120 22550 12190
rect 22620 12120 22760 12190
rect 22830 12120 22880 12190
rect 22950 12120 23090 12190
rect 23160 12120 23210 12190
rect 23280 12120 23420 12190
rect 23490 12120 23540 12190
rect 23610 12120 23750 12190
rect 23820 12120 23870 12190
rect 23940 12120 24080 12190
rect 24150 12120 24200 12190
rect 24270 12120 24300 12190
rect 21300 12110 24300 12120
rect 18870 12090 24300 12110
rect 11690 12070 11930 12090
rect 12020 12070 12260 12090
rect 12350 12070 12590 12090
rect 12680 12070 12920 12090
rect 13010 12070 13250 12090
rect 13340 12070 13580 12090
rect 13670 12070 13910 12090
rect 14000 12070 14240 12090
rect 14330 12070 14570 12090
rect 14660 12070 14900 12090
rect 14990 12070 15230 12090
rect 15320 12070 15560 12090
rect 15650 12070 15890 12090
rect 15980 12070 16220 12090
rect 16310 12070 16550 12090
rect 16640 12070 16880 12090
rect 19080 12070 19320 12090
rect 19410 12070 19650 12090
rect 19740 12070 19980 12090
rect 20070 12070 20310 12090
rect 20400 12070 20640 12090
rect 20730 12070 20970 12090
rect 21060 12070 21300 12090
rect 21390 12070 21630 12090
rect 21720 12070 21960 12090
rect 22050 12070 22290 12090
rect 22380 12070 22620 12090
rect 22710 12070 22950 12090
rect 23040 12070 23280 12090
rect 23370 12070 23610 12090
rect 23700 12070 23940 12090
rect 24030 12070 24270 12090
<< via1 >>
rect 11690 17490 11760 17560
rect 11810 17490 11880 17560
rect 12020 17490 12090 17560
rect 12140 17490 12210 17560
rect 12350 17490 12420 17560
rect 12470 17490 12540 17560
rect 12680 17490 12750 17560
rect 12800 17490 12870 17560
rect 13010 17490 13080 17560
rect 13130 17490 13200 17560
rect 13340 17490 13410 17560
rect 13460 17490 13530 17560
rect 13670 17490 13740 17560
rect 13790 17490 13860 17560
rect 14000 17490 14070 17560
rect 14120 17490 14190 17560
rect 14330 17490 14400 17560
rect 14450 17490 14520 17560
rect 14660 17500 14730 17570
rect 14780 17500 14850 17570
rect 14990 17500 15060 17570
rect 15110 17500 15180 17570
rect 15320 17500 15390 17570
rect 15440 17500 15510 17570
rect 15650 17490 15720 17560
rect 15770 17490 15840 17560
rect 15980 17490 16050 17560
rect 16100 17490 16170 17560
rect 16310 17490 16380 17560
rect 16430 17490 16500 17560
rect 16640 17490 16710 17560
rect 16760 17490 16830 17560
rect 11690 17370 11760 17440
rect 11810 17370 11880 17440
rect 12020 17370 12090 17440
rect 12140 17370 12210 17440
rect 12350 17370 12420 17440
rect 12470 17370 12540 17440
rect 12680 17370 12750 17440
rect 12800 17370 12870 17440
rect 13010 17370 13080 17440
rect 13130 17370 13200 17440
rect 13340 17370 13410 17440
rect 13460 17370 13530 17440
rect 13670 17370 13740 17440
rect 13790 17370 13860 17440
rect 14000 17370 14070 17440
rect 14120 17370 14190 17440
rect 14330 17370 14400 17440
rect 14450 17370 14520 17440
rect 14660 17380 14730 17450
rect 14780 17380 14850 17450
rect 14990 17380 15060 17450
rect 15110 17380 15180 17450
rect 15320 17380 15390 17450
rect 15440 17380 15510 17450
rect 15650 17370 15720 17440
rect 15770 17370 15840 17440
rect 15980 17370 16050 17440
rect 16100 17370 16170 17440
rect 16310 17370 16380 17440
rect 16430 17370 16500 17440
rect 16640 17370 16710 17440
rect 16760 17370 16830 17440
rect 19130 17490 19200 17560
rect 19250 17490 19320 17560
rect 19460 17490 19530 17560
rect 19580 17490 19650 17560
rect 19790 17490 19860 17560
rect 19910 17490 19980 17560
rect 20120 17490 20190 17560
rect 20240 17490 20310 17560
rect 20450 17500 20520 17570
rect 20570 17500 20640 17570
rect 20780 17500 20850 17570
rect 20900 17500 20970 17570
rect 21110 17500 21180 17570
rect 21230 17500 21300 17570
rect 21440 17490 21510 17560
rect 21560 17490 21630 17560
rect 21770 17490 21840 17560
rect 21890 17490 21960 17560
rect 22100 17490 22170 17560
rect 22220 17490 22290 17560
rect 22430 17490 22500 17560
rect 22550 17490 22620 17560
rect 22760 17490 22830 17560
rect 22880 17490 22950 17560
rect 23090 17490 23160 17560
rect 23210 17490 23280 17560
rect 23420 17490 23490 17560
rect 23540 17490 23610 17560
rect 23750 17490 23820 17560
rect 23870 17490 23940 17560
rect 24080 17490 24150 17560
rect 24200 17490 24270 17560
rect 19130 17370 19200 17440
rect 19250 17370 19320 17440
rect 19460 17370 19530 17440
rect 19580 17370 19650 17440
rect 19790 17370 19860 17440
rect 19910 17370 19980 17440
rect 20120 17370 20190 17440
rect 20240 17370 20310 17440
rect 20450 17380 20520 17450
rect 20570 17380 20640 17450
rect 20780 17380 20850 17450
rect 20900 17380 20970 17450
rect 21110 17380 21180 17450
rect 21230 17380 21300 17450
rect 21440 17370 21510 17440
rect 21560 17370 21630 17440
rect 21770 17370 21840 17440
rect 21890 17370 21960 17440
rect 22100 17370 22170 17440
rect 22220 17370 22290 17440
rect 22430 17370 22500 17440
rect 22550 17370 22620 17440
rect 22760 17370 22830 17440
rect 22880 17370 22950 17440
rect 23090 17370 23160 17440
rect 23210 17370 23280 17440
rect 23420 17370 23490 17440
rect 23540 17370 23610 17440
rect 23750 17370 23820 17440
rect 23870 17370 23940 17440
rect 24080 17370 24150 17440
rect 24200 17370 24270 17440
rect 11650 15930 11710 15990
rect 11740 15930 11800 15990
rect 11830 15930 11890 15990
rect 11920 15930 11980 15990
rect 12010 15930 12070 15990
rect 12100 15930 12160 15990
rect 12190 15930 12250 15990
rect 12280 15930 12340 15990
rect 12370 15930 12430 15990
rect 12460 15930 12520 15990
rect 12550 15930 12610 15990
rect 12640 15930 12700 15990
rect 12730 15930 12790 15990
rect 12820 15930 12880 15990
rect 12910 15930 12970 15990
rect 13000 15930 13060 15990
rect 13090 15930 13150 15990
rect 13180 15930 13240 15990
rect 13270 15930 13330 15990
rect 13360 15930 13420 15990
rect 13450 15930 13510 15990
rect 13540 15930 13600 15990
rect 13630 15930 13690 15990
rect 13720 15930 13780 15990
rect 13810 15930 13870 15990
rect 13900 15930 13960 15990
rect 13990 15930 14050 15990
rect 14080 15930 14140 15990
rect 14170 15930 14230 15990
rect 14260 15930 14320 15990
rect 14350 15930 14410 15990
rect 14440 15930 14500 15990
rect 14530 15930 14590 15990
rect 14620 15930 14680 15990
rect 14710 15930 14770 15990
rect 14800 15930 14860 15990
rect 14890 15930 14950 15990
rect 14980 15930 15040 15990
rect 15070 15930 15130 15990
rect 15160 15930 15220 15990
rect 15250 15930 15310 15990
rect 15340 15930 15400 15990
rect 15430 15930 15490 15990
rect 15520 15930 15580 15990
rect 15610 15930 15670 15990
rect 15700 15930 15760 15990
rect 15790 15930 15850 15990
rect 15880 15930 15940 15990
rect 15970 15930 16030 15990
rect 16060 15930 16120 15990
rect 16150 15930 16210 15990
rect 16240 15930 16300 15990
rect 16330 15930 16390 15990
rect 16420 15930 16480 15990
rect 16510 15930 16570 15990
rect 16600 15930 16660 15990
rect 16690 15930 16750 15990
rect 16780 15930 16840 15990
rect 16870 15930 16930 15990
rect 16960 15930 17020 15990
rect 17050 15930 17110 15990
rect 17740 15980 17810 16070
rect 17840 15980 17910 16070
rect 17940 15980 18010 16070
rect 18040 15980 18110 16070
rect 18140 15980 18210 16070
rect 11650 15840 11710 15900
rect 11740 15840 11800 15900
rect 11830 15840 11890 15900
rect 11920 15840 11980 15900
rect 12010 15840 12070 15900
rect 12100 15840 12160 15900
rect 12190 15840 12250 15900
rect 12280 15840 12340 15900
rect 12370 15840 12430 15900
rect 12460 15840 12520 15900
rect 12550 15840 12610 15900
rect 12640 15840 12700 15900
rect 12730 15840 12790 15900
rect 12820 15840 12880 15900
rect 12910 15840 12970 15900
rect 13000 15840 13060 15900
rect 13090 15840 13150 15900
rect 13180 15840 13240 15900
rect 13270 15840 13330 15900
rect 13360 15840 13420 15900
rect 13450 15840 13510 15900
rect 13540 15840 13600 15900
rect 13630 15840 13690 15900
rect 13720 15840 13780 15900
rect 13810 15840 13870 15900
rect 13900 15840 13960 15900
rect 13990 15840 14050 15900
rect 14080 15840 14140 15900
rect 14170 15840 14230 15900
rect 14260 15840 14320 15900
rect 14350 15840 14410 15900
rect 14440 15840 14500 15900
rect 14530 15840 14590 15900
rect 14620 15840 14680 15900
rect 14710 15840 14770 15900
rect 14800 15840 14860 15900
rect 14890 15840 14950 15900
rect 14980 15840 15040 15900
rect 15070 15840 15130 15900
rect 15160 15840 15220 15900
rect 15250 15840 15310 15900
rect 15340 15840 15400 15900
rect 15430 15840 15490 15900
rect 15520 15840 15580 15900
rect 15610 15840 15670 15900
rect 15700 15840 15760 15900
rect 15790 15840 15850 15900
rect 15880 15840 15940 15900
rect 15970 15840 16030 15900
rect 16060 15840 16120 15900
rect 16150 15840 16210 15900
rect 16240 15840 16300 15900
rect 16330 15840 16390 15900
rect 16420 15840 16480 15900
rect 16510 15840 16570 15900
rect 16600 15840 16660 15900
rect 16690 15840 16750 15900
rect 16780 15840 16840 15900
rect 16870 15840 16930 15900
rect 16960 15840 17020 15900
rect 17050 15840 17110 15900
rect 17740 15850 17810 15940
rect 17840 15850 17910 15940
rect 17940 15850 18010 15940
rect 18040 15850 18110 15940
rect 18140 15850 18210 15940
rect 19030 15930 19090 15990
rect 19120 15930 19180 15990
rect 19210 15930 19270 15990
rect 19300 15930 19360 15990
rect 19390 15930 19450 15990
rect 19480 15930 19540 15990
rect 19570 15930 19630 15990
rect 19660 15930 19720 15990
rect 19750 15930 19810 15990
rect 19840 15930 19900 15990
rect 19930 15930 19990 15990
rect 20020 15930 20080 15990
rect 20110 15930 20170 15990
rect 20200 15930 20260 15990
rect 20290 15930 20350 15990
rect 20380 15930 20440 15990
rect 20470 15930 20530 15990
rect 20560 15930 20620 15990
rect 20650 15930 20710 15990
rect 20740 15930 20800 15990
rect 20830 15930 20890 15990
rect 20920 15930 20980 15990
rect 21010 15930 21070 15990
rect 21100 15930 21160 15990
rect 21190 15930 21250 15990
rect 21280 15930 21340 15990
rect 21370 15930 21430 15990
rect 21460 15930 21520 15990
rect 21550 15930 21610 15990
rect 21640 15930 21700 15990
rect 21730 15930 21790 15990
rect 21820 15930 21880 15990
rect 21910 15930 21970 15990
rect 22000 15930 22060 15990
rect 22090 15930 22150 15990
rect 22180 15930 22240 15990
rect 22270 15930 22330 15990
rect 22360 15930 22420 15990
rect 22450 15930 22510 15990
rect 22540 15930 22600 15990
rect 22630 15930 22690 15990
rect 22720 15930 22780 15990
rect 22810 15930 22870 15990
rect 22900 15930 22960 15990
rect 22990 15930 23050 15990
rect 23080 15930 23140 15990
rect 23170 15930 23230 15990
rect 23260 15930 23320 15990
rect 23350 15930 23410 15990
rect 23440 15930 23500 15990
rect 23530 15930 23590 15990
rect 23620 15930 23680 15990
rect 23710 15930 23770 15990
rect 23800 15930 23860 15990
rect 23890 15930 23950 15990
rect 23980 15930 24040 15990
rect 24070 15930 24130 15990
rect 24160 15930 24220 15990
rect 24250 15930 24310 15990
rect 19030 15840 19090 15900
rect 19120 15840 19180 15900
rect 19210 15840 19270 15900
rect 19300 15840 19360 15900
rect 19390 15840 19450 15900
rect 19480 15840 19540 15900
rect 19570 15840 19630 15900
rect 19660 15840 19720 15900
rect 19750 15840 19810 15900
rect 19840 15840 19900 15900
rect 19930 15840 19990 15900
rect 20020 15840 20080 15900
rect 20110 15840 20170 15900
rect 20200 15840 20260 15900
rect 20290 15840 20350 15900
rect 20380 15840 20440 15900
rect 20470 15840 20530 15900
rect 20560 15840 20620 15900
rect 20650 15840 20710 15900
rect 20740 15840 20800 15900
rect 20830 15840 20890 15900
rect 20920 15840 20980 15900
rect 21010 15840 21070 15900
rect 21100 15840 21160 15900
rect 21190 15840 21250 15900
rect 21280 15840 21340 15900
rect 21370 15840 21430 15900
rect 21460 15840 21520 15900
rect 21550 15840 21610 15900
rect 21640 15840 21700 15900
rect 21730 15840 21790 15900
rect 21820 15840 21880 15900
rect 21910 15840 21970 15900
rect 22000 15840 22060 15900
rect 22090 15840 22150 15900
rect 22180 15840 22240 15900
rect 22270 15840 22330 15900
rect 22360 15840 22420 15900
rect 22450 15840 22510 15900
rect 22540 15840 22600 15900
rect 22630 15840 22690 15900
rect 22720 15840 22780 15900
rect 22810 15840 22870 15900
rect 22900 15840 22960 15900
rect 22990 15840 23050 15900
rect 23080 15840 23140 15900
rect 23170 15840 23230 15900
rect 23260 15840 23320 15900
rect 23350 15840 23410 15900
rect 23440 15840 23500 15900
rect 23530 15840 23590 15900
rect 23620 15840 23680 15900
rect 23710 15840 23770 15900
rect 23800 15840 23860 15900
rect 23890 15840 23950 15900
rect 23980 15840 24040 15900
rect 24070 15840 24130 15900
rect 24160 15840 24220 15900
rect 24250 15840 24310 15900
rect 11650 13800 11710 13860
rect 11740 13800 11800 13860
rect 11830 13800 11890 13860
rect 11920 13800 11980 13860
rect 12010 13800 12070 13860
rect 12100 13800 12160 13860
rect 12190 13800 12250 13860
rect 12280 13800 12340 13860
rect 12370 13800 12430 13860
rect 12460 13800 12520 13860
rect 12550 13800 12610 13860
rect 12640 13800 12700 13860
rect 12730 13800 12790 13860
rect 12820 13800 12880 13860
rect 12910 13800 12970 13860
rect 13000 13800 13060 13860
rect 13090 13800 13150 13860
rect 13180 13800 13240 13860
rect 13270 13800 13330 13860
rect 13360 13800 13420 13860
rect 13450 13800 13510 13860
rect 13540 13800 13600 13860
rect 13630 13800 13690 13860
rect 13720 13800 13780 13860
rect 13810 13800 13870 13860
rect 13900 13800 13960 13860
rect 13990 13800 14050 13860
rect 14080 13800 14140 13860
rect 14170 13800 14230 13860
rect 14260 13800 14320 13860
rect 14350 13800 14410 13860
rect 14440 13800 14500 13860
rect 14530 13800 14590 13860
rect 14620 13800 14680 13860
rect 14710 13800 14770 13860
rect 14800 13800 14860 13860
rect 14890 13800 14950 13860
rect 14980 13800 15040 13860
rect 15070 13800 15130 13860
rect 15160 13800 15220 13860
rect 15250 13800 15310 13860
rect 15340 13800 15400 13860
rect 15430 13800 15490 13860
rect 15520 13800 15580 13860
rect 15610 13800 15670 13860
rect 15700 13800 15760 13860
rect 15790 13800 15850 13860
rect 15880 13800 15940 13860
rect 15970 13800 16030 13860
rect 16060 13800 16120 13860
rect 16150 13800 16210 13860
rect 16240 13800 16300 13860
rect 16330 13800 16390 13860
rect 16420 13800 16480 13860
rect 16510 13800 16570 13860
rect 16600 13800 16660 13860
rect 16690 13800 16750 13860
rect 16780 13800 16840 13860
rect 16870 13800 16930 13860
rect 11650 13710 11710 13770
rect 11740 13710 11800 13770
rect 11830 13710 11890 13770
rect 11920 13710 11980 13770
rect 12010 13710 12070 13770
rect 12100 13710 12160 13770
rect 12190 13710 12250 13770
rect 12280 13710 12340 13770
rect 12370 13710 12430 13770
rect 12460 13710 12520 13770
rect 12550 13710 12610 13770
rect 12640 13710 12700 13770
rect 12730 13710 12790 13770
rect 12820 13710 12880 13770
rect 12910 13710 12970 13770
rect 13000 13710 13060 13770
rect 13090 13710 13150 13770
rect 13180 13710 13240 13770
rect 13270 13710 13330 13770
rect 13360 13710 13420 13770
rect 13450 13710 13510 13770
rect 13540 13710 13600 13770
rect 13630 13710 13690 13770
rect 13720 13710 13780 13770
rect 13810 13710 13870 13770
rect 13900 13710 13960 13770
rect 13990 13710 14050 13770
rect 14080 13710 14140 13770
rect 14170 13710 14230 13770
rect 14260 13710 14320 13770
rect 14350 13710 14410 13770
rect 14440 13710 14500 13770
rect 14530 13710 14590 13770
rect 14620 13710 14680 13770
rect 14710 13710 14770 13770
rect 14800 13710 14860 13770
rect 14890 13710 14950 13770
rect 14980 13710 15040 13770
rect 15070 13710 15130 13770
rect 15160 13710 15220 13770
rect 15250 13710 15310 13770
rect 15340 13710 15400 13770
rect 15430 13710 15490 13770
rect 15520 13710 15580 13770
rect 15610 13710 15670 13770
rect 15700 13710 15760 13770
rect 15790 13710 15850 13770
rect 15880 13710 15940 13770
rect 15970 13710 16030 13770
rect 16060 13710 16120 13770
rect 16150 13710 16210 13770
rect 16240 13710 16300 13770
rect 16330 13710 16390 13770
rect 16420 13710 16480 13770
rect 16510 13710 16570 13770
rect 16600 13710 16660 13770
rect 16690 13710 16750 13770
rect 16780 13710 16840 13770
rect 16870 13710 16930 13770
rect 17740 13760 17810 13850
rect 17840 13760 17910 13850
rect 17940 13760 18010 13850
rect 18040 13760 18110 13850
rect 18140 13760 18210 13850
rect 18850 13800 18910 13860
rect 18940 13800 19000 13860
rect 19030 13800 19090 13860
rect 19120 13800 19180 13860
rect 19210 13800 19270 13860
rect 19300 13800 19360 13860
rect 19390 13800 19450 13860
rect 19480 13800 19540 13860
rect 19570 13800 19630 13860
rect 19660 13800 19720 13860
rect 19750 13800 19810 13860
rect 19840 13800 19900 13860
rect 19930 13800 19990 13860
rect 20020 13800 20080 13860
rect 20110 13800 20170 13860
rect 20200 13800 20260 13860
rect 20290 13800 20350 13860
rect 20380 13800 20440 13860
rect 20470 13800 20530 13860
rect 20560 13800 20620 13860
rect 20650 13800 20710 13860
rect 20740 13800 20800 13860
rect 20830 13800 20890 13860
rect 20920 13800 20980 13860
rect 21010 13800 21070 13860
rect 21100 13800 21160 13860
rect 21190 13800 21250 13860
rect 21280 13800 21340 13860
rect 21370 13800 21430 13860
rect 21460 13800 21520 13860
rect 21550 13800 21610 13860
rect 21640 13800 21700 13860
rect 21730 13800 21790 13860
rect 21820 13800 21880 13860
rect 21910 13800 21970 13860
rect 22000 13800 22060 13860
rect 22090 13800 22150 13860
rect 22180 13800 22240 13860
rect 22270 13800 22330 13860
rect 22360 13800 22420 13860
rect 22450 13800 22510 13860
rect 22540 13800 22600 13860
rect 22630 13800 22690 13860
rect 22720 13800 22780 13860
rect 22810 13800 22870 13860
rect 22900 13800 22960 13860
rect 22990 13800 23050 13860
rect 23080 13800 23140 13860
rect 23170 13800 23230 13860
rect 23260 13800 23320 13860
rect 23350 13800 23410 13860
rect 23440 13800 23500 13860
rect 23530 13800 23590 13860
rect 23620 13800 23680 13860
rect 23710 13800 23770 13860
rect 23800 13800 23860 13860
rect 23890 13800 23950 13860
rect 23980 13800 24040 13860
rect 24070 13800 24130 13860
rect 24160 13800 24220 13860
rect 24250 13800 24310 13860
rect 17740 13630 17810 13720
rect 17840 13630 17910 13720
rect 17940 13630 18010 13720
rect 18040 13630 18110 13720
rect 18140 13630 18210 13720
rect 18850 13710 18910 13770
rect 18940 13710 19000 13770
rect 19030 13710 19090 13770
rect 19120 13710 19180 13770
rect 19210 13710 19270 13770
rect 19300 13710 19360 13770
rect 19390 13710 19450 13770
rect 19480 13710 19540 13770
rect 19570 13710 19630 13770
rect 19660 13710 19720 13770
rect 19750 13710 19810 13770
rect 19840 13710 19900 13770
rect 19930 13710 19990 13770
rect 20020 13710 20080 13770
rect 20110 13710 20170 13770
rect 20200 13710 20260 13770
rect 20290 13710 20350 13770
rect 20380 13710 20440 13770
rect 20470 13710 20530 13770
rect 20560 13710 20620 13770
rect 20650 13710 20710 13770
rect 20740 13710 20800 13770
rect 20830 13710 20890 13770
rect 20920 13710 20980 13770
rect 21010 13710 21070 13770
rect 21100 13710 21160 13770
rect 21190 13710 21250 13770
rect 21280 13710 21340 13770
rect 21370 13710 21430 13770
rect 21460 13710 21520 13770
rect 21550 13710 21610 13770
rect 21640 13710 21700 13770
rect 21730 13710 21790 13770
rect 21820 13710 21880 13770
rect 21910 13710 21970 13770
rect 22000 13710 22060 13770
rect 22090 13710 22150 13770
rect 22180 13710 22240 13770
rect 22270 13710 22330 13770
rect 22360 13710 22420 13770
rect 22450 13710 22510 13770
rect 22540 13710 22600 13770
rect 22630 13710 22690 13770
rect 22720 13710 22780 13770
rect 22810 13710 22870 13770
rect 22900 13710 22960 13770
rect 22990 13710 23050 13770
rect 23080 13710 23140 13770
rect 23170 13710 23230 13770
rect 23260 13710 23320 13770
rect 23350 13710 23410 13770
rect 23440 13710 23500 13770
rect 23530 13710 23590 13770
rect 23620 13710 23680 13770
rect 23710 13710 23770 13770
rect 23800 13710 23860 13770
rect 23890 13710 23950 13770
rect 23980 13710 24040 13770
rect 24070 13710 24130 13770
rect 24160 13710 24220 13770
rect 24250 13710 24310 13770
rect 11690 12240 11760 12310
rect 11810 12240 11880 12310
rect 12020 12240 12090 12310
rect 12140 12240 12210 12310
rect 12350 12240 12420 12310
rect 12470 12240 12540 12310
rect 12680 12240 12750 12310
rect 12800 12240 12870 12310
rect 13010 12240 13080 12310
rect 13130 12240 13200 12310
rect 13340 12240 13410 12310
rect 13460 12240 13530 12310
rect 13670 12240 13740 12310
rect 13790 12240 13860 12310
rect 14000 12240 14070 12310
rect 14120 12240 14190 12310
rect 14330 12240 14400 12310
rect 14450 12240 14520 12310
rect 14660 12230 14730 12300
rect 14780 12230 14850 12300
rect 14990 12230 15060 12300
rect 15110 12230 15180 12300
rect 15320 12230 15390 12300
rect 15440 12230 15510 12300
rect 15650 12240 15720 12310
rect 15770 12240 15840 12310
rect 15980 12240 16050 12310
rect 16100 12240 16170 12310
rect 16310 12240 16380 12310
rect 16430 12240 16500 12310
rect 16640 12240 16710 12310
rect 16760 12240 16830 12310
rect 11690 12120 11760 12190
rect 11810 12120 11880 12190
rect 12020 12120 12090 12190
rect 12140 12120 12210 12190
rect 12350 12120 12420 12190
rect 12470 12120 12540 12190
rect 12680 12120 12750 12190
rect 12800 12120 12870 12190
rect 13010 12120 13080 12190
rect 13130 12120 13200 12190
rect 13340 12120 13410 12190
rect 13460 12120 13530 12190
rect 13670 12120 13740 12190
rect 13790 12120 13860 12190
rect 14000 12120 14070 12190
rect 14120 12120 14190 12190
rect 14330 12120 14400 12190
rect 14450 12120 14520 12190
rect 14660 12110 14730 12180
rect 14780 12110 14850 12180
rect 14990 12110 15060 12180
rect 15110 12110 15180 12180
rect 15320 12110 15390 12180
rect 15440 12110 15510 12180
rect 15650 12120 15720 12190
rect 15770 12120 15840 12190
rect 15980 12120 16050 12190
rect 16100 12120 16170 12190
rect 16310 12120 16380 12190
rect 16430 12120 16500 12190
rect 16640 12120 16710 12190
rect 16760 12120 16830 12190
rect 19130 12240 19200 12310
rect 19250 12240 19320 12310
rect 19460 12240 19530 12310
rect 19580 12240 19650 12310
rect 19790 12240 19860 12310
rect 19910 12240 19980 12310
rect 20120 12240 20190 12310
rect 20240 12240 20310 12310
rect 20450 12230 20520 12300
rect 20570 12230 20640 12300
rect 20780 12230 20850 12300
rect 20900 12230 20970 12300
rect 21110 12230 21180 12300
rect 21230 12230 21300 12300
rect 21440 12240 21510 12310
rect 21560 12240 21630 12310
rect 21770 12240 21840 12310
rect 21890 12240 21960 12310
rect 22100 12240 22170 12310
rect 22220 12240 22290 12310
rect 22430 12240 22500 12310
rect 22550 12240 22620 12310
rect 22760 12240 22830 12310
rect 22880 12240 22950 12310
rect 23090 12240 23160 12310
rect 23210 12240 23280 12310
rect 23420 12240 23490 12310
rect 23540 12240 23610 12310
rect 23750 12240 23820 12310
rect 23870 12240 23940 12310
rect 24080 12240 24150 12310
rect 24200 12240 24270 12310
rect 19130 12120 19200 12190
rect 19250 12120 19320 12190
rect 19460 12120 19530 12190
rect 19580 12120 19650 12190
rect 19790 12120 19860 12190
rect 19910 12120 19980 12190
rect 20120 12120 20190 12190
rect 20240 12120 20310 12190
rect 20450 12110 20520 12180
rect 20570 12110 20640 12180
rect 20780 12110 20850 12180
rect 20900 12110 20970 12180
rect 21110 12110 21180 12180
rect 21230 12110 21300 12180
rect 21440 12120 21510 12190
rect 21560 12120 21630 12190
rect 21770 12120 21840 12190
rect 21890 12120 21960 12190
rect 22100 12120 22170 12190
rect 22220 12120 22290 12190
rect 22430 12120 22500 12190
rect 22550 12120 22620 12190
rect 22760 12120 22830 12190
rect 22880 12120 22950 12190
rect 23090 12120 23160 12190
rect 23210 12120 23280 12190
rect 23420 12120 23490 12190
rect 23540 12120 23610 12190
rect 23750 12120 23820 12190
rect 23870 12120 23940 12190
rect 24080 12120 24150 12190
rect 24200 12120 24270 12190
<< metal2 >>
rect 11690 17590 11930 17610
rect 12020 17590 12260 17610
rect 12350 17590 12590 17610
rect 12680 17590 12920 17610
rect 13010 17590 13250 17610
rect 13340 17590 13580 17610
rect 13670 17590 13910 17610
rect 14000 17590 14240 17610
rect 14330 17590 14570 17610
rect 14660 17590 14900 17610
rect 14990 17590 15230 17610
rect 15320 17590 15560 17610
rect 15650 17590 15890 17610
rect 15980 17590 16220 17610
rect 16310 17590 16550 17610
rect 16640 17590 16880 17610
rect 19080 17590 19320 17610
rect 19410 17590 19650 17610
rect 19740 17590 19980 17610
rect 20070 17590 20310 17610
rect 20400 17590 20640 17610
rect 20730 17590 20970 17610
rect 21060 17590 21300 17610
rect 21390 17590 21630 17610
rect 21720 17590 21960 17610
rect 22050 17590 22290 17610
rect 22380 17590 22620 17610
rect 22710 17590 22950 17610
rect 23040 17590 23280 17610
rect 23370 17590 23610 17610
rect 23700 17590 23940 17610
rect 24030 17590 24270 17610
rect 11660 17570 17090 17590
rect 11660 17560 14660 17570
rect 11660 17490 11690 17560
rect 11760 17490 11810 17560
rect 11880 17490 12020 17560
rect 12090 17490 12140 17560
rect 12210 17490 12350 17560
rect 12420 17490 12470 17560
rect 12540 17490 12680 17560
rect 12750 17490 12800 17560
rect 12870 17490 13010 17560
rect 13080 17490 13130 17560
rect 13200 17490 13340 17560
rect 13410 17490 13460 17560
rect 13530 17490 13670 17560
rect 13740 17490 13790 17560
rect 13860 17490 14000 17560
rect 14070 17490 14120 17560
rect 14190 17490 14330 17560
rect 14400 17490 14450 17560
rect 14520 17500 14660 17560
rect 14730 17500 14780 17570
rect 14850 17500 14990 17570
rect 15060 17500 15110 17570
rect 15180 17500 15320 17570
rect 15390 17500 15440 17570
rect 15510 17560 17090 17570
rect 15510 17500 15650 17560
rect 14520 17490 15650 17500
rect 15720 17490 15770 17560
rect 15840 17490 15980 17560
rect 16050 17490 16100 17560
rect 16170 17490 16310 17560
rect 16380 17490 16430 17560
rect 16500 17490 16640 17560
rect 16710 17490 16760 17560
rect 16830 17490 17090 17560
rect 11660 17450 17090 17490
rect 11660 17440 14660 17450
rect 11660 17370 11690 17440
rect 11760 17370 11810 17440
rect 11880 17370 12020 17440
rect 12090 17370 12140 17440
rect 12210 17370 12350 17440
rect 12420 17370 12470 17440
rect 12540 17370 12680 17440
rect 12750 17370 12800 17440
rect 12870 17370 13010 17440
rect 13080 17370 13130 17440
rect 13200 17370 13340 17440
rect 13410 17370 13460 17440
rect 13530 17370 13670 17440
rect 13740 17370 13790 17440
rect 13860 17370 14000 17440
rect 14070 17370 14120 17440
rect 14190 17370 14330 17440
rect 14400 17370 14450 17440
rect 14520 17380 14660 17440
rect 14730 17380 14780 17450
rect 14850 17380 14990 17450
rect 15060 17380 15110 17450
rect 15180 17380 15320 17450
rect 15390 17380 15440 17450
rect 15510 17440 17090 17450
rect 15510 17380 15650 17440
rect 14520 17370 15650 17380
rect 15720 17370 15770 17440
rect 15840 17370 15980 17440
rect 16050 17370 16100 17440
rect 16170 17370 16310 17440
rect 16380 17370 16430 17440
rect 16500 17370 16640 17440
rect 16710 17370 16760 17440
rect 16830 17370 17090 17440
rect 11660 17340 17090 17370
rect 18870 17570 24300 17590
rect 18870 17560 20450 17570
rect 18870 17490 19130 17560
rect 19200 17490 19250 17560
rect 19320 17490 19460 17560
rect 19530 17490 19580 17560
rect 19650 17490 19790 17560
rect 19860 17490 19910 17560
rect 19980 17490 20120 17560
rect 20190 17490 20240 17560
rect 20310 17500 20450 17560
rect 20520 17500 20570 17570
rect 20640 17500 20780 17570
rect 20850 17500 20900 17570
rect 20970 17500 21110 17570
rect 21180 17500 21230 17570
rect 21300 17560 24300 17570
rect 21300 17500 21440 17560
rect 20310 17490 21440 17500
rect 21510 17490 21560 17560
rect 21630 17490 21770 17560
rect 21840 17490 21890 17560
rect 21960 17490 22100 17560
rect 22170 17490 22220 17560
rect 22290 17490 22430 17560
rect 22500 17490 22550 17560
rect 22620 17490 22760 17560
rect 22830 17490 22880 17560
rect 22950 17490 23090 17560
rect 23160 17490 23210 17560
rect 23280 17490 23420 17560
rect 23490 17490 23540 17560
rect 23610 17490 23750 17560
rect 23820 17490 23870 17560
rect 23940 17490 24080 17560
rect 24150 17490 24200 17560
rect 24270 17490 24300 17560
rect 18870 17450 24300 17490
rect 18870 17440 20450 17450
rect 18870 17370 19130 17440
rect 19200 17370 19250 17440
rect 19320 17370 19460 17440
rect 19530 17370 19580 17440
rect 19650 17370 19790 17440
rect 19860 17370 19910 17440
rect 19980 17370 20120 17440
rect 20190 17370 20240 17440
rect 20310 17380 20450 17440
rect 20520 17380 20570 17450
rect 20640 17380 20780 17450
rect 20850 17380 20900 17450
rect 20970 17380 21110 17450
rect 21180 17380 21230 17450
rect 21300 17440 24300 17450
rect 21300 17380 21440 17440
rect 20310 17370 21440 17380
rect 21510 17370 21560 17440
rect 21630 17370 21770 17440
rect 21840 17370 21890 17440
rect 21960 17370 22100 17440
rect 22170 17370 22220 17440
rect 22290 17370 22430 17440
rect 22500 17370 22550 17440
rect 22620 17370 22760 17440
rect 22830 17370 22880 17440
rect 22950 17370 23090 17440
rect 23160 17370 23210 17440
rect 23280 17370 23420 17440
rect 23490 17370 23540 17440
rect 23610 17370 23750 17440
rect 23820 17370 23870 17440
rect 23940 17370 24080 17440
rect 24150 17370 24200 17440
rect 24270 17370 24300 17440
rect 18870 17340 24300 17370
rect 17690 16070 18260 16100
rect 17690 16000 17740 16070
rect 11630 15990 17740 16000
rect 11630 15930 11650 15990
rect 11710 15930 11740 15990
rect 11800 15930 11830 15990
rect 11890 15930 11920 15990
rect 11980 15930 12010 15990
rect 12070 15930 12100 15990
rect 12160 15930 12190 15990
rect 12250 15930 12280 15990
rect 12340 15930 12370 15990
rect 12430 15930 12460 15990
rect 12520 15930 12550 15990
rect 12610 15930 12640 15990
rect 12700 15930 12730 15990
rect 12790 15930 12820 15990
rect 12880 15930 12910 15990
rect 12970 15930 13000 15990
rect 13060 15930 13090 15990
rect 13150 15930 13180 15990
rect 13240 15930 13270 15990
rect 13330 15930 13360 15990
rect 13420 15930 13450 15990
rect 13510 15930 13540 15990
rect 13600 15930 13630 15990
rect 13690 15930 13720 15990
rect 13780 15930 13810 15990
rect 13870 15930 13900 15990
rect 13960 15930 13990 15990
rect 14050 15930 14080 15990
rect 14140 15930 14170 15990
rect 14230 15930 14260 15990
rect 14320 15930 14350 15990
rect 14410 15930 14440 15990
rect 14500 15930 14530 15990
rect 14590 15930 14620 15990
rect 14680 15930 14710 15990
rect 14770 15930 14800 15990
rect 14860 15930 14890 15990
rect 14950 15930 14980 15990
rect 15040 15930 15070 15990
rect 15130 15930 15160 15990
rect 15220 15930 15250 15990
rect 15310 15930 15340 15990
rect 15400 15930 15430 15990
rect 15490 15930 15520 15990
rect 15580 15930 15610 15990
rect 15670 15930 15700 15990
rect 15760 15930 15790 15990
rect 15850 15930 15880 15990
rect 15940 15930 15970 15990
rect 16030 15930 16060 15990
rect 16120 15930 16150 15990
rect 16210 15930 16240 15990
rect 16300 15930 16330 15990
rect 16390 15930 16420 15990
rect 16480 15930 16510 15990
rect 16570 15930 16600 15990
rect 16660 15930 16690 15990
rect 16750 15930 16780 15990
rect 16840 15930 16870 15990
rect 16930 15930 16960 15990
rect 17020 15930 17050 15990
rect 17110 15980 17740 15990
rect 17810 15980 17840 16070
rect 17910 15980 17940 16070
rect 18010 15980 18040 16070
rect 18110 15980 18140 16070
rect 18210 15980 18260 16070
rect 17110 15940 18260 15980
rect 17110 15930 17740 15940
rect 11630 15900 17740 15930
rect 11630 15840 11650 15900
rect 11710 15840 11740 15900
rect 11800 15840 11830 15900
rect 11890 15840 11920 15900
rect 11980 15840 12010 15900
rect 12070 15840 12100 15900
rect 12160 15840 12190 15900
rect 12250 15840 12280 15900
rect 12340 15840 12370 15900
rect 12430 15840 12460 15900
rect 12520 15840 12550 15900
rect 12610 15840 12640 15900
rect 12700 15840 12730 15900
rect 12790 15840 12820 15900
rect 12880 15840 12910 15900
rect 12970 15840 13000 15900
rect 13060 15840 13090 15900
rect 13150 15840 13180 15900
rect 13240 15840 13270 15900
rect 13330 15840 13360 15900
rect 13420 15840 13450 15900
rect 13510 15840 13540 15900
rect 13600 15840 13630 15900
rect 13690 15840 13720 15900
rect 13780 15840 13810 15900
rect 13870 15840 13900 15900
rect 13960 15840 13990 15900
rect 14050 15840 14080 15900
rect 14140 15840 14170 15900
rect 14230 15840 14260 15900
rect 14320 15840 14350 15900
rect 14410 15840 14440 15900
rect 14500 15840 14530 15900
rect 14590 15840 14620 15900
rect 14680 15840 14710 15900
rect 14770 15840 14800 15900
rect 14860 15840 14890 15900
rect 14950 15840 14980 15900
rect 15040 15840 15070 15900
rect 15130 15840 15160 15900
rect 15220 15840 15250 15900
rect 15310 15840 15340 15900
rect 15400 15840 15430 15900
rect 15490 15840 15520 15900
rect 15580 15840 15610 15900
rect 15670 15840 15700 15900
rect 15760 15840 15790 15900
rect 15850 15840 15880 15900
rect 15940 15840 15970 15900
rect 16030 15840 16060 15900
rect 16120 15840 16150 15900
rect 16210 15840 16240 15900
rect 16300 15840 16330 15900
rect 16390 15840 16420 15900
rect 16480 15840 16510 15900
rect 16570 15840 16600 15900
rect 16660 15840 16690 15900
rect 16750 15840 16780 15900
rect 16840 15840 16870 15900
rect 16930 15840 16960 15900
rect 17020 15840 17050 15900
rect 17110 15850 17740 15900
rect 17810 15850 17840 15940
rect 17910 15850 17940 15940
rect 18010 15850 18040 15940
rect 18110 15850 18140 15940
rect 18210 15850 18260 15940
rect 17110 15840 18260 15850
rect 11630 15820 18260 15840
rect 18980 15990 24330 16000
rect 18980 15930 19030 15990
rect 19090 15930 19120 15990
rect 19180 15930 19210 15990
rect 19270 15930 19300 15990
rect 19360 15930 19390 15990
rect 19450 15930 19480 15990
rect 19540 15930 19570 15990
rect 19630 15930 19660 15990
rect 19720 15930 19750 15990
rect 19810 15930 19840 15990
rect 19900 15930 19930 15990
rect 19990 15930 20020 15990
rect 20080 15930 20110 15990
rect 20170 15930 20200 15990
rect 20260 15930 20290 15990
rect 20350 15930 20380 15990
rect 20440 15930 20470 15990
rect 20530 15930 20560 15990
rect 20620 15930 20650 15990
rect 20710 15930 20740 15990
rect 20800 15930 20830 15990
rect 20890 15930 20920 15990
rect 20980 15930 21010 15990
rect 21070 15930 21100 15990
rect 21160 15930 21190 15990
rect 21250 15930 21280 15990
rect 21340 15930 21370 15990
rect 21430 15930 21460 15990
rect 21520 15930 21550 15990
rect 21610 15930 21640 15990
rect 21700 15930 21730 15990
rect 21790 15930 21820 15990
rect 21880 15930 21910 15990
rect 21970 15930 22000 15990
rect 22060 15930 22090 15990
rect 22150 15930 22180 15990
rect 22240 15930 22270 15990
rect 22330 15930 22360 15990
rect 22420 15930 22450 15990
rect 22510 15930 22540 15990
rect 22600 15930 22630 15990
rect 22690 15930 22720 15990
rect 22780 15930 22810 15990
rect 22870 15930 22900 15990
rect 22960 15930 22990 15990
rect 23050 15930 23080 15990
rect 23140 15930 23170 15990
rect 23230 15930 23260 15990
rect 23320 15930 23350 15990
rect 23410 15930 23440 15990
rect 23500 15930 23530 15990
rect 23590 15930 23620 15990
rect 23680 15930 23710 15990
rect 23770 15930 23800 15990
rect 23860 15930 23890 15990
rect 23950 15930 23980 15990
rect 24040 15930 24070 15990
rect 24130 15930 24160 15990
rect 24220 15930 24250 15990
rect 24310 15930 24330 15990
rect 18980 15900 24330 15930
rect 18980 15840 19030 15900
rect 19090 15840 19120 15900
rect 19180 15840 19210 15900
rect 19270 15840 19300 15900
rect 19360 15840 19390 15900
rect 19450 15840 19480 15900
rect 19540 15840 19570 15900
rect 19630 15840 19660 15900
rect 19720 15840 19750 15900
rect 19810 15840 19840 15900
rect 19900 15840 19930 15900
rect 19990 15840 20020 15900
rect 20080 15840 20110 15900
rect 20170 15840 20200 15900
rect 20260 15840 20290 15900
rect 20350 15840 20380 15900
rect 20440 15840 20470 15900
rect 20530 15840 20560 15900
rect 20620 15840 20650 15900
rect 20710 15840 20740 15900
rect 20800 15840 20830 15900
rect 20890 15840 20920 15900
rect 20980 15840 21010 15900
rect 21070 15840 21100 15900
rect 21160 15840 21190 15900
rect 21250 15840 21280 15900
rect 21340 15840 21370 15900
rect 21430 15840 21460 15900
rect 21520 15840 21550 15900
rect 21610 15840 21640 15900
rect 21700 15840 21730 15900
rect 21790 15840 21820 15900
rect 21880 15840 21910 15900
rect 21970 15840 22000 15900
rect 22060 15840 22090 15900
rect 22150 15840 22180 15900
rect 22240 15840 22270 15900
rect 22330 15840 22360 15900
rect 22420 15840 22450 15900
rect 22510 15840 22540 15900
rect 22600 15840 22630 15900
rect 22690 15840 22720 15900
rect 22780 15840 22810 15900
rect 22870 15840 22900 15900
rect 22960 15840 22990 15900
rect 23050 15840 23080 15900
rect 23140 15840 23170 15900
rect 23230 15840 23260 15900
rect 23320 15840 23350 15900
rect 23410 15840 23440 15900
rect 23500 15840 23530 15900
rect 23590 15840 23620 15900
rect 23680 15840 23710 15900
rect 23770 15840 23800 15900
rect 23860 15840 23890 15900
rect 23950 15840 23980 15900
rect 24040 15840 24070 15900
rect 24130 15840 24160 15900
rect 24220 15840 24250 15900
rect 24310 15840 24330 15900
rect 18980 15820 24330 15840
rect 11630 13860 16980 13880
rect 11630 13800 11650 13860
rect 11710 13800 11740 13860
rect 11800 13800 11830 13860
rect 11890 13800 11920 13860
rect 11980 13800 12010 13860
rect 12070 13800 12100 13860
rect 12160 13800 12190 13860
rect 12250 13800 12280 13860
rect 12340 13800 12370 13860
rect 12430 13800 12460 13860
rect 12520 13800 12550 13860
rect 12610 13800 12640 13860
rect 12700 13800 12730 13860
rect 12790 13800 12820 13860
rect 12880 13800 12910 13860
rect 12970 13800 13000 13860
rect 13060 13800 13090 13860
rect 13150 13800 13180 13860
rect 13240 13800 13270 13860
rect 13330 13800 13360 13860
rect 13420 13800 13450 13860
rect 13510 13800 13540 13860
rect 13600 13800 13630 13860
rect 13690 13800 13720 13860
rect 13780 13800 13810 13860
rect 13870 13800 13900 13860
rect 13960 13800 13990 13860
rect 14050 13800 14080 13860
rect 14140 13800 14170 13860
rect 14230 13800 14260 13860
rect 14320 13800 14350 13860
rect 14410 13800 14440 13860
rect 14500 13800 14530 13860
rect 14590 13800 14620 13860
rect 14680 13800 14710 13860
rect 14770 13800 14800 13860
rect 14860 13800 14890 13860
rect 14950 13800 14980 13860
rect 15040 13800 15070 13860
rect 15130 13800 15160 13860
rect 15220 13800 15250 13860
rect 15310 13800 15340 13860
rect 15400 13800 15430 13860
rect 15490 13800 15520 13860
rect 15580 13800 15610 13860
rect 15670 13800 15700 13860
rect 15760 13800 15790 13860
rect 15850 13800 15880 13860
rect 15940 13800 15970 13860
rect 16030 13800 16060 13860
rect 16120 13800 16150 13860
rect 16210 13800 16240 13860
rect 16300 13800 16330 13860
rect 16390 13800 16420 13860
rect 16480 13800 16510 13860
rect 16570 13800 16600 13860
rect 16660 13800 16690 13860
rect 16750 13800 16780 13860
rect 16840 13800 16870 13860
rect 16930 13800 16980 13860
rect 11630 13770 16980 13800
rect 11630 13710 11650 13770
rect 11710 13710 11740 13770
rect 11800 13710 11830 13770
rect 11890 13710 11920 13770
rect 11980 13710 12010 13770
rect 12070 13710 12100 13770
rect 12160 13710 12190 13770
rect 12250 13710 12280 13770
rect 12340 13710 12370 13770
rect 12430 13710 12460 13770
rect 12520 13710 12550 13770
rect 12610 13710 12640 13770
rect 12700 13710 12730 13770
rect 12790 13710 12820 13770
rect 12880 13710 12910 13770
rect 12970 13710 13000 13770
rect 13060 13710 13090 13770
rect 13150 13710 13180 13770
rect 13240 13710 13270 13770
rect 13330 13710 13360 13770
rect 13420 13710 13450 13770
rect 13510 13710 13540 13770
rect 13600 13710 13630 13770
rect 13690 13710 13720 13770
rect 13780 13710 13810 13770
rect 13870 13710 13900 13770
rect 13960 13710 13990 13770
rect 14050 13710 14080 13770
rect 14140 13710 14170 13770
rect 14230 13710 14260 13770
rect 14320 13710 14350 13770
rect 14410 13710 14440 13770
rect 14500 13710 14530 13770
rect 14590 13710 14620 13770
rect 14680 13710 14710 13770
rect 14770 13710 14800 13770
rect 14860 13710 14890 13770
rect 14950 13710 14980 13770
rect 15040 13710 15070 13770
rect 15130 13710 15160 13770
rect 15220 13710 15250 13770
rect 15310 13710 15340 13770
rect 15400 13710 15430 13770
rect 15490 13710 15520 13770
rect 15580 13710 15610 13770
rect 15670 13710 15700 13770
rect 15760 13710 15790 13770
rect 15850 13710 15880 13770
rect 15940 13710 15970 13770
rect 16030 13710 16060 13770
rect 16120 13710 16150 13770
rect 16210 13710 16240 13770
rect 16300 13710 16330 13770
rect 16390 13710 16420 13770
rect 16480 13710 16510 13770
rect 16570 13710 16600 13770
rect 16660 13710 16690 13770
rect 16750 13710 16780 13770
rect 16840 13710 16870 13770
rect 16930 13710 16980 13770
rect 11630 13700 16980 13710
rect 17690 13860 24330 13880
rect 17690 13850 18850 13860
rect 17690 13760 17740 13850
rect 17810 13760 17840 13850
rect 17910 13760 17940 13850
rect 18010 13760 18040 13850
rect 18110 13760 18140 13850
rect 18210 13800 18850 13850
rect 18910 13800 18940 13860
rect 19000 13800 19030 13860
rect 19090 13800 19120 13860
rect 19180 13800 19210 13860
rect 19270 13800 19300 13860
rect 19360 13800 19390 13860
rect 19450 13800 19480 13860
rect 19540 13800 19570 13860
rect 19630 13800 19660 13860
rect 19720 13800 19750 13860
rect 19810 13800 19840 13860
rect 19900 13800 19930 13860
rect 19990 13800 20020 13860
rect 20080 13800 20110 13860
rect 20170 13800 20200 13860
rect 20260 13800 20290 13860
rect 20350 13800 20380 13860
rect 20440 13800 20470 13860
rect 20530 13800 20560 13860
rect 20620 13800 20650 13860
rect 20710 13800 20740 13860
rect 20800 13800 20830 13860
rect 20890 13800 20920 13860
rect 20980 13800 21010 13860
rect 21070 13800 21100 13860
rect 21160 13800 21190 13860
rect 21250 13800 21280 13860
rect 21340 13800 21370 13860
rect 21430 13800 21460 13860
rect 21520 13800 21550 13860
rect 21610 13800 21640 13860
rect 21700 13800 21730 13860
rect 21790 13800 21820 13860
rect 21880 13800 21910 13860
rect 21970 13800 22000 13860
rect 22060 13800 22090 13860
rect 22150 13800 22180 13860
rect 22240 13800 22270 13860
rect 22330 13800 22360 13860
rect 22420 13800 22450 13860
rect 22510 13800 22540 13860
rect 22600 13800 22630 13860
rect 22690 13800 22720 13860
rect 22780 13800 22810 13860
rect 22870 13800 22900 13860
rect 22960 13800 22990 13860
rect 23050 13800 23080 13860
rect 23140 13800 23170 13860
rect 23230 13800 23260 13860
rect 23320 13800 23350 13860
rect 23410 13800 23440 13860
rect 23500 13800 23530 13860
rect 23590 13800 23620 13860
rect 23680 13800 23710 13860
rect 23770 13800 23800 13860
rect 23860 13800 23890 13860
rect 23950 13800 23980 13860
rect 24040 13800 24070 13860
rect 24130 13800 24160 13860
rect 24220 13800 24250 13860
rect 24310 13800 24330 13860
rect 18210 13770 24330 13800
rect 18210 13760 18850 13770
rect 17690 13720 18850 13760
rect 17690 13630 17740 13720
rect 17810 13630 17840 13720
rect 17910 13630 17940 13720
rect 18010 13630 18040 13720
rect 18110 13630 18140 13720
rect 18210 13710 18850 13720
rect 18910 13710 18940 13770
rect 19000 13710 19030 13770
rect 19090 13710 19120 13770
rect 19180 13710 19210 13770
rect 19270 13710 19300 13770
rect 19360 13710 19390 13770
rect 19450 13710 19480 13770
rect 19540 13710 19570 13770
rect 19630 13710 19660 13770
rect 19720 13710 19750 13770
rect 19810 13710 19840 13770
rect 19900 13710 19930 13770
rect 19990 13710 20020 13770
rect 20080 13710 20110 13770
rect 20170 13710 20200 13770
rect 20260 13710 20290 13770
rect 20350 13710 20380 13770
rect 20440 13710 20470 13770
rect 20530 13710 20560 13770
rect 20620 13710 20650 13770
rect 20710 13710 20740 13770
rect 20800 13710 20830 13770
rect 20890 13710 20920 13770
rect 20980 13710 21010 13770
rect 21070 13710 21100 13770
rect 21160 13710 21190 13770
rect 21250 13710 21280 13770
rect 21340 13710 21370 13770
rect 21430 13710 21460 13770
rect 21520 13710 21550 13770
rect 21610 13710 21640 13770
rect 21700 13710 21730 13770
rect 21790 13710 21820 13770
rect 21880 13710 21910 13770
rect 21970 13710 22000 13770
rect 22060 13710 22090 13770
rect 22150 13710 22180 13770
rect 22240 13710 22270 13770
rect 22330 13710 22360 13770
rect 22420 13710 22450 13770
rect 22510 13710 22540 13770
rect 22600 13710 22630 13770
rect 22690 13710 22720 13770
rect 22780 13710 22810 13770
rect 22870 13710 22900 13770
rect 22960 13710 22990 13770
rect 23050 13710 23080 13770
rect 23140 13710 23170 13770
rect 23230 13710 23260 13770
rect 23320 13710 23350 13770
rect 23410 13710 23440 13770
rect 23500 13710 23530 13770
rect 23590 13710 23620 13770
rect 23680 13710 23710 13770
rect 23770 13710 23800 13770
rect 23860 13710 23890 13770
rect 23950 13710 23980 13770
rect 24040 13710 24070 13770
rect 24130 13710 24160 13770
rect 24220 13710 24250 13770
rect 24310 13710 24330 13770
rect 18210 13700 24330 13710
rect 18210 13630 18260 13700
rect 17690 13600 18260 13630
rect 11660 12310 17090 12340
rect 11660 12240 11690 12310
rect 11760 12240 11810 12310
rect 11880 12240 12020 12310
rect 12090 12240 12140 12310
rect 12210 12240 12350 12310
rect 12420 12240 12470 12310
rect 12540 12240 12680 12310
rect 12750 12240 12800 12310
rect 12870 12240 13010 12310
rect 13080 12240 13130 12310
rect 13200 12240 13340 12310
rect 13410 12240 13460 12310
rect 13530 12240 13670 12310
rect 13740 12240 13790 12310
rect 13860 12240 14000 12310
rect 14070 12240 14120 12310
rect 14190 12240 14330 12310
rect 14400 12240 14450 12310
rect 14520 12300 15650 12310
rect 14520 12240 14660 12300
rect 11660 12230 14660 12240
rect 14730 12230 14780 12300
rect 14850 12230 14990 12300
rect 15060 12230 15110 12300
rect 15180 12230 15320 12300
rect 15390 12230 15440 12300
rect 15510 12240 15650 12300
rect 15720 12240 15770 12310
rect 15840 12240 15980 12310
rect 16050 12240 16100 12310
rect 16170 12240 16310 12310
rect 16380 12240 16430 12310
rect 16500 12240 16640 12310
rect 16710 12240 16760 12310
rect 16830 12240 17090 12310
rect 15510 12230 17090 12240
rect 11660 12190 17090 12230
rect 11660 12120 11690 12190
rect 11760 12120 11810 12190
rect 11880 12120 12020 12190
rect 12090 12120 12140 12190
rect 12210 12120 12350 12190
rect 12420 12120 12470 12190
rect 12540 12120 12680 12190
rect 12750 12120 12800 12190
rect 12870 12120 13010 12190
rect 13080 12120 13130 12190
rect 13200 12120 13340 12190
rect 13410 12120 13460 12190
rect 13530 12120 13670 12190
rect 13740 12120 13790 12190
rect 13860 12120 14000 12190
rect 14070 12120 14120 12190
rect 14190 12120 14330 12190
rect 14400 12120 14450 12190
rect 14520 12180 15650 12190
rect 14520 12120 14660 12180
rect 11660 12110 14660 12120
rect 14730 12110 14780 12180
rect 14850 12110 14990 12180
rect 15060 12110 15110 12180
rect 15180 12110 15320 12180
rect 15390 12110 15440 12180
rect 15510 12120 15650 12180
rect 15720 12120 15770 12190
rect 15840 12120 15980 12190
rect 16050 12120 16100 12190
rect 16170 12120 16310 12190
rect 16380 12120 16430 12190
rect 16500 12120 16640 12190
rect 16710 12120 16760 12190
rect 16830 12120 17090 12190
rect 15510 12110 17090 12120
rect 11660 12090 17090 12110
rect 18870 12310 24300 12340
rect 18870 12240 19130 12310
rect 19200 12240 19250 12310
rect 19320 12240 19460 12310
rect 19530 12240 19580 12310
rect 19650 12240 19790 12310
rect 19860 12240 19910 12310
rect 19980 12240 20120 12310
rect 20190 12240 20240 12310
rect 20310 12300 21440 12310
rect 20310 12240 20450 12300
rect 18870 12230 20450 12240
rect 20520 12230 20570 12300
rect 20640 12230 20780 12300
rect 20850 12230 20900 12300
rect 20970 12230 21110 12300
rect 21180 12230 21230 12300
rect 21300 12240 21440 12300
rect 21510 12240 21560 12310
rect 21630 12240 21770 12310
rect 21840 12240 21890 12310
rect 21960 12240 22100 12310
rect 22170 12240 22220 12310
rect 22290 12240 22430 12310
rect 22500 12240 22550 12310
rect 22620 12240 22760 12310
rect 22830 12240 22880 12310
rect 22950 12240 23090 12310
rect 23160 12240 23210 12310
rect 23280 12240 23420 12310
rect 23490 12240 23540 12310
rect 23610 12240 23750 12310
rect 23820 12240 23870 12310
rect 23940 12240 24080 12310
rect 24150 12240 24200 12310
rect 24270 12240 24300 12310
rect 21300 12230 24300 12240
rect 18870 12190 24300 12230
rect 18870 12120 19130 12190
rect 19200 12120 19250 12190
rect 19320 12120 19460 12190
rect 19530 12120 19580 12190
rect 19650 12120 19790 12190
rect 19860 12120 19910 12190
rect 19980 12120 20120 12190
rect 20190 12120 20240 12190
rect 20310 12180 21440 12190
rect 20310 12120 20450 12180
rect 18870 12110 20450 12120
rect 20520 12110 20570 12180
rect 20640 12110 20780 12180
rect 20850 12110 20900 12180
rect 20970 12110 21110 12180
rect 21180 12110 21230 12180
rect 21300 12120 21440 12180
rect 21510 12120 21560 12190
rect 21630 12120 21770 12190
rect 21840 12120 21890 12190
rect 21960 12120 22100 12190
rect 22170 12120 22220 12190
rect 22290 12120 22430 12190
rect 22500 12120 22550 12190
rect 22620 12120 22760 12190
rect 22830 12120 22880 12190
rect 22950 12120 23090 12190
rect 23160 12120 23210 12190
rect 23280 12120 23420 12190
rect 23490 12120 23540 12190
rect 23610 12120 23750 12190
rect 23820 12120 23870 12190
rect 23940 12120 24080 12190
rect 24150 12120 24200 12190
rect 24270 12120 24300 12190
rect 21300 12110 24300 12120
rect 18870 12090 24300 12110
rect 11690 12070 11930 12090
rect 12020 12070 12260 12090
rect 12350 12070 12590 12090
rect 12680 12070 12920 12090
rect 13010 12070 13250 12090
rect 13340 12070 13580 12090
rect 13670 12070 13910 12090
rect 14000 12070 14240 12090
rect 14330 12070 14570 12090
rect 14660 12070 14900 12090
rect 14990 12070 15230 12090
rect 15320 12070 15560 12090
rect 15650 12070 15890 12090
rect 15980 12070 16220 12090
rect 16310 12070 16550 12090
rect 16640 12070 16880 12090
rect 19080 12070 19320 12090
rect 19410 12070 19650 12090
rect 19740 12070 19980 12090
rect 20070 12070 20310 12090
rect 20400 12070 20640 12090
rect 20730 12070 20970 12090
rect 21060 12070 21300 12090
rect 21390 12070 21630 12090
rect 21720 12070 21960 12090
rect 22050 12070 22290 12090
rect 22380 12070 22620 12090
rect 22710 12070 22950 12090
rect 23040 12070 23280 12090
rect 23370 12070 23610 12090
rect 23700 12070 23940 12090
rect 24030 12070 24270 12090
<< via2 >>
rect 11690 17490 11760 17560
rect 11810 17490 11880 17560
rect 12020 17490 12090 17560
rect 12140 17490 12210 17560
rect 12350 17490 12420 17560
rect 12470 17490 12540 17560
rect 12680 17490 12750 17560
rect 12800 17490 12870 17560
rect 13010 17490 13080 17560
rect 13130 17490 13200 17560
rect 13340 17490 13410 17560
rect 13460 17490 13530 17560
rect 13670 17490 13740 17560
rect 13790 17490 13860 17560
rect 14000 17490 14070 17560
rect 14120 17490 14190 17560
rect 14330 17490 14400 17560
rect 14450 17490 14520 17560
rect 14660 17500 14730 17570
rect 14780 17500 14850 17570
rect 14990 17500 15060 17570
rect 15110 17500 15180 17570
rect 15320 17500 15390 17570
rect 15440 17500 15510 17570
rect 15650 17490 15720 17560
rect 15770 17490 15840 17560
rect 15980 17490 16050 17560
rect 16100 17490 16170 17560
rect 16310 17490 16380 17560
rect 16430 17490 16500 17560
rect 16640 17490 16710 17560
rect 16760 17490 16830 17560
rect 11690 17370 11760 17440
rect 11810 17370 11880 17440
rect 12020 17370 12090 17440
rect 12140 17370 12210 17440
rect 12350 17370 12420 17440
rect 12470 17370 12540 17440
rect 12680 17370 12750 17440
rect 12800 17370 12870 17440
rect 13010 17370 13080 17440
rect 13130 17370 13200 17440
rect 13340 17370 13410 17440
rect 13460 17370 13530 17440
rect 13670 17370 13740 17440
rect 13790 17370 13860 17440
rect 14000 17370 14070 17440
rect 14120 17370 14190 17440
rect 14330 17370 14400 17440
rect 14450 17370 14520 17440
rect 14660 17380 14730 17450
rect 14780 17380 14850 17450
rect 14990 17380 15060 17450
rect 15110 17380 15180 17450
rect 15320 17380 15390 17450
rect 15440 17380 15510 17450
rect 15650 17370 15720 17440
rect 15770 17370 15840 17440
rect 15980 17370 16050 17440
rect 16100 17370 16170 17440
rect 16310 17370 16380 17440
rect 16430 17370 16500 17440
rect 16640 17370 16710 17440
rect 16760 17370 16830 17440
rect 19130 17490 19200 17560
rect 19250 17490 19320 17560
rect 19460 17490 19530 17560
rect 19580 17490 19650 17560
rect 19790 17490 19860 17560
rect 19910 17490 19980 17560
rect 20120 17490 20190 17560
rect 20240 17490 20310 17560
rect 20450 17500 20520 17570
rect 20570 17500 20640 17570
rect 20780 17500 20850 17570
rect 20900 17500 20970 17570
rect 21110 17500 21180 17570
rect 21230 17500 21300 17570
rect 21440 17490 21510 17560
rect 21560 17490 21630 17560
rect 21770 17490 21840 17560
rect 21890 17490 21960 17560
rect 22100 17490 22170 17560
rect 22220 17490 22290 17560
rect 22430 17490 22500 17560
rect 22550 17490 22620 17560
rect 22760 17490 22830 17560
rect 22880 17490 22950 17560
rect 23090 17490 23160 17560
rect 23210 17490 23280 17560
rect 23420 17490 23490 17560
rect 23540 17490 23610 17560
rect 23750 17490 23820 17560
rect 23870 17490 23940 17560
rect 24080 17490 24150 17560
rect 24200 17490 24270 17560
rect 19130 17370 19200 17440
rect 19250 17370 19320 17440
rect 19460 17370 19530 17440
rect 19580 17370 19650 17440
rect 19790 17370 19860 17440
rect 19910 17370 19980 17440
rect 20120 17370 20190 17440
rect 20240 17370 20310 17440
rect 20450 17380 20520 17450
rect 20570 17380 20640 17450
rect 20780 17380 20850 17450
rect 20900 17380 20970 17450
rect 21110 17380 21180 17450
rect 21230 17380 21300 17450
rect 21440 17370 21510 17440
rect 21560 17370 21630 17440
rect 21770 17370 21840 17440
rect 21890 17370 21960 17440
rect 22100 17370 22170 17440
rect 22220 17370 22290 17440
rect 22430 17370 22500 17440
rect 22550 17370 22620 17440
rect 22760 17370 22830 17440
rect 22880 17370 22950 17440
rect 23090 17370 23160 17440
rect 23210 17370 23280 17440
rect 23420 17370 23490 17440
rect 23540 17370 23610 17440
rect 23750 17370 23820 17440
rect 23870 17370 23940 17440
rect 24080 17370 24150 17440
rect 24200 17370 24270 17440
rect 11650 15930 11710 15990
rect 11740 15930 11800 15990
rect 11830 15930 11890 15990
rect 11920 15930 11980 15990
rect 12010 15930 12070 15990
rect 12100 15930 12160 15990
rect 12190 15930 12250 15990
rect 12280 15930 12340 15990
rect 12370 15930 12430 15990
rect 12460 15930 12520 15990
rect 12550 15930 12610 15990
rect 12640 15930 12700 15990
rect 12730 15930 12790 15990
rect 12820 15930 12880 15990
rect 12910 15930 12970 15990
rect 13000 15930 13060 15990
rect 13090 15930 13150 15990
rect 13180 15930 13240 15990
rect 13270 15930 13330 15990
rect 13360 15930 13420 15990
rect 13450 15930 13510 15990
rect 13540 15930 13600 15990
rect 13630 15930 13690 15990
rect 13720 15930 13780 15990
rect 13810 15930 13870 15990
rect 13900 15930 13960 15990
rect 13990 15930 14050 15990
rect 14080 15930 14140 15990
rect 14170 15930 14230 15990
rect 14260 15930 14320 15990
rect 14350 15930 14410 15990
rect 14440 15930 14500 15990
rect 14530 15930 14590 15990
rect 14620 15930 14680 15990
rect 14710 15930 14770 15990
rect 14800 15930 14860 15990
rect 14890 15930 14950 15990
rect 14980 15930 15040 15990
rect 15070 15930 15130 15990
rect 15160 15930 15220 15990
rect 15250 15930 15310 15990
rect 15340 15930 15400 15990
rect 15430 15930 15490 15990
rect 15520 15930 15580 15990
rect 15610 15930 15670 15990
rect 15700 15930 15760 15990
rect 15790 15930 15850 15990
rect 15880 15930 15940 15990
rect 15970 15930 16030 15990
rect 16060 15930 16120 15990
rect 16150 15930 16210 15990
rect 16240 15930 16300 15990
rect 16330 15930 16390 15990
rect 16420 15930 16480 15990
rect 16510 15930 16570 15990
rect 16600 15930 16660 15990
rect 16690 15930 16750 15990
rect 16780 15930 16840 15990
rect 16870 15930 16930 15990
rect 16960 15930 17020 15990
rect 17050 15930 17110 15990
rect 17740 15980 17810 16070
rect 17840 15980 17910 16070
rect 17940 15980 18010 16070
rect 18040 15980 18110 16070
rect 18140 15980 18210 16070
rect 11650 15840 11710 15900
rect 11740 15840 11800 15900
rect 11830 15840 11890 15900
rect 11920 15840 11980 15900
rect 12010 15840 12070 15900
rect 12100 15840 12160 15900
rect 12190 15840 12250 15900
rect 12280 15840 12340 15900
rect 12370 15840 12430 15900
rect 12460 15840 12520 15900
rect 12550 15840 12610 15900
rect 12640 15840 12700 15900
rect 12730 15840 12790 15900
rect 12820 15840 12880 15900
rect 12910 15840 12970 15900
rect 13000 15840 13060 15900
rect 13090 15840 13150 15900
rect 13180 15840 13240 15900
rect 13270 15840 13330 15900
rect 13360 15840 13420 15900
rect 13450 15840 13510 15900
rect 13540 15840 13600 15900
rect 13630 15840 13690 15900
rect 13720 15840 13780 15900
rect 13810 15840 13870 15900
rect 13900 15840 13960 15900
rect 13990 15840 14050 15900
rect 14080 15840 14140 15900
rect 14170 15840 14230 15900
rect 14260 15840 14320 15900
rect 14350 15840 14410 15900
rect 14440 15840 14500 15900
rect 14530 15840 14590 15900
rect 14620 15840 14680 15900
rect 14710 15840 14770 15900
rect 14800 15840 14860 15900
rect 14890 15840 14950 15900
rect 14980 15840 15040 15900
rect 15070 15840 15130 15900
rect 15160 15840 15220 15900
rect 15250 15840 15310 15900
rect 15340 15840 15400 15900
rect 15430 15840 15490 15900
rect 15520 15840 15580 15900
rect 15610 15840 15670 15900
rect 15700 15840 15760 15900
rect 15790 15840 15850 15900
rect 15880 15840 15940 15900
rect 15970 15840 16030 15900
rect 16060 15840 16120 15900
rect 16150 15840 16210 15900
rect 16240 15840 16300 15900
rect 16330 15840 16390 15900
rect 16420 15840 16480 15900
rect 16510 15840 16570 15900
rect 16600 15840 16660 15900
rect 16690 15840 16750 15900
rect 16780 15840 16840 15900
rect 16870 15840 16930 15900
rect 16960 15840 17020 15900
rect 17050 15840 17110 15900
rect 17740 15850 17810 15940
rect 17840 15850 17910 15940
rect 17940 15850 18010 15940
rect 18040 15850 18110 15940
rect 18140 15850 18210 15940
rect 19030 15930 19090 15990
rect 19120 15930 19180 15990
rect 19210 15930 19270 15990
rect 19300 15930 19360 15990
rect 19390 15930 19450 15990
rect 19480 15930 19540 15990
rect 19570 15930 19630 15990
rect 19660 15930 19720 15990
rect 19750 15930 19810 15990
rect 19840 15930 19900 15990
rect 19930 15930 19990 15990
rect 20020 15930 20080 15990
rect 20110 15930 20170 15990
rect 20200 15930 20260 15990
rect 20290 15930 20350 15990
rect 20380 15930 20440 15990
rect 20470 15930 20530 15990
rect 20560 15930 20620 15990
rect 20650 15930 20710 15990
rect 20740 15930 20800 15990
rect 20830 15930 20890 15990
rect 20920 15930 20980 15990
rect 21010 15930 21070 15990
rect 21100 15930 21160 15990
rect 21190 15930 21250 15990
rect 21280 15930 21340 15990
rect 21370 15930 21430 15990
rect 21460 15930 21520 15990
rect 21550 15930 21610 15990
rect 21640 15930 21700 15990
rect 21730 15930 21790 15990
rect 21820 15930 21880 15990
rect 21910 15930 21970 15990
rect 22000 15930 22060 15990
rect 22090 15930 22150 15990
rect 22180 15930 22240 15990
rect 22270 15930 22330 15990
rect 22360 15930 22420 15990
rect 22450 15930 22510 15990
rect 22540 15930 22600 15990
rect 22630 15930 22690 15990
rect 22720 15930 22780 15990
rect 22810 15930 22870 15990
rect 22900 15930 22960 15990
rect 22990 15930 23050 15990
rect 23080 15930 23140 15990
rect 23170 15930 23230 15990
rect 23260 15930 23320 15990
rect 23350 15930 23410 15990
rect 23440 15930 23500 15990
rect 23530 15930 23590 15990
rect 23620 15930 23680 15990
rect 23710 15930 23770 15990
rect 23800 15930 23860 15990
rect 23890 15930 23950 15990
rect 23980 15930 24040 15990
rect 24070 15930 24130 15990
rect 24160 15930 24220 15990
rect 24250 15930 24310 15990
rect 19030 15840 19090 15900
rect 19120 15840 19180 15900
rect 19210 15840 19270 15900
rect 19300 15840 19360 15900
rect 19390 15840 19450 15900
rect 19480 15840 19540 15900
rect 19570 15840 19630 15900
rect 19660 15840 19720 15900
rect 19750 15840 19810 15900
rect 19840 15840 19900 15900
rect 19930 15840 19990 15900
rect 20020 15840 20080 15900
rect 20110 15840 20170 15900
rect 20200 15840 20260 15900
rect 20290 15840 20350 15900
rect 20380 15840 20440 15900
rect 20470 15840 20530 15900
rect 20560 15840 20620 15900
rect 20650 15840 20710 15900
rect 20740 15840 20800 15900
rect 20830 15840 20890 15900
rect 20920 15840 20980 15900
rect 21010 15840 21070 15900
rect 21100 15840 21160 15900
rect 21190 15840 21250 15900
rect 21280 15840 21340 15900
rect 21370 15840 21430 15900
rect 21460 15840 21520 15900
rect 21550 15840 21610 15900
rect 21640 15840 21700 15900
rect 21730 15840 21790 15900
rect 21820 15840 21880 15900
rect 21910 15840 21970 15900
rect 22000 15840 22060 15900
rect 22090 15840 22150 15900
rect 22180 15840 22240 15900
rect 22270 15840 22330 15900
rect 22360 15840 22420 15900
rect 22450 15840 22510 15900
rect 22540 15840 22600 15900
rect 22630 15840 22690 15900
rect 22720 15840 22780 15900
rect 22810 15840 22870 15900
rect 22900 15840 22960 15900
rect 22990 15840 23050 15900
rect 23080 15840 23140 15900
rect 23170 15840 23230 15900
rect 23260 15840 23320 15900
rect 23350 15840 23410 15900
rect 23440 15840 23500 15900
rect 23530 15840 23590 15900
rect 23620 15840 23680 15900
rect 23710 15840 23770 15900
rect 23800 15840 23860 15900
rect 23890 15840 23950 15900
rect 23980 15840 24040 15900
rect 24070 15840 24130 15900
rect 24160 15840 24220 15900
rect 24250 15840 24310 15900
rect 11650 13800 11710 13860
rect 11740 13800 11800 13860
rect 11830 13800 11890 13860
rect 11920 13800 11980 13860
rect 12010 13800 12070 13860
rect 12100 13800 12160 13860
rect 12190 13800 12250 13860
rect 12280 13800 12340 13860
rect 12370 13800 12430 13860
rect 12460 13800 12520 13860
rect 12550 13800 12610 13860
rect 12640 13800 12700 13860
rect 12730 13800 12790 13860
rect 12820 13800 12880 13860
rect 12910 13800 12970 13860
rect 13000 13800 13060 13860
rect 13090 13800 13150 13860
rect 13180 13800 13240 13860
rect 13270 13800 13330 13860
rect 13360 13800 13420 13860
rect 13450 13800 13510 13860
rect 13540 13800 13600 13860
rect 13630 13800 13690 13860
rect 13720 13800 13780 13860
rect 13810 13800 13870 13860
rect 13900 13800 13960 13860
rect 13990 13800 14050 13860
rect 14080 13800 14140 13860
rect 14170 13800 14230 13860
rect 14260 13800 14320 13860
rect 14350 13800 14410 13860
rect 14440 13800 14500 13860
rect 14530 13800 14590 13860
rect 14620 13800 14680 13860
rect 14710 13800 14770 13860
rect 14800 13800 14860 13860
rect 14890 13800 14950 13860
rect 14980 13800 15040 13860
rect 15070 13800 15130 13860
rect 15160 13800 15220 13860
rect 15250 13800 15310 13860
rect 15340 13800 15400 13860
rect 15430 13800 15490 13860
rect 15520 13800 15580 13860
rect 15610 13800 15670 13860
rect 15700 13800 15760 13860
rect 15790 13800 15850 13860
rect 15880 13800 15940 13860
rect 15970 13800 16030 13860
rect 16060 13800 16120 13860
rect 16150 13800 16210 13860
rect 16240 13800 16300 13860
rect 16330 13800 16390 13860
rect 16420 13800 16480 13860
rect 16510 13800 16570 13860
rect 16600 13800 16660 13860
rect 16690 13800 16750 13860
rect 16780 13800 16840 13860
rect 16870 13800 16930 13860
rect 11650 13710 11710 13770
rect 11740 13710 11800 13770
rect 11830 13710 11890 13770
rect 11920 13710 11980 13770
rect 12010 13710 12070 13770
rect 12100 13710 12160 13770
rect 12190 13710 12250 13770
rect 12280 13710 12340 13770
rect 12370 13710 12430 13770
rect 12460 13710 12520 13770
rect 12550 13710 12610 13770
rect 12640 13710 12700 13770
rect 12730 13710 12790 13770
rect 12820 13710 12880 13770
rect 12910 13710 12970 13770
rect 13000 13710 13060 13770
rect 13090 13710 13150 13770
rect 13180 13710 13240 13770
rect 13270 13710 13330 13770
rect 13360 13710 13420 13770
rect 13450 13710 13510 13770
rect 13540 13710 13600 13770
rect 13630 13710 13690 13770
rect 13720 13710 13780 13770
rect 13810 13710 13870 13770
rect 13900 13710 13960 13770
rect 13990 13710 14050 13770
rect 14080 13710 14140 13770
rect 14170 13710 14230 13770
rect 14260 13710 14320 13770
rect 14350 13710 14410 13770
rect 14440 13710 14500 13770
rect 14530 13710 14590 13770
rect 14620 13710 14680 13770
rect 14710 13710 14770 13770
rect 14800 13710 14860 13770
rect 14890 13710 14950 13770
rect 14980 13710 15040 13770
rect 15070 13710 15130 13770
rect 15160 13710 15220 13770
rect 15250 13710 15310 13770
rect 15340 13710 15400 13770
rect 15430 13710 15490 13770
rect 15520 13710 15580 13770
rect 15610 13710 15670 13770
rect 15700 13710 15760 13770
rect 15790 13710 15850 13770
rect 15880 13710 15940 13770
rect 15970 13710 16030 13770
rect 16060 13710 16120 13770
rect 16150 13710 16210 13770
rect 16240 13710 16300 13770
rect 16330 13710 16390 13770
rect 16420 13710 16480 13770
rect 16510 13710 16570 13770
rect 16600 13710 16660 13770
rect 16690 13710 16750 13770
rect 16780 13710 16840 13770
rect 16870 13710 16930 13770
rect 17740 13760 17810 13850
rect 17840 13760 17910 13850
rect 17940 13760 18010 13850
rect 18040 13760 18110 13850
rect 18140 13760 18210 13850
rect 18850 13800 18910 13860
rect 18940 13800 19000 13860
rect 19030 13800 19090 13860
rect 19120 13800 19180 13860
rect 19210 13800 19270 13860
rect 19300 13800 19360 13860
rect 19390 13800 19450 13860
rect 19480 13800 19540 13860
rect 19570 13800 19630 13860
rect 19660 13800 19720 13860
rect 19750 13800 19810 13860
rect 19840 13800 19900 13860
rect 19930 13800 19990 13860
rect 20020 13800 20080 13860
rect 20110 13800 20170 13860
rect 20200 13800 20260 13860
rect 20290 13800 20350 13860
rect 20380 13800 20440 13860
rect 20470 13800 20530 13860
rect 20560 13800 20620 13860
rect 20650 13800 20710 13860
rect 20740 13800 20800 13860
rect 20830 13800 20890 13860
rect 20920 13800 20980 13860
rect 21010 13800 21070 13860
rect 21100 13800 21160 13860
rect 21190 13800 21250 13860
rect 21280 13800 21340 13860
rect 21370 13800 21430 13860
rect 21460 13800 21520 13860
rect 21550 13800 21610 13860
rect 21640 13800 21700 13860
rect 21730 13800 21790 13860
rect 21820 13800 21880 13860
rect 21910 13800 21970 13860
rect 22000 13800 22060 13860
rect 22090 13800 22150 13860
rect 22180 13800 22240 13860
rect 22270 13800 22330 13860
rect 22360 13800 22420 13860
rect 22450 13800 22510 13860
rect 22540 13800 22600 13860
rect 22630 13800 22690 13860
rect 22720 13800 22780 13860
rect 22810 13800 22870 13860
rect 22900 13800 22960 13860
rect 22990 13800 23050 13860
rect 23080 13800 23140 13860
rect 23170 13800 23230 13860
rect 23260 13800 23320 13860
rect 23350 13800 23410 13860
rect 23440 13800 23500 13860
rect 23530 13800 23590 13860
rect 23620 13800 23680 13860
rect 23710 13800 23770 13860
rect 23800 13800 23860 13860
rect 23890 13800 23950 13860
rect 23980 13800 24040 13860
rect 24070 13800 24130 13860
rect 24160 13800 24220 13860
rect 24250 13800 24310 13860
rect 17740 13630 17810 13720
rect 17840 13630 17910 13720
rect 17940 13630 18010 13720
rect 18040 13630 18110 13720
rect 18140 13630 18210 13720
rect 18850 13710 18910 13770
rect 18940 13710 19000 13770
rect 19030 13710 19090 13770
rect 19120 13710 19180 13770
rect 19210 13710 19270 13770
rect 19300 13710 19360 13770
rect 19390 13710 19450 13770
rect 19480 13710 19540 13770
rect 19570 13710 19630 13770
rect 19660 13710 19720 13770
rect 19750 13710 19810 13770
rect 19840 13710 19900 13770
rect 19930 13710 19990 13770
rect 20020 13710 20080 13770
rect 20110 13710 20170 13770
rect 20200 13710 20260 13770
rect 20290 13710 20350 13770
rect 20380 13710 20440 13770
rect 20470 13710 20530 13770
rect 20560 13710 20620 13770
rect 20650 13710 20710 13770
rect 20740 13710 20800 13770
rect 20830 13710 20890 13770
rect 20920 13710 20980 13770
rect 21010 13710 21070 13770
rect 21100 13710 21160 13770
rect 21190 13710 21250 13770
rect 21280 13710 21340 13770
rect 21370 13710 21430 13770
rect 21460 13710 21520 13770
rect 21550 13710 21610 13770
rect 21640 13710 21700 13770
rect 21730 13710 21790 13770
rect 21820 13710 21880 13770
rect 21910 13710 21970 13770
rect 22000 13710 22060 13770
rect 22090 13710 22150 13770
rect 22180 13710 22240 13770
rect 22270 13710 22330 13770
rect 22360 13710 22420 13770
rect 22450 13710 22510 13770
rect 22540 13710 22600 13770
rect 22630 13710 22690 13770
rect 22720 13710 22780 13770
rect 22810 13710 22870 13770
rect 22900 13710 22960 13770
rect 22990 13710 23050 13770
rect 23080 13710 23140 13770
rect 23170 13710 23230 13770
rect 23260 13710 23320 13770
rect 23350 13710 23410 13770
rect 23440 13710 23500 13770
rect 23530 13710 23590 13770
rect 23620 13710 23680 13770
rect 23710 13710 23770 13770
rect 23800 13710 23860 13770
rect 23890 13710 23950 13770
rect 23980 13710 24040 13770
rect 24070 13710 24130 13770
rect 24160 13710 24220 13770
rect 24250 13710 24310 13770
rect 11690 12240 11760 12310
rect 11810 12240 11880 12310
rect 12020 12240 12090 12310
rect 12140 12240 12210 12310
rect 12350 12240 12420 12310
rect 12470 12240 12540 12310
rect 12680 12240 12750 12310
rect 12800 12240 12870 12310
rect 13010 12240 13080 12310
rect 13130 12240 13200 12310
rect 13340 12240 13410 12310
rect 13460 12240 13530 12310
rect 13670 12240 13740 12310
rect 13790 12240 13860 12310
rect 14000 12240 14070 12310
rect 14120 12240 14190 12310
rect 14330 12240 14400 12310
rect 14450 12240 14520 12310
rect 14660 12230 14730 12300
rect 14780 12230 14850 12300
rect 14990 12230 15060 12300
rect 15110 12230 15180 12300
rect 15320 12230 15390 12300
rect 15440 12230 15510 12300
rect 15650 12240 15720 12310
rect 15770 12240 15840 12310
rect 15980 12240 16050 12310
rect 16100 12240 16170 12310
rect 16310 12240 16380 12310
rect 16430 12240 16500 12310
rect 16640 12240 16710 12310
rect 16760 12240 16830 12310
rect 11690 12120 11760 12190
rect 11810 12120 11880 12190
rect 12020 12120 12090 12190
rect 12140 12120 12210 12190
rect 12350 12120 12420 12190
rect 12470 12120 12540 12190
rect 12680 12120 12750 12190
rect 12800 12120 12870 12190
rect 13010 12120 13080 12190
rect 13130 12120 13200 12190
rect 13340 12120 13410 12190
rect 13460 12120 13530 12190
rect 13670 12120 13740 12190
rect 13790 12120 13860 12190
rect 14000 12120 14070 12190
rect 14120 12120 14190 12190
rect 14330 12120 14400 12190
rect 14450 12120 14520 12190
rect 14660 12110 14730 12180
rect 14780 12110 14850 12180
rect 14990 12110 15060 12180
rect 15110 12110 15180 12180
rect 15320 12110 15390 12180
rect 15440 12110 15510 12180
rect 15650 12120 15720 12190
rect 15770 12120 15840 12190
rect 15980 12120 16050 12190
rect 16100 12120 16170 12190
rect 16310 12120 16380 12190
rect 16430 12120 16500 12190
rect 16640 12120 16710 12190
rect 16760 12120 16830 12190
rect 19130 12240 19200 12310
rect 19250 12240 19320 12310
rect 19460 12240 19530 12310
rect 19580 12240 19650 12310
rect 19790 12240 19860 12310
rect 19910 12240 19980 12310
rect 20120 12240 20190 12310
rect 20240 12240 20310 12310
rect 20450 12230 20520 12300
rect 20570 12230 20640 12300
rect 20780 12230 20850 12300
rect 20900 12230 20970 12300
rect 21110 12230 21180 12300
rect 21230 12230 21300 12300
rect 21440 12240 21510 12310
rect 21560 12240 21630 12310
rect 21770 12240 21840 12310
rect 21890 12240 21960 12310
rect 22100 12240 22170 12310
rect 22220 12240 22290 12310
rect 22430 12240 22500 12310
rect 22550 12240 22620 12310
rect 22760 12240 22830 12310
rect 22880 12240 22950 12310
rect 23090 12240 23160 12310
rect 23210 12240 23280 12310
rect 23420 12240 23490 12310
rect 23540 12240 23610 12310
rect 23750 12240 23820 12310
rect 23870 12240 23940 12310
rect 24080 12240 24150 12310
rect 24200 12240 24270 12310
rect 19130 12120 19200 12190
rect 19250 12120 19320 12190
rect 19460 12120 19530 12190
rect 19580 12120 19650 12190
rect 19790 12120 19860 12190
rect 19910 12120 19980 12190
rect 20120 12120 20190 12190
rect 20240 12120 20310 12190
rect 20450 12110 20520 12180
rect 20570 12110 20640 12180
rect 20780 12110 20850 12180
rect 20900 12110 20970 12180
rect 21110 12110 21180 12180
rect 21230 12110 21300 12180
rect 21440 12120 21510 12190
rect 21560 12120 21630 12190
rect 21770 12120 21840 12190
rect 21890 12120 21960 12190
rect 22100 12120 22170 12190
rect 22220 12120 22290 12190
rect 22430 12120 22500 12190
rect 22550 12120 22620 12190
rect 22760 12120 22830 12190
rect 22880 12120 22950 12190
rect 23090 12120 23160 12190
rect 23210 12120 23280 12190
rect 23420 12120 23490 12190
rect 23540 12120 23610 12190
rect 23750 12120 23820 12190
rect 23870 12120 23940 12190
rect 24080 12120 24150 12190
rect 24200 12120 24270 12190
<< metal3 >>
rect 11690 17590 11930 17610
rect 12020 17590 12260 17610
rect 12350 17590 12590 17610
rect 12680 17590 12920 17610
rect 13010 17590 13250 17610
rect 13340 17590 13580 17610
rect 13670 17590 13910 17610
rect 14000 17590 14240 17610
rect 14330 17590 14570 17610
rect 14660 17590 14900 17610
rect 14990 17590 15230 17610
rect 15320 17590 15560 17610
rect 15650 17590 15890 17610
rect 15980 17590 16220 17610
rect 16310 17590 16550 17610
rect 16640 17590 16880 17610
rect 19080 17590 19320 17610
rect 19410 17590 19650 17610
rect 19740 17590 19980 17610
rect 20070 17590 20310 17610
rect 20400 17590 20640 17610
rect 20730 17590 20970 17610
rect 21060 17590 21300 17610
rect 21390 17590 21630 17610
rect 21720 17590 21960 17610
rect 22050 17590 22290 17610
rect 22380 17590 22620 17610
rect 22710 17590 22950 17610
rect 23040 17590 23280 17610
rect 23370 17590 23610 17610
rect 23700 17590 23940 17610
rect 24030 17590 24270 17610
rect 11660 17570 17090 17590
rect 11660 17560 14660 17570
rect 11660 17490 11690 17560
rect 11760 17490 11810 17560
rect 11880 17490 12020 17560
rect 12090 17490 12140 17560
rect 12210 17490 12350 17560
rect 12420 17490 12470 17560
rect 12540 17490 12680 17560
rect 12750 17490 12800 17560
rect 12870 17490 13010 17560
rect 13080 17490 13130 17560
rect 13200 17490 13340 17560
rect 13410 17490 13460 17560
rect 13530 17490 13670 17560
rect 13740 17490 13790 17560
rect 13860 17490 14000 17560
rect 14070 17490 14120 17560
rect 14190 17490 14330 17560
rect 14400 17490 14450 17560
rect 14520 17500 14660 17560
rect 14730 17500 14780 17570
rect 14850 17500 14990 17570
rect 15060 17500 15110 17570
rect 15180 17500 15320 17570
rect 15390 17500 15440 17570
rect 15510 17560 17090 17570
rect 15510 17500 15650 17560
rect 14520 17490 15650 17500
rect 15720 17490 15770 17560
rect 15840 17490 15980 17560
rect 16050 17490 16100 17560
rect 16170 17490 16310 17560
rect 16380 17490 16430 17560
rect 16500 17490 16640 17560
rect 16710 17490 16760 17560
rect 16830 17490 17090 17560
rect 11660 17450 17090 17490
rect 11660 17440 14660 17450
rect 11660 17370 11690 17440
rect 11760 17370 11810 17440
rect 11880 17370 12020 17440
rect 12090 17370 12140 17440
rect 12210 17370 12350 17440
rect 12420 17370 12470 17440
rect 12540 17370 12680 17440
rect 12750 17370 12800 17440
rect 12870 17370 13010 17440
rect 13080 17370 13130 17440
rect 13200 17370 13340 17440
rect 13410 17370 13460 17440
rect 13530 17370 13670 17440
rect 13740 17370 13790 17440
rect 13860 17370 14000 17440
rect 14070 17370 14120 17440
rect 14190 17370 14330 17440
rect 14400 17370 14450 17440
rect 14520 17380 14660 17440
rect 14730 17380 14780 17450
rect 14850 17380 14990 17450
rect 15060 17380 15110 17450
rect 15180 17380 15320 17450
rect 15390 17380 15440 17450
rect 15510 17440 17090 17450
rect 15510 17380 15650 17440
rect 14520 17370 15650 17380
rect 15720 17370 15770 17440
rect 15840 17370 15980 17440
rect 16050 17370 16100 17440
rect 16170 17370 16310 17440
rect 16380 17370 16430 17440
rect 16500 17370 16640 17440
rect 16710 17370 16760 17440
rect 16830 17370 17090 17440
rect 11660 17340 17090 17370
rect 18870 17570 24300 17590
rect 18870 17560 20450 17570
rect 18870 17490 19130 17560
rect 19200 17490 19250 17560
rect 19320 17490 19460 17560
rect 19530 17490 19580 17560
rect 19650 17490 19790 17560
rect 19860 17490 19910 17560
rect 19980 17490 20120 17560
rect 20190 17490 20240 17560
rect 20310 17500 20450 17560
rect 20520 17500 20570 17570
rect 20640 17500 20780 17570
rect 20850 17500 20900 17570
rect 20970 17500 21110 17570
rect 21180 17500 21230 17570
rect 21300 17560 24300 17570
rect 21300 17500 21440 17560
rect 20310 17490 21440 17500
rect 21510 17490 21560 17560
rect 21630 17490 21770 17560
rect 21840 17490 21890 17560
rect 21960 17490 22100 17560
rect 22170 17490 22220 17560
rect 22290 17490 22430 17560
rect 22500 17490 22550 17560
rect 22620 17490 22760 17560
rect 22830 17490 22880 17560
rect 22950 17490 23090 17560
rect 23160 17490 23210 17560
rect 23280 17490 23420 17560
rect 23490 17490 23540 17560
rect 23610 17490 23750 17560
rect 23820 17490 23870 17560
rect 23940 17490 24080 17560
rect 24150 17490 24200 17560
rect 24270 17490 24300 17560
rect 18870 17450 24300 17490
rect 18870 17440 20450 17450
rect 18870 17370 19130 17440
rect 19200 17370 19250 17440
rect 19320 17370 19460 17440
rect 19530 17370 19580 17440
rect 19650 17370 19790 17440
rect 19860 17370 19910 17440
rect 19980 17370 20120 17440
rect 20190 17370 20240 17440
rect 20310 17380 20450 17440
rect 20520 17380 20570 17450
rect 20640 17380 20780 17450
rect 20850 17380 20900 17450
rect 20970 17380 21110 17450
rect 21180 17380 21230 17450
rect 21300 17440 24300 17450
rect 21300 17380 21440 17440
rect 20310 17370 21440 17380
rect 21510 17370 21560 17440
rect 21630 17370 21770 17440
rect 21840 17370 21890 17440
rect 21960 17370 22100 17440
rect 22170 17370 22220 17440
rect 22290 17370 22430 17440
rect 22500 17370 22550 17440
rect 22620 17370 22760 17440
rect 22830 17370 22880 17440
rect 22950 17370 23090 17440
rect 23160 17370 23210 17440
rect 23280 17370 23420 17440
rect 23490 17370 23540 17440
rect 23610 17370 23750 17440
rect 23820 17370 23870 17440
rect 23940 17370 24080 17440
rect 24150 17370 24200 17440
rect 24270 17370 24300 17440
rect 18870 17340 24300 17370
rect 17690 16070 18260 16100
rect 17690 16000 17740 16070
rect 11630 15990 17740 16000
rect 11630 15930 11650 15990
rect 11710 15930 11740 15990
rect 11800 15930 11830 15990
rect 11890 15930 11920 15990
rect 11980 15930 12010 15990
rect 12070 15930 12100 15990
rect 12160 15930 12190 15990
rect 12250 15930 12280 15990
rect 12340 15930 12370 15990
rect 12430 15930 12460 15990
rect 12520 15930 12550 15990
rect 12610 15930 12640 15990
rect 12700 15930 12730 15990
rect 12790 15930 12820 15990
rect 12880 15930 12910 15990
rect 12970 15930 13000 15990
rect 13060 15930 13090 15990
rect 13150 15930 13180 15990
rect 13240 15930 13270 15990
rect 13330 15930 13360 15990
rect 13420 15930 13450 15990
rect 13510 15930 13540 15990
rect 13600 15930 13630 15990
rect 13690 15930 13720 15990
rect 13780 15930 13810 15990
rect 13870 15930 13900 15990
rect 13960 15930 13990 15990
rect 14050 15930 14080 15990
rect 14140 15930 14170 15990
rect 14230 15930 14260 15990
rect 14320 15930 14350 15990
rect 14410 15930 14440 15990
rect 14500 15930 14530 15990
rect 14590 15930 14620 15990
rect 14680 15930 14710 15990
rect 14770 15930 14800 15990
rect 14860 15930 14890 15990
rect 14950 15930 14980 15990
rect 15040 15930 15070 15990
rect 15130 15930 15160 15990
rect 15220 15930 15250 15990
rect 15310 15930 15340 15990
rect 15400 15930 15430 15990
rect 15490 15930 15520 15990
rect 15580 15930 15610 15990
rect 15670 15930 15700 15990
rect 15760 15930 15790 15990
rect 15850 15930 15880 15990
rect 15940 15930 15970 15990
rect 16030 15930 16060 15990
rect 16120 15930 16150 15990
rect 16210 15930 16240 15990
rect 16300 15930 16330 15990
rect 16390 15930 16420 15990
rect 16480 15930 16510 15990
rect 16570 15930 16600 15990
rect 16660 15930 16690 15990
rect 16750 15930 16780 15990
rect 16840 15930 16870 15990
rect 16930 15930 16960 15990
rect 17020 15930 17050 15990
rect 17110 15980 17740 15990
rect 17810 15980 17840 16070
rect 17910 15980 17940 16070
rect 18010 15980 18040 16070
rect 18110 15980 18140 16070
rect 18210 15980 18260 16070
rect 17110 15940 18260 15980
rect 17110 15930 17740 15940
rect 11630 15900 17740 15930
rect 11630 15840 11650 15900
rect 11710 15840 11740 15900
rect 11800 15840 11830 15900
rect 11890 15840 11920 15900
rect 11980 15840 12010 15900
rect 12070 15840 12100 15900
rect 12160 15840 12190 15900
rect 12250 15840 12280 15900
rect 12340 15840 12370 15900
rect 12430 15840 12460 15900
rect 12520 15840 12550 15900
rect 12610 15840 12640 15900
rect 12700 15840 12730 15900
rect 12790 15840 12820 15900
rect 12880 15840 12910 15900
rect 12970 15840 13000 15900
rect 13060 15840 13090 15900
rect 13150 15840 13180 15900
rect 13240 15840 13270 15900
rect 13330 15840 13360 15900
rect 13420 15840 13450 15900
rect 13510 15840 13540 15900
rect 13600 15840 13630 15900
rect 13690 15840 13720 15900
rect 13780 15840 13810 15900
rect 13870 15840 13900 15900
rect 13960 15840 13990 15900
rect 14050 15840 14080 15900
rect 14140 15840 14170 15900
rect 14230 15840 14260 15900
rect 14320 15840 14350 15900
rect 14410 15840 14440 15900
rect 14500 15840 14530 15900
rect 14590 15840 14620 15900
rect 14680 15840 14710 15900
rect 14770 15840 14800 15900
rect 14860 15840 14890 15900
rect 14950 15840 14980 15900
rect 15040 15840 15070 15900
rect 15130 15840 15160 15900
rect 15220 15840 15250 15900
rect 15310 15840 15340 15900
rect 15400 15840 15430 15900
rect 15490 15840 15520 15900
rect 15580 15840 15610 15900
rect 15670 15840 15700 15900
rect 15760 15840 15790 15900
rect 15850 15840 15880 15900
rect 15940 15840 15970 15900
rect 16030 15840 16060 15900
rect 16120 15840 16150 15900
rect 16210 15840 16240 15900
rect 16300 15840 16330 15900
rect 16390 15840 16420 15900
rect 16480 15840 16510 15900
rect 16570 15840 16600 15900
rect 16660 15840 16690 15900
rect 16750 15840 16780 15900
rect 16840 15840 16870 15900
rect 16930 15840 16960 15900
rect 17020 15840 17050 15900
rect 17110 15850 17740 15900
rect 17810 15850 17840 15940
rect 17910 15850 17940 15940
rect 18010 15850 18040 15940
rect 18110 15850 18140 15940
rect 18210 15850 18260 15940
rect 17110 15840 18260 15850
rect 11630 15820 18260 15840
rect 18980 15990 24330 16000
rect 18980 15930 19030 15990
rect 19090 15930 19120 15990
rect 19180 15930 19210 15990
rect 19270 15930 19300 15990
rect 19360 15930 19390 15990
rect 19450 15930 19480 15990
rect 19540 15930 19570 15990
rect 19630 15930 19660 15990
rect 19720 15930 19750 15990
rect 19810 15930 19840 15990
rect 19900 15930 19930 15990
rect 19990 15930 20020 15990
rect 20080 15930 20110 15990
rect 20170 15930 20200 15990
rect 20260 15930 20290 15990
rect 20350 15930 20380 15990
rect 20440 15930 20470 15990
rect 20530 15930 20560 15990
rect 20620 15930 20650 15990
rect 20710 15930 20740 15990
rect 20800 15930 20830 15990
rect 20890 15930 20920 15990
rect 20980 15930 21010 15990
rect 21070 15930 21100 15990
rect 21160 15930 21190 15990
rect 21250 15930 21280 15990
rect 21340 15930 21370 15990
rect 21430 15930 21460 15990
rect 21520 15930 21550 15990
rect 21610 15930 21640 15990
rect 21700 15930 21730 15990
rect 21790 15930 21820 15990
rect 21880 15930 21910 15990
rect 21970 15930 22000 15990
rect 22060 15930 22090 15990
rect 22150 15930 22180 15990
rect 22240 15930 22270 15990
rect 22330 15930 22360 15990
rect 22420 15930 22450 15990
rect 22510 15930 22540 15990
rect 22600 15930 22630 15990
rect 22690 15930 22720 15990
rect 22780 15930 22810 15990
rect 22870 15930 22900 15990
rect 22960 15930 22990 15990
rect 23050 15930 23080 15990
rect 23140 15930 23170 15990
rect 23230 15930 23260 15990
rect 23320 15930 23350 15990
rect 23410 15930 23440 15990
rect 23500 15930 23530 15990
rect 23590 15930 23620 15990
rect 23680 15930 23710 15990
rect 23770 15930 23800 15990
rect 23860 15930 23890 15990
rect 23950 15930 23980 15990
rect 24040 15930 24070 15990
rect 24130 15930 24160 15990
rect 24220 15930 24250 15990
rect 24310 15930 24330 15990
rect 18980 15900 24330 15930
rect 18980 15840 19030 15900
rect 19090 15840 19120 15900
rect 19180 15840 19210 15900
rect 19270 15840 19300 15900
rect 19360 15840 19390 15900
rect 19450 15840 19480 15900
rect 19540 15840 19570 15900
rect 19630 15840 19660 15900
rect 19720 15840 19750 15900
rect 19810 15840 19840 15900
rect 19900 15840 19930 15900
rect 19990 15840 20020 15900
rect 20080 15840 20110 15900
rect 20170 15840 20200 15900
rect 20260 15840 20290 15900
rect 20350 15840 20380 15900
rect 20440 15840 20470 15900
rect 20530 15840 20560 15900
rect 20620 15840 20650 15900
rect 20710 15840 20740 15900
rect 20800 15840 20830 15900
rect 20890 15840 20920 15900
rect 20980 15840 21010 15900
rect 21070 15840 21100 15900
rect 21160 15840 21190 15900
rect 21250 15840 21280 15900
rect 21340 15840 21370 15900
rect 21430 15840 21460 15900
rect 21520 15840 21550 15900
rect 21610 15840 21640 15900
rect 21700 15840 21730 15900
rect 21790 15840 21820 15900
rect 21880 15840 21910 15900
rect 21970 15840 22000 15900
rect 22060 15840 22090 15900
rect 22150 15840 22180 15900
rect 22240 15840 22270 15900
rect 22330 15840 22360 15900
rect 22420 15840 22450 15900
rect 22510 15840 22540 15900
rect 22600 15840 22630 15900
rect 22690 15840 22720 15900
rect 22780 15840 22810 15900
rect 22870 15840 22900 15900
rect 22960 15840 22990 15900
rect 23050 15840 23080 15900
rect 23140 15840 23170 15900
rect 23230 15840 23260 15900
rect 23320 15840 23350 15900
rect 23410 15840 23440 15900
rect 23500 15840 23530 15900
rect 23590 15840 23620 15900
rect 23680 15840 23710 15900
rect 23770 15840 23800 15900
rect 23860 15840 23890 15900
rect 23950 15840 23980 15900
rect 24040 15840 24070 15900
rect 24130 15840 24160 15900
rect 24220 15840 24250 15900
rect 24310 15840 24330 15900
rect 11630 13860 16980 15820
rect 18980 13880 24330 15840
rect 11630 13800 11650 13860
rect 11710 13800 11740 13860
rect 11800 13800 11830 13860
rect 11890 13800 11920 13860
rect 11980 13800 12010 13860
rect 12070 13800 12100 13860
rect 12160 13800 12190 13860
rect 12250 13800 12280 13860
rect 12340 13800 12370 13860
rect 12430 13800 12460 13860
rect 12520 13800 12550 13860
rect 12610 13800 12640 13860
rect 12700 13800 12730 13860
rect 12790 13800 12820 13860
rect 12880 13800 12910 13860
rect 12970 13800 13000 13860
rect 13060 13800 13090 13860
rect 13150 13800 13180 13860
rect 13240 13800 13270 13860
rect 13330 13800 13360 13860
rect 13420 13800 13450 13860
rect 13510 13800 13540 13860
rect 13600 13800 13630 13860
rect 13690 13800 13720 13860
rect 13780 13800 13810 13860
rect 13870 13800 13900 13860
rect 13960 13800 13990 13860
rect 14050 13800 14080 13860
rect 14140 13800 14170 13860
rect 14230 13800 14260 13860
rect 14320 13800 14350 13860
rect 14410 13800 14440 13860
rect 14500 13800 14530 13860
rect 14590 13800 14620 13860
rect 14680 13800 14710 13860
rect 14770 13800 14800 13860
rect 14860 13800 14890 13860
rect 14950 13800 14980 13860
rect 15040 13800 15070 13860
rect 15130 13800 15160 13860
rect 15220 13800 15250 13860
rect 15310 13800 15340 13860
rect 15400 13800 15430 13860
rect 15490 13800 15520 13860
rect 15580 13800 15610 13860
rect 15670 13800 15700 13860
rect 15760 13800 15790 13860
rect 15850 13800 15880 13860
rect 15940 13800 15970 13860
rect 16030 13800 16060 13860
rect 16120 13800 16150 13860
rect 16210 13800 16240 13860
rect 16300 13800 16330 13860
rect 16390 13800 16420 13860
rect 16480 13800 16510 13860
rect 16570 13800 16600 13860
rect 16660 13800 16690 13860
rect 16750 13800 16780 13860
rect 16840 13800 16870 13860
rect 16930 13800 16980 13860
rect 11630 13770 16980 13800
rect 11630 13710 11650 13770
rect 11710 13710 11740 13770
rect 11800 13710 11830 13770
rect 11890 13710 11920 13770
rect 11980 13710 12010 13770
rect 12070 13710 12100 13770
rect 12160 13710 12190 13770
rect 12250 13710 12280 13770
rect 12340 13710 12370 13770
rect 12430 13710 12460 13770
rect 12520 13710 12550 13770
rect 12610 13710 12640 13770
rect 12700 13710 12730 13770
rect 12790 13710 12820 13770
rect 12880 13710 12910 13770
rect 12970 13710 13000 13770
rect 13060 13710 13090 13770
rect 13150 13710 13180 13770
rect 13240 13710 13270 13770
rect 13330 13710 13360 13770
rect 13420 13710 13450 13770
rect 13510 13710 13540 13770
rect 13600 13710 13630 13770
rect 13690 13710 13720 13770
rect 13780 13710 13810 13770
rect 13870 13710 13900 13770
rect 13960 13710 13990 13770
rect 14050 13710 14080 13770
rect 14140 13710 14170 13770
rect 14230 13710 14260 13770
rect 14320 13710 14350 13770
rect 14410 13710 14440 13770
rect 14500 13710 14530 13770
rect 14590 13710 14620 13770
rect 14680 13710 14710 13770
rect 14770 13710 14800 13770
rect 14860 13710 14890 13770
rect 14950 13710 14980 13770
rect 15040 13710 15070 13770
rect 15130 13710 15160 13770
rect 15220 13710 15250 13770
rect 15310 13710 15340 13770
rect 15400 13710 15430 13770
rect 15490 13710 15520 13770
rect 15580 13710 15610 13770
rect 15670 13710 15700 13770
rect 15760 13710 15790 13770
rect 15850 13710 15880 13770
rect 15940 13710 15970 13770
rect 16030 13710 16060 13770
rect 16120 13710 16150 13770
rect 16210 13710 16240 13770
rect 16300 13710 16330 13770
rect 16390 13710 16420 13770
rect 16480 13710 16510 13770
rect 16570 13710 16600 13770
rect 16660 13710 16690 13770
rect 16750 13710 16780 13770
rect 16840 13710 16870 13770
rect 16930 13710 16980 13770
rect 11630 13700 16980 13710
rect 17690 13860 24330 13880
rect 17690 13850 18850 13860
rect 17690 13760 17740 13850
rect 17810 13760 17840 13850
rect 17910 13760 17940 13850
rect 18010 13760 18040 13850
rect 18110 13760 18140 13850
rect 18210 13800 18850 13850
rect 18910 13800 18940 13860
rect 19000 13800 19030 13860
rect 19090 13800 19120 13860
rect 19180 13800 19210 13860
rect 19270 13800 19300 13860
rect 19360 13800 19390 13860
rect 19450 13800 19480 13860
rect 19540 13800 19570 13860
rect 19630 13800 19660 13860
rect 19720 13800 19750 13860
rect 19810 13800 19840 13860
rect 19900 13800 19930 13860
rect 19990 13800 20020 13860
rect 20080 13800 20110 13860
rect 20170 13800 20200 13860
rect 20260 13800 20290 13860
rect 20350 13800 20380 13860
rect 20440 13800 20470 13860
rect 20530 13800 20560 13860
rect 20620 13800 20650 13860
rect 20710 13800 20740 13860
rect 20800 13800 20830 13860
rect 20890 13800 20920 13860
rect 20980 13800 21010 13860
rect 21070 13800 21100 13860
rect 21160 13800 21190 13860
rect 21250 13800 21280 13860
rect 21340 13800 21370 13860
rect 21430 13800 21460 13860
rect 21520 13800 21550 13860
rect 21610 13800 21640 13860
rect 21700 13800 21730 13860
rect 21790 13800 21820 13860
rect 21880 13800 21910 13860
rect 21970 13800 22000 13860
rect 22060 13800 22090 13860
rect 22150 13800 22180 13860
rect 22240 13800 22270 13860
rect 22330 13800 22360 13860
rect 22420 13800 22450 13860
rect 22510 13800 22540 13860
rect 22600 13800 22630 13860
rect 22690 13800 22720 13860
rect 22780 13800 22810 13860
rect 22870 13800 22900 13860
rect 22960 13800 22990 13860
rect 23050 13800 23080 13860
rect 23140 13800 23170 13860
rect 23230 13800 23260 13860
rect 23320 13800 23350 13860
rect 23410 13800 23440 13860
rect 23500 13800 23530 13860
rect 23590 13800 23620 13860
rect 23680 13800 23710 13860
rect 23770 13800 23800 13860
rect 23860 13800 23890 13860
rect 23950 13800 23980 13860
rect 24040 13800 24070 13860
rect 24130 13800 24160 13860
rect 24220 13800 24250 13860
rect 24310 13800 24330 13860
rect 18210 13770 24330 13800
rect 18210 13760 18850 13770
rect 17690 13720 18850 13760
rect 17690 13630 17740 13720
rect 17810 13630 17840 13720
rect 17910 13630 17940 13720
rect 18010 13630 18040 13720
rect 18110 13630 18140 13720
rect 18210 13710 18850 13720
rect 18910 13710 18940 13770
rect 19000 13710 19030 13770
rect 19090 13710 19120 13770
rect 19180 13710 19210 13770
rect 19270 13710 19300 13770
rect 19360 13710 19390 13770
rect 19450 13710 19480 13770
rect 19540 13710 19570 13770
rect 19630 13710 19660 13770
rect 19720 13710 19750 13770
rect 19810 13710 19840 13770
rect 19900 13710 19930 13770
rect 19990 13710 20020 13770
rect 20080 13710 20110 13770
rect 20170 13710 20200 13770
rect 20260 13710 20290 13770
rect 20350 13710 20380 13770
rect 20440 13710 20470 13770
rect 20530 13710 20560 13770
rect 20620 13710 20650 13770
rect 20710 13710 20740 13770
rect 20800 13710 20830 13770
rect 20890 13710 20920 13770
rect 20980 13710 21010 13770
rect 21070 13710 21100 13770
rect 21160 13710 21190 13770
rect 21250 13710 21280 13770
rect 21340 13710 21370 13770
rect 21430 13710 21460 13770
rect 21520 13710 21550 13770
rect 21610 13710 21640 13770
rect 21700 13710 21730 13770
rect 21790 13710 21820 13770
rect 21880 13710 21910 13770
rect 21970 13710 22000 13770
rect 22060 13710 22090 13770
rect 22150 13710 22180 13770
rect 22240 13710 22270 13770
rect 22330 13710 22360 13770
rect 22420 13710 22450 13770
rect 22510 13710 22540 13770
rect 22600 13710 22630 13770
rect 22690 13710 22720 13770
rect 22780 13710 22810 13770
rect 22870 13710 22900 13770
rect 22960 13710 22990 13770
rect 23050 13710 23080 13770
rect 23140 13710 23170 13770
rect 23230 13710 23260 13770
rect 23320 13710 23350 13770
rect 23410 13710 23440 13770
rect 23500 13710 23530 13770
rect 23590 13710 23620 13770
rect 23680 13710 23710 13770
rect 23770 13710 23800 13770
rect 23860 13710 23890 13770
rect 23950 13710 23980 13770
rect 24040 13710 24070 13770
rect 24130 13710 24160 13770
rect 24220 13710 24250 13770
rect 24310 13710 24330 13770
rect 18210 13700 24330 13710
rect 18210 13630 18260 13700
rect 17690 13600 18260 13630
rect 11660 12310 17090 12340
rect 11660 12240 11690 12310
rect 11760 12240 11810 12310
rect 11880 12240 12020 12310
rect 12090 12240 12140 12310
rect 12210 12240 12350 12310
rect 12420 12240 12470 12310
rect 12540 12240 12680 12310
rect 12750 12240 12800 12310
rect 12870 12240 13010 12310
rect 13080 12240 13130 12310
rect 13200 12240 13340 12310
rect 13410 12240 13460 12310
rect 13530 12240 13670 12310
rect 13740 12240 13790 12310
rect 13860 12240 14000 12310
rect 14070 12240 14120 12310
rect 14190 12240 14330 12310
rect 14400 12240 14450 12310
rect 14520 12300 15650 12310
rect 14520 12240 14660 12300
rect 11660 12230 14660 12240
rect 14730 12230 14780 12300
rect 14850 12230 14990 12300
rect 15060 12230 15110 12300
rect 15180 12230 15320 12300
rect 15390 12230 15440 12300
rect 15510 12240 15650 12300
rect 15720 12240 15770 12310
rect 15840 12240 15980 12310
rect 16050 12240 16100 12310
rect 16170 12240 16310 12310
rect 16380 12240 16430 12310
rect 16500 12240 16640 12310
rect 16710 12240 16760 12310
rect 16830 12240 17090 12310
rect 15510 12230 17090 12240
rect 11660 12190 17090 12230
rect 11660 12120 11690 12190
rect 11760 12120 11810 12190
rect 11880 12120 12020 12190
rect 12090 12120 12140 12190
rect 12210 12120 12350 12190
rect 12420 12120 12470 12190
rect 12540 12120 12680 12190
rect 12750 12120 12800 12190
rect 12870 12120 13010 12190
rect 13080 12120 13130 12190
rect 13200 12120 13340 12190
rect 13410 12120 13460 12190
rect 13530 12120 13670 12190
rect 13740 12120 13790 12190
rect 13860 12120 14000 12190
rect 14070 12120 14120 12190
rect 14190 12120 14330 12190
rect 14400 12120 14450 12190
rect 14520 12180 15650 12190
rect 14520 12120 14660 12180
rect 11660 12110 14660 12120
rect 14730 12110 14780 12180
rect 14850 12110 14990 12180
rect 15060 12110 15110 12180
rect 15180 12110 15320 12180
rect 15390 12110 15440 12180
rect 15510 12120 15650 12180
rect 15720 12120 15770 12190
rect 15840 12120 15980 12190
rect 16050 12120 16100 12190
rect 16170 12120 16310 12190
rect 16380 12120 16430 12190
rect 16500 12120 16640 12190
rect 16710 12120 16760 12190
rect 16830 12120 17090 12190
rect 15510 12110 17090 12120
rect 11660 12090 17090 12110
rect 18870 12310 24300 12340
rect 18870 12240 19130 12310
rect 19200 12240 19250 12310
rect 19320 12240 19460 12310
rect 19530 12240 19580 12310
rect 19650 12240 19790 12310
rect 19860 12240 19910 12310
rect 19980 12240 20120 12310
rect 20190 12240 20240 12310
rect 20310 12300 21440 12310
rect 20310 12240 20450 12300
rect 18870 12230 20450 12240
rect 20520 12230 20570 12300
rect 20640 12230 20780 12300
rect 20850 12230 20900 12300
rect 20970 12230 21110 12300
rect 21180 12230 21230 12300
rect 21300 12240 21440 12300
rect 21510 12240 21560 12310
rect 21630 12240 21770 12310
rect 21840 12240 21890 12310
rect 21960 12240 22100 12310
rect 22170 12240 22220 12310
rect 22290 12240 22430 12310
rect 22500 12240 22550 12310
rect 22620 12240 22760 12310
rect 22830 12240 22880 12310
rect 22950 12240 23090 12310
rect 23160 12240 23210 12310
rect 23280 12240 23420 12310
rect 23490 12240 23540 12310
rect 23610 12240 23750 12310
rect 23820 12240 23870 12310
rect 23940 12240 24080 12310
rect 24150 12240 24200 12310
rect 24270 12240 24300 12310
rect 21300 12230 24300 12240
rect 18870 12190 24300 12230
rect 18870 12120 19130 12190
rect 19200 12120 19250 12190
rect 19320 12120 19460 12190
rect 19530 12120 19580 12190
rect 19650 12120 19790 12190
rect 19860 12120 19910 12190
rect 19980 12120 20120 12190
rect 20190 12120 20240 12190
rect 20310 12180 21440 12190
rect 20310 12120 20450 12180
rect 18870 12110 20450 12120
rect 20520 12110 20570 12180
rect 20640 12110 20780 12180
rect 20850 12110 20900 12180
rect 20970 12110 21110 12180
rect 21180 12110 21230 12180
rect 21300 12120 21440 12180
rect 21510 12120 21560 12190
rect 21630 12120 21770 12190
rect 21840 12120 21890 12190
rect 21960 12120 22100 12190
rect 22170 12120 22220 12190
rect 22290 12120 22430 12190
rect 22500 12120 22550 12190
rect 22620 12120 22760 12190
rect 22830 12120 22880 12190
rect 22950 12120 23090 12190
rect 23160 12120 23210 12190
rect 23280 12120 23420 12190
rect 23490 12120 23540 12190
rect 23610 12120 23750 12190
rect 23820 12120 23870 12190
rect 23940 12120 24080 12190
rect 24150 12120 24200 12190
rect 24270 12120 24300 12190
rect 21300 12110 24300 12120
rect 18870 12090 24300 12110
rect 11690 12070 11930 12090
rect 12020 12070 12260 12090
rect 12350 12070 12590 12090
rect 12680 12070 12920 12090
rect 13010 12070 13250 12090
rect 13340 12070 13580 12090
rect 13670 12070 13910 12090
rect 14000 12070 14240 12090
rect 14330 12070 14570 12090
rect 14660 12070 14900 12090
rect 14990 12070 15230 12090
rect 15320 12070 15560 12090
rect 15650 12070 15890 12090
rect 15980 12070 16220 12090
rect 16310 12070 16550 12090
rect 16640 12070 16880 12090
rect 19080 12070 19320 12090
rect 19410 12070 19650 12090
rect 19740 12070 19980 12090
rect 20070 12070 20310 12090
rect 20400 12070 20640 12090
rect 20730 12070 20970 12090
rect 21060 12070 21300 12090
rect 21390 12070 21630 12090
rect 21720 12070 21960 12090
rect 22050 12070 22290 12090
rect 22380 12070 22620 12090
rect 22710 12070 22950 12090
rect 23040 12070 23280 12090
rect 23370 12070 23610 12090
rect 23700 12070 23940 12090
rect 24030 12070 24270 12090
<< via3 >>
rect 11690 17490 11760 17560
rect 11810 17490 11880 17560
rect 12020 17490 12090 17560
rect 12140 17490 12210 17560
rect 12350 17490 12420 17560
rect 12470 17490 12540 17560
rect 12680 17490 12750 17560
rect 12800 17490 12870 17560
rect 13010 17490 13080 17560
rect 13130 17490 13200 17560
rect 13340 17490 13410 17560
rect 13460 17490 13530 17560
rect 13670 17490 13740 17560
rect 13790 17490 13860 17560
rect 14000 17490 14070 17560
rect 14120 17490 14190 17560
rect 14330 17490 14400 17560
rect 14450 17490 14520 17560
rect 14660 17500 14730 17570
rect 14780 17500 14850 17570
rect 14990 17500 15060 17570
rect 15110 17500 15180 17570
rect 15320 17500 15390 17570
rect 15440 17500 15510 17570
rect 15650 17490 15720 17560
rect 15770 17490 15840 17560
rect 15980 17490 16050 17560
rect 16100 17490 16170 17560
rect 16310 17490 16380 17560
rect 16430 17490 16500 17560
rect 16640 17490 16710 17560
rect 16760 17490 16830 17560
rect 11690 17370 11760 17440
rect 11810 17370 11880 17440
rect 12020 17370 12090 17440
rect 12140 17370 12210 17440
rect 12350 17370 12420 17440
rect 12470 17370 12540 17440
rect 12680 17370 12750 17440
rect 12800 17370 12870 17440
rect 13010 17370 13080 17440
rect 13130 17370 13200 17440
rect 13340 17370 13410 17440
rect 13460 17370 13530 17440
rect 13670 17370 13740 17440
rect 13790 17370 13860 17440
rect 14000 17370 14070 17440
rect 14120 17370 14190 17440
rect 14330 17370 14400 17440
rect 14450 17370 14520 17440
rect 14660 17380 14730 17450
rect 14780 17380 14850 17450
rect 14990 17380 15060 17450
rect 15110 17380 15180 17450
rect 15320 17380 15390 17450
rect 15440 17380 15510 17450
rect 15650 17370 15720 17440
rect 15770 17370 15840 17440
rect 15980 17370 16050 17440
rect 16100 17370 16170 17440
rect 16310 17370 16380 17440
rect 16430 17370 16500 17440
rect 16640 17370 16710 17440
rect 16760 17370 16830 17440
rect 19130 17490 19200 17560
rect 19250 17490 19320 17560
rect 19460 17490 19530 17560
rect 19580 17490 19650 17560
rect 19790 17490 19860 17560
rect 19910 17490 19980 17560
rect 20120 17490 20190 17560
rect 20240 17490 20310 17560
rect 20450 17500 20520 17570
rect 20570 17500 20640 17570
rect 20780 17500 20850 17570
rect 20900 17500 20970 17570
rect 21110 17500 21180 17570
rect 21230 17500 21300 17570
rect 21440 17490 21510 17560
rect 21560 17490 21630 17560
rect 21770 17490 21840 17560
rect 21890 17490 21960 17560
rect 22100 17490 22170 17560
rect 22220 17490 22290 17560
rect 22430 17490 22500 17560
rect 22550 17490 22620 17560
rect 22760 17490 22830 17560
rect 22880 17490 22950 17560
rect 23090 17490 23160 17560
rect 23210 17490 23280 17560
rect 23420 17490 23490 17560
rect 23540 17490 23610 17560
rect 23750 17490 23820 17560
rect 23870 17490 23940 17560
rect 24080 17490 24150 17560
rect 24200 17490 24270 17560
rect 19130 17370 19200 17440
rect 19250 17370 19320 17440
rect 19460 17370 19530 17440
rect 19580 17370 19650 17440
rect 19790 17370 19860 17440
rect 19910 17370 19980 17440
rect 20120 17370 20190 17440
rect 20240 17370 20310 17440
rect 20450 17380 20520 17450
rect 20570 17380 20640 17450
rect 20780 17380 20850 17450
rect 20900 17380 20970 17450
rect 21110 17380 21180 17450
rect 21230 17380 21300 17450
rect 21440 17370 21510 17440
rect 21560 17370 21630 17440
rect 21770 17370 21840 17440
rect 21890 17370 21960 17440
rect 22100 17370 22170 17440
rect 22220 17370 22290 17440
rect 22430 17370 22500 17440
rect 22550 17370 22620 17440
rect 22760 17370 22830 17440
rect 22880 17370 22950 17440
rect 23090 17370 23160 17440
rect 23210 17370 23280 17440
rect 23420 17370 23490 17440
rect 23540 17370 23610 17440
rect 23750 17370 23820 17440
rect 23870 17370 23940 17440
rect 24080 17370 24150 17440
rect 24200 17370 24270 17440
rect 17740 15980 17810 16070
rect 17840 15980 17910 16070
rect 17940 15980 18010 16070
rect 18040 15980 18110 16070
rect 18140 15980 18210 16070
rect 17740 15850 17810 15940
rect 17840 15850 17910 15940
rect 17940 15850 18010 15940
rect 18040 15850 18110 15940
rect 18140 15850 18210 15940
rect 17740 13760 17810 13850
rect 17840 13760 17910 13850
rect 17940 13760 18010 13850
rect 18040 13760 18110 13850
rect 18140 13760 18210 13850
rect 17740 13630 17810 13720
rect 17840 13630 17910 13720
rect 17940 13630 18010 13720
rect 18040 13630 18110 13720
rect 18140 13630 18210 13720
rect 11690 12240 11760 12310
rect 11810 12240 11880 12310
rect 12020 12240 12090 12310
rect 12140 12240 12210 12310
rect 12350 12240 12420 12310
rect 12470 12240 12540 12310
rect 12680 12240 12750 12310
rect 12800 12240 12870 12310
rect 13010 12240 13080 12310
rect 13130 12240 13200 12310
rect 13340 12240 13410 12310
rect 13460 12240 13530 12310
rect 13670 12240 13740 12310
rect 13790 12240 13860 12310
rect 14000 12240 14070 12310
rect 14120 12240 14190 12310
rect 14330 12240 14400 12310
rect 14450 12240 14520 12310
rect 14660 12230 14730 12300
rect 14780 12230 14850 12300
rect 14990 12230 15060 12300
rect 15110 12230 15180 12300
rect 15320 12230 15390 12300
rect 15440 12230 15510 12300
rect 15650 12240 15720 12310
rect 15770 12240 15840 12310
rect 15980 12240 16050 12310
rect 16100 12240 16170 12310
rect 16310 12240 16380 12310
rect 16430 12240 16500 12310
rect 16640 12240 16710 12310
rect 16760 12240 16830 12310
rect 11690 12120 11760 12190
rect 11810 12120 11880 12190
rect 12020 12120 12090 12190
rect 12140 12120 12210 12190
rect 12350 12120 12420 12190
rect 12470 12120 12540 12190
rect 12680 12120 12750 12190
rect 12800 12120 12870 12190
rect 13010 12120 13080 12190
rect 13130 12120 13200 12190
rect 13340 12120 13410 12190
rect 13460 12120 13530 12190
rect 13670 12120 13740 12190
rect 13790 12120 13860 12190
rect 14000 12120 14070 12190
rect 14120 12120 14190 12190
rect 14330 12120 14400 12190
rect 14450 12120 14520 12190
rect 14660 12110 14730 12180
rect 14780 12110 14850 12180
rect 14990 12110 15060 12180
rect 15110 12110 15180 12180
rect 15320 12110 15390 12180
rect 15440 12110 15510 12180
rect 15650 12120 15720 12190
rect 15770 12120 15840 12190
rect 15980 12120 16050 12190
rect 16100 12120 16170 12190
rect 16310 12120 16380 12190
rect 16430 12120 16500 12190
rect 16640 12120 16710 12190
rect 16760 12120 16830 12190
rect 19130 12240 19200 12310
rect 19250 12240 19320 12310
rect 19460 12240 19530 12310
rect 19580 12240 19650 12310
rect 19790 12240 19860 12310
rect 19910 12240 19980 12310
rect 20120 12240 20190 12310
rect 20240 12240 20310 12310
rect 20450 12230 20520 12300
rect 20570 12230 20640 12300
rect 20780 12230 20850 12300
rect 20900 12230 20970 12300
rect 21110 12230 21180 12300
rect 21230 12230 21300 12300
rect 21440 12240 21510 12310
rect 21560 12240 21630 12310
rect 21770 12240 21840 12310
rect 21890 12240 21960 12310
rect 22100 12240 22170 12310
rect 22220 12240 22290 12310
rect 22430 12240 22500 12310
rect 22550 12240 22620 12310
rect 22760 12240 22830 12310
rect 22880 12240 22950 12310
rect 23090 12240 23160 12310
rect 23210 12240 23280 12310
rect 23420 12240 23490 12310
rect 23540 12240 23610 12310
rect 23750 12240 23820 12310
rect 23870 12240 23940 12310
rect 24080 12240 24150 12310
rect 24200 12240 24270 12310
rect 19130 12120 19200 12190
rect 19250 12120 19320 12190
rect 19460 12120 19530 12190
rect 19580 12120 19650 12190
rect 19790 12120 19860 12190
rect 19910 12120 19980 12190
rect 20120 12120 20190 12190
rect 20240 12120 20310 12190
rect 20450 12110 20520 12180
rect 20570 12110 20640 12180
rect 20780 12110 20850 12180
rect 20900 12110 20970 12180
rect 21110 12110 21180 12180
rect 21230 12110 21300 12180
rect 21440 12120 21510 12190
rect 21560 12120 21630 12190
rect 21770 12120 21840 12190
rect 21890 12120 21960 12190
rect 22100 12120 22170 12190
rect 22220 12120 22290 12190
rect 22430 12120 22500 12190
rect 22550 12120 22620 12190
rect 22760 12120 22830 12190
rect 22880 12120 22950 12190
rect 23090 12120 23160 12190
rect 23210 12120 23280 12190
rect 23420 12120 23490 12190
rect 23540 12120 23610 12190
rect 23750 12120 23820 12190
rect 23870 12120 23940 12190
rect 24080 12120 24150 12190
rect 24200 12120 24270 12190
<< metal4 >>
rect 17180 17660 18780 18230
rect 11660 17610 17090 17660
rect 11660 17370 11690 17610
rect 11930 17370 12020 17610
rect 12260 17370 12350 17610
rect 12590 17370 12680 17610
rect 12920 17370 13010 17610
rect 13250 17370 13340 17610
rect 13580 17370 13670 17610
rect 13910 17370 14000 17610
rect 14240 17370 14330 17610
rect 14570 17370 14660 17610
rect 14900 17370 14990 17610
rect 15230 17370 15320 17610
rect 15560 17370 15650 17610
rect 15890 17370 15980 17610
rect 16220 17370 16310 17610
rect 16550 17370 16640 17610
rect 16880 17370 17090 17610
rect 11660 17340 17090 17370
rect 17180 17340 18790 17660
rect 18870 17610 24300 17660
rect 18870 17370 19080 17610
rect 19320 17370 19410 17610
rect 19650 17370 19740 17610
rect 19980 17370 20070 17610
rect 20310 17370 20400 17610
rect 20640 17370 20730 17610
rect 20970 17370 21060 17610
rect 21300 17370 21390 17610
rect 21630 17370 21720 17610
rect 21960 17370 22050 17610
rect 22290 17370 22380 17610
rect 22620 17370 22710 17610
rect 22950 17370 23040 17610
rect 23280 17370 23370 17610
rect 23610 17370 23700 17610
rect 23940 17370 24030 17610
rect 24270 17370 24300 17610
rect 18870 17340 24300 17370
rect 17180 16070 18780 17340
rect 17180 15980 17740 16070
rect 17810 15980 17840 16070
rect 17910 15980 17940 16070
rect 18010 15980 18040 16070
rect 18110 15980 18140 16070
rect 18210 15980 18780 16070
rect 17180 15940 18780 15980
rect 17180 15850 17740 15940
rect 17810 15850 17840 15940
rect 17910 15850 17940 15940
rect 18010 15850 18040 15940
rect 18110 15850 18140 15940
rect 18210 15850 18780 15940
rect 17180 15820 18780 15850
rect 17180 15810 17690 15820
rect 18260 15810 18780 15820
rect 17180 13850 18780 13880
rect 17180 13760 17740 13850
rect 17810 13760 17840 13850
rect 17910 13760 17940 13850
rect 18010 13760 18040 13850
rect 18110 13760 18140 13850
rect 18210 13760 18780 13850
rect 17180 13720 18780 13760
rect 17180 13630 17740 13720
rect 17810 13630 17840 13720
rect 17910 13630 17940 13720
rect 18010 13630 18040 13720
rect 18110 13630 18140 13720
rect 18210 13630 18780 13720
rect 17180 12340 18780 13630
rect 11660 12310 17090 12340
rect 11660 12070 11690 12310
rect 11930 12070 12020 12310
rect 12260 12070 12350 12310
rect 12590 12070 12680 12310
rect 12920 12070 13010 12310
rect 13250 12070 13340 12310
rect 13580 12070 13670 12310
rect 13910 12070 14000 12310
rect 14240 12070 14330 12310
rect 14570 12070 14660 12310
rect 14900 12070 14990 12310
rect 15230 12070 15320 12310
rect 15560 12070 15650 12310
rect 15890 12070 15980 12310
rect 16220 12070 16310 12310
rect 16550 12070 16640 12310
rect 16880 12070 17090 12310
rect 11660 12020 17090 12070
rect 17180 12020 18800 12340
rect 18870 12310 24300 12340
rect 18870 12070 19080 12310
rect 19320 12070 19410 12310
rect 19650 12070 19740 12310
rect 19980 12070 20070 12310
rect 20310 12070 20400 12310
rect 20640 12070 20730 12310
rect 20970 12070 21060 12310
rect 21300 12070 21390 12310
rect 21630 12070 21720 12310
rect 21960 12070 22050 12310
rect 22290 12070 22380 12310
rect 22620 12070 22710 12310
rect 22950 12070 23040 12310
rect 23280 12070 23370 12310
rect 23610 12070 23700 12310
rect 23940 12070 24030 12310
rect 24270 12070 24300 12310
rect 18870 12020 24300 12070
rect 17180 11470 18780 12020
<< via4 >>
rect 11690 17560 11930 17610
rect 11690 17490 11760 17560
rect 11760 17490 11810 17560
rect 11810 17490 11880 17560
rect 11880 17490 11930 17560
rect 11690 17440 11930 17490
rect 11690 17370 11760 17440
rect 11760 17370 11810 17440
rect 11810 17370 11880 17440
rect 11880 17370 11930 17440
rect 12020 17560 12260 17610
rect 12020 17490 12090 17560
rect 12090 17490 12140 17560
rect 12140 17490 12210 17560
rect 12210 17490 12260 17560
rect 12020 17440 12260 17490
rect 12020 17370 12090 17440
rect 12090 17370 12140 17440
rect 12140 17370 12210 17440
rect 12210 17370 12260 17440
rect 12350 17560 12590 17610
rect 12350 17490 12420 17560
rect 12420 17490 12470 17560
rect 12470 17490 12540 17560
rect 12540 17490 12590 17560
rect 12350 17440 12590 17490
rect 12350 17370 12420 17440
rect 12420 17370 12470 17440
rect 12470 17370 12540 17440
rect 12540 17370 12590 17440
rect 12680 17560 12920 17610
rect 12680 17490 12750 17560
rect 12750 17490 12800 17560
rect 12800 17490 12870 17560
rect 12870 17490 12920 17560
rect 12680 17440 12920 17490
rect 12680 17370 12750 17440
rect 12750 17370 12800 17440
rect 12800 17370 12870 17440
rect 12870 17370 12920 17440
rect 13010 17560 13250 17610
rect 13010 17490 13080 17560
rect 13080 17490 13130 17560
rect 13130 17490 13200 17560
rect 13200 17490 13250 17560
rect 13010 17440 13250 17490
rect 13010 17370 13080 17440
rect 13080 17370 13130 17440
rect 13130 17370 13200 17440
rect 13200 17370 13250 17440
rect 13340 17560 13580 17610
rect 13340 17490 13410 17560
rect 13410 17490 13460 17560
rect 13460 17490 13530 17560
rect 13530 17490 13580 17560
rect 13340 17440 13580 17490
rect 13340 17370 13410 17440
rect 13410 17370 13460 17440
rect 13460 17370 13530 17440
rect 13530 17370 13580 17440
rect 13670 17560 13910 17610
rect 13670 17490 13740 17560
rect 13740 17490 13790 17560
rect 13790 17490 13860 17560
rect 13860 17490 13910 17560
rect 13670 17440 13910 17490
rect 13670 17370 13740 17440
rect 13740 17370 13790 17440
rect 13790 17370 13860 17440
rect 13860 17370 13910 17440
rect 14000 17560 14240 17610
rect 14000 17490 14070 17560
rect 14070 17490 14120 17560
rect 14120 17490 14190 17560
rect 14190 17490 14240 17560
rect 14000 17440 14240 17490
rect 14000 17370 14070 17440
rect 14070 17370 14120 17440
rect 14120 17370 14190 17440
rect 14190 17370 14240 17440
rect 14330 17560 14570 17610
rect 14330 17490 14400 17560
rect 14400 17490 14450 17560
rect 14450 17490 14520 17560
rect 14520 17490 14570 17560
rect 14330 17440 14570 17490
rect 14330 17370 14400 17440
rect 14400 17370 14450 17440
rect 14450 17370 14520 17440
rect 14520 17370 14570 17440
rect 14660 17570 14900 17610
rect 14660 17500 14730 17570
rect 14730 17500 14780 17570
rect 14780 17500 14850 17570
rect 14850 17500 14900 17570
rect 14660 17450 14900 17500
rect 14660 17380 14730 17450
rect 14730 17380 14780 17450
rect 14780 17380 14850 17450
rect 14850 17380 14900 17450
rect 14660 17370 14900 17380
rect 14990 17570 15230 17610
rect 14990 17500 15060 17570
rect 15060 17500 15110 17570
rect 15110 17500 15180 17570
rect 15180 17500 15230 17570
rect 14990 17450 15230 17500
rect 14990 17380 15060 17450
rect 15060 17380 15110 17450
rect 15110 17380 15180 17450
rect 15180 17380 15230 17450
rect 14990 17370 15230 17380
rect 15320 17570 15560 17610
rect 15320 17500 15390 17570
rect 15390 17500 15440 17570
rect 15440 17500 15510 17570
rect 15510 17500 15560 17570
rect 15320 17450 15560 17500
rect 15320 17380 15390 17450
rect 15390 17380 15440 17450
rect 15440 17380 15510 17450
rect 15510 17380 15560 17450
rect 15320 17370 15560 17380
rect 15650 17560 15890 17610
rect 15650 17490 15720 17560
rect 15720 17490 15770 17560
rect 15770 17490 15840 17560
rect 15840 17490 15890 17560
rect 15650 17440 15890 17490
rect 15650 17370 15720 17440
rect 15720 17370 15770 17440
rect 15770 17370 15840 17440
rect 15840 17370 15890 17440
rect 15980 17560 16220 17610
rect 15980 17490 16050 17560
rect 16050 17490 16100 17560
rect 16100 17490 16170 17560
rect 16170 17490 16220 17560
rect 15980 17440 16220 17490
rect 15980 17370 16050 17440
rect 16050 17370 16100 17440
rect 16100 17370 16170 17440
rect 16170 17370 16220 17440
rect 16310 17560 16550 17610
rect 16310 17490 16380 17560
rect 16380 17490 16430 17560
rect 16430 17490 16500 17560
rect 16500 17490 16550 17560
rect 16310 17440 16550 17490
rect 16310 17370 16380 17440
rect 16380 17370 16430 17440
rect 16430 17370 16500 17440
rect 16500 17370 16550 17440
rect 16640 17560 16880 17610
rect 16640 17490 16710 17560
rect 16710 17490 16760 17560
rect 16760 17490 16830 17560
rect 16830 17490 16880 17560
rect 16640 17440 16880 17490
rect 16640 17370 16710 17440
rect 16710 17370 16760 17440
rect 16760 17370 16830 17440
rect 16830 17370 16880 17440
rect 19080 17560 19320 17610
rect 19080 17490 19130 17560
rect 19130 17490 19200 17560
rect 19200 17490 19250 17560
rect 19250 17490 19320 17560
rect 19080 17440 19320 17490
rect 19080 17370 19130 17440
rect 19130 17370 19200 17440
rect 19200 17370 19250 17440
rect 19250 17370 19320 17440
rect 19410 17560 19650 17610
rect 19410 17490 19460 17560
rect 19460 17490 19530 17560
rect 19530 17490 19580 17560
rect 19580 17490 19650 17560
rect 19410 17440 19650 17490
rect 19410 17370 19460 17440
rect 19460 17370 19530 17440
rect 19530 17370 19580 17440
rect 19580 17370 19650 17440
rect 19740 17560 19980 17610
rect 19740 17490 19790 17560
rect 19790 17490 19860 17560
rect 19860 17490 19910 17560
rect 19910 17490 19980 17560
rect 19740 17440 19980 17490
rect 19740 17370 19790 17440
rect 19790 17370 19860 17440
rect 19860 17370 19910 17440
rect 19910 17370 19980 17440
rect 20070 17560 20310 17610
rect 20070 17490 20120 17560
rect 20120 17490 20190 17560
rect 20190 17490 20240 17560
rect 20240 17490 20310 17560
rect 20070 17440 20310 17490
rect 20070 17370 20120 17440
rect 20120 17370 20190 17440
rect 20190 17370 20240 17440
rect 20240 17370 20310 17440
rect 20400 17570 20640 17610
rect 20400 17500 20450 17570
rect 20450 17500 20520 17570
rect 20520 17500 20570 17570
rect 20570 17500 20640 17570
rect 20400 17450 20640 17500
rect 20400 17380 20450 17450
rect 20450 17380 20520 17450
rect 20520 17380 20570 17450
rect 20570 17380 20640 17450
rect 20400 17370 20640 17380
rect 20730 17570 20970 17610
rect 20730 17500 20780 17570
rect 20780 17500 20850 17570
rect 20850 17500 20900 17570
rect 20900 17500 20970 17570
rect 20730 17450 20970 17500
rect 20730 17380 20780 17450
rect 20780 17380 20850 17450
rect 20850 17380 20900 17450
rect 20900 17380 20970 17450
rect 20730 17370 20970 17380
rect 21060 17570 21300 17610
rect 21060 17500 21110 17570
rect 21110 17500 21180 17570
rect 21180 17500 21230 17570
rect 21230 17500 21300 17570
rect 21060 17450 21300 17500
rect 21060 17380 21110 17450
rect 21110 17380 21180 17450
rect 21180 17380 21230 17450
rect 21230 17380 21300 17450
rect 21060 17370 21300 17380
rect 21390 17560 21630 17610
rect 21390 17490 21440 17560
rect 21440 17490 21510 17560
rect 21510 17490 21560 17560
rect 21560 17490 21630 17560
rect 21390 17440 21630 17490
rect 21390 17370 21440 17440
rect 21440 17370 21510 17440
rect 21510 17370 21560 17440
rect 21560 17370 21630 17440
rect 21720 17560 21960 17610
rect 21720 17490 21770 17560
rect 21770 17490 21840 17560
rect 21840 17490 21890 17560
rect 21890 17490 21960 17560
rect 21720 17440 21960 17490
rect 21720 17370 21770 17440
rect 21770 17370 21840 17440
rect 21840 17370 21890 17440
rect 21890 17370 21960 17440
rect 22050 17560 22290 17610
rect 22050 17490 22100 17560
rect 22100 17490 22170 17560
rect 22170 17490 22220 17560
rect 22220 17490 22290 17560
rect 22050 17440 22290 17490
rect 22050 17370 22100 17440
rect 22100 17370 22170 17440
rect 22170 17370 22220 17440
rect 22220 17370 22290 17440
rect 22380 17560 22620 17610
rect 22380 17490 22430 17560
rect 22430 17490 22500 17560
rect 22500 17490 22550 17560
rect 22550 17490 22620 17560
rect 22380 17440 22620 17490
rect 22380 17370 22430 17440
rect 22430 17370 22500 17440
rect 22500 17370 22550 17440
rect 22550 17370 22620 17440
rect 22710 17560 22950 17610
rect 22710 17490 22760 17560
rect 22760 17490 22830 17560
rect 22830 17490 22880 17560
rect 22880 17490 22950 17560
rect 22710 17440 22950 17490
rect 22710 17370 22760 17440
rect 22760 17370 22830 17440
rect 22830 17370 22880 17440
rect 22880 17370 22950 17440
rect 23040 17560 23280 17610
rect 23040 17490 23090 17560
rect 23090 17490 23160 17560
rect 23160 17490 23210 17560
rect 23210 17490 23280 17560
rect 23040 17440 23280 17490
rect 23040 17370 23090 17440
rect 23090 17370 23160 17440
rect 23160 17370 23210 17440
rect 23210 17370 23280 17440
rect 23370 17560 23610 17610
rect 23370 17490 23420 17560
rect 23420 17490 23490 17560
rect 23490 17490 23540 17560
rect 23540 17490 23610 17560
rect 23370 17440 23610 17490
rect 23370 17370 23420 17440
rect 23420 17370 23490 17440
rect 23490 17370 23540 17440
rect 23540 17370 23610 17440
rect 23700 17560 23940 17610
rect 23700 17490 23750 17560
rect 23750 17490 23820 17560
rect 23820 17490 23870 17560
rect 23870 17490 23940 17560
rect 23700 17440 23940 17490
rect 23700 17370 23750 17440
rect 23750 17370 23820 17440
rect 23820 17370 23870 17440
rect 23870 17370 23940 17440
rect 24030 17560 24270 17610
rect 24030 17490 24080 17560
rect 24080 17490 24150 17560
rect 24150 17490 24200 17560
rect 24200 17490 24270 17560
rect 24030 17440 24270 17490
rect 24030 17370 24080 17440
rect 24080 17370 24150 17440
rect 24150 17370 24200 17440
rect 24200 17370 24270 17440
rect 11690 12240 11760 12310
rect 11760 12240 11810 12310
rect 11810 12240 11880 12310
rect 11880 12240 11930 12310
rect 11690 12190 11930 12240
rect 11690 12120 11760 12190
rect 11760 12120 11810 12190
rect 11810 12120 11880 12190
rect 11880 12120 11930 12190
rect 11690 12070 11930 12120
rect 12020 12240 12090 12310
rect 12090 12240 12140 12310
rect 12140 12240 12210 12310
rect 12210 12240 12260 12310
rect 12020 12190 12260 12240
rect 12020 12120 12090 12190
rect 12090 12120 12140 12190
rect 12140 12120 12210 12190
rect 12210 12120 12260 12190
rect 12020 12070 12260 12120
rect 12350 12240 12420 12310
rect 12420 12240 12470 12310
rect 12470 12240 12540 12310
rect 12540 12240 12590 12310
rect 12350 12190 12590 12240
rect 12350 12120 12420 12190
rect 12420 12120 12470 12190
rect 12470 12120 12540 12190
rect 12540 12120 12590 12190
rect 12350 12070 12590 12120
rect 12680 12240 12750 12310
rect 12750 12240 12800 12310
rect 12800 12240 12870 12310
rect 12870 12240 12920 12310
rect 12680 12190 12920 12240
rect 12680 12120 12750 12190
rect 12750 12120 12800 12190
rect 12800 12120 12870 12190
rect 12870 12120 12920 12190
rect 12680 12070 12920 12120
rect 13010 12240 13080 12310
rect 13080 12240 13130 12310
rect 13130 12240 13200 12310
rect 13200 12240 13250 12310
rect 13010 12190 13250 12240
rect 13010 12120 13080 12190
rect 13080 12120 13130 12190
rect 13130 12120 13200 12190
rect 13200 12120 13250 12190
rect 13010 12070 13250 12120
rect 13340 12240 13410 12310
rect 13410 12240 13460 12310
rect 13460 12240 13530 12310
rect 13530 12240 13580 12310
rect 13340 12190 13580 12240
rect 13340 12120 13410 12190
rect 13410 12120 13460 12190
rect 13460 12120 13530 12190
rect 13530 12120 13580 12190
rect 13340 12070 13580 12120
rect 13670 12240 13740 12310
rect 13740 12240 13790 12310
rect 13790 12240 13860 12310
rect 13860 12240 13910 12310
rect 13670 12190 13910 12240
rect 13670 12120 13740 12190
rect 13740 12120 13790 12190
rect 13790 12120 13860 12190
rect 13860 12120 13910 12190
rect 13670 12070 13910 12120
rect 14000 12240 14070 12310
rect 14070 12240 14120 12310
rect 14120 12240 14190 12310
rect 14190 12240 14240 12310
rect 14000 12190 14240 12240
rect 14000 12120 14070 12190
rect 14070 12120 14120 12190
rect 14120 12120 14190 12190
rect 14190 12120 14240 12190
rect 14000 12070 14240 12120
rect 14330 12240 14400 12310
rect 14400 12240 14450 12310
rect 14450 12240 14520 12310
rect 14520 12240 14570 12310
rect 14330 12190 14570 12240
rect 14330 12120 14400 12190
rect 14400 12120 14450 12190
rect 14450 12120 14520 12190
rect 14520 12120 14570 12190
rect 14330 12070 14570 12120
rect 14660 12300 14900 12310
rect 14660 12230 14730 12300
rect 14730 12230 14780 12300
rect 14780 12230 14850 12300
rect 14850 12230 14900 12300
rect 14660 12180 14900 12230
rect 14660 12110 14730 12180
rect 14730 12110 14780 12180
rect 14780 12110 14850 12180
rect 14850 12110 14900 12180
rect 14660 12070 14900 12110
rect 14990 12300 15230 12310
rect 14990 12230 15060 12300
rect 15060 12230 15110 12300
rect 15110 12230 15180 12300
rect 15180 12230 15230 12300
rect 14990 12180 15230 12230
rect 14990 12110 15060 12180
rect 15060 12110 15110 12180
rect 15110 12110 15180 12180
rect 15180 12110 15230 12180
rect 14990 12070 15230 12110
rect 15320 12300 15560 12310
rect 15320 12230 15390 12300
rect 15390 12230 15440 12300
rect 15440 12230 15510 12300
rect 15510 12230 15560 12300
rect 15320 12180 15560 12230
rect 15320 12110 15390 12180
rect 15390 12110 15440 12180
rect 15440 12110 15510 12180
rect 15510 12110 15560 12180
rect 15320 12070 15560 12110
rect 15650 12240 15720 12310
rect 15720 12240 15770 12310
rect 15770 12240 15840 12310
rect 15840 12240 15890 12310
rect 15650 12190 15890 12240
rect 15650 12120 15720 12190
rect 15720 12120 15770 12190
rect 15770 12120 15840 12190
rect 15840 12120 15890 12190
rect 15650 12070 15890 12120
rect 15980 12240 16050 12310
rect 16050 12240 16100 12310
rect 16100 12240 16170 12310
rect 16170 12240 16220 12310
rect 15980 12190 16220 12240
rect 15980 12120 16050 12190
rect 16050 12120 16100 12190
rect 16100 12120 16170 12190
rect 16170 12120 16220 12190
rect 15980 12070 16220 12120
rect 16310 12240 16380 12310
rect 16380 12240 16430 12310
rect 16430 12240 16500 12310
rect 16500 12240 16550 12310
rect 16310 12190 16550 12240
rect 16310 12120 16380 12190
rect 16380 12120 16430 12190
rect 16430 12120 16500 12190
rect 16500 12120 16550 12190
rect 16310 12070 16550 12120
rect 16640 12240 16710 12310
rect 16710 12240 16760 12310
rect 16760 12240 16830 12310
rect 16830 12240 16880 12310
rect 16640 12190 16880 12240
rect 16640 12120 16710 12190
rect 16710 12120 16760 12190
rect 16760 12120 16830 12190
rect 16830 12120 16880 12190
rect 16640 12070 16880 12120
rect 19080 12240 19130 12310
rect 19130 12240 19200 12310
rect 19200 12240 19250 12310
rect 19250 12240 19320 12310
rect 19080 12190 19320 12240
rect 19080 12120 19130 12190
rect 19130 12120 19200 12190
rect 19200 12120 19250 12190
rect 19250 12120 19320 12190
rect 19080 12070 19320 12120
rect 19410 12240 19460 12310
rect 19460 12240 19530 12310
rect 19530 12240 19580 12310
rect 19580 12240 19650 12310
rect 19410 12190 19650 12240
rect 19410 12120 19460 12190
rect 19460 12120 19530 12190
rect 19530 12120 19580 12190
rect 19580 12120 19650 12190
rect 19410 12070 19650 12120
rect 19740 12240 19790 12310
rect 19790 12240 19860 12310
rect 19860 12240 19910 12310
rect 19910 12240 19980 12310
rect 19740 12190 19980 12240
rect 19740 12120 19790 12190
rect 19790 12120 19860 12190
rect 19860 12120 19910 12190
rect 19910 12120 19980 12190
rect 19740 12070 19980 12120
rect 20070 12240 20120 12310
rect 20120 12240 20190 12310
rect 20190 12240 20240 12310
rect 20240 12240 20310 12310
rect 20070 12190 20310 12240
rect 20070 12120 20120 12190
rect 20120 12120 20190 12190
rect 20190 12120 20240 12190
rect 20240 12120 20310 12190
rect 20070 12070 20310 12120
rect 20400 12300 20640 12310
rect 20400 12230 20450 12300
rect 20450 12230 20520 12300
rect 20520 12230 20570 12300
rect 20570 12230 20640 12300
rect 20400 12180 20640 12230
rect 20400 12110 20450 12180
rect 20450 12110 20520 12180
rect 20520 12110 20570 12180
rect 20570 12110 20640 12180
rect 20400 12070 20640 12110
rect 20730 12300 20970 12310
rect 20730 12230 20780 12300
rect 20780 12230 20850 12300
rect 20850 12230 20900 12300
rect 20900 12230 20970 12300
rect 20730 12180 20970 12230
rect 20730 12110 20780 12180
rect 20780 12110 20850 12180
rect 20850 12110 20900 12180
rect 20900 12110 20970 12180
rect 20730 12070 20970 12110
rect 21060 12300 21300 12310
rect 21060 12230 21110 12300
rect 21110 12230 21180 12300
rect 21180 12230 21230 12300
rect 21230 12230 21300 12300
rect 21060 12180 21300 12230
rect 21060 12110 21110 12180
rect 21110 12110 21180 12180
rect 21180 12110 21230 12180
rect 21230 12110 21300 12180
rect 21060 12070 21300 12110
rect 21390 12240 21440 12310
rect 21440 12240 21510 12310
rect 21510 12240 21560 12310
rect 21560 12240 21630 12310
rect 21390 12190 21630 12240
rect 21390 12120 21440 12190
rect 21440 12120 21510 12190
rect 21510 12120 21560 12190
rect 21560 12120 21630 12190
rect 21390 12070 21630 12120
rect 21720 12240 21770 12310
rect 21770 12240 21840 12310
rect 21840 12240 21890 12310
rect 21890 12240 21960 12310
rect 21720 12190 21960 12240
rect 21720 12120 21770 12190
rect 21770 12120 21840 12190
rect 21840 12120 21890 12190
rect 21890 12120 21960 12190
rect 21720 12070 21960 12120
rect 22050 12240 22100 12310
rect 22100 12240 22170 12310
rect 22170 12240 22220 12310
rect 22220 12240 22290 12310
rect 22050 12190 22290 12240
rect 22050 12120 22100 12190
rect 22100 12120 22170 12190
rect 22170 12120 22220 12190
rect 22220 12120 22290 12190
rect 22050 12070 22290 12120
rect 22380 12240 22430 12310
rect 22430 12240 22500 12310
rect 22500 12240 22550 12310
rect 22550 12240 22620 12310
rect 22380 12190 22620 12240
rect 22380 12120 22430 12190
rect 22430 12120 22500 12190
rect 22500 12120 22550 12190
rect 22550 12120 22620 12190
rect 22380 12070 22620 12120
rect 22710 12240 22760 12310
rect 22760 12240 22830 12310
rect 22830 12240 22880 12310
rect 22880 12240 22950 12310
rect 22710 12190 22950 12240
rect 22710 12120 22760 12190
rect 22760 12120 22830 12190
rect 22830 12120 22880 12190
rect 22880 12120 22950 12190
rect 22710 12070 22950 12120
rect 23040 12240 23090 12310
rect 23090 12240 23160 12310
rect 23160 12240 23210 12310
rect 23210 12240 23280 12310
rect 23040 12190 23280 12240
rect 23040 12120 23090 12190
rect 23090 12120 23160 12190
rect 23160 12120 23210 12190
rect 23210 12120 23280 12190
rect 23040 12070 23280 12120
rect 23370 12240 23420 12310
rect 23420 12240 23490 12310
rect 23490 12240 23540 12310
rect 23540 12240 23610 12310
rect 23370 12190 23610 12240
rect 23370 12120 23420 12190
rect 23420 12120 23490 12190
rect 23490 12120 23540 12190
rect 23540 12120 23610 12190
rect 23370 12070 23610 12120
rect 23700 12240 23750 12310
rect 23750 12240 23820 12310
rect 23820 12240 23870 12310
rect 23870 12240 23940 12310
rect 23700 12190 23940 12240
rect 23700 12120 23750 12190
rect 23750 12120 23820 12190
rect 23820 12120 23870 12190
rect 23870 12120 23940 12190
rect 23700 12070 23940 12120
rect 24030 12240 24080 12310
rect 24080 12240 24150 12310
rect 24150 12240 24200 12310
rect 24200 12240 24270 12310
rect 24030 12190 24270 12240
rect 24030 12120 24080 12190
rect 24080 12120 24150 12190
rect 24150 12120 24200 12190
rect 24200 12120 24270 12190
rect 24030 12070 24270 12120
<< metal5 >>
rect 11660 17610 24300 17660
rect 11660 17370 11690 17610
rect 11930 17370 12020 17610
rect 12260 17370 12350 17610
rect 12590 17370 12680 17610
rect 12920 17370 13010 17610
rect 13250 17370 13340 17610
rect 13580 17370 13670 17610
rect 13910 17370 14000 17610
rect 14240 17370 14330 17610
rect 14570 17370 14660 17610
rect 14900 17370 14990 17610
rect 15230 17370 15320 17610
rect 15560 17370 15650 17610
rect 15890 17370 15980 17610
rect 16220 17370 16310 17610
rect 16550 17370 16640 17610
rect 16880 17370 19080 17610
rect 19320 17370 19410 17610
rect 19650 17370 19740 17610
rect 19980 17370 20070 17610
rect 20310 17370 20400 17610
rect 20640 17370 20730 17610
rect 20970 17370 21060 17610
rect 21300 17370 21390 17610
rect 21630 17370 21720 17610
rect 21960 17370 22050 17610
rect 22290 17370 22380 17610
rect 22620 17370 22710 17610
rect 22950 17370 23040 17610
rect 23280 17370 23370 17610
rect 23610 17370 23700 17610
rect 23940 17370 24030 17610
rect 24270 17370 24300 17610
rect 11660 17340 24300 17370
rect 11660 12310 24300 12340
rect 11660 12070 11690 12310
rect 11930 12070 12020 12310
rect 12260 12070 12350 12310
rect 12590 12070 12680 12310
rect 12920 12070 13010 12310
rect 13250 12070 13340 12310
rect 13580 12070 13670 12310
rect 13910 12070 14000 12310
rect 14240 12070 14330 12310
rect 14570 12070 14660 12310
rect 14900 12070 14990 12310
rect 15230 12070 15320 12310
rect 15560 12070 15650 12310
rect 15890 12070 15980 12310
rect 16220 12070 16310 12310
rect 16550 12070 16640 12310
rect 16880 12070 19080 12310
rect 19320 12070 19410 12310
rect 19650 12070 19740 12310
rect 19980 12070 20070 12310
rect 20310 12070 20400 12310
rect 20640 12070 20730 12310
rect 20970 12070 21060 12310
rect 21300 12070 21390 12310
rect 21630 12070 21720 12310
rect 21960 12070 22050 12310
rect 22290 12070 22380 12310
rect 22620 12070 22710 12310
rect 22950 12070 23040 12310
rect 23280 12070 23370 12310
rect 23610 12070 23700 12310
rect 23940 12070 24030 12310
rect 24270 12070 24300 12310
rect 11660 12020 24300 12070
<< comment >>
rect 11570 16320 11630 16350
rect 24330 16320 24390 16350
rect 11570 13350 11630 13380
rect 24330 13350 24390 13380
<< labels >>
rlabel metal4 17450 11600 17450 11600 1 out
port 1 n
rlabel metal4 17450 18150 17450 18150 1 in
port 2 n
rlabel metal5 16990 17630 16990 17630 1 VDD
port 3 n
rlabel metal5 17090 12040 17090 12040 1 GND
port 4 n
<< end >>
